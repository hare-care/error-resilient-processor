magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< dnwell >>
rect 626 9736 14336 36182
<< nwell >>
rect 517 35918 14447 36293
rect 517 10000 832 35918
rect 1593 30774 13423 31518
rect 1593 27622 2336 30774
rect 12680 27622 13423 30774
rect 1593 26878 13423 27622
rect 14072 10000 14447 35918
rect 517 9625 14447 10000
<< pwell >>
rect 219 36363 14750 36600
rect 219 9554 456 36363
rect 1122 34548 13870 34720
rect 1122 10388 1294 34548
rect 13698 10388 13870 34548
rect 1122 10216 13870 10388
rect 14513 9554 14750 36363
rect 219 9317 14750 9554
<< mvpsubdiff >>
rect 245 36498 14724 36574
rect 245 36464 532 36498
rect 566 36464 600 36498
rect 634 36464 668 36498
rect 702 36464 736 36498
rect 770 36464 804 36498
rect 838 36464 872 36498
rect 906 36464 940 36498
rect 974 36464 1008 36498
rect 1042 36464 1076 36498
rect 1110 36464 1144 36498
rect 1178 36464 1212 36498
rect 1246 36464 1280 36498
rect 1314 36464 1348 36498
rect 1382 36464 1416 36498
rect 1450 36464 1484 36498
rect 1518 36464 1552 36498
rect 1586 36464 1620 36498
rect 1654 36464 1688 36498
rect 1722 36464 1756 36498
rect 1790 36464 1824 36498
rect 1858 36464 1892 36498
rect 1926 36464 1960 36498
rect 1994 36464 2028 36498
rect 2062 36464 2096 36498
rect 2130 36464 2164 36498
rect 2198 36464 2232 36498
rect 2266 36464 2300 36498
rect 2334 36464 2368 36498
rect 2402 36464 2436 36498
rect 2470 36464 2504 36498
rect 2538 36464 2572 36498
rect 2606 36464 2640 36498
rect 2674 36464 2708 36498
rect 2742 36464 2776 36498
rect 2810 36464 2844 36498
rect 2878 36464 2912 36498
rect 2946 36464 2980 36498
rect 3014 36464 3048 36498
rect 3082 36464 3116 36498
rect 3150 36464 3184 36498
rect 3218 36464 3252 36498
rect 3286 36464 3320 36498
rect 3354 36464 3388 36498
rect 3422 36464 3456 36498
rect 3490 36464 3524 36498
rect 3558 36464 3592 36498
rect 3626 36464 3660 36498
rect 3694 36464 3728 36498
rect 3762 36464 3796 36498
rect 3830 36464 3864 36498
rect 3898 36464 3932 36498
rect 3966 36464 4000 36498
rect 4034 36464 4068 36498
rect 4102 36464 4136 36498
rect 4170 36464 4204 36498
rect 4238 36464 4272 36498
rect 4306 36464 4340 36498
rect 4374 36464 4408 36498
rect 4442 36464 4476 36498
rect 4510 36464 4544 36498
rect 4578 36464 4612 36498
rect 4646 36464 4680 36498
rect 4714 36464 4748 36498
rect 4782 36464 4816 36498
rect 4850 36464 4884 36498
rect 4918 36464 4952 36498
rect 4986 36464 5020 36498
rect 5054 36464 5088 36498
rect 5122 36464 5156 36498
rect 5190 36464 5224 36498
rect 5258 36464 5292 36498
rect 5326 36464 5360 36498
rect 5394 36464 5428 36498
rect 5462 36464 5496 36498
rect 5530 36464 5564 36498
rect 5598 36464 5632 36498
rect 5666 36464 5700 36498
rect 5734 36464 5768 36498
rect 5802 36464 5836 36498
rect 5870 36464 5904 36498
rect 5938 36464 5972 36498
rect 6006 36464 6040 36498
rect 6074 36464 6108 36498
rect 6142 36464 6176 36498
rect 6210 36464 6244 36498
rect 6278 36464 6312 36498
rect 6346 36464 6380 36498
rect 6414 36464 6448 36498
rect 6482 36464 6516 36498
rect 6550 36464 6584 36498
rect 6618 36464 6652 36498
rect 6686 36464 6720 36498
rect 6754 36464 6788 36498
rect 6822 36464 6856 36498
rect 6890 36464 6924 36498
rect 6958 36464 6992 36498
rect 7026 36464 7060 36498
rect 7094 36464 7128 36498
rect 7162 36464 7196 36498
rect 7230 36464 7264 36498
rect 7298 36464 7332 36498
rect 7366 36464 7400 36498
rect 7434 36464 7468 36498
rect 7502 36464 7536 36498
rect 7570 36464 7604 36498
rect 7638 36464 7672 36498
rect 7706 36464 7740 36498
rect 7774 36464 7808 36498
rect 7842 36464 7876 36498
rect 7910 36464 7944 36498
rect 7978 36464 8012 36498
rect 8046 36464 8080 36498
rect 8114 36464 8148 36498
rect 8182 36464 8216 36498
rect 8250 36464 8284 36498
rect 8318 36464 8352 36498
rect 8386 36464 8420 36498
rect 8454 36464 8488 36498
rect 8522 36464 8556 36498
rect 8590 36464 8624 36498
rect 8658 36464 8692 36498
rect 8726 36464 8760 36498
rect 8794 36464 8828 36498
rect 8862 36464 8896 36498
rect 8930 36464 8964 36498
rect 8998 36464 9032 36498
rect 9066 36464 9100 36498
rect 9134 36464 9168 36498
rect 9202 36464 9236 36498
rect 9270 36464 9304 36498
rect 9338 36464 9372 36498
rect 9406 36464 9440 36498
rect 9474 36464 9508 36498
rect 9542 36464 9576 36498
rect 9610 36464 9644 36498
rect 9678 36464 9712 36498
rect 9746 36464 9780 36498
rect 9814 36464 9848 36498
rect 9882 36464 9916 36498
rect 9950 36464 9984 36498
rect 10018 36464 10052 36498
rect 10086 36464 10120 36498
rect 10154 36464 10188 36498
rect 10222 36464 10256 36498
rect 10290 36464 10324 36498
rect 10358 36464 10392 36498
rect 10426 36464 10460 36498
rect 10494 36464 10528 36498
rect 10562 36464 10596 36498
rect 10630 36464 10664 36498
rect 10698 36464 10732 36498
rect 10766 36464 10800 36498
rect 10834 36464 10868 36498
rect 10902 36464 10936 36498
rect 10970 36464 11004 36498
rect 11038 36464 11072 36498
rect 11106 36464 11140 36498
rect 11174 36464 11208 36498
rect 11242 36464 11276 36498
rect 11310 36464 11344 36498
rect 11378 36464 11412 36498
rect 11446 36464 11480 36498
rect 11514 36464 11548 36498
rect 11582 36464 11616 36498
rect 11650 36464 11684 36498
rect 11718 36464 11752 36498
rect 11786 36464 11820 36498
rect 11854 36464 11888 36498
rect 11922 36464 11956 36498
rect 11990 36464 12024 36498
rect 12058 36464 12092 36498
rect 12126 36464 12160 36498
rect 12194 36464 12228 36498
rect 12262 36464 12296 36498
rect 12330 36464 12364 36498
rect 12398 36464 12432 36498
rect 12466 36464 12500 36498
rect 12534 36464 12568 36498
rect 12602 36464 12636 36498
rect 12670 36464 12704 36498
rect 12738 36464 12772 36498
rect 12806 36464 12840 36498
rect 12874 36464 12908 36498
rect 12942 36464 12976 36498
rect 13010 36464 13044 36498
rect 13078 36464 13112 36498
rect 13146 36464 13180 36498
rect 13214 36464 13248 36498
rect 13282 36464 13316 36498
rect 13350 36464 13384 36498
rect 13418 36464 13452 36498
rect 13486 36464 13520 36498
rect 13554 36464 13588 36498
rect 13622 36464 13656 36498
rect 13690 36464 13724 36498
rect 13758 36464 13792 36498
rect 13826 36464 13860 36498
rect 13894 36464 13928 36498
rect 13962 36464 13996 36498
rect 14030 36464 14064 36498
rect 14098 36464 14132 36498
rect 14166 36464 14200 36498
rect 14234 36464 14268 36498
rect 14302 36464 14336 36498
rect 14370 36464 14404 36498
rect 14438 36464 14472 36498
rect 14506 36464 14724 36498
rect 245 36389 14724 36464
rect 245 36311 430 36389
rect 245 36277 317 36311
rect 351 36277 430 36311
rect 245 36243 430 36277
rect 245 36209 317 36243
rect 351 36209 430 36243
rect 14539 36309 14724 36389
rect 14539 36275 14611 36309
rect 14645 36275 14724 36309
rect 14539 36241 14724 36275
rect 245 36175 430 36209
rect 245 36141 317 36175
rect 351 36141 430 36175
rect 245 36107 430 36141
rect 245 36073 317 36107
rect 351 36073 430 36107
rect 245 36039 430 36073
rect 245 36005 317 36039
rect 351 36005 430 36039
rect 245 35971 430 36005
rect 245 35937 317 35971
rect 351 35937 430 35971
rect 245 35903 430 35937
rect 245 35869 317 35903
rect 351 35869 430 35903
rect 245 35835 430 35869
rect 245 35801 317 35835
rect 351 35801 430 35835
rect 245 35767 430 35801
rect 245 35733 317 35767
rect 351 35733 430 35767
rect 245 35699 430 35733
rect 245 35665 317 35699
rect 351 35665 430 35699
rect 245 35631 430 35665
rect 245 35597 317 35631
rect 351 35597 430 35631
rect 245 35563 430 35597
rect 245 35529 317 35563
rect 351 35529 430 35563
rect 245 35495 430 35529
rect 245 35461 317 35495
rect 351 35461 430 35495
rect 245 35427 430 35461
rect 245 35393 317 35427
rect 351 35393 430 35427
rect 245 35359 430 35393
rect 245 35325 317 35359
rect 351 35325 430 35359
rect 245 35291 430 35325
rect 245 35257 317 35291
rect 351 35257 430 35291
rect 245 35223 430 35257
rect 245 35189 317 35223
rect 351 35189 430 35223
rect 245 35155 430 35189
rect 245 35121 317 35155
rect 351 35121 430 35155
rect 245 35087 430 35121
rect 245 35053 317 35087
rect 351 35053 430 35087
rect 245 35019 430 35053
rect 245 34985 317 35019
rect 351 34985 430 35019
rect 245 34951 430 34985
rect 245 34917 317 34951
rect 351 34917 430 34951
rect 245 34883 430 34917
rect 245 34849 317 34883
rect 351 34849 430 34883
rect 245 34815 430 34849
rect 245 34781 317 34815
rect 351 34781 430 34815
rect 245 34747 430 34781
rect 245 34713 317 34747
rect 351 34713 430 34747
rect 245 34679 430 34713
rect 245 34645 317 34679
rect 351 34645 430 34679
rect 245 34611 430 34645
rect 245 34577 317 34611
rect 351 34577 430 34611
rect 245 34543 430 34577
rect 245 34509 317 34543
rect 351 34509 430 34543
rect 245 34475 430 34509
rect 245 34441 317 34475
rect 351 34441 430 34475
rect 245 34407 430 34441
rect 245 34373 317 34407
rect 351 34373 430 34407
rect 245 34339 430 34373
rect 245 34305 317 34339
rect 351 34305 430 34339
rect 245 34271 430 34305
rect 245 34237 317 34271
rect 351 34237 430 34271
rect 245 34203 430 34237
rect 245 34169 317 34203
rect 351 34169 430 34203
rect 245 34135 430 34169
rect 245 34101 317 34135
rect 351 34101 430 34135
rect 245 34067 430 34101
rect 245 34033 317 34067
rect 351 34033 430 34067
rect 245 33999 430 34033
rect 245 33965 317 33999
rect 351 33965 430 33999
rect 245 33931 430 33965
rect 245 33897 317 33931
rect 351 33897 430 33931
rect 245 33863 430 33897
rect 245 33829 317 33863
rect 351 33829 430 33863
rect 245 33795 430 33829
rect 245 33761 317 33795
rect 351 33761 430 33795
rect 245 33727 430 33761
rect 245 33693 317 33727
rect 351 33693 430 33727
rect 245 33659 430 33693
rect 245 33625 317 33659
rect 351 33625 430 33659
rect 245 33591 430 33625
rect 245 33557 317 33591
rect 351 33557 430 33591
rect 245 33523 430 33557
rect 245 33489 317 33523
rect 351 33489 430 33523
rect 245 33455 430 33489
rect 245 33421 317 33455
rect 351 33421 430 33455
rect 245 33387 430 33421
rect 245 33353 317 33387
rect 351 33353 430 33387
rect 245 33319 430 33353
rect 245 33285 317 33319
rect 351 33285 430 33319
rect 245 33251 430 33285
rect 245 33217 317 33251
rect 351 33217 430 33251
rect 245 33183 430 33217
rect 245 33149 317 33183
rect 351 33149 430 33183
rect 245 33115 430 33149
rect 245 33081 317 33115
rect 351 33081 430 33115
rect 245 33047 430 33081
rect 245 33013 317 33047
rect 351 33013 430 33047
rect 245 32979 430 33013
rect 245 32945 317 32979
rect 351 32945 430 32979
rect 245 32911 430 32945
rect 245 32877 317 32911
rect 351 32877 430 32911
rect 245 32843 430 32877
rect 245 32809 317 32843
rect 351 32809 430 32843
rect 245 32775 430 32809
rect 245 32741 317 32775
rect 351 32741 430 32775
rect 245 32707 430 32741
rect 245 32673 317 32707
rect 351 32673 430 32707
rect 245 32639 430 32673
rect 245 32605 317 32639
rect 351 32605 430 32639
rect 245 32571 430 32605
rect 245 32537 317 32571
rect 351 32537 430 32571
rect 245 32503 430 32537
rect 245 32469 317 32503
rect 351 32469 430 32503
rect 245 32435 430 32469
rect 245 32401 317 32435
rect 351 32401 430 32435
rect 245 32367 430 32401
rect 245 32333 317 32367
rect 351 32333 430 32367
rect 245 32299 430 32333
rect 245 32265 317 32299
rect 351 32265 430 32299
rect 245 32231 430 32265
rect 245 32197 317 32231
rect 351 32197 430 32231
rect 245 32163 430 32197
rect 245 32129 317 32163
rect 351 32129 430 32163
rect 245 32095 430 32129
rect 245 32061 317 32095
rect 351 32061 430 32095
rect 245 32027 430 32061
rect 245 31993 317 32027
rect 351 31993 430 32027
rect 245 31959 430 31993
rect 245 31925 317 31959
rect 351 31925 430 31959
rect 245 31891 430 31925
rect 245 31857 317 31891
rect 351 31857 430 31891
rect 245 31823 430 31857
rect 245 31789 317 31823
rect 351 31789 430 31823
rect 245 31755 430 31789
rect 245 31721 317 31755
rect 351 31721 430 31755
rect 245 31687 430 31721
rect 245 31653 317 31687
rect 351 31653 430 31687
rect 245 31619 430 31653
rect 245 31585 317 31619
rect 351 31585 430 31619
rect 245 31551 430 31585
rect 245 31517 317 31551
rect 351 31517 430 31551
rect 245 31483 430 31517
rect 245 31449 317 31483
rect 351 31449 430 31483
rect 245 31415 430 31449
rect 245 31381 317 31415
rect 351 31381 430 31415
rect 245 31347 430 31381
rect 245 31313 317 31347
rect 351 31313 430 31347
rect 245 31279 430 31313
rect 245 31245 317 31279
rect 351 31245 430 31279
rect 245 31211 430 31245
rect 245 31177 317 31211
rect 351 31177 430 31211
rect 245 31143 430 31177
rect 245 31109 317 31143
rect 351 31109 430 31143
rect 245 31075 430 31109
rect 245 31041 317 31075
rect 351 31041 430 31075
rect 245 31007 430 31041
rect 245 30973 317 31007
rect 351 30973 430 31007
rect 245 30939 430 30973
rect 245 30905 317 30939
rect 351 30905 430 30939
rect 245 30871 430 30905
rect 245 30837 317 30871
rect 351 30837 430 30871
rect 245 30803 430 30837
rect 245 30769 317 30803
rect 351 30769 430 30803
rect 245 30735 430 30769
rect 245 30701 317 30735
rect 351 30701 430 30735
rect 245 30667 430 30701
rect 245 30633 317 30667
rect 351 30633 430 30667
rect 245 30599 430 30633
rect 245 30565 317 30599
rect 351 30565 430 30599
rect 245 30531 430 30565
rect 245 30497 317 30531
rect 351 30497 430 30531
rect 245 30463 430 30497
rect 245 30429 317 30463
rect 351 30429 430 30463
rect 245 30395 430 30429
rect 245 30361 317 30395
rect 351 30361 430 30395
rect 245 30327 430 30361
rect 245 30293 317 30327
rect 351 30293 430 30327
rect 245 30259 430 30293
rect 245 30225 317 30259
rect 351 30225 430 30259
rect 245 30191 430 30225
rect 245 30157 317 30191
rect 351 30157 430 30191
rect 245 30123 430 30157
rect 245 30089 317 30123
rect 351 30089 430 30123
rect 245 30055 430 30089
rect 245 30021 317 30055
rect 351 30021 430 30055
rect 245 29987 430 30021
rect 245 29953 317 29987
rect 351 29953 430 29987
rect 245 29919 430 29953
rect 245 29885 317 29919
rect 351 29885 430 29919
rect 245 29851 430 29885
rect 245 29817 317 29851
rect 351 29817 430 29851
rect 245 29783 430 29817
rect 245 29749 317 29783
rect 351 29749 430 29783
rect 245 29715 430 29749
rect 245 29681 317 29715
rect 351 29681 430 29715
rect 245 29647 430 29681
rect 245 29613 317 29647
rect 351 29613 430 29647
rect 245 29579 430 29613
rect 245 29545 317 29579
rect 351 29545 430 29579
rect 245 29511 430 29545
rect 245 29477 317 29511
rect 351 29477 430 29511
rect 245 29443 430 29477
rect 245 29409 317 29443
rect 351 29409 430 29443
rect 245 29375 430 29409
rect 245 29341 317 29375
rect 351 29341 430 29375
rect 245 29307 430 29341
rect 245 29273 317 29307
rect 351 29273 430 29307
rect 245 29239 430 29273
rect 245 29205 317 29239
rect 351 29205 430 29239
rect 245 29171 430 29205
rect 245 29137 317 29171
rect 351 29137 430 29171
rect 245 29103 430 29137
rect 245 29069 317 29103
rect 351 29069 430 29103
rect 245 29035 430 29069
rect 245 29001 317 29035
rect 351 29001 430 29035
rect 245 28967 430 29001
rect 245 28933 317 28967
rect 351 28933 430 28967
rect 245 28899 430 28933
rect 245 28865 317 28899
rect 351 28865 430 28899
rect 245 28831 430 28865
rect 245 28797 317 28831
rect 351 28797 430 28831
rect 245 28763 430 28797
rect 245 28729 317 28763
rect 351 28729 430 28763
rect 245 28695 430 28729
rect 245 28661 317 28695
rect 351 28661 430 28695
rect 245 28627 430 28661
rect 245 28593 317 28627
rect 351 28593 430 28627
rect 245 28559 430 28593
rect 245 28525 317 28559
rect 351 28525 430 28559
rect 245 28491 430 28525
rect 245 28457 317 28491
rect 351 28457 430 28491
rect 245 28423 430 28457
rect 245 28389 317 28423
rect 351 28389 430 28423
rect 245 28355 430 28389
rect 245 28321 317 28355
rect 351 28321 430 28355
rect 245 28287 430 28321
rect 245 28253 317 28287
rect 351 28253 430 28287
rect 245 28219 430 28253
rect 245 28185 317 28219
rect 351 28185 430 28219
rect 245 28151 430 28185
rect 245 28117 317 28151
rect 351 28117 430 28151
rect 245 28083 430 28117
rect 245 28049 317 28083
rect 351 28049 430 28083
rect 245 28015 430 28049
rect 245 27981 317 28015
rect 351 27981 430 28015
rect 245 27947 430 27981
rect 245 27913 317 27947
rect 351 27913 430 27947
rect 245 27879 430 27913
rect 245 27845 317 27879
rect 351 27845 430 27879
rect 245 27811 430 27845
rect 245 27777 317 27811
rect 351 27777 430 27811
rect 245 27743 430 27777
rect 245 27709 317 27743
rect 351 27709 430 27743
rect 245 27675 430 27709
rect 245 27641 317 27675
rect 351 27641 430 27675
rect 245 27607 430 27641
rect 245 27573 317 27607
rect 351 27573 430 27607
rect 245 27539 430 27573
rect 245 27505 317 27539
rect 351 27505 430 27539
rect 245 27471 430 27505
rect 245 27437 317 27471
rect 351 27437 430 27471
rect 245 27403 430 27437
rect 245 27369 317 27403
rect 351 27369 430 27403
rect 245 27335 430 27369
rect 245 27301 317 27335
rect 351 27301 430 27335
rect 245 27267 430 27301
rect 245 27233 317 27267
rect 351 27233 430 27267
rect 245 27199 430 27233
rect 245 27165 317 27199
rect 351 27165 430 27199
rect 245 27131 430 27165
rect 245 27097 317 27131
rect 351 27097 430 27131
rect 245 27063 430 27097
rect 245 27029 317 27063
rect 351 27029 430 27063
rect 245 26995 430 27029
rect 245 26961 317 26995
rect 351 26961 430 26995
rect 245 26927 430 26961
rect 245 26893 317 26927
rect 351 26893 430 26927
rect 245 26859 430 26893
rect 245 26825 317 26859
rect 351 26825 430 26859
rect 245 26791 430 26825
rect 245 26757 317 26791
rect 351 26757 430 26791
rect 245 26723 430 26757
rect 245 26689 317 26723
rect 351 26689 430 26723
rect 245 26655 430 26689
rect 245 26621 317 26655
rect 351 26621 430 26655
rect 245 26587 430 26621
rect 245 26553 317 26587
rect 351 26553 430 26587
rect 245 26519 430 26553
rect 245 26485 317 26519
rect 351 26485 430 26519
rect 245 26451 430 26485
rect 245 26417 317 26451
rect 351 26417 430 26451
rect 245 26383 430 26417
rect 245 26349 317 26383
rect 351 26349 430 26383
rect 245 26315 430 26349
rect 245 26281 317 26315
rect 351 26281 430 26315
rect 245 26247 430 26281
rect 245 26213 317 26247
rect 351 26213 430 26247
rect 245 26179 430 26213
rect 245 26145 317 26179
rect 351 26145 430 26179
rect 245 26111 430 26145
rect 245 26077 317 26111
rect 351 26077 430 26111
rect 245 26043 430 26077
rect 245 26009 317 26043
rect 351 26009 430 26043
rect 245 25975 430 26009
rect 245 25941 317 25975
rect 351 25941 430 25975
rect 245 25907 430 25941
rect 245 25873 317 25907
rect 351 25873 430 25907
rect 245 25839 430 25873
rect 245 25805 317 25839
rect 351 25805 430 25839
rect 245 25771 430 25805
rect 245 25737 317 25771
rect 351 25737 430 25771
rect 245 25703 430 25737
rect 245 25669 317 25703
rect 351 25669 430 25703
rect 245 25635 430 25669
rect 245 25601 317 25635
rect 351 25601 430 25635
rect 245 25567 430 25601
rect 245 25533 317 25567
rect 351 25533 430 25567
rect 245 25499 430 25533
rect 245 25465 317 25499
rect 351 25465 430 25499
rect 245 25431 430 25465
rect 245 25397 317 25431
rect 351 25397 430 25431
rect 245 25363 430 25397
rect 245 25329 317 25363
rect 351 25329 430 25363
rect 245 25295 430 25329
rect 245 25261 317 25295
rect 351 25261 430 25295
rect 245 25227 430 25261
rect 245 25193 317 25227
rect 351 25193 430 25227
rect 245 25159 430 25193
rect 245 25125 317 25159
rect 351 25125 430 25159
rect 245 25091 430 25125
rect 245 25057 317 25091
rect 351 25057 430 25091
rect 245 25023 430 25057
rect 245 24989 317 25023
rect 351 24989 430 25023
rect 245 24955 430 24989
rect 245 24921 317 24955
rect 351 24921 430 24955
rect 245 24887 430 24921
rect 245 24853 317 24887
rect 351 24853 430 24887
rect 245 24819 430 24853
rect 245 24785 317 24819
rect 351 24785 430 24819
rect 245 24751 430 24785
rect 245 24717 317 24751
rect 351 24717 430 24751
rect 245 24683 430 24717
rect 245 24649 317 24683
rect 351 24649 430 24683
rect 245 24615 430 24649
rect 245 24581 317 24615
rect 351 24581 430 24615
rect 245 24547 430 24581
rect 245 24513 317 24547
rect 351 24513 430 24547
rect 245 24479 430 24513
rect 245 24445 317 24479
rect 351 24445 430 24479
rect 245 24411 430 24445
rect 245 24377 317 24411
rect 351 24377 430 24411
rect 245 24343 430 24377
rect 245 24309 317 24343
rect 351 24309 430 24343
rect 245 24275 430 24309
rect 245 24241 317 24275
rect 351 24241 430 24275
rect 245 24207 430 24241
rect 245 24173 317 24207
rect 351 24173 430 24207
rect 245 24139 430 24173
rect 245 24105 317 24139
rect 351 24105 430 24139
rect 245 24071 430 24105
rect 245 24037 317 24071
rect 351 24037 430 24071
rect 245 24003 430 24037
rect 245 23969 317 24003
rect 351 23969 430 24003
rect 245 23935 430 23969
rect 245 23901 317 23935
rect 351 23901 430 23935
rect 245 23867 430 23901
rect 245 23833 317 23867
rect 351 23833 430 23867
rect 245 23799 430 23833
rect 245 23765 317 23799
rect 351 23765 430 23799
rect 245 23731 430 23765
rect 245 23697 317 23731
rect 351 23697 430 23731
rect 245 23663 430 23697
rect 245 23629 317 23663
rect 351 23629 430 23663
rect 245 23595 430 23629
rect 245 23561 317 23595
rect 351 23561 430 23595
rect 245 23527 430 23561
rect 245 23493 317 23527
rect 351 23493 430 23527
rect 245 23459 430 23493
rect 245 23425 317 23459
rect 351 23425 430 23459
rect 245 23391 430 23425
rect 245 23357 317 23391
rect 351 23357 430 23391
rect 245 23323 430 23357
rect 245 23289 317 23323
rect 351 23289 430 23323
rect 245 23255 430 23289
rect 245 23221 317 23255
rect 351 23221 430 23255
rect 245 23187 430 23221
rect 245 23153 317 23187
rect 351 23153 430 23187
rect 245 23119 430 23153
rect 245 23085 317 23119
rect 351 23085 430 23119
rect 245 23051 430 23085
rect 245 23017 317 23051
rect 351 23017 430 23051
rect 245 22983 430 23017
rect 245 22949 317 22983
rect 351 22949 430 22983
rect 245 22915 430 22949
rect 245 22881 317 22915
rect 351 22881 430 22915
rect 245 22847 430 22881
rect 245 22813 317 22847
rect 351 22813 430 22847
rect 245 22779 430 22813
rect 245 22745 317 22779
rect 351 22745 430 22779
rect 245 22711 430 22745
rect 245 22677 317 22711
rect 351 22677 430 22711
rect 245 22643 430 22677
rect 245 22609 317 22643
rect 351 22609 430 22643
rect 245 22575 430 22609
rect 245 22541 317 22575
rect 351 22541 430 22575
rect 245 22507 430 22541
rect 245 22473 317 22507
rect 351 22473 430 22507
rect 245 22439 430 22473
rect 245 22405 317 22439
rect 351 22405 430 22439
rect 245 22371 430 22405
rect 245 22337 317 22371
rect 351 22337 430 22371
rect 245 22303 430 22337
rect 245 22269 317 22303
rect 351 22269 430 22303
rect 245 22235 430 22269
rect 245 22201 317 22235
rect 351 22201 430 22235
rect 245 22167 430 22201
rect 245 22133 317 22167
rect 351 22133 430 22167
rect 245 22099 430 22133
rect 245 22065 317 22099
rect 351 22065 430 22099
rect 245 22031 430 22065
rect 245 21997 317 22031
rect 351 21997 430 22031
rect 245 21963 430 21997
rect 245 21929 317 21963
rect 351 21929 430 21963
rect 245 21895 430 21929
rect 245 21861 317 21895
rect 351 21861 430 21895
rect 245 21827 430 21861
rect 245 21793 317 21827
rect 351 21793 430 21827
rect 245 21759 430 21793
rect 245 21725 317 21759
rect 351 21725 430 21759
rect 245 21691 430 21725
rect 245 21657 317 21691
rect 351 21657 430 21691
rect 245 21623 430 21657
rect 245 21589 317 21623
rect 351 21589 430 21623
rect 245 21555 430 21589
rect 245 21521 317 21555
rect 351 21521 430 21555
rect 245 21487 430 21521
rect 245 21453 317 21487
rect 351 21453 430 21487
rect 245 21419 430 21453
rect 245 21385 317 21419
rect 351 21385 430 21419
rect 245 21351 430 21385
rect 245 21317 317 21351
rect 351 21317 430 21351
rect 245 21283 430 21317
rect 245 21249 317 21283
rect 351 21249 430 21283
rect 245 21215 430 21249
rect 245 21181 317 21215
rect 351 21181 430 21215
rect 245 21147 430 21181
rect 245 21113 317 21147
rect 351 21113 430 21147
rect 245 21079 430 21113
rect 245 21045 317 21079
rect 351 21045 430 21079
rect 245 21011 430 21045
rect 245 20977 317 21011
rect 351 20977 430 21011
rect 245 20943 430 20977
rect 245 20909 317 20943
rect 351 20909 430 20943
rect 245 20875 430 20909
rect 245 20841 317 20875
rect 351 20841 430 20875
rect 245 20807 430 20841
rect 245 20773 317 20807
rect 351 20773 430 20807
rect 245 20739 430 20773
rect 245 20705 317 20739
rect 351 20705 430 20739
rect 245 20671 430 20705
rect 245 20637 317 20671
rect 351 20637 430 20671
rect 245 20603 430 20637
rect 245 20569 317 20603
rect 351 20569 430 20603
rect 245 20535 430 20569
rect 245 20501 317 20535
rect 351 20501 430 20535
rect 245 20467 430 20501
rect 245 20433 317 20467
rect 351 20433 430 20467
rect 245 20399 430 20433
rect 245 20365 317 20399
rect 351 20365 430 20399
rect 245 20331 430 20365
rect 245 20297 317 20331
rect 351 20297 430 20331
rect 245 20263 430 20297
rect 245 20229 317 20263
rect 351 20229 430 20263
rect 245 20195 430 20229
rect 245 20161 317 20195
rect 351 20161 430 20195
rect 245 20127 430 20161
rect 245 20093 317 20127
rect 351 20093 430 20127
rect 245 20059 430 20093
rect 245 20025 317 20059
rect 351 20025 430 20059
rect 245 19991 430 20025
rect 245 19957 317 19991
rect 351 19957 430 19991
rect 245 19923 430 19957
rect 245 19889 317 19923
rect 351 19889 430 19923
rect 245 19855 430 19889
rect 245 19821 317 19855
rect 351 19821 430 19855
rect 245 19787 430 19821
rect 245 19753 317 19787
rect 351 19753 430 19787
rect 245 19719 430 19753
rect 245 19685 317 19719
rect 351 19685 430 19719
rect 245 19651 430 19685
rect 245 19617 317 19651
rect 351 19617 430 19651
rect 245 19583 430 19617
rect 245 19549 317 19583
rect 351 19549 430 19583
rect 245 19515 430 19549
rect 245 19481 317 19515
rect 351 19481 430 19515
rect 245 19447 430 19481
rect 245 19413 317 19447
rect 351 19413 430 19447
rect 245 19379 430 19413
rect 245 19345 317 19379
rect 351 19345 430 19379
rect 245 19311 430 19345
rect 245 19277 317 19311
rect 351 19277 430 19311
rect 245 19243 430 19277
rect 245 19209 317 19243
rect 351 19209 430 19243
rect 245 19175 430 19209
rect 245 19141 317 19175
rect 351 19141 430 19175
rect 245 19107 430 19141
rect 245 19073 317 19107
rect 351 19073 430 19107
rect 245 19039 430 19073
rect 245 19005 317 19039
rect 351 19005 430 19039
rect 245 18971 430 19005
rect 245 18937 317 18971
rect 351 18937 430 18971
rect 245 18903 430 18937
rect 245 18869 317 18903
rect 351 18869 430 18903
rect 245 18835 430 18869
rect 245 18801 317 18835
rect 351 18801 430 18835
rect 245 18767 430 18801
rect 245 18733 317 18767
rect 351 18733 430 18767
rect 245 18699 430 18733
rect 245 18665 317 18699
rect 351 18665 430 18699
rect 245 18631 430 18665
rect 245 18597 317 18631
rect 351 18597 430 18631
rect 245 18563 430 18597
rect 245 18529 317 18563
rect 351 18529 430 18563
rect 245 18495 430 18529
rect 245 18461 317 18495
rect 351 18461 430 18495
rect 245 18427 430 18461
rect 245 18393 317 18427
rect 351 18393 430 18427
rect 245 18359 430 18393
rect 245 18325 317 18359
rect 351 18325 430 18359
rect 245 18291 430 18325
rect 245 18257 317 18291
rect 351 18257 430 18291
rect 245 18223 430 18257
rect 245 18189 317 18223
rect 351 18189 430 18223
rect 245 18155 430 18189
rect 245 18121 317 18155
rect 351 18121 430 18155
rect 245 18087 430 18121
rect 245 18053 317 18087
rect 351 18053 430 18087
rect 245 18019 430 18053
rect 245 17985 317 18019
rect 351 17985 430 18019
rect 245 17951 430 17985
rect 245 17917 317 17951
rect 351 17917 430 17951
rect 245 17883 430 17917
rect 245 17849 317 17883
rect 351 17849 430 17883
rect 245 17815 430 17849
rect 245 17781 317 17815
rect 351 17781 430 17815
rect 245 17747 430 17781
rect 245 17713 317 17747
rect 351 17713 430 17747
rect 245 17679 430 17713
rect 245 17645 317 17679
rect 351 17645 430 17679
rect 245 17611 430 17645
rect 245 17577 317 17611
rect 351 17577 430 17611
rect 245 17543 430 17577
rect 245 17509 317 17543
rect 351 17509 430 17543
rect 245 17475 430 17509
rect 245 17441 317 17475
rect 351 17441 430 17475
rect 245 17407 430 17441
rect 245 17373 317 17407
rect 351 17373 430 17407
rect 245 17339 430 17373
rect 245 17305 317 17339
rect 351 17305 430 17339
rect 245 17271 430 17305
rect 245 17237 317 17271
rect 351 17237 430 17271
rect 245 17203 430 17237
rect 245 17169 317 17203
rect 351 17169 430 17203
rect 245 17135 430 17169
rect 245 17101 317 17135
rect 351 17101 430 17135
rect 245 17067 430 17101
rect 245 17033 317 17067
rect 351 17033 430 17067
rect 245 16999 430 17033
rect 245 16965 317 16999
rect 351 16965 430 16999
rect 245 16931 430 16965
rect 245 16897 317 16931
rect 351 16897 430 16931
rect 245 16863 430 16897
rect 245 16829 317 16863
rect 351 16829 430 16863
rect 245 16795 430 16829
rect 245 16761 317 16795
rect 351 16761 430 16795
rect 245 16727 430 16761
rect 245 16693 317 16727
rect 351 16693 430 16727
rect 245 16659 430 16693
rect 245 16625 317 16659
rect 351 16625 430 16659
rect 245 16591 430 16625
rect 245 16557 317 16591
rect 351 16557 430 16591
rect 245 16523 430 16557
rect 245 16489 317 16523
rect 351 16489 430 16523
rect 245 16455 430 16489
rect 245 16421 317 16455
rect 351 16421 430 16455
rect 245 16387 430 16421
rect 245 16353 317 16387
rect 351 16353 430 16387
rect 245 16319 430 16353
rect 245 16285 317 16319
rect 351 16285 430 16319
rect 245 16251 430 16285
rect 245 16217 317 16251
rect 351 16217 430 16251
rect 245 16183 430 16217
rect 245 16149 317 16183
rect 351 16149 430 16183
rect 245 16115 430 16149
rect 245 16081 317 16115
rect 351 16081 430 16115
rect 245 16047 430 16081
rect 245 16013 317 16047
rect 351 16013 430 16047
rect 245 15979 430 16013
rect 245 15945 317 15979
rect 351 15945 430 15979
rect 245 15911 430 15945
rect 245 15877 317 15911
rect 351 15877 430 15911
rect 245 15843 430 15877
rect 245 15809 317 15843
rect 351 15809 430 15843
rect 245 15775 430 15809
rect 245 15741 317 15775
rect 351 15741 430 15775
rect 245 15707 430 15741
rect 245 15673 317 15707
rect 351 15673 430 15707
rect 245 15639 430 15673
rect 245 15605 317 15639
rect 351 15605 430 15639
rect 245 15571 430 15605
rect 245 15537 317 15571
rect 351 15537 430 15571
rect 245 15503 430 15537
rect 245 15469 317 15503
rect 351 15469 430 15503
rect 245 15435 430 15469
rect 245 15401 317 15435
rect 351 15401 430 15435
rect 245 15367 430 15401
rect 245 15333 317 15367
rect 351 15333 430 15367
rect 245 15299 430 15333
rect 245 15265 317 15299
rect 351 15265 430 15299
rect 245 15231 430 15265
rect 245 15197 317 15231
rect 351 15197 430 15231
rect 245 15163 430 15197
rect 245 15129 317 15163
rect 351 15129 430 15163
rect 245 15095 430 15129
rect 245 15061 317 15095
rect 351 15061 430 15095
rect 245 15027 430 15061
rect 245 14993 317 15027
rect 351 14993 430 15027
rect 245 14959 430 14993
rect 245 14925 317 14959
rect 351 14925 430 14959
rect 245 14891 430 14925
rect 245 14857 317 14891
rect 351 14857 430 14891
rect 245 14823 430 14857
rect 245 14789 317 14823
rect 351 14789 430 14823
rect 245 14755 430 14789
rect 245 14721 317 14755
rect 351 14721 430 14755
rect 245 14687 430 14721
rect 245 14653 317 14687
rect 351 14653 430 14687
rect 245 14619 430 14653
rect 245 14585 317 14619
rect 351 14585 430 14619
rect 245 14551 430 14585
rect 245 14517 317 14551
rect 351 14517 430 14551
rect 245 14483 430 14517
rect 245 14449 317 14483
rect 351 14449 430 14483
rect 245 14415 430 14449
rect 245 14381 317 14415
rect 351 14381 430 14415
rect 245 14347 430 14381
rect 245 14313 317 14347
rect 351 14313 430 14347
rect 245 14279 430 14313
rect 245 14245 317 14279
rect 351 14245 430 14279
rect 245 14211 430 14245
rect 245 14177 317 14211
rect 351 14177 430 14211
rect 245 14143 430 14177
rect 245 14109 317 14143
rect 351 14109 430 14143
rect 245 14075 430 14109
rect 245 14041 317 14075
rect 351 14041 430 14075
rect 245 14007 430 14041
rect 245 13973 317 14007
rect 351 13973 430 14007
rect 245 13939 430 13973
rect 245 13905 317 13939
rect 351 13905 430 13939
rect 245 13871 430 13905
rect 245 13837 317 13871
rect 351 13837 430 13871
rect 245 13803 430 13837
rect 245 13769 317 13803
rect 351 13769 430 13803
rect 245 13735 430 13769
rect 245 13701 317 13735
rect 351 13701 430 13735
rect 245 13667 430 13701
rect 245 13633 317 13667
rect 351 13633 430 13667
rect 245 13599 430 13633
rect 245 13565 317 13599
rect 351 13565 430 13599
rect 245 13531 430 13565
rect 245 13497 317 13531
rect 351 13497 430 13531
rect 245 13463 430 13497
rect 245 13429 317 13463
rect 351 13429 430 13463
rect 245 13395 430 13429
rect 245 13361 317 13395
rect 351 13361 430 13395
rect 245 13327 430 13361
rect 245 13293 317 13327
rect 351 13293 430 13327
rect 245 13259 430 13293
rect 245 13225 317 13259
rect 351 13225 430 13259
rect 245 13191 430 13225
rect 245 13157 317 13191
rect 351 13157 430 13191
rect 245 13123 430 13157
rect 245 13089 317 13123
rect 351 13089 430 13123
rect 245 13055 430 13089
rect 245 13021 317 13055
rect 351 13021 430 13055
rect 245 12987 430 13021
rect 245 12953 317 12987
rect 351 12953 430 12987
rect 245 12919 430 12953
rect 245 12885 317 12919
rect 351 12885 430 12919
rect 245 12851 430 12885
rect 245 12817 317 12851
rect 351 12817 430 12851
rect 245 12783 430 12817
rect 245 12749 317 12783
rect 351 12749 430 12783
rect 245 12715 430 12749
rect 245 12681 317 12715
rect 351 12681 430 12715
rect 245 12647 430 12681
rect 245 12613 317 12647
rect 351 12613 430 12647
rect 245 12579 430 12613
rect 245 12545 317 12579
rect 351 12545 430 12579
rect 245 12511 430 12545
rect 245 12477 317 12511
rect 351 12477 430 12511
rect 245 12443 430 12477
rect 245 12409 317 12443
rect 351 12409 430 12443
rect 245 12375 430 12409
rect 245 12341 317 12375
rect 351 12341 430 12375
rect 245 12307 430 12341
rect 245 12273 317 12307
rect 351 12273 430 12307
rect 245 12239 430 12273
rect 245 12205 317 12239
rect 351 12205 430 12239
rect 245 12171 430 12205
rect 245 12137 317 12171
rect 351 12137 430 12171
rect 245 12103 430 12137
rect 245 12069 317 12103
rect 351 12069 430 12103
rect 245 12035 430 12069
rect 245 12001 317 12035
rect 351 12001 430 12035
rect 245 11967 430 12001
rect 245 11933 317 11967
rect 351 11933 430 11967
rect 245 11899 430 11933
rect 245 11865 317 11899
rect 351 11865 430 11899
rect 245 11831 430 11865
rect 245 11797 317 11831
rect 351 11797 430 11831
rect 245 11763 430 11797
rect 245 11729 317 11763
rect 351 11729 430 11763
rect 245 11695 430 11729
rect 245 11661 317 11695
rect 351 11661 430 11695
rect 245 11627 430 11661
rect 245 11593 317 11627
rect 351 11593 430 11627
rect 245 11559 430 11593
rect 245 11525 317 11559
rect 351 11525 430 11559
rect 245 11491 430 11525
rect 245 11457 317 11491
rect 351 11457 430 11491
rect 245 11423 430 11457
rect 245 11389 317 11423
rect 351 11389 430 11423
rect 245 11355 430 11389
rect 245 11321 317 11355
rect 351 11321 430 11355
rect 245 11287 430 11321
rect 245 11253 317 11287
rect 351 11253 430 11287
rect 245 11219 430 11253
rect 245 11185 317 11219
rect 351 11185 430 11219
rect 245 11151 430 11185
rect 245 11117 317 11151
rect 351 11117 430 11151
rect 245 11083 430 11117
rect 245 11049 317 11083
rect 351 11049 430 11083
rect 245 11015 430 11049
rect 245 10981 317 11015
rect 351 10981 430 11015
rect 245 10947 430 10981
rect 245 10913 317 10947
rect 351 10913 430 10947
rect 245 10879 430 10913
rect 245 10845 317 10879
rect 351 10845 430 10879
rect 245 10811 430 10845
rect 245 10777 317 10811
rect 351 10777 430 10811
rect 245 10743 430 10777
rect 245 10709 317 10743
rect 351 10709 430 10743
rect 245 10675 430 10709
rect 245 10641 317 10675
rect 351 10641 430 10675
rect 245 10607 430 10641
rect 245 10573 317 10607
rect 351 10573 430 10607
rect 245 10539 430 10573
rect 245 10505 317 10539
rect 351 10505 430 10539
rect 245 10471 430 10505
rect 245 10437 317 10471
rect 351 10437 430 10471
rect 245 10403 430 10437
rect 245 10369 317 10403
rect 351 10369 430 10403
rect 245 10335 430 10369
rect 245 10301 317 10335
rect 351 10301 430 10335
rect 245 10267 430 10301
rect 245 10233 317 10267
rect 351 10233 430 10267
rect 245 10199 430 10233
rect 245 10165 317 10199
rect 351 10165 430 10199
rect 245 10131 430 10165
rect 245 10097 317 10131
rect 351 10097 430 10131
rect 245 10063 430 10097
rect 245 10029 317 10063
rect 351 10029 430 10063
rect 245 9995 430 10029
rect 245 9961 317 9995
rect 351 9961 430 9995
rect 245 9927 430 9961
rect 245 9893 317 9927
rect 351 9893 430 9927
rect 245 9859 430 9893
rect 245 9825 317 9859
rect 351 9825 430 9859
rect 245 9791 430 9825
rect 245 9757 317 9791
rect 351 9757 430 9791
rect 245 9723 430 9757
rect 245 9689 317 9723
rect 351 9689 430 9723
rect 1148 34650 13844 34694
rect 1148 34616 1327 34650
rect 1361 34616 1395 34650
rect 1429 34616 1463 34650
rect 1497 34616 1531 34650
rect 1565 34616 1599 34650
rect 1633 34616 1667 34650
rect 1701 34616 1735 34650
rect 1769 34616 1803 34650
rect 1837 34616 1871 34650
rect 1905 34616 1939 34650
rect 1973 34616 2007 34650
rect 2041 34616 2075 34650
rect 2109 34616 2143 34650
rect 2177 34616 2211 34650
rect 2245 34616 2279 34650
rect 2313 34616 2347 34650
rect 2381 34616 2415 34650
rect 2449 34616 2483 34650
rect 2517 34616 2551 34650
rect 2585 34616 2619 34650
rect 2653 34616 2687 34650
rect 2721 34616 2755 34650
rect 2789 34616 2823 34650
rect 2857 34616 2891 34650
rect 2925 34616 2959 34650
rect 2993 34616 3027 34650
rect 3061 34616 3095 34650
rect 3129 34616 3163 34650
rect 3197 34616 3231 34650
rect 3265 34616 3299 34650
rect 3333 34616 3367 34650
rect 3401 34616 3435 34650
rect 3469 34616 3503 34650
rect 3537 34616 3571 34650
rect 3605 34616 3639 34650
rect 3673 34616 3707 34650
rect 3741 34616 3775 34650
rect 3809 34616 3843 34650
rect 3877 34616 3911 34650
rect 3945 34616 3979 34650
rect 4013 34616 4047 34650
rect 4081 34616 4115 34650
rect 4149 34616 4183 34650
rect 4217 34616 4251 34650
rect 4285 34616 4319 34650
rect 4353 34616 4387 34650
rect 4421 34616 4455 34650
rect 4489 34616 4523 34650
rect 4557 34616 4591 34650
rect 4625 34616 4659 34650
rect 4693 34616 4727 34650
rect 4761 34616 4795 34650
rect 4829 34616 4863 34650
rect 4897 34616 4931 34650
rect 4965 34616 4999 34650
rect 5033 34616 5067 34650
rect 5101 34616 5135 34650
rect 5169 34616 5203 34650
rect 5237 34616 5271 34650
rect 5305 34616 5339 34650
rect 5373 34616 5407 34650
rect 5441 34616 5475 34650
rect 5509 34616 5543 34650
rect 5577 34616 5611 34650
rect 5645 34616 5679 34650
rect 5713 34616 5747 34650
rect 5781 34616 5815 34650
rect 5849 34616 5883 34650
rect 5917 34616 5951 34650
rect 5985 34616 6019 34650
rect 6053 34616 6087 34650
rect 6121 34616 6155 34650
rect 6189 34616 6223 34650
rect 6257 34616 6291 34650
rect 6325 34616 6359 34650
rect 6393 34616 6427 34650
rect 6461 34616 6495 34650
rect 6529 34616 6563 34650
rect 6597 34616 6631 34650
rect 6665 34616 6699 34650
rect 6733 34616 6767 34650
rect 6801 34616 6835 34650
rect 6869 34616 6903 34650
rect 6937 34616 6971 34650
rect 7005 34616 7039 34650
rect 7073 34616 7107 34650
rect 7141 34616 7175 34650
rect 7209 34616 7243 34650
rect 7277 34616 7311 34650
rect 7345 34616 7379 34650
rect 7413 34616 7447 34650
rect 7481 34616 7515 34650
rect 7549 34616 7583 34650
rect 7617 34616 7651 34650
rect 7685 34616 7719 34650
rect 7753 34616 7787 34650
rect 7821 34616 7855 34650
rect 7889 34616 7923 34650
rect 7957 34616 7991 34650
rect 8025 34616 8059 34650
rect 8093 34616 8127 34650
rect 8161 34616 8195 34650
rect 8229 34616 8263 34650
rect 8297 34616 8331 34650
rect 8365 34616 8399 34650
rect 8433 34616 8467 34650
rect 8501 34616 8535 34650
rect 8569 34616 8603 34650
rect 8637 34616 8671 34650
rect 8705 34616 8739 34650
rect 8773 34616 8807 34650
rect 8841 34616 8875 34650
rect 8909 34616 8943 34650
rect 8977 34616 9011 34650
rect 9045 34616 9079 34650
rect 9113 34616 9147 34650
rect 9181 34616 9215 34650
rect 9249 34616 9283 34650
rect 9317 34616 9351 34650
rect 9385 34616 9419 34650
rect 9453 34616 9487 34650
rect 9521 34616 9555 34650
rect 9589 34616 9623 34650
rect 9657 34616 9691 34650
rect 9725 34616 9759 34650
rect 9793 34616 9827 34650
rect 9861 34616 9895 34650
rect 9929 34616 9963 34650
rect 9997 34616 10031 34650
rect 10065 34616 10099 34650
rect 10133 34616 10167 34650
rect 10201 34616 10235 34650
rect 10269 34616 10303 34650
rect 10337 34616 10371 34650
rect 10405 34616 10439 34650
rect 10473 34616 10507 34650
rect 10541 34616 10575 34650
rect 10609 34616 10643 34650
rect 10677 34616 10711 34650
rect 10745 34616 10779 34650
rect 10813 34616 10847 34650
rect 10881 34616 10915 34650
rect 10949 34616 10983 34650
rect 11017 34616 11051 34650
rect 11085 34616 11119 34650
rect 11153 34616 11187 34650
rect 11221 34616 11255 34650
rect 11289 34616 11323 34650
rect 11357 34616 11391 34650
rect 11425 34616 11459 34650
rect 11493 34616 11527 34650
rect 11561 34616 11595 34650
rect 11629 34616 11663 34650
rect 11697 34616 11731 34650
rect 11765 34616 11799 34650
rect 11833 34616 11867 34650
rect 11901 34616 11935 34650
rect 11969 34616 12003 34650
rect 12037 34616 12071 34650
rect 12105 34616 12139 34650
rect 12173 34616 12207 34650
rect 12241 34616 12275 34650
rect 12309 34616 12343 34650
rect 12377 34616 12411 34650
rect 12445 34616 12479 34650
rect 12513 34616 12547 34650
rect 12581 34616 12615 34650
rect 12649 34616 12683 34650
rect 12717 34616 12751 34650
rect 12785 34616 12819 34650
rect 12853 34616 12887 34650
rect 12921 34616 12955 34650
rect 12989 34616 13023 34650
rect 13057 34616 13091 34650
rect 13125 34616 13159 34650
rect 13193 34616 13227 34650
rect 13261 34616 13295 34650
rect 13329 34616 13363 34650
rect 13397 34616 13431 34650
rect 13465 34616 13499 34650
rect 13533 34616 13567 34650
rect 13601 34616 13635 34650
rect 13669 34616 13844 34650
rect 1148 34574 13844 34616
rect 1148 34521 1268 34574
rect 1148 34487 1192 34521
rect 1226 34487 1268 34521
rect 1148 34453 1268 34487
rect 1148 34419 1192 34453
rect 1226 34419 1268 34453
rect 1148 34385 1268 34419
rect 1148 34351 1192 34385
rect 1226 34351 1268 34385
rect 1148 34317 1268 34351
rect 1148 34283 1192 34317
rect 1226 34283 1268 34317
rect 1148 34249 1268 34283
rect 1148 34215 1192 34249
rect 1226 34215 1268 34249
rect 1148 34181 1268 34215
rect 1148 34147 1192 34181
rect 1226 34147 1268 34181
rect 1148 34113 1268 34147
rect 1148 34079 1192 34113
rect 1226 34079 1268 34113
rect 1148 34045 1268 34079
rect 1148 34011 1192 34045
rect 1226 34011 1268 34045
rect 1148 33977 1268 34011
rect 1148 33943 1192 33977
rect 1226 33943 1268 33977
rect 1148 33909 1268 33943
rect 1148 33875 1192 33909
rect 1226 33875 1268 33909
rect 1148 33841 1268 33875
rect 1148 33807 1192 33841
rect 1226 33807 1268 33841
rect 1148 33773 1268 33807
rect 1148 33739 1192 33773
rect 1226 33739 1268 33773
rect 1148 33705 1268 33739
rect 1148 33671 1192 33705
rect 1226 33671 1268 33705
rect 1148 33637 1268 33671
rect 1148 33603 1192 33637
rect 1226 33603 1268 33637
rect 1148 33569 1268 33603
rect 1148 33535 1192 33569
rect 1226 33535 1268 33569
rect 1148 33501 1268 33535
rect 1148 33467 1192 33501
rect 1226 33467 1268 33501
rect 1148 33433 1268 33467
rect 1148 33399 1192 33433
rect 1226 33399 1268 33433
rect 1148 33365 1268 33399
rect 1148 33331 1192 33365
rect 1226 33331 1268 33365
rect 1148 33297 1268 33331
rect 1148 33263 1192 33297
rect 1226 33263 1268 33297
rect 1148 33229 1268 33263
rect 1148 33195 1192 33229
rect 1226 33195 1268 33229
rect 1148 33161 1268 33195
rect 1148 33127 1192 33161
rect 1226 33127 1268 33161
rect 1148 33093 1268 33127
rect 1148 33059 1192 33093
rect 1226 33059 1268 33093
rect 1148 33025 1268 33059
rect 1148 32991 1192 33025
rect 1226 32991 1268 33025
rect 1148 32957 1268 32991
rect 1148 32923 1192 32957
rect 1226 32923 1268 32957
rect 1148 32889 1268 32923
rect 1148 32855 1192 32889
rect 1226 32855 1268 32889
rect 1148 32821 1268 32855
rect 1148 32787 1192 32821
rect 1226 32787 1268 32821
rect 1148 32753 1268 32787
rect 1148 32719 1192 32753
rect 1226 32719 1268 32753
rect 1148 32685 1268 32719
rect 1148 32651 1192 32685
rect 1226 32651 1268 32685
rect 1148 32617 1268 32651
rect 1148 32583 1192 32617
rect 1226 32583 1268 32617
rect 1148 32549 1268 32583
rect 1148 32515 1192 32549
rect 1226 32515 1268 32549
rect 1148 32481 1268 32515
rect 1148 32447 1192 32481
rect 1226 32447 1268 32481
rect 1148 32413 1268 32447
rect 1148 32379 1192 32413
rect 1226 32379 1268 32413
rect 1148 32345 1268 32379
rect 1148 32311 1192 32345
rect 1226 32311 1268 32345
rect 1148 32277 1268 32311
rect 1148 32243 1192 32277
rect 1226 32243 1268 32277
rect 1148 32209 1268 32243
rect 1148 32175 1192 32209
rect 1226 32175 1268 32209
rect 1148 32141 1268 32175
rect 1148 32107 1192 32141
rect 1226 32107 1268 32141
rect 1148 32073 1268 32107
rect 1148 32039 1192 32073
rect 1226 32039 1268 32073
rect 1148 32005 1268 32039
rect 1148 31971 1192 32005
rect 1226 31971 1268 32005
rect 1148 31937 1268 31971
rect 1148 31903 1192 31937
rect 1226 31903 1268 31937
rect 1148 31869 1268 31903
rect 1148 31835 1192 31869
rect 1226 31835 1268 31869
rect 1148 31801 1268 31835
rect 1148 31767 1192 31801
rect 1226 31767 1268 31801
rect 1148 31733 1268 31767
rect 1148 31699 1192 31733
rect 1226 31699 1268 31733
rect 1148 31665 1268 31699
rect 1148 31631 1192 31665
rect 1226 31631 1268 31665
rect 1148 31597 1268 31631
rect 1148 31563 1192 31597
rect 1226 31563 1268 31597
rect 1148 31529 1268 31563
rect 1148 31495 1192 31529
rect 1226 31495 1268 31529
rect 1148 31461 1268 31495
rect 1148 31427 1192 31461
rect 1226 31427 1268 31461
rect 1148 31393 1268 31427
rect 1148 31359 1192 31393
rect 1226 31359 1268 31393
rect 13724 34534 13844 34574
rect 13724 34500 13768 34534
rect 13802 34500 13844 34534
rect 13724 34466 13844 34500
rect 13724 34432 13768 34466
rect 13802 34432 13844 34466
rect 13724 34398 13844 34432
rect 13724 34364 13768 34398
rect 13802 34364 13844 34398
rect 13724 34330 13844 34364
rect 13724 34296 13768 34330
rect 13802 34296 13844 34330
rect 13724 34262 13844 34296
rect 13724 34228 13768 34262
rect 13802 34228 13844 34262
rect 13724 34194 13844 34228
rect 13724 34160 13768 34194
rect 13802 34160 13844 34194
rect 13724 34126 13844 34160
rect 13724 34092 13768 34126
rect 13802 34092 13844 34126
rect 13724 34058 13844 34092
rect 13724 34024 13768 34058
rect 13802 34024 13844 34058
rect 13724 33990 13844 34024
rect 13724 33956 13768 33990
rect 13802 33956 13844 33990
rect 13724 33922 13844 33956
rect 13724 33888 13768 33922
rect 13802 33888 13844 33922
rect 13724 33854 13844 33888
rect 13724 33820 13768 33854
rect 13802 33820 13844 33854
rect 13724 33786 13844 33820
rect 13724 33752 13768 33786
rect 13802 33752 13844 33786
rect 13724 33718 13844 33752
rect 13724 33684 13768 33718
rect 13802 33684 13844 33718
rect 13724 33650 13844 33684
rect 13724 33616 13768 33650
rect 13802 33616 13844 33650
rect 13724 33582 13844 33616
rect 13724 33548 13768 33582
rect 13802 33548 13844 33582
rect 13724 33514 13844 33548
rect 13724 33480 13768 33514
rect 13802 33480 13844 33514
rect 13724 33446 13844 33480
rect 13724 33412 13768 33446
rect 13802 33412 13844 33446
rect 13724 33378 13844 33412
rect 13724 33344 13768 33378
rect 13802 33344 13844 33378
rect 13724 33310 13844 33344
rect 13724 33276 13768 33310
rect 13802 33276 13844 33310
rect 13724 33242 13844 33276
rect 13724 33208 13768 33242
rect 13802 33208 13844 33242
rect 13724 33174 13844 33208
rect 13724 33140 13768 33174
rect 13802 33140 13844 33174
rect 13724 33106 13844 33140
rect 13724 33072 13768 33106
rect 13802 33072 13844 33106
rect 13724 33038 13844 33072
rect 13724 33004 13768 33038
rect 13802 33004 13844 33038
rect 13724 32970 13844 33004
rect 13724 32936 13768 32970
rect 13802 32936 13844 32970
rect 13724 32902 13844 32936
rect 13724 32868 13768 32902
rect 13802 32868 13844 32902
rect 13724 32834 13844 32868
rect 13724 32800 13768 32834
rect 13802 32800 13844 32834
rect 13724 32766 13844 32800
rect 13724 32732 13768 32766
rect 13802 32732 13844 32766
rect 13724 32698 13844 32732
rect 13724 32664 13768 32698
rect 13802 32664 13844 32698
rect 13724 32630 13844 32664
rect 13724 32596 13768 32630
rect 13802 32596 13844 32630
rect 13724 32562 13844 32596
rect 13724 32528 13768 32562
rect 13802 32528 13844 32562
rect 13724 32494 13844 32528
rect 13724 32460 13768 32494
rect 13802 32460 13844 32494
rect 13724 32426 13844 32460
rect 13724 32392 13768 32426
rect 13802 32392 13844 32426
rect 13724 32358 13844 32392
rect 13724 32324 13768 32358
rect 13802 32324 13844 32358
rect 13724 32290 13844 32324
rect 13724 32256 13768 32290
rect 13802 32256 13844 32290
rect 13724 32222 13844 32256
rect 13724 32188 13768 32222
rect 13802 32188 13844 32222
rect 13724 32154 13844 32188
rect 13724 32120 13768 32154
rect 13802 32120 13844 32154
rect 13724 32086 13844 32120
rect 13724 32052 13768 32086
rect 13802 32052 13844 32086
rect 13724 32018 13844 32052
rect 13724 31984 13768 32018
rect 13802 31984 13844 32018
rect 13724 31950 13844 31984
rect 13724 31916 13768 31950
rect 13802 31916 13844 31950
rect 13724 31882 13844 31916
rect 13724 31848 13768 31882
rect 13802 31848 13844 31882
rect 13724 31814 13844 31848
rect 13724 31780 13768 31814
rect 13802 31780 13844 31814
rect 13724 31746 13844 31780
rect 13724 31712 13768 31746
rect 13802 31712 13844 31746
rect 13724 31678 13844 31712
rect 13724 31644 13768 31678
rect 13802 31644 13844 31678
rect 13724 31610 13844 31644
rect 13724 31576 13768 31610
rect 13802 31576 13844 31610
rect 13724 31542 13844 31576
rect 13724 31508 13768 31542
rect 13802 31508 13844 31542
rect 13724 31474 13844 31508
rect 13724 31440 13768 31474
rect 13802 31440 13844 31474
rect 13724 31406 13844 31440
rect 1148 31325 1268 31359
rect 1148 31291 1192 31325
rect 1226 31291 1268 31325
rect 1148 31257 1268 31291
rect 1148 31223 1192 31257
rect 1226 31223 1268 31257
rect 1148 31189 1268 31223
rect 1148 31155 1192 31189
rect 1226 31155 1268 31189
rect 1148 31121 1268 31155
rect 1148 31087 1192 31121
rect 1226 31087 1268 31121
rect 1148 31053 1268 31087
rect 1148 31019 1192 31053
rect 1226 31019 1268 31053
rect 1148 30985 1268 31019
rect 1148 30951 1192 30985
rect 1226 30951 1268 30985
rect 1148 30917 1268 30951
rect 1148 30883 1192 30917
rect 1226 30883 1268 30917
rect 1148 30849 1268 30883
rect 1148 30815 1192 30849
rect 1226 30815 1268 30849
rect 1148 30781 1268 30815
rect 1148 30747 1192 30781
rect 1226 30747 1268 30781
rect 1148 30713 1268 30747
rect 1148 30679 1192 30713
rect 1226 30679 1268 30713
rect 1148 30645 1268 30679
rect 1148 30611 1192 30645
rect 1226 30611 1268 30645
rect 1148 30577 1268 30611
rect 1148 30543 1192 30577
rect 1226 30543 1268 30577
rect 1148 30509 1268 30543
rect 1148 30475 1192 30509
rect 1226 30475 1268 30509
rect 1148 30441 1268 30475
rect 1148 30407 1192 30441
rect 1226 30407 1268 30441
rect 1148 30373 1268 30407
rect 1148 30339 1192 30373
rect 1226 30339 1268 30373
rect 1148 30305 1268 30339
rect 1148 30271 1192 30305
rect 1226 30271 1268 30305
rect 1148 30237 1268 30271
rect 1148 30203 1192 30237
rect 1226 30203 1268 30237
rect 1148 30169 1268 30203
rect 1148 30135 1192 30169
rect 1226 30135 1268 30169
rect 1148 30101 1268 30135
rect 1148 30067 1192 30101
rect 1226 30067 1268 30101
rect 1148 30033 1268 30067
rect 1148 29999 1192 30033
rect 1226 29999 1268 30033
rect 1148 29965 1268 29999
rect 1148 29931 1192 29965
rect 1226 29931 1268 29965
rect 1148 29897 1268 29931
rect 1148 29863 1192 29897
rect 1226 29863 1268 29897
rect 1148 29829 1268 29863
rect 1148 29795 1192 29829
rect 1226 29795 1268 29829
rect 1148 29761 1268 29795
rect 1148 29727 1192 29761
rect 1226 29727 1268 29761
rect 1148 29693 1268 29727
rect 1148 29659 1192 29693
rect 1226 29659 1268 29693
rect 1148 29625 1268 29659
rect 1148 29591 1192 29625
rect 1226 29591 1268 29625
rect 1148 29557 1268 29591
rect 1148 29523 1192 29557
rect 1226 29523 1268 29557
rect 1148 29489 1268 29523
rect 1148 29455 1192 29489
rect 1226 29455 1268 29489
rect 1148 29421 1268 29455
rect 1148 29387 1192 29421
rect 1226 29387 1268 29421
rect 1148 29353 1268 29387
rect 1148 29319 1192 29353
rect 1226 29319 1268 29353
rect 1148 29285 1268 29319
rect 1148 29251 1192 29285
rect 1226 29251 1268 29285
rect 1148 29217 1268 29251
rect 1148 29183 1192 29217
rect 1226 29183 1268 29217
rect 1148 29149 1268 29183
rect 1148 29115 1192 29149
rect 1226 29115 1268 29149
rect 1148 29081 1268 29115
rect 1148 29047 1192 29081
rect 1226 29047 1268 29081
rect 1148 29013 1268 29047
rect 1148 28979 1192 29013
rect 1226 28979 1268 29013
rect 1148 28945 1268 28979
rect 1148 28911 1192 28945
rect 1226 28911 1268 28945
rect 1148 28877 1268 28911
rect 1148 28843 1192 28877
rect 1226 28843 1268 28877
rect 1148 28809 1268 28843
rect 1148 28775 1192 28809
rect 1226 28775 1268 28809
rect 1148 28741 1268 28775
rect 1148 28707 1192 28741
rect 1226 28707 1268 28741
rect 1148 28673 1268 28707
rect 1148 28639 1192 28673
rect 1226 28639 1268 28673
rect 1148 28605 1268 28639
rect 1148 28571 1192 28605
rect 1226 28571 1268 28605
rect 1148 28537 1268 28571
rect 1148 28503 1192 28537
rect 1226 28503 1268 28537
rect 1148 28469 1268 28503
rect 1148 28435 1192 28469
rect 1226 28435 1268 28469
rect 1148 28401 1268 28435
rect 1148 28367 1192 28401
rect 1226 28367 1268 28401
rect 1148 28333 1268 28367
rect 1148 28299 1192 28333
rect 1226 28299 1268 28333
rect 1148 28265 1268 28299
rect 1148 28231 1192 28265
rect 1226 28231 1268 28265
rect 1148 28197 1268 28231
rect 1148 28163 1192 28197
rect 1226 28163 1268 28197
rect 1148 28129 1268 28163
rect 1148 28095 1192 28129
rect 1226 28095 1268 28129
rect 1148 28061 1268 28095
rect 1148 28027 1192 28061
rect 1226 28027 1268 28061
rect 1148 27993 1268 28027
rect 1148 27959 1192 27993
rect 1226 27959 1268 27993
rect 1148 27925 1268 27959
rect 1148 27891 1192 27925
rect 1226 27891 1268 27925
rect 1148 27857 1268 27891
rect 1148 27823 1192 27857
rect 1226 27823 1268 27857
rect 1148 27789 1268 27823
rect 1148 27755 1192 27789
rect 1226 27755 1268 27789
rect 1148 27721 1268 27755
rect 1148 27687 1192 27721
rect 1226 27687 1268 27721
rect 1148 27653 1268 27687
rect 1148 27619 1192 27653
rect 1226 27619 1268 27653
rect 1148 27585 1268 27619
rect 1148 27551 1192 27585
rect 1226 27551 1268 27585
rect 1148 27517 1268 27551
rect 1148 27483 1192 27517
rect 1226 27483 1268 27517
rect 1148 27449 1268 27483
rect 1148 27415 1192 27449
rect 1226 27415 1268 27449
rect 1148 27381 1268 27415
rect 1148 27347 1192 27381
rect 1226 27347 1268 27381
rect 1148 27313 1268 27347
rect 1148 27279 1192 27313
rect 1226 27279 1268 27313
rect 1148 27245 1268 27279
rect 1148 27211 1192 27245
rect 1226 27211 1268 27245
rect 1148 27177 1268 27211
rect 1148 27143 1192 27177
rect 1226 27143 1268 27177
rect 1148 27109 1268 27143
rect 1148 27075 1192 27109
rect 1226 27075 1268 27109
rect 1148 27041 1268 27075
rect 1148 27007 1192 27041
rect 1226 27007 1268 27041
rect 13724 31372 13768 31406
rect 13802 31372 13844 31406
rect 13724 31338 13844 31372
rect 13724 31304 13768 31338
rect 13802 31304 13844 31338
rect 13724 31270 13844 31304
rect 13724 31236 13768 31270
rect 13802 31236 13844 31270
rect 13724 31202 13844 31236
rect 13724 31168 13768 31202
rect 13802 31168 13844 31202
rect 13724 31134 13844 31168
rect 13724 31100 13768 31134
rect 13802 31100 13844 31134
rect 13724 31066 13844 31100
rect 13724 31032 13768 31066
rect 13802 31032 13844 31066
rect 13724 30998 13844 31032
rect 13724 30964 13768 30998
rect 13802 30964 13844 30998
rect 13724 30930 13844 30964
rect 13724 30896 13768 30930
rect 13802 30896 13844 30930
rect 13724 30862 13844 30896
rect 13724 30828 13768 30862
rect 13802 30828 13844 30862
rect 13724 30794 13844 30828
rect 13724 30760 13768 30794
rect 13802 30760 13844 30794
rect 13724 30726 13844 30760
rect 13724 30692 13768 30726
rect 13802 30692 13844 30726
rect 13724 30658 13844 30692
rect 13724 30624 13768 30658
rect 13802 30624 13844 30658
rect 13724 30590 13844 30624
rect 13724 30556 13768 30590
rect 13802 30556 13844 30590
rect 13724 30522 13844 30556
rect 13724 30488 13768 30522
rect 13802 30488 13844 30522
rect 13724 30454 13844 30488
rect 13724 30420 13768 30454
rect 13802 30420 13844 30454
rect 13724 30386 13844 30420
rect 13724 30352 13768 30386
rect 13802 30352 13844 30386
rect 13724 30318 13844 30352
rect 13724 30284 13768 30318
rect 13802 30284 13844 30318
rect 13724 30250 13844 30284
rect 13724 30216 13768 30250
rect 13802 30216 13844 30250
rect 13724 30182 13844 30216
rect 13724 30148 13768 30182
rect 13802 30148 13844 30182
rect 13724 30114 13844 30148
rect 13724 30080 13768 30114
rect 13802 30080 13844 30114
rect 13724 30046 13844 30080
rect 13724 30012 13768 30046
rect 13802 30012 13844 30046
rect 13724 29978 13844 30012
rect 13724 29944 13768 29978
rect 13802 29944 13844 29978
rect 13724 29910 13844 29944
rect 13724 29876 13768 29910
rect 13802 29876 13844 29910
rect 13724 29842 13844 29876
rect 13724 29808 13768 29842
rect 13802 29808 13844 29842
rect 13724 29774 13844 29808
rect 13724 29740 13768 29774
rect 13802 29740 13844 29774
rect 13724 29706 13844 29740
rect 13724 29672 13768 29706
rect 13802 29672 13844 29706
rect 13724 29638 13844 29672
rect 13724 29604 13768 29638
rect 13802 29604 13844 29638
rect 13724 29570 13844 29604
rect 13724 29536 13768 29570
rect 13802 29536 13844 29570
rect 13724 29502 13844 29536
rect 13724 29468 13768 29502
rect 13802 29468 13844 29502
rect 13724 29434 13844 29468
rect 13724 29400 13768 29434
rect 13802 29400 13844 29434
rect 13724 29366 13844 29400
rect 13724 29332 13768 29366
rect 13802 29332 13844 29366
rect 13724 29298 13844 29332
rect 13724 29264 13768 29298
rect 13802 29264 13844 29298
rect 13724 29230 13844 29264
rect 13724 29196 13768 29230
rect 13802 29196 13844 29230
rect 13724 29162 13844 29196
rect 13724 29128 13768 29162
rect 13802 29128 13844 29162
rect 13724 29094 13844 29128
rect 13724 29060 13768 29094
rect 13802 29060 13844 29094
rect 13724 29026 13844 29060
rect 13724 28992 13768 29026
rect 13802 28992 13844 29026
rect 13724 28958 13844 28992
rect 13724 28924 13768 28958
rect 13802 28924 13844 28958
rect 13724 28890 13844 28924
rect 13724 28856 13768 28890
rect 13802 28856 13844 28890
rect 13724 28822 13844 28856
rect 13724 28788 13768 28822
rect 13802 28788 13844 28822
rect 13724 28754 13844 28788
rect 13724 28720 13768 28754
rect 13802 28720 13844 28754
rect 13724 28686 13844 28720
rect 13724 28652 13768 28686
rect 13802 28652 13844 28686
rect 13724 28618 13844 28652
rect 13724 28584 13768 28618
rect 13802 28584 13844 28618
rect 13724 28550 13844 28584
rect 13724 28516 13768 28550
rect 13802 28516 13844 28550
rect 13724 28482 13844 28516
rect 13724 28448 13768 28482
rect 13802 28448 13844 28482
rect 13724 28414 13844 28448
rect 13724 28380 13768 28414
rect 13802 28380 13844 28414
rect 13724 28346 13844 28380
rect 13724 28312 13768 28346
rect 13802 28312 13844 28346
rect 13724 28278 13844 28312
rect 13724 28244 13768 28278
rect 13802 28244 13844 28278
rect 13724 28210 13844 28244
rect 13724 28176 13768 28210
rect 13802 28176 13844 28210
rect 13724 28142 13844 28176
rect 13724 28108 13768 28142
rect 13802 28108 13844 28142
rect 13724 28074 13844 28108
rect 13724 28040 13768 28074
rect 13802 28040 13844 28074
rect 13724 28006 13844 28040
rect 13724 27972 13768 28006
rect 13802 27972 13844 28006
rect 13724 27938 13844 27972
rect 13724 27904 13768 27938
rect 13802 27904 13844 27938
rect 13724 27870 13844 27904
rect 13724 27836 13768 27870
rect 13802 27836 13844 27870
rect 13724 27802 13844 27836
rect 13724 27768 13768 27802
rect 13802 27768 13844 27802
rect 13724 27734 13844 27768
rect 13724 27700 13768 27734
rect 13802 27700 13844 27734
rect 13724 27666 13844 27700
rect 13724 27632 13768 27666
rect 13802 27632 13844 27666
rect 13724 27598 13844 27632
rect 13724 27564 13768 27598
rect 13802 27564 13844 27598
rect 13724 27530 13844 27564
rect 13724 27496 13768 27530
rect 13802 27496 13844 27530
rect 13724 27462 13844 27496
rect 13724 27428 13768 27462
rect 13802 27428 13844 27462
rect 13724 27394 13844 27428
rect 13724 27360 13768 27394
rect 13802 27360 13844 27394
rect 13724 27326 13844 27360
rect 13724 27292 13768 27326
rect 13802 27292 13844 27326
rect 13724 27258 13844 27292
rect 13724 27224 13768 27258
rect 13802 27224 13844 27258
rect 13724 27190 13844 27224
rect 13724 27156 13768 27190
rect 13802 27156 13844 27190
rect 13724 27122 13844 27156
rect 13724 27088 13768 27122
rect 13802 27088 13844 27122
rect 13724 27054 13844 27088
rect 13724 27020 13768 27054
rect 13802 27020 13844 27054
rect 1148 26973 1268 27007
rect 1148 26939 1192 26973
rect 1226 26939 1268 26973
rect 1148 26905 1268 26939
rect 1148 26871 1192 26905
rect 1226 26871 1268 26905
rect 1148 26837 1268 26871
rect 1148 26803 1192 26837
rect 1226 26803 1268 26837
rect 1148 26769 1268 26803
rect 1148 26735 1192 26769
rect 1226 26735 1268 26769
rect 1148 26701 1268 26735
rect 1148 26667 1192 26701
rect 1226 26667 1268 26701
rect 1148 26633 1268 26667
rect 1148 26599 1192 26633
rect 1226 26599 1268 26633
rect 1148 26565 1268 26599
rect 1148 26531 1192 26565
rect 1226 26531 1268 26565
rect 1148 26497 1268 26531
rect 1148 26463 1192 26497
rect 1226 26463 1268 26497
rect 1148 26429 1268 26463
rect 1148 26395 1192 26429
rect 1226 26395 1268 26429
rect 1148 26361 1268 26395
rect 1148 26327 1192 26361
rect 1226 26327 1268 26361
rect 1148 26293 1268 26327
rect 1148 26259 1192 26293
rect 1226 26259 1268 26293
rect 1148 26225 1268 26259
rect 1148 26191 1192 26225
rect 1226 26191 1268 26225
rect 1148 26157 1268 26191
rect 1148 26123 1192 26157
rect 1226 26123 1268 26157
rect 1148 26089 1268 26123
rect 1148 26055 1192 26089
rect 1226 26055 1268 26089
rect 1148 26021 1268 26055
rect 1148 25987 1192 26021
rect 1226 25987 1268 26021
rect 1148 25953 1268 25987
rect 1148 25919 1192 25953
rect 1226 25919 1268 25953
rect 1148 25885 1268 25919
rect 1148 25851 1192 25885
rect 1226 25851 1268 25885
rect 1148 25817 1268 25851
rect 1148 25783 1192 25817
rect 1226 25783 1268 25817
rect 1148 25749 1268 25783
rect 1148 25715 1192 25749
rect 1226 25715 1268 25749
rect 1148 25681 1268 25715
rect 1148 25647 1192 25681
rect 1226 25647 1268 25681
rect 1148 25613 1268 25647
rect 1148 25579 1192 25613
rect 1226 25579 1268 25613
rect 1148 25545 1268 25579
rect 1148 25511 1192 25545
rect 1226 25511 1268 25545
rect 1148 25477 1268 25511
rect 1148 25443 1192 25477
rect 1226 25443 1268 25477
rect 1148 25409 1268 25443
rect 1148 25375 1192 25409
rect 1226 25375 1268 25409
rect 1148 25341 1268 25375
rect 1148 25307 1192 25341
rect 1226 25307 1268 25341
rect 1148 25273 1268 25307
rect 1148 25239 1192 25273
rect 1226 25239 1268 25273
rect 1148 25205 1268 25239
rect 1148 25171 1192 25205
rect 1226 25171 1268 25205
rect 1148 25137 1268 25171
rect 1148 25103 1192 25137
rect 1226 25103 1268 25137
rect 1148 25069 1268 25103
rect 1148 25035 1192 25069
rect 1226 25035 1268 25069
rect 1148 25001 1268 25035
rect 1148 24967 1192 25001
rect 1226 24967 1268 25001
rect 1148 24933 1268 24967
rect 1148 24899 1192 24933
rect 1226 24899 1268 24933
rect 1148 24865 1268 24899
rect 1148 24831 1192 24865
rect 1226 24831 1268 24865
rect 1148 24797 1268 24831
rect 1148 24763 1192 24797
rect 1226 24763 1268 24797
rect 1148 24729 1268 24763
rect 1148 24695 1192 24729
rect 1226 24695 1268 24729
rect 1148 24661 1268 24695
rect 1148 24627 1192 24661
rect 1226 24627 1268 24661
rect 1148 24593 1268 24627
rect 1148 24559 1192 24593
rect 1226 24559 1268 24593
rect 1148 24525 1268 24559
rect 1148 24491 1192 24525
rect 1226 24491 1268 24525
rect 1148 24457 1268 24491
rect 1148 24423 1192 24457
rect 1226 24423 1268 24457
rect 1148 24389 1268 24423
rect 1148 24355 1192 24389
rect 1226 24355 1268 24389
rect 1148 24321 1268 24355
rect 1148 24287 1192 24321
rect 1226 24287 1268 24321
rect 1148 24253 1268 24287
rect 1148 24219 1192 24253
rect 1226 24219 1268 24253
rect 1148 24185 1268 24219
rect 1148 24151 1192 24185
rect 1226 24151 1268 24185
rect 1148 24117 1268 24151
rect 1148 24083 1192 24117
rect 1226 24083 1268 24117
rect 1148 24049 1268 24083
rect 1148 24015 1192 24049
rect 1226 24015 1268 24049
rect 1148 23981 1268 24015
rect 1148 23947 1192 23981
rect 1226 23947 1268 23981
rect 1148 23913 1268 23947
rect 1148 23879 1192 23913
rect 1226 23879 1268 23913
rect 1148 23845 1268 23879
rect 1148 23811 1192 23845
rect 1226 23811 1268 23845
rect 1148 23777 1268 23811
rect 1148 23743 1192 23777
rect 1226 23743 1268 23777
rect 1148 23709 1268 23743
rect 1148 23675 1192 23709
rect 1226 23675 1268 23709
rect 1148 23641 1268 23675
rect 1148 23607 1192 23641
rect 1226 23607 1268 23641
rect 1148 23573 1268 23607
rect 1148 23539 1192 23573
rect 1226 23539 1268 23573
rect 1148 23505 1268 23539
rect 1148 23471 1192 23505
rect 1226 23471 1268 23505
rect 1148 23437 1268 23471
rect 1148 23403 1192 23437
rect 1226 23403 1268 23437
rect 1148 23369 1268 23403
rect 1148 23335 1192 23369
rect 1226 23335 1268 23369
rect 1148 23301 1268 23335
rect 1148 23267 1192 23301
rect 1226 23267 1268 23301
rect 1148 23233 1268 23267
rect 1148 23199 1192 23233
rect 1226 23199 1268 23233
rect 1148 23165 1268 23199
rect 1148 23131 1192 23165
rect 1226 23131 1268 23165
rect 1148 23097 1268 23131
rect 1148 23063 1192 23097
rect 1226 23063 1268 23097
rect 1148 23029 1268 23063
rect 1148 22995 1192 23029
rect 1226 22995 1268 23029
rect 1148 22961 1268 22995
rect 1148 22927 1192 22961
rect 1226 22927 1268 22961
rect 1148 22893 1268 22927
rect 1148 22859 1192 22893
rect 1226 22859 1268 22893
rect 1148 22825 1268 22859
rect 1148 22791 1192 22825
rect 1226 22791 1268 22825
rect 1148 22757 1268 22791
rect 1148 22723 1192 22757
rect 1226 22723 1268 22757
rect 1148 22689 1268 22723
rect 1148 22655 1192 22689
rect 1226 22655 1268 22689
rect 1148 22621 1268 22655
rect 1148 22587 1192 22621
rect 1226 22587 1268 22621
rect 1148 22553 1268 22587
rect 1148 22519 1192 22553
rect 1226 22519 1268 22553
rect 1148 22485 1268 22519
rect 1148 22451 1192 22485
rect 1226 22451 1268 22485
rect 1148 22417 1268 22451
rect 1148 22383 1192 22417
rect 1226 22383 1268 22417
rect 1148 22349 1268 22383
rect 1148 22315 1192 22349
rect 1226 22315 1268 22349
rect 1148 22281 1268 22315
rect 1148 22247 1192 22281
rect 1226 22247 1268 22281
rect 1148 22213 1268 22247
rect 1148 22179 1192 22213
rect 1226 22179 1268 22213
rect 1148 22145 1268 22179
rect 1148 22111 1192 22145
rect 1226 22111 1268 22145
rect 1148 22077 1268 22111
rect 1148 22043 1192 22077
rect 1226 22043 1268 22077
rect 1148 22009 1268 22043
rect 1148 21975 1192 22009
rect 1226 21975 1268 22009
rect 1148 21941 1268 21975
rect 1148 21907 1192 21941
rect 1226 21907 1268 21941
rect 1148 21873 1268 21907
rect 1148 21839 1192 21873
rect 1226 21839 1268 21873
rect 1148 21805 1268 21839
rect 1148 21771 1192 21805
rect 1226 21771 1268 21805
rect 1148 21737 1268 21771
rect 1148 21703 1192 21737
rect 1226 21703 1268 21737
rect 1148 21669 1268 21703
rect 1148 21635 1192 21669
rect 1226 21635 1268 21669
rect 1148 21601 1268 21635
rect 1148 21567 1192 21601
rect 1226 21567 1268 21601
rect 1148 21533 1268 21567
rect 1148 21499 1192 21533
rect 1226 21499 1268 21533
rect 1148 21465 1268 21499
rect 1148 21431 1192 21465
rect 1226 21431 1268 21465
rect 1148 21397 1268 21431
rect 1148 21363 1192 21397
rect 1226 21363 1268 21397
rect 1148 21329 1268 21363
rect 1148 21295 1192 21329
rect 1226 21295 1268 21329
rect 1148 21261 1268 21295
rect 1148 21227 1192 21261
rect 1226 21227 1268 21261
rect 1148 21193 1268 21227
rect 1148 21159 1192 21193
rect 1226 21159 1268 21193
rect 1148 21125 1268 21159
rect 1148 21091 1192 21125
rect 1226 21091 1268 21125
rect 1148 21057 1268 21091
rect 1148 21023 1192 21057
rect 1226 21023 1268 21057
rect 1148 20989 1268 21023
rect 1148 20955 1192 20989
rect 1226 20955 1268 20989
rect 1148 20921 1268 20955
rect 1148 20887 1192 20921
rect 1226 20887 1268 20921
rect 1148 20853 1268 20887
rect 1148 20819 1192 20853
rect 1226 20819 1268 20853
rect 1148 20785 1268 20819
rect 1148 20751 1192 20785
rect 1226 20751 1268 20785
rect 1148 20717 1268 20751
rect 1148 20683 1192 20717
rect 1226 20683 1268 20717
rect 1148 20649 1268 20683
rect 1148 20615 1192 20649
rect 1226 20615 1268 20649
rect 1148 20581 1268 20615
rect 1148 20547 1192 20581
rect 1226 20547 1268 20581
rect 1148 20513 1268 20547
rect 1148 20479 1192 20513
rect 1226 20479 1268 20513
rect 1148 20445 1268 20479
rect 1148 20411 1192 20445
rect 1226 20411 1268 20445
rect 1148 20377 1268 20411
rect 1148 20343 1192 20377
rect 1226 20343 1268 20377
rect 1148 20309 1268 20343
rect 1148 20275 1192 20309
rect 1226 20275 1268 20309
rect 1148 20241 1268 20275
rect 1148 20207 1192 20241
rect 1226 20207 1268 20241
rect 1148 20173 1268 20207
rect 1148 20139 1192 20173
rect 1226 20139 1268 20173
rect 1148 20105 1268 20139
rect 1148 20071 1192 20105
rect 1226 20071 1268 20105
rect 1148 20037 1268 20071
rect 1148 20003 1192 20037
rect 1226 20003 1268 20037
rect 1148 19969 1268 20003
rect 1148 19935 1192 19969
rect 1226 19935 1268 19969
rect 1148 19901 1268 19935
rect 1148 19867 1192 19901
rect 1226 19867 1268 19901
rect 1148 19833 1268 19867
rect 1148 19799 1192 19833
rect 1226 19799 1268 19833
rect 1148 19765 1268 19799
rect 1148 19731 1192 19765
rect 1226 19731 1268 19765
rect 1148 19697 1268 19731
rect 1148 19663 1192 19697
rect 1226 19663 1268 19697
rect 1148 19629 1268 19663
rect 1148 19595 1192 19629
rect 1226 19595 1268 19629
rect 1148 19561 1268 19595
rect 1148 19527 1192 19561
rect 1226 19527 1268 19561
rect 1148 19493 1268 19527
rect 1148 19459 1192 19493
rect 1226 19459 1268 19493
rect 1148 19425 1268 19459
rect 1148 19391 1192 19425
rect 1226 19391 1268 19425
rect 1148 19357 1268 19391
rect 1148 19323 1192 19357
rect 1226 19323 1268 19357
rect 1148 19289 1268 19323
rect 1148 19255 1192 19289
rect 1226 19255 1268 19289
rect 1148 19221 1268 19255
rect 1148 19187 1192 19221
rect 1226 19187 1268 19221
rect 1148 19153 1268 19187
rect 1148 19119 1192 19153
rect 1226 19119 1268 19153
rect 1148 19085 1268 19119
rect 1148 19051 1192 19085
rect 1226 19051 1268 19085
rect 1148 19017 1268 19051
rect 1148 18983 1192 19017
rect 1226 18983 1268 19017
rect 1148 18949 1268 18983
rect 1148 18915 1192 18949
rect 1226 18915 1268 18949
rect 1148 18881 1268 18915
rect 1148 18847 1192 18881
rect 1226 18847 1268 18881
rect 1148 18813 1268 18847
rect 1148 18779 1192 18813
rect 1226 18779 1268 18813
rect 1148 18745 1268 18779
rect 1148 18711 1192 18745
rect 1226 18711 1268 18745
rect 1148 18677 1268 18711
rect 1148 18643 1192 18677
rect 1226 18643 1268 18677
rect 1148 18609 1268 18643
rect 1148 18575 1192 18609
rect 1226 18575 1268 18609
rect 1148 18541 1268 18575
rect 1148 18507 1192 18541
rect 1226 18507 1268 18541
rect 1148 18473 1268 18507
rect 1148 18439 1192 18473
rect 1226 18439 1268 18473
rect 1148 18405 1268 18439
rect 1148 18371 1192 18405
rect 1226 18371 1268 18405
rect 1148 18337 1268 18371
rect 1148 18303 1192 18337
rect 1226 18303 1268 18337
rect 1148 18269 1268 18303
rect 1148 18235 1192 18269
rect 1226 18235 1268 18269
rect 1148 18201 1268 18235
rect 1148 18167 1192 18201
rect 1226 18167 1268 18201
rect 1148 18133 1268 18167
rect 1148 18099 1192 18133
rect 1226 18099 1268 18133
rect 1148 18065 1268 18099
rect 1148 18031 1192 18065
rect 1226 18031 1268 18065
rect 1148 17997 1268 18031
rect 1148 17963 1192 17997
rect 1226 17963 1268 17997
rect 1148 17929 1268 17963
rect 1148 17895 1192 17929
rect 1226 17895 1268 17929
rect 1148 17861 1268 17895
rect 1148 17827 1192 17861
rect 1226 17827 1268 17861
rect 1148 17793 1268 17827
rect 1148 17759 1192 17793
rect 1226 17759 1268 17793
rect 1148 17725 1268 17759
rect 1148 17691 1192 17725
rect 1226 17691 1268 17725
rect 1148 17657 1268 17691
rect 1148 17623 1192 17657
rect 1226 17623 1268 17657
rect 1148 17589 1268 17623
rect 1148 17555 1192 17589
rect 1226 17555 1268 17589
rect 1148 17521 1268 17555
rect 1148 17487 1192 17521
rect 1226 17487 1268 17521
rect 1148 17453 1268 17487
rect 1148 17419 1192 17453
rect 1226 17419 1268 17453
rect 1148 17385 1268 17419
rect 1148 17351 1192 17385
rect 1226 17351 1268 17385
rect 1148 17317 1268 17351
rect 1148 17283 1192 17317
rect 1226 17283 1268 17317
rect 1148 17249 1268 17283
rect 1148 17215 1192 17249
rect 1226 17215 1268 17249
rect 1148 17181 1268 17215
rect 1148 17147 1192 17181
rect 1226 17147 1268 17181
rect 1148 17113 1268 17147
rect 1148 17079 1192 17113
rect 1226 17079 1268 17113
rect 1148 17045 1268 17079
rect 1148 17011 1192 17045
rect 1226 17011 1268 17045
rect 1148 16977 1268 17011
rect 1148 16943 1192 16977
rect 1226 16943 1268 16977
rect 1148 16909 1268 16943
rect 1148 16875 1192 16909
rect 1226 16875 1268 16909
rect 1148 16841 1268 16875
rect 1148 16807 1192 16841
rect 1226 16807 1268 16841
rect 1148 16773 1268 16807
rect 1148 16739 1192 16773
rect 1226 16739 1268 16773
rect 1148 16705 1268 16739
rect 1148 16671 1192 16705
rect 1226 16671 1268 16705
rect 1148 16637 1268 16671
rect 1148 16603 1192 16637
rect 1226 16603 1268 16637
rect 1148 16569 1268 16603
rect 1148 16535 1192 16569
rect 1226 16535 1268 16569
rect 1148 16501 1268 16535
rect 1148 16467 1192 16501
rect 1226 16467 1268 16501
rect 1148 16433 1268 16467
rect 1148 16399 1192 16433
rect 1226 16399 1268 16433
rect 1148 16365 1268 16399
rect 1148 16331 1192 16365
rect 1226 16331 1268 16365
rect 1148 16297 1268 16331
rect 1148 16263 1192 16297
rect 1226 16263 1268 16297
rect 1148 16229 1268 16263
rect 1148 16195 1192 16229
rect 1226 16195 1268 16229
rect 1148 16161 1268 16195
rect 1148 16127 1192 16161
rect 1226 16127 1268 16161
rect 1148 16093 1268 16127
rect 1148 16059 1192 16093
rect 1226 16059 1268 16093
rect 1148 16025 1268 16059
rect 1148 15991 1192 16025
rect 1226 15991 1268 16025
rect 1148 15957 1268 15991
rect 1148 15923 1192 15957
rect 1226 15923 1268 15957
rect 1148 15889 1268 15923
rect 1148 15855 1192 15889
rect 1226 15855 1268 15889
rect 1148 15821 1268 15855
rect 1148 15787 1192 15821
rect 1226 15787 1268 15821
rect 1148 15753 1268 15787
rect 1148 15719 1192 15753
rect 1226 15719 1268 15753
rect 1148 15685 1268 15719
rect 1148 15651 1192 15685
rect 1226 15651 1268 15685
rect 1148 15617 1268 15651
rect 1148 15583 1192 15617
rect 1226 15583 1268 15617
rect 1148 15549 1268 15583
rect 1148 15515 1192 15549
rect 1226 15515 1268 15549
rect 1148 15481 1268 15515
rect 1148 15447 1192 15481
rect 1226 15447 1268 15481
rect 1148 15413 1268 15447
rect 1148 15379 1192 15413
rect 1226 15379 1268 15413
rect 1148 15345 1268 15379
rect 1148 15311 1192 15345
rect 1226 15311 1268 15345
rect 1148 15277 1268 15311
rect 1148 15243 1192 15277
rect 1226 15243 1268 15277
rect 1148 15209 1268 15243
rect 1148 15175 1192 15209
rect 1226 15175 1268 15209
rect 1148 15141 1268 15175
rect 1148 15107 1192 15141
rect 1226 15107 1268 15141
rect 1148 15073 1268 15107
rect 1148 15039 1192 15073
rect 1226 15039 1268 15073
rect 1148 15005 1268 15039
rect 1148 14971 1192 15005
rect 1226 14971 1268 15005
rect 1148 14937 1268 14971
rect 1148 14903 1192 14937
rect 1226 14903 1268 14937
rect 1148 14869 1268 14903
rect 1148 14835 1192 14869
rect 1226 14835 1268 14869
rect 1148 14801 1268 14835
rect 1148 14767 1192 14801
rect 1226 14767 1268 14801
rect 1148 14733 1268 14767
rect 1148 14699 1192 14733
rect 1226 14699 1268 14733
rect 1148 14665 1268 14699
rect 1148 14631 1192 14665
rect 1226 14631 1268 14665
rect 1148 14597 1268 14631
rect 1148 14563 1192 14597
rect 1226 14563 1268 14597
rect 1148 14529 1268 14563
rect 1148 14495 1192 14529
rect 1226 14495 1268 14529
rect 1148 14461 1268 14495
rect 1148 14427 1192 14461
rect 1226 14427 1268 14461
rect 1148 14393 1268 14427
rect 1148 14359 1192 14393
rect 1226 14359 1268 14393
rect 1148 14325 1268 14359
rect 1148 14291 1192 14325
rect 1226 14291 1268 14325
rect 1148 14257 1268 14291
rect 1148 14223 1192 14257
rect 1226 14223 1268 14257
rect 1148 14189 1268 14223
rect 1148 14155 1192 14189
rect 1226 14155 1268 14189
rect 1148 14121 1268 14155
rect 1148 14087 1192 14121
rect 1226 14087 1268 14121
rect 1148 14053 1268 14087
rect 1148 14019 1192 14053
rect 1226 14019 1268 14053
rect 1148 13985 1268 14019
rect 1148 13951 1192 13985
rect 1226 13951 1268 13985
rect 1148 13917 1268 13951
rect 1148 13883 1192 13917
rect 1226 13883 1268 13917
rect 1148 13849 1268 13883
rect 1148 13815 1192 13849
rect 1226 13815 1268 13849
rect 1148 13781 1268 13815
rect 1148 13747 1192 13781
rect 1226 13747 1268 13781
rect 1148 13713 1268 13747
rect 1148 13679 1192 13713
rect 1226 13679 1268 13713
rect 1148 13645 1268 13679
rect 1148 13611 1192 13645
rect 1226 13611 1268 13645
rect 1148 13577 1268 13611
rect 1148 13543 1192 13577
rect 1226 13543 1268 13577
rect 1148 13509 1268 13543
rect 1148 13475 1192 13509
rect 1226 13475 1268 13509
rect 1148 13441 1268 13475
rect 1148 13407 1192 13441
rect 1226 13407 1268 13441
rect 1148 13373 1268 13407
rect 1148 13339 1192 13373
rect 1226 13339 1268 13373
rect 1148 13305 1268 13339
rect 1148 13271 1192 13305
rect 1226 13271 1268 13305
rect 1148 13237 1268 13271
rect 1148 13203 1192 13237
rect 1226 13203 1268 13237
rect 1148 13169 1268 13203
rect 1148 13135 1192 13169
rect 1226 13135 1268 13169
rect 1148 13101 1268 13135
rect 1148 13067 1192 13101
rect 1226 13067 1268 13101
rect 1148 13033 1268 13067
rect 1148 12999 1192 13033
rect 1226 12999 1268 13033
rect 1148 12965 1268 12999
rect 1148 12931 1192 12965
rect 1226 12931 1268 12965
rect 1148 12897 1268 12931
rect 1148 12863 1192 12897
rect 1226 12863 1268 12897
rect 1148 12829 1268 12863
rect 1148 12795 1192 12829
rect 1226 12795 1268 12829
rect 1148 12761 1268 12795
rect 1148 12727 1192 12761
rect 1226 12727 1268 12761
rect 1148 12693 1268 12727
rect 1148 12659 1192 12693
rect 1226 12659 1268 12693
rect 1148 12625 1268 12659
rect 1148 12591 1192 12625
rect 1226 12591 1268 12625
rect 1148 12557 1268 12591
rect 1148 12523 1192 12557
rect 1226 12523 1268 12557
rect 1148 12489 1268 12523
rect 1148 12455 1192 12489
rect 1226 12455 1268 12489
rect 1148 12421 1268 12455
rect 1148 12387 1192 12421
rect 1226 12387 1268 12421
rect 1148 12353 1268 12387
rect 1148 12319 1192 12353
rect 1226 12319 1268 12353
rect 1148 12285 1268 12319
rect 1148 12251 1192 12285
rect 1226 12251 1268 12285
rect 1148 12217 1268 12251
rect 1148 12183 1192 12217
rect 1226 12183 1268 12217
rect 1148 12149 1268 12183
rect 1148 12115 1192 12149
rect 1226 12115 1268 12149
rect 1148 12081 1268 12115
rect 1148 12047 1192 12081
rect 1226 12047 1268 12081
rect 1148 12013 1268 12047
rect 1148 11979 1192 12013
rect 1226 11979 1268 12013
rect 1148 11945 1268 11979
rect 1148 11911 1192 11945
rect 1226 11911 1268 11945
rect 1148 11877 1268 11911
rect 1148 11843 1192 11877
rect 1226 11843 1268 11877
rect 1148 11809 1268 11843
rect 1148 11775 1192 11809
rect 1226 11775 1268 11809
rect 1148 11741 1268 11775
rect 1148 11707 1192 11741
rect 1226 11707 1268 11741
rect 1148 11673 1268 11707
rect 1148 11639 1192 11673
rect 1226 11639 1268 11673
rect 1148 11605 1268 11639
rect 1148 11571 1192 11605
rect 1226 11571 1268 11605
rect 1148 11537 1268 11571
rect 1148 11503 1192 11537
rect 1226 11503 1268 11537
rect 1148 11469 1268 11503
rect 1148 11435 1192 11469
rect 1226 11435 1268 11469
rect 1148 11401 1268 11435
rect 1148 11367 1192 11401
rect 1226 11367 1268 11401
rect 1148 11333 1268 11367
rect 1148 11299 1192 11333
rect 1226 11299 1268 11333
rect 1148 11265 1268 11299
rect 1148 11231 1192 11265
rect 1226 11231 1268 11265
rect 1148 11197 1268 11231
rect 1148 11163 1192 11197
rect 1226 11163 1268 11197
rect 1148 11129 1268 11163
rect 1148 11095 1192 11129
rect 1226 11095 1268 11129
rect 1148 11061 1268 11095
rect 1148 11027 1192 11061
rect 1226 11027 1268 11061
rect 1148 10993 1268 11027
rect 1148 10959 1192 10993
rect 1226 10959 1268 10993
rect 1148 10925 1268 10959
rect 1148 10891 1192 10925
rect 1226 10891 1268 10925
rect 1148 10857 1268 10891
rect 1148 10823 1192 10857
rect 1226 10823 1268 10857
rect 1148 10789 1268 10823
rect 1148 10755 1192 10789
rect 1226 10755 1268 10789
rect 1148 10721 1268 10755
rect 1148 10687 1192 10721
rect 1226 10687 1268 10721
rect 1148 10653 1268 10687
rect 1148 10619 1192 10653
rect 1226 10619 1268 10653
rect 1148 10585 1268 10619
rect 1148 10551 1192 10585
rect 1226 10551 1268 10585
rect 1148 10517 1268 10551
rect 1148 10483 1192 10517
rect 1226 10483 1268 10517
rect 1148 10449 1268 10483
rect 1148 10415 1192 10449
rect 1226 10415 1268 10449
rect 1148 10362 1268 10415
rect 13724 26986 13844 27020
rect 13724 26952 13768 26986
rect 13802 26952 13844 26986
rect 13724 26918 13844 26952
rect 13724 26884 13768 26918
rect 13802 26884 13844 26918
rect 13724 26850 13844 26884
rect 13724 26816 13768 26850
rect 13802 26816 13844 26850
rect 13724 26782 13844 26816
rect 13724 26748 13768 26782
rect 13802 26748 13844 26782
rect 13724 26714 13844 26748
rect 13724 26680 13768 26714
rect 13802 26680 13844 26714
rect 13724 26646 13844 26680
rect 13724 26612 13768 26646
rect 13802 26612 13844 26646
rect 13724 26578 13844 26612
rect 13724 26544 13768 26578
rect 13802 26544 13844 26578
rect 13724 26510 13844 26544
rect 13724 26476 13768 26510
rect 13802 26476 13844 26510
rect 13724 26442 13844 26476
rect 13724 26408 13768 26442
rect 13802 26408 13844 26442
rect 13724 26374 13844 26408
rect 13724 26340 13768 26374
rect 13802 26340 13844 26374
rect 13724 26306 13844 26340
rect 13724 26272 13768 26306
rect 13802 26272 13844 26306
rect 13724 26238 13844 26272
rect 13724 26204 13768 26238
rect 13802 26204 13844 26238
rect 13724 26170 13844 26204
rect 13724 26136 13768 26170
rect 13802 26136 13844 26170
rect 13724 26102 13844 26136
rect 13724 26068 13768 26102
rect 13802 26068 13844 26102
rect 13724 26034 13844 26068
rect 13724 26000 13768 26034
rect 13802 26000 13844 26034
rect 13724 25966 13844 26000
rect 13724 25932 13768 25966
rect 13802 25932 13844 25966
rect 13724 25898 13844 25932
rect 13724 25864 13768 25898
rect 13802 25864 13844 25898
rect 13724 25830 13844 25864
rect 13724 25796 13768 25830
rect 13802 25796 13844 25830
rect 13724 25762 13844 25796
rect 13724 25728 13768 25762
rect 13802 25728 13844 25762
rect 13724 25694 13844 25728
rect 13724 25660 13768 25694
rect 13802 25660 13844 25694
rect 13724 25626 13844 25660
rect 13724 25592 13768 25626
rect 13802 25592 13844 25626
rect 13724 25558 13844 25592
rect 13724 25524 13768 25558
rect 13802 25524 13844 25558
rect 13724 25490 13844 25524
rect 13724 25456 13768 25490
rect 13802 25456 13844 25490
rect 13724 25422 13844 25456
rect 13724 25388 13768 25422
rect 13802 25388 13844 25422
rect 13724 25354 13844 25388
rect 13724 25320 13768 25354
rect 13802 25320 13844 25354
rect 13724 25286 13844 25320
rect 13724 25252 13768 25286
rect 13802 25252 13844 25286
rect 13724 25218 13844 25252
rect 13724 25184 13768 25218
rect 13802 25184 13844 25218
rect 13724 25150 13844 25184
rect 13724 25116 13768 25150
rect 13802 25116 13844 25150
rect 13724 25082 13844 25116
rect 13724 25048 13768 25082
rect 13802 25048 13844 25082
rect 13724 25014 13844 25048
rect 13724 24980 13768 25014
rect 13802 24980 13844 25014
rect 13724 24946 13844 24980
rect 13724 24912 13768 24946
rect 13802 24912 13844 24946
rect 13724 24878 13844 24912
rect 13724 24844 13768 24878
rect 13802 24844 13844 24878
rect 13724 24810 13844 24844
rect 13724 24776 13768 24810
rect 13802 24776 13844 24810
rect 13724 24742 13844 24776
rect 13724 24708 13768 24742
rect 13802 24708 13844 24742
rect 13724 24674 13844 24708
rect 13724 24640 13768 24674
rect 13802 24640 13844 24674
rect 13724 24606 13844 24640
rect 13724 24572 13768 24606
rect 13802 24572 13844 24606
rect 13724 24538 13844 24572
rect 13724 24504 13768 24538
rect 13802 24504 13844 24538
rect 13724 24470 13844 24504
rect 13724 24436 13768 24470
rect 13802 24436 13844 24470
rect 13724 24402 13844 24436
rect 13724 24368 13768 24402
rect 13802 24368 13844 24402
rect 13724 24334 13844 24368
rect 13724 24300 13768 24334
rect 13802 24300 13844 24334
rect 13724 24266 13844 24300
rect 13724 24232 13768 24266
rect 13802 24232 13844 24266
rect 13724 24198 13844 24232
rect 13724 24164 13768 24198
rect 13802 24164 13844 24198
rect 13724 24130 13844 24164
rect 13724 24096 13768 24130
rect 13802 24096 13844 24130
rect 13724 24062 13844 24096
rect 13724 24028 13768 24062
rect 13802 24028 13844 24062
rect 13724 23994 13844 24028
rect 13724 23960 13768 23994
rect 13802 23960 13844 23994
rect 13724 23926 13844 23960
rect 13724 23892 13768 23926
rect 13802 23892 13844 23926
rect 13724 23858 13844 23892
rect 13724 23824 13768 23858
rect 13802 23824 13844 23858
rect 13724 23790 13844 23824
rect 13724 23756 13768 23790
rect 13802 23756 13844 23790
rect 13724 23722 13844 23756
rect 13724 23688 13768 23722
rect 13802 23688 13844 23722
rect 13724 23654 13844 23688
rect 13724 23620 13768 23654
rect 13802 23620 13844 23654
rect 13724 23586 13844 23620
rect 13724 23552 13768 23586
rect 13802 23552 13844 23586
rect 13724 23518 13844 23552
rect 13724 23484 13768 23518
rect 13802 23484 13844 23518
rect 13724 23450 13844 23484
rect 13724 23416 13768 23450
rect 13802 23416 13844 23450
rect 13724 23382 13844 23416
rect 13724 23348 13768 23382
rect 13802 23348 13844 23382
rect 13724 23314 13844 23348
rect 13724 23280 13768 23314
rect 13802 23280 13844 23314
rect 13724 23246 13844 23280
rect 13724 23212 13768 23246
rect 13802 23212 13844 23246
rect 13724 23178 13844 23212
rect 13724 23144 13768 23178
rect 13802 23144 13844 23178
rect 13724 23110 13844 23144
rect 13724 23076 13768 23110
rect 13802 23076 13844 23110
rect 13724 23042 13844 23076
rect 13724 23008 13768 23042
rect 13802 23008 13844 23042
rect 13724 22974 13844 23008
rect 13724 22940 13768 22974
rect 13802 22940 13844 22974
rect 13724 22906 13844 22940
rect 13724 22872 13768 22906
rect 13802 22872 13844 22906
rect 13724 22838 13844 22872
rect 13724 22804 13768 22838
rect 13802 22804 13844 22838
rect 13724 22770 13844 22804
rect 13724 22736 13768 22770
rect 13802 22736 13844 22770
rect 13724 22702 13844 22736
rect 13724 22668 13768 22702
rect 13802 22668 13844 22702
rect 13724 22634 13844 22668
rect 13724 22600 13768 22634
rect 13802 22600 13844 22634
rect 13724 22566 13844 22600
rect 13724 22532 13768 22566
rect 13802 22532 13844 22566
rect 13724 22498 13844 22532
rect 13724 22464 13768 22498
rect 13802 22464 13844 22498
rect 13724 22430 13844 22464
rect 13724 22396 13768 22430
rect 13802 22396 13844 22430
rect 13724 22362 13844 22396
rect 13724 22328 13768 22362
rect 13802 22328 13844 22362
rect 13724 22294 13844 22328
rect 13724 22260 13768 22294
rect 13802 22260 13844 22294
rect 13724 22226 13844 22260
rect 13724 22192 13768 22226
rect 13802 22192 13844 22226
rect 13724 22158 13844 22192
rect 13724 22124 13768 22158
rect 13802 22124 13844 22158
rect 13724 22090 13844 22124
rect 13724 22056 13768 22090
rect 13802 22056 13844 22090
rect 13724 22022 13844 22056
rect 13724 21988 13768 22022
rect 13802 21988 13844 22022
rect 13724 21954 13844 21988
rect 13724 21920 13768 21954
rect 13802 21920 13844 21954
rect 13724 21886 13844 21920
rect 13724 21852 13768 21886
rect 13802 21852 13844 21886
rect 13724 21818 13844 21852
rect 13724 21784 13768 21818
rect 13802 21784 13844 21818
rect 13724 21750 13844 21784
rect 13724 21716 13768 21750
rect 13802 21716 13844 21750
rect 13724 21682 13844 21716
rect 13724 21648 13768 21682
rect 13802 21648 13844 21682
rect 13724 21614 13844 21648
rect 13724 21580 13768 21614
rect 13802 21580 13844 21614
rect 13724 21546 13844 21580
rect 13724 21512 13768 21546
rect 13802 21512 13844 21546
rect 13724 21478 13844 21512
rect 13724 21444 13768 21478
rect 13802 21444 13844 21478
rect 13724 21410 13844 21444
rect 13724 21376 13768 21410
rect 13802 21376 13844 21410
rect 13724 21342 13844 21376
rect 13724 21308 13768 21342
rect 13802 21308 13844 21342
rect 13724 21274 13844 21308
rect 13724 21240 13768 21274
rect 13802 21240 13844 21274
rect 13724 21206 13844 21240
rect 13724 21172 13768 21206
rect 13802 21172 13844 21206
rect 13724 21138 13844 21172
rect 13724 21104 13768 21138
rect 13802 21104 13844 21138
rect 13724 21070 13844 21104
rect 13724 21036 13768 21070
rect 13802 21036 13844 21070
rect 13724 21002 13844 21036
rect 13724 20968 13768 21002
rect 13802 20968 13844 21002
rect 13724 20934 13844 20968
rect 13724 20900 13768 20934
rect 13802 20900 13844 20934
rect 13724 20866 13844 20900
rect 13724 20832 13768 20866
rect 13802 20832 13844 20866
rect 13724 20798 13844 20832
rect 13724 20764 13768 20798
rect 13802 20764 13844 20798
rect 13724 20730 13844 20764
rect 13724 20696 13768 20730
rect 13802 20696 13844 20730
rect 13724 20662 13844 20696
rect 13724 20628 13768 20662
rect 13802 20628 13844 20662
rect 13724 20594 13844 20628
rect 13724 20560 13768 20594
rect 13802 20560 13844 20594
rect 13724 20526 13844 20560
rect 13724 20492 13768 20526
rect 13802 20492 13844 20526
rect 13724 20458 13844 20492
rect 13724 20424 13768 20458
rect 13802 20424 13844 20458
rect 13724 20390 13844 20424
rect 13724 20356 13768 20390
rect 13802 20356 13844 20390
rect 13724 20322 13844 20356
rect 13724 20288 13768 20322
rect 13802 20288 13844 20322
rect 13724 20254 13844 20288
rect 13724 20220 13768 20254
rect 13802 20220 13844 20254
rect 13724 20186 13844 20220
rect 13724 20152 13768 20186
rect 13802 20152 13844 20186
rect 13724 20118 13844 20152
rect 13724 20084 13768 20118
rect 13802 20084 13844 20118
rect 13724 20050 13844 20084
rect 13724 20016 13768 20050
rect 13802 20016 13844 20050
rect 13724 19982 13844 20016
rect 13724 19948 13768 19982
rect 13802 19948 13844 19982
rect 13724 19914 13844 19948
rect 13724 19880 13768 19914
rect 13802 19880 13844 19914
rect 13724 19846 13844 19880
rect 13724 19812 13768 19846
rect 13802 19812 13844 19846
rect 13724 19778 13844 19812
rect 13724 19744 13768 19778
rect 13802 19744 13844 19778
rect 13724 19710 13844 19744
rect 13724 19676 13768 19710
rect 13802 19676 13844 19710
rect 13724 19642 13844 19676
rect 13724 19608 13768 19642
rect 13802 19608 13844 19642
rect 13724 19574 13844 19608
rect 13724 19540 13768 19574
rect 13802 19540 13844 19574
rect 13724 19506 13844 19540
rect 13724 19472 13768 19506
rect 13802 19472 13844 19506
rect 13724 19438 13844 19472
rect 13724 19404 13768 19438
rect 13802 19404 13844 19438
rect 13724 19370 13844 19404
rect 13724 19336 13768 19370
rect 13802 19336 13844 19370
rect 13724 19302 13844 19336
rect 13724 19268 13768 19302
rect 13802 19268 13844 19302
rect 13724 19234 13844 19268
rect 13724 19200 13768 19234
rect 13802 19200 13844 19234
rect 13724 19166 13844 19200
rect 13724 19132 13768 19166
rect 13802 19132 13844 19166
rect 13724 19098 13844 19132
rect 13724 19064 13768 19098
rect 13802 19064 13844 19098
rect 13724 19030 13844 19064
rect 13724 18996 13768 19030
rect 13802 18996 13844 19030
rect 13724 18962 13844 18996
rect 13724 18928 13768 18962
rect 13802 18928 13844 18962
rect 13724 18894 13844 18928
rect 13724 18860 13768 18894
rect 13802 18860 13844 18894
rect 13724 18826 13844 18860
rect 13724 18792 13768 18826
rect 13802 18792 13844 18826
rect 13724 18758 13844 18792
rect 13724 18724 13768 18758
rect 13802 18724 13844 18758
rect 13724 18690 13844 18724
rect 13724 18656 13768 18690
rect 13802 18656 13844 18690
rect 13724 18622 13844 18656
rect 13724 18588 13768 18622
rect 13802 18588 13844 18622
rect 13724 18554 13844 18588
rect 13724 18520 13768 18554
rect 13802 18520 13844 18554
rect 13724 18486 13844 18520
rect 13724 18452 13768 18486
rect 13802 18452 13844 18486
rect 13724 18418 13844 18452
rect 13724 18384 13768 18418
rect 13802 18384 13844 18418
rect 13724 18350 13844 18384
rect 13724 18316 13768 18350
rect 13802 18316 13844 18350
rect 13724 18282 13844 18316
rect 13724 18248 13768 18282
rect 13802 18248 13844 18282
rect 13724 18214 13844 18248
rect 13724 18180 13768 18214
rect 13802 18180 13844 18214
rect 13724 18146 13844 18180
rect 13724 18112 13768 18146
rect 13802 18112 13844 18146
rect 13724 18078 13844 18112
rect 13724 18044 13768 18078
rect 13802 18044 13844 18078
rect 13724 18010 13844 18044
rect 13724 17976 13768 18010
rect 13802 17976 13844 18010
rect 13724 17942 13844 17976
rect 13724 17908 13768 17942
rect 13802 17908 13844 17942
rect 13724 17874 13844 17908
rect 13724 17840 13768 17874
rect 13802 17840 13844 17874
rect 13724 17806 13844 17840
rect 13724 17772 13768 17806
rect 13802 17772 13844 17806
rect 13724 17738 13844 17772
rect 13724 17704 13768 17738
rect 13802 17704 13844 17738
rect 13724 17670 13844 17704
rect 13724 17636 13768 17670
rect 13802 17636 13844 17670
rect 13724 17602 13844 17636
rect 13724 17568 13768 17602
rect 13802 17568 13844 17602
rect 13724 17534 13844 17568
rect 13724 17500 13768 17534
rect 13802 17500 13844 17534
rect 13724 17466 13844 17500
rect 13724 17432 13768 17466
rect 13802 17432 13844 17466
rect 13724 17398 13844 17432
rect 13724 17364 13768 17398
rect 13802 17364 13844 17398
rect 13724 17330 13844 17364
rect 13724 17296 13768 17330
rect 13802 17296 13844 17330
rect 13724 17262 13844 17296
rect 13724 17228 13768 17262
rect 13802 17228 13844 17262
rect 13724 17194 13844 17228
rect 13724 17160 13768 17194
rect 13802 17160 13844 17194
rect 13724 17126 13844 17160
rect 13724 17092 13768 17126
rect 13802 17092 13844 17126
rect 13724 17058 13844 17092
rect 13724 17024 13768 17058
rect 13802 17024 13844 17058
rect 13724 16990 13844 17024
rect 13724 16956 13768 16990
rect 13802 16956 13844 16990
rect 13724 16922 13844 16956
rect 13724 16888 13768 16922
rect 13802 16888 13844 16922
rect 13724 16854 13844 16888
rect 13724 16820 13768 16854
rect 13802 16820 13844 16854
rect 13724 16786 13844 16820
rect 13724 16752 13768 16786
rect 13802 16752 13844 16786
rect 13724 16718 13844 16752
rect 13724 16684 13768 16718
rect 13802 16684 13844 16718
rect 13724 16650 13844 16684
rect 13724 16616 13768 16650
rect 13802 16616 13844 16650
rect 13724 16582 13844 16616
rect 13724 16548 13768 16582
rect 13802 16548 13844 16582
rect 13724 16514 13844 16548
rect 13724 16480 13768 16514
rect 13802 16480 13844 16514
rect 13724 16446 13844 16480
rect 13724 16412 13768 16446
rect 13802 16412 13844 16446
rect 13724 16378 13844 16412
rect 13724 16344 13768 16378
rect 13802 16344 13844 16378
rect 13724 16310 13844 16344
rect 13724 16276 13768 16310
rect 13802 16276 13844 16310
rect 13724 16242 13844 16276
rect 13724 16208 13768 16242
rect 13802 16208 13844 16242
rect 13724 16174 13844 16208
rect 13724 16140 13768 16174
rect 13802 16140 13844 16174
rect 13724 16106 13844 16140
rect 13724 16072 13768 16106
rect 13802 16072 13844 16106
rect 13724 16038 13844 16072
rect 13724 16004 13768 16038
rect 13802 16004 13844 16038
rect 13724 15970 13844 16004
rect 13724 15936 13768 15970
rect 13802 15936 13844 15970
rect 13724 15902 13844 15936
rect 13724 15868 13768 15902
rect 13802 15868 13844 15902
rect 13724 15834 13844 15868
rect 13724 15800 13768 15834
rect 13802 15800 13844 15834
rect 13724 15766 13844 15800
rect 13724 15732 13768 15766
rect 13802 15732 13844 15766
rect 13724 15698 13844 15732
rect 13724 15664 13768 15698
rect 13802 15664 13844 15698
rect 13724 15630 13844 15664
rect 13724 15596 13768 15630
rect 13802 15596 13844 15630
rect 13724 15562 13844 15596
rect 13724 15528 13768 15562
rect 13802 15528 13844 15562
rect 13724 15494 13844 15528
rect 13724 15460 13768 15494
rect 13802 15460 13844 15494
rect 13724 15426 13844 15460
rect 13724 15392 13768 15426
rect 13802 15392 13844 15426
rect 13724 15358 13844 15392
rect 13724 15324 13768 15358
rect 13802 15324 13844 15358
rect 13724 15290 13844 15324
rect 13724 15256 13768 15290
rect 13802 15256 13844 15290
rect 13724 15222 13844 15256
rect 13724 15188 13768 15222
rect 13802 15188 13844 15222
rect 13724 15154 13844 15188
rect 13724 15120 13768 15154
rect 13802 15120 13844 15154
rect 13724 15086 13844 15120
rect 13724 15052 13768 15086
rect 13802 15052 13844 15086
rect 13724 15018 13844 15052
rect 13724 14984 13768 15018
rect 13802 14984 13844 15018
rect 13724 14950 13844 14984
rect 13724 14916 13768 14950
rect 13802 14916 13844 14950
rect 13724 14882 13844 14916
rect 13724 14848 13768 14882
rect 13802 14848 13844 14882
rect 13724 14814 13844 14848
rect 13724 14780 13768 14814
rect 13802 14780 13844 14814
rect 13724 14746 13844 14780
rect 13724 14712 13768 14746
rect 13802 14712 13844 14746
rect 13724 14678 13844 14712
rect 13724 14644 13768 14678
rect 13802 14644 13844 14678
rect 13724 14610 13844 14644
rect 13724 14576 13768 14610
rect 13802 14576 13844 14610
rect 13724 14542 13844 14576
rect 13724 14508 13768 14542
rect 13802 14508 13844 14542
rect 13724 14474 13844 14508
rect 13724 14440 13768 14474
rect 13802 14440 13844 14474
rect 13724 14406 13844 14440
rect 13724 14372 13768 14406
rect 13802 14372 13844 14406
rect 13724 14338 13844 14372
rect 13724 14304 13768 14338
rect 13802 14304 13844 14338
rect 13724 14270 13844 14304
rect 13724 14236 13768 14270
rect 13802 14236 13844 14270
rect 13724 14202 13844 14236
rect 13724 14168 13768 14202
rect 13802 14168 13844 14202
rect 13724 14134 13844 14168
rect 13724 14100 13768 14134
rect 13802 14100 13844 14134
rect 13724 14066 13844 14100
rect 13724 14032 13768 14066
rect 13802 14032 13844 14066
rect 13724 13998 13844 14032
rect 13724 13964 13768 13998
rect 13802 13964 13844 13998
rect 13724 13930 13844 13964
rect 13724 13896 13768 13930
rect 13802 13896 13844 13930
rect 13724 13862 13844 13896
rect 13724 13828 13768 13862
rect 13802 13828 13844 13862
rect 13724 13794 13844 13828
rect 13724 13760 13768 13794
rect 13802 13760 13844 13794
rect 13724 13726 13844 13760
rect 13724 13692 13768 13726
rect 13802 13692 13844 13726
rect 13724 13658 13844 13692
rect 13724 13624 13768 13658
rect 13802 13624 13844 13658
rect 13724 13590 13844 13624
rect 13724 13556 13768 13590
rect 13802 13556 13844 13590
rect 13724 13522 13844 13556
rect 13724 13488 13768 13522
rect 13802 13488 13844 13522
rect 13724 13454 13844 13488
rect 13724 13420 13768 13454
rect 13802 13420 13844 13454
rect 13724 13386 13844 13420
rect 13724 13352 13768 13386
rect 13802 13352 13844 13386
rect 13724 13318 13844 13352
rect 13724 13284 13768 13318
rect 13802 13284 13844 13318
rect 13724 13250 13844 13284
rect 13724 13216 13768 13250
rect 13802 13216 13844 13250
rect 13724 13182 13844 13216
rect 13724 13148 13768 13182
rect 13802 13148 13844 13182
rect 13724 13114 13844 13148
rect 13724 13080 13768 13114
rect 13802 13080 13844 13114
rect 13724 13046 13844 13080
rect 13724 13012 13768 13046
rect 13802 13012 13844 13046
rect 13724 12978 13844 13012
rect 13724 12944 13768 12978
rect 13802 12944 13844 12978
rect 13724 12910 13844 12944
rect 13724 12876 13768 12910
rect 13802 12876 13844 12910
rect 13724 12842 13844 12876
rect 13724 12808 13768 12842
rect 13802 12808 13844 12842
rect 13724 12774 13844 12808
rect 13724 12740 13768 12774
rect 13802 12740 13844 12774
rect 13724 12706 13844 12740
rect 13724 12672 13768 12706
rect 13802 12672 13844 12706
rect 13724 12638 13844 12672
rect 13724 12604 13768 12638
rect 13802 12604 13844 12638
rect 13724 12570 13844 12604
rect 13724 12536 13768 12570
rect 13802 12536 13844 12570
rect 13724 12502 13844 12536
rect 13724 12468 13768 12502
rect 13802 12468 13844 12502
rect 13724 12434 13844 12468
rect 13724 12400 13768 12434
rect 13802 12400 13844 12434
rect 13724 12366 13844 12400
rect 13724 12332 13768 12366
rect 13802 12332 13844 12366
rect 13724 12298 13844 12332
rect 13724 12264 13768 12298
rect 13802 12264 13844 12298
rect 13724 12230 13844 12264
rect 13724 12196 13768 12230
rect 13802 12196 13844 12230
rect 13724 12162 13844 12196
rect 13724 12128 13768 12162
rect 13802 12128 13844 12162
rect 13724 12094 13844 12128
rect 13724 12060 13768 12094
rect 13802 12060 13844 12094
rect 13724 12026 13844 12060
rect 13724 11992 13768 12026
rect 13802 11992 13844 12026
rect 13724 11958 13844 11992
rect 13724 11924 13768 11958
rect 13802 11924 13844 11958
rect 13724 11890 13844 11924
rect 13724 11856 13768 11890
rect 13802 11856 13844 11890
rect 13724 11822 13844 11856
rect 13724 11788 13768 11822
rect 13802 11788 13844 11822
rect 13724 11754 13844 11788
rect 13724 11720 13768 11754
rect 13802 11720 13844 11754
rect 13724 11686 13844 11720
rect 13724 11652 13768 11686
rect 13802 11652 13844 11686
rect 13724 11618 13844 11652
rect 13724 11584 13768 11618
rect 13802 11584 13844 11618
rect 13724 11550 13844 11584
rect 13724 11516 13768 11550
rect 13802 11516 13844 11550
rect 13724 11482 13844 11516
rect 13724 11448 13768 11482
rect 13802 11448 13844 11482
rect 13724 11414 13844 11448
rect 13724 11380 13768 11414
rect 13802 11380 13844 11414
rect 13724 11346 13844 11380
rect 13724 11312 13768 11346
rect 13802 11312 13844 11346
rect 13724 11278 13844 11312
rect 13724 11244 13768 11278
rect 13802 11244 13844 11278
rect 13724 11210 13844 11244
rect 13724 11176 13768 11210
rect 13802 11176 13844 11210
rect 13724 11142 13844 11176
rect 13724 11108 13768 11142
rect 13802 11108 13844 11142
rect 13724 11074 13844 11108
rect 13724 11040 13768 11074
rect 13802 11040 13844 11074
rect 13724 11006 13844 11040
rect 13724 10972 13768 11006
rect 13802 10972 13844 11006
rect 13724 10938 13844 10972
rect 13724 10904 13768 10938
rect 13802 10904 13844 10938
rect 13724 10870 13844 10904
rect 13724 10836 13768 10870
rect 13802 10836 13844 10870
rect 13724 10802 13844 10836
rect 13724 10768 13768 10802
rect 13802 10768 13844 10802
rect 13724 10734 13844 10768
rect 13724 10700 13768 10734
rect 13802 10700 13844 10734
rect 13724 10666 13844 10700
rect 13724 10632 13768 10666
rect 13802 10632 13844 10666
rect 13724 10598 13844 10632
rect 13724 10564 13768 10598
rect 13802 10564 13844 10598
rect 13724 10530 13844 10564
rect 13724 10496 13768 10530
rect 13802 10496 13844 10530
rect 13724 10462 13844 10496
rect 13724 10428 13768 10462
rect 13802 10428 13844 10462
rect 13724 10394 13844 10428
rect 13724 10362 13768 10394
rect 1148 10360 13768 10362
rect 13802 10360 13844 10394
rect 1148 10318 13844 10360
rect 1148 10284 1329 10318
rect 1363 10284 1397 10318
rect 1431 10284 1465 10318
rect 1499 10284 1533 10318
rect 1567 10284 1601 10318
rect 1635 10284 1669 10318
rect 1703 10284 1737 10318
rect 1771 10284 1805 10318
rect 1839 10284 1873 10318
rect 1907 10284 1941 10318
rect 1975 10284 2009 10318
rect 2043 10284 2077 10318
rect 2111 10284 2145 10318
rect 2179 10284 2213 10318
rect 2247 10284 2281 10318
rect 2315 10284 2349 10318
rect 2383 10284 2417 10318
rect 2451 10284 2485 10318
rect 2519 10284 2553 10318
rect 2587 10284 2621 10318
rect 2655 10284 2689 10318
rect 2723 10284 2757 10318
rect 2791 10284 2825 10318
rect 2859 10284 2893 10318
rect 2927 10284 2961 10318
rect 2995 10284 3029 10318
rect 3063 10284 3097 10318
rect 3131 10284 3165 10318
rect 3199 10284 3233 10318
rect 3267 10284 3301 10318
rect 3335 10284 3369 10318
rect 3403 10284 3437 10318
rect 3471 10284 3505 10318
rect 3539 10284 3573 10318
rect 3607 10284 3641 10318
rect 3675 10284 3709 10318
rect 3743 10284 3777 10318
rect 3811 10284 3845 10318
rect 3879 10284 3913 10318
rect 3947 10284 3981 10318
rect 4015 10284 4049 10318
rect 4083 10284 4117 10318
rect 4151 10284 4185 10318
rect 4219 10284 4253 10318
rect 4287 10284 4321 10318
rect 4355 10284 4389 10318
rect 4423 10284 4457 10318
rect 4491 10284 4525 10318
rect 4559 10284 4593 10318
rect 4627 10284 4661 10318
rect 4695 10284 4729 10318
rect 4763 10284 4797 10318
rect 4831 10284 4865 10318
rect 4899 10284 4933 10318
rect 4967 10284 5001 10318
rect 5035 10284 5069 10318
rect 5103 10284 5137 10318
rect 5171 10284 5205 10318
rect 5239 10284 5273 10318
rect 5307 10284 5341 10318
rect 5375 10284 5409 10318
rect 5443 10284 5477 10318
rect 5511 10284 5545 10318
rect 5579 10284 5613 10318
rect 5647 10284 5681 10318
rect 5715 10284 5749 10318
rect 5783 10284 5817 10318
rect 5851 10284 5885 10318
rect 5919 10284 5953 10318
rect 5987 10284 6021 10318
rect 6055 10284 6089 10318
rect 6123 10284 6157 10318
rect 6191 10284 6225 10318
rect 6259 10284 6293 10318
rect 6327 10284 6361 10318
rect 6395 10284 6429 10318
rect 6463 10284 6497 10318
rect 6531 10284 6565 10318
rect 6599 10284 6633 10318
rect 6667 10284 6701 10318
rect 6735 10284 6769 10318
rect 6803 10284 6837 10318
rect 6871 10284 6905 10318
rect 6939 10284 6973 10318
rect 7007 10284 7041 10318
rect 7075 10284 7109 10318
rect 7143 10284 7177 10318
rect 7211 10284 7245 10318
rect 7279 10284 7313 10318
rect 7347 10284 7381 10318
rect 7415 10284 7449 10318
rect 7483 10284 7517 10318
rect 7551 10284 7585 10318
rect 7619 10284 7653 10318
rect 7687 10284 7721 10318
rect 7755 10284 7789 10318
rect 7823 10284 7857 10318
rect 7891 10284 7925 10318
rect 7959 10284 7993 10318
rect 8027 10284 8061 10318
rect 8095 10284 8129 10318
rect 8163 10284 8197 10318
rect 8231 10284 8265 10318
rect 8299 10284 8333 10318
rect 8367 10284 8401 10318
rect 8435 10284 8469 10318
rect 8503 10284 8537 10318
rect 8571 10284 8605 10318
rect 8639 10284 8673 10318
rect 8707 10284 8741 10318
rect 8775 10284 8809 10318
rect 8843 10284 8877 10318
rect 8911 10284 8945 10318
rect 8979 10284 9013 10318
rect 9047 10284 9081 10318
rect 9115 10284 9149 10318
rect 9183 10284 9217 10318
rect 9251 10284 9285 10318
rect 9319 10284 9353 10318
rect 9387 10284 9421 10318
rect 9455 10284 9489 10318
rect 9523 10284 9557 10318
rect 9591 10284 9625 10318
rect 9659 10284 9693 10318
rect 9727 10284 9761 10318
rect 9795 10284 9829 10318
rect 9863 10284 9897 10318
rect 9931 10284 9965 10318
rect 9999 10284 10033 10318
rect 10067 10284 10101 10318
rect 10135 10284 10169 10318
rect 10203 10284 10237 10318
rect 10271 10284 10305 10318
rect 10339 10284 10373 10318
rect 10407 10284 10441 10318
rect 10475 10284 10509 10318
rect 10543 10284 10577 10318
rect 10611 10284 10645 10318
rect 10679 10284 10713 10318
rect 10747 10284 10781 10318
rect 10815 10284 10849 10318
rect 10883 10284 10917 10318
rect 10951 10284 10985 10318
rect 11019 10284 11053 10318
rect 11087 10284 11121 10318
rect 11155 10284 11189 10318
rect 11223 10284 11257 10318
rect 11291 10284 11325 10318
rect 11359 10284 11393 10318
rect 11427 10284 11461 10318
rect 11495 10284 11529 10318
rect 11563 10284 11597 10318
rect 11631 10284 11665 10318
rect 11699 10284 11733 10318
rect 11767 10284 11801 10318
rect 11835 10284 11869 10318
rect 11903 10284 11937 10318
rect 11971 10284 12005 10318
rect 12039 10284 12073 10318
rect 12107 10284 12141 10318
rect 12175 10284 12209 10318
rect 12243 10284 12277 10318
rect 12311 10284 12345 10318
rect 12379 10284 12413 10318
rect 12447 10284 12481 10318
rect 12515 10284 12549 10318
rect 12583 10284 12617 10318
rect 12651 10284 12685 10318
rect 12719 10284 12753 10318
rect 12787 10284 12821 10318
rect 12855 10284 12889 10318
rect 12923 10284 12957 10318
rect 12991 10284 13025 10318
rect 13059 10284 13093 10318
rect 13127 10284 13161 10318
rect 13195 10284 13229 10318
rect 13263 10284 13297 10318
rect 13331 10284 13365 10318
rect 13399 10284 13433 10318
rect 13467 10284 13501 10318
rect 13535 10284 13569 10318
rect 13603 10284 13637 10318
rect 13671 10284 13844 10318
rect 1148 10242 13844 10284
rect 14539 36207 14611 36241
rect 14645 36207 14724 36241
rect 14539 36173 14724 36207
rect 14539 36139 14611 36173
rect 14645 36139 14724 36173
rect 14539 36105 14724 36139
rect 14539 36071 14611 36105
rect 14645 36071 14724 36105
rect 14539 36037 14724 36071
rect 14539 36003 14611 36037
rect 14645 36003 14724 36037
rect 14539 35969 14724 36003
rect 14539 35935 14611 35969
rect 14645 35935 14724 35969
rect 14539 35901 14724 35935
rect 14539 35867 14611 35901
rect 14645 35867 14724 35901
rect 14539 35833 14724 35867
rect 14539 35799 14611 35833
rect 14645 35799 14724 35833
rect 14539 35765 14724 35799
rect 14539 35731 14611 35765
rect 14645 35731 14724 35765
rect 14539 35697 14724 35731
rect 14539 35663 14611 35697
rect 14645 35663 14724 35697
rect 14539 35629 14724 35663
rect 14539 35595 14611 35629
rect 14645 35595 14724 35629
rect 14539 35561 14724 35595
rect 14539 35527 14611 35561
rect 14645 35527 14724 35561
rect 14539 35493 14724 35527
rect 14539 35459 14611 35493
rect 14645 35459 14724 35493
rect 14539 35425 14724 35459
rect 14539 35391 14611 35425
rect 14645 35391 14724 35425
rect 14539 35357 14724 35391
rect 14539 35323 14611 35357
rect 14645 35323 14724 35357
rect 14539 35289 14724 35323
rect 14539 35255 14611 35289
rect 14645 35255 14724 35289
rect 14539 35221 14724 35255
rect 14539 35187 14611 35221
rect 14645 35187 14724 35221
rect 14539 35153 14724 35187
rect 14539 35119 14611 35153
rect 14645 35119 14724 35153
rect 14539 35085 14724 35119
rect 14539 35051 14611 35085
rect 14645 35051 14724 35085
rect 14539 35017 14724 35051
rect 14539 34983 14611 35017
rect 14645 34983 14724 35017
rect 14539 34949 14724 34983
rect 14539 34915 14611 34949
rect 14645 34915 14724 34949
rect 14539 34881 14724 34915
rect 14539 34847 14611 34881
rect 14645 34847 14724 34881
rect 14539 34813 14724 34847
rect 14539 34779 14611 34813
rect 14645 34779 14724 34813
rect 14539 34745 14724 34779
rect 14539 34711 14611 34745
rect 14645 34711 14724 34745
rect 14539 34677 14724 34711
rect 14539 34643 14611 34677
rect 14645 34643 14724 34677
rect 14539 34609 14724 34643
rect 14539 34575 14611 34609
rect 14645 34575 14724 34609
rect 14539 34541 14724 34575
rect 14539 34507 14611 34541
rect 14645 34507 14724 34541
rect 14539 34473 14724 34507
rect 14539 34439 14611 34473
rect 14645 34439 14724 34473
rect 14539 34405 14724 34439
rect 14539 34371 14611 34405
rect 14645 34371 14724 34405
rect 14539 34337 14724 34371
rect 14539 34303 14611 34337
rect 14645 34303 14724 34337
rect 14539 34269 14724 34303
rect 14539 34235 14611 34269
rect 14645 34235 14724 34269
rect 14539 34201 14724 34235
rect 14539 34167 14611 34201
rect 14645 34167 14724 34201
rect 14539 34133 14724 34167
rect 14539 34099 14611 34133
rect 14645 34099 14724 34133
rect 14539 34065 14724 34099
rect 14539 34031 14611 34065
rect 14645 34031 14724 34065
rect 14539 33997 14724 34031
rect 14539 33963 14611 33997
rect 14645 33963 14724 33997
rect 14539 33929 14724 33963
rect 14539 33895 14611 33929
rect 14645 33895 14724 33929
rect 14539 33861 14724 33895
rect 14539 33827 14611 33861
rect 14645 33827 14724 33861
rect 14539 33793 14724 33827
rect 14539 33759 14611 33793
rect 14645 33759 14724 33793
rect 14539 33725 14724 33759
rect 14539 33691 14611 33725
rect 14645 33691 14724 33725
rect 14539 33657 14724 33691
rect 14539 33623 14611 33657
rect 14645 33623 14724 33657
rect 14539 33589 14724 33623
rect 14539 33555 14611 33589
rect 14645 33555 14724 33589
rect 14539 33521 14724 33555
rect 14539 33487 14611 33521
rect 14645 33487 14724 33521
rect 14539 33453 14724 33487
rect 14539 33419 14611 33453
rect 14645 33419 14724 33453
rect 14539 33385 14724 33419
rect 14539 33351 14611 33385
rect 14645 33351 14724 33385
rect 14539 33317 14724 33351
rect 14539 33283 14611 33317
rect 14645 33283 14724 33317
rect 14539 33249 14724 33283
rect 14539 33215 14611 33249
rect 14645 33215 14724 33249
rect 14539 33181 14724 33215
rect 14539 33147 14611 33181
rect 14645 33147 14724 33181
rect 14539 33113 14724 33147
rect 14539 33079 14611 33113
rect 14645 33079 14724 33113
rect 14539 33045 14724 33079
rect 14539 33011 14611 33045
rect 14645 33011 14724 33045
rect 14539 32977 14724 33011
rect 14539 32943 14611 32977
rect 14645 32943 14724 32977
rect 14539 32909 14724 32943
rect 14539 32875 14611 32909
rect 14645 32875 14724 32909
rect 14539 32841 14724 32875
rect 14539 32807 14611 32841
rect 14645 32807 14724 32841
rect 14539 32773 14724 32807
rect 14539 32739 14611 32773
rect 14645 32739 14724 32773
rect 14539 32705 14724 32739
rect 14539 32671 14611 32705
rect 14645 32671 14724 32705
rect 14539 32637 14724 32671
rect 14539 32603 14611 32637
rect 14645 32603 14724 32637
rect 14539 32569 14724 32603
rect 14539 32535 14611 32569
rect 14645 32535 14724 32569
rect 14539 32501 14724 32535
rect 14539 32467 14611 32501
rect 14645 32467 14724 32501
rect 14539 32433 14724 32467
rect 14539 32399 14611 32433
rect 14645 32399 14724 32433
rect 14539 32365 14724 32399
rect 14539 32331 14611 32365
rect 14645 32331 14724 32365
rect 14539 32297 14724 32331
rect 14539 32263 14611 32297
rect 14645 32263 14724 32297
rect 14539 32229 14724 32263
rect 14539 32195 14611 32229
rect 14645 32195 14724 32229
rect 14539 32161 14724 32195
rect 14539 32127 14611 32161
rect 14645 32127 14724 32161
rect 14539 32093 14724 32127
rect 14539 32059 14611 32093
rect 14645 32059 14724 32093
rect 14539 32025 14724 32059
rect 14539 31991 14611 32025
rect 14645 31991 14724 32025
rect 14539 31957 14724 31991
rect 14539 31923 14611 31957
rect 14645 31923 14724 31957
rect 14539 31889 14724 31923
rect 14539 31855 14611 31889
rect 14645 31855 14724 31889
rect 14539 31821 14724 31855
rect 14539 31787 14611 31821
rect 14645 31787 14724 31821
rect 14539 31753 14724 31787
rect 14539 31719 14611 31753
rect 14645 31719 14724 31753
rect 14539 31685 14724 31719
rect 14539 31651 14611 31685
rect 14645 31651 14724 31685
rect 14539 31617 14724 31651
rect 14539 31583 14611 31617
rect 14645 31583 14724 31617
rect 14539 31549 14724 31583
rect 14539 31515 14611 31549
rect 14645 31515 14724 31549
rect 14539 31481 14724 31515
rect 14539 31447 14611 31481
rect 14645 31447 14724 31481
rect 14539 31413 14724 31447
rect 14539 31379 14611 31413
rect 14645 31379 14724 31413
rect 14539 31345 14724 31379
rect 14539 31311 14611 31345
rect 14645 31311 14724 31345
rect 14539 31277 14724 31311
rect 14539 31243 14611 31277
rect 14645 31243 14724 31277
rect 14539 31209 14724 31243
rect 14539 31175 14611 31209
rect 14645 31175 14724 31209
rect 14539 31141 14724 31175
rect 14539 31107 14611 31141
rect 14645 31107 14724 31141
rect 14539 31073 14724 31107
rect 14539 31039 14611 31073
rect 14645 31039 14724 31073
rect 14539 31005 14724 31039
rect 14539 30971 14611 31005
rect 14645 30971 14724 31005
rect 14539 30937 14724 30971
rect 14539 30903 14611 30937
rect 14645 30903 14724 30937
rect 14539 30869 14724 30903
rect 14539 30835 14611 30869
rect 14645 30835 14724 30869
rect 14539 30801 14724 30835
rect 14539 30767 14611 30801
rect 14645 30767 14724 30801
rect 14539 30733 14724 30767
rect 14539 30699 14611 30733
rect 14645 30699 14724 30733
rect 14539 30665 14724 30699
rect 14539 30631 14611 30665
rect 14645 30631 14724 30665
rect 14539 30597 14724 30631
rect 14539 30563 14611 30597
rect 14645 30563 14724 30597
rect 14539 30529 14724 30563
rect 14539 30495 14611 30529
rect 14645 30495 14724 30529
rect 14539 30461 14724 30495
rect 14539 30427 14611 30461
rect 14645 30427 14724 30461
rect 14539 30393 14724 30427
rect 14539 30359 14611 30393
rect 14645 30359 14724 30393
rect 14539 30325 14724 30359
rect 14539 30291 14611 30325
rect 14645 30291 14724 30325
rect 14539 30257 14724 30291
rect 14539 30223 14611 30257
rect 14645 30223 14724 30257
rect 14539 30189 14724 30223
rect 14539 30155 14611 30189
rect 14645 30155 14724 30189
rect 14539 30121 14724 30155
rect 14539 30087 14611 30121
rect 14645 30087 14724 30121
rect 14539 30053 14724 30087
rect 14539 30019 14611 30053
rect 14645 30019 14724 30053
rect 14539 29985 14724 30019
rect 14539 29951 14611 29985
rect 14645 29951 14724 29985
rect 14539 29917 14724 29951
rect 14539 29883 14611 29917
rect 14645 29883 14724 29917
rect 14539 29849 14724 29883
rect 14539 29815 14611 29849
rect 14645 29815 14724 29849
rect 14539 29781 14724 29815
rect 14539 29747 14611 29781
rect 14645 29747 14724 29781
rect 14539 29713 14724 29747
rect 14539 29679 14611 29713
rect 14645 29679 14724 29713
rect 14539 29645 14724 29679
rect 14539 29611 14611 29645
rect 14645 29611 14724 29645
rect 14539 29577 14724 29611
rect 14539 29543 14611 29577
rect 14645 29543 14724 29577
rect 14539 29509 14724 29543
rect 14539 29475 14611 29509
rect 14645 29475 14724 29509
rect 14539 29441 14724 29475
rect 14539 29407 14611 29441
rect 14645 29407 14724 29441
rect 14539 29373 14724 29407
rect 14539 29339 14611 29373
rect 14645 29339 14724 29373
rect 14539 29305 14724 29339
rect 14539 29271 14611 29305
rect 14645 29271 14724 29305
rect 14539 29237 14724 29271
rect 14539 29203 14611 29237
rect 14645 29203 14724 29237
rect 14539 29169 14724 29203
rect 14539 29135 14611 29169
rect 14645 29135 14724 29169
rect 14539 29101 14724 29135
rect 14539 29067 14611 29101
rect 14645 29067 14724 29101
rect 14539 29033 14724 29067
rect 14539 28999 14611 29033
rect 14645 28999 14724 29033
rect 14539 28965 14724 28999
rect 14539 28931 14611 28965
rect 14645 28931 14724 28965
rect 14539 28897 14724 28931
rect 14539 28863 14611 28897
rect 14645 28863 14724 28897
rect 14539 28829 14724 28863
rect 14539 28795 14611 28829
rect 14645 28795 14724 28829
rect 14539 28761 14724 28795
rect 14539 28727 14611 28761
rect 14645 28727 14724 28761
rect 14539 28693 14724 28727
rect 14539 28659 14611 28693
rect 14645 28659 14724 28693
rect 14539 28625 14724 28659
rect 14539 28591 14611 28625
rect 14645 28591 14724 28625
rect 14539 28557 14724 28591
rect 14539 28523 14611 28557
rect 14645 28523 14724 28557
rect 14539 28489 14724 28523
rect 14539 28455 14611 28489
rect 14645 28455 14724 28489
rect 14539 28421 14724 28455
rect 14539 28387 14611 28421
rect 14645 28387 14724 28421
rect 14539 28353 14724 28387
rect 14539 28319 14611 28353
rect 14645 28319 14724 28353
rect 14539 28285 14724 28319
rect 14539 28251 14611 28285
rect 14645 28251 14724 28285
rect 14539 28217 14724 28251
rect 14539 28183 14611 28217
rect 14645 28183 14724 28217
rect 14539 28149 14724 28183
rect 14539 28115 14611 28149
rect 14645 28115 14724 28149
rect 14539 28081 14724 28115
rect 14539 28047 14611 28081
rect 14645 28047 14724 28081
rect 14539 28013 14724 28047
rect 14539 27979 14611 28013
rect 14645 27979 14724 28013
rect 14539 27945 14724 27979
rect 14539 27911 14611 27945
rect 14645 27911 14724 27945
rect 14539 27877 14724 27911
rect 14539 27843 14611 27877
rect 14645 27843 14724 27877
rect 14539 27809 14724 27843
rect 14539 27775 14611 27809
rect 14645 27775 14724 27809
rect 14539 27741 14724 27775
rect 14539 27707 14611 27741
rect 14645 27707 14724 27741
rect 14539 27673 14724 27707
rect 14539 27639 14611 27673
rect 14645 27639 14724 27673
rect 14539 27605 14724 27639
rect 14539 27571 14611 27605
rect 14645 27571 14724 27605
rect 14539 27537 14724 27571
rect 14539 27503 14611 27537
rect 14645 27503 14724 27537
rect 14539 27469 14724 27503
rect 14539 27435 14611 27469
rect 14645 27435 14724 27469
rect 14539 27401 14724 27435
rect 14539 27367 14611 27401
rect 14645 27367 14724 27401
rect 14539 27333 14724 27367
rect 14539 27299 14611 27333
rect 14645 27299 14724 27333
rect 14539 27265 14724 27299
rect 14539 27231 14611 27265
rect 14645 27231 14724 27265
rect 14539 27197 14724 27231
rect 14539 27163 14611 27197
rect 14645 27163 14724 27197
rect 14539 27129 14724 27163
rect 14539 27095 14611 27129
rect 14645 27095 14724 27129
rect 14539 27061 14724 27095
rect 14539 27027 14611 27061
rect 14645 27027 14724 27061
rect 14539 26993 14724 27027
rect 14539 26959 14611 26993
rect 14645 26959 14724 26993
rect 14539 26925 14724 26959
rect 14539 26891 14611 26925
rect 14645 26891 14724 26925
rect 14539 26857 14724 26891
rect 14539 26823 14611 26857
rect 14645 26823 14724 26857
rect 14539 26789 14724 26823
rect 14539 26755 14611 26789
rect 14645 26755 14724 26789
rect 14539 26721 14724 26755
rect 14539 26687 14611 26721
rect 14645 26687 14724 26721
rect 14539 26653 14724 26687
rect 14539 26619 14611 26653
rect 14645 26619 14724 26653
rect 14539 26585 14724 26619
rect 14539 26551 14611 26585
rect 14645 26551 14724 26585
rect 14539 26517 14724 26551
rect 14539 26483 14611 26517
rect 14645 26483 14724 26517
rect 14539 26449 14724 26483
rect 14539 26415 14611 26449
rect 14645 26415 14724 26449
rect 14539 26381 14724 26415
rect 14539 26347 14611 26381
rect 14645 26347 14724 26381
rect 14539 26313 14724 26347
rect 14539 26279 14611 26313
rect 14645 26279 14724 26313
rect 14539 26245 14724 26279
rect 14539 26211 14611 26245
rect 14645 26211 14724 26245
rect 14539 26177 14724 26211
rect 14539 26143 14611 26177
rect 14645 26143 14724 26177
rect 14539 26109 14724 26143
rect 14539 26075 14611 26109
rect 14645 26075 14724 26109
rect 14539 26041 14724 26075
rect 14539 26007 14611 26041
rect 14645 26007 14724 26041
rect 14539 25973 14724 26007
rect 14539 25939 14611 25973
rect 14645 25939 14724 25973
rect 14539 25905 14724 25939
rect 14539 25871 14611 25905
rect 14645 25871 14724 25905
rect 14539 25837 14724 25871
rect 14539 25803 14611 25837
rect 14645 25803 14724 25837
rect 14539 25769 14724 25803
rect 14539 25735 14611 25769
rect 14645 25735 14724 25769
rect 14539 25701 14724 25735
rect 14539 25667 14611 25701
rect 14645 25667 14724 25701
rect 14539 25633 14724 25667
rect 14539 25599 14611 25633
rect 14645 25599 14724 25633
rect 14539 25565 14724 25599
rect 14539 25531 14611 25565
rect 14645 25531 14724 25565
rect 14539 25497 14724 25531
rect 14539 25463 14611 25497
rect 14645 25463 14724 25497
rect 14539 25429 14724 25463
rect 14539 25395 14611 25429
rect 14645 25395 14724 25429
rect 14539 25361 14724 25395
rect 14539 25327 14611 25361
rect 14645 25327 14724 25361
rect 14539 25293 14724 25327
rect 14539 25259 14611 25293
rect 14645 25259 14724 25293
rect 14539 25225 14724 25259
rect 14539 25191 14611 25225
rect 14645 25191 14724 25225
rect 14539 25157 14724 25191
rect 14539 25123 14611 25157
rect 14645 25123 14724 25157
rect 14539 25089 14724 25123
rect 14539 25055 14611 25089
rect 14645 25055 14724 25089
rect 14539 25021 14724 25055
rect 14539 24987 14611 25021
rect 14645 24987 14724 25021
rect 14539 24953 14724 24987
rect 14539 24919 14611 24953
rect 14645 24919 14724 24953
rect 14539 24885 14724 24919
rect 14539 24851 14611 24885
rect 14645 24851 14724 24885
rect 14539 24817 14724 24851
rect 14539 24783 14611 24817
rect 14645 24783 14724 24817
rect 14539 24749 14724 24783
rect 14539 24715 14611 24749
rect 14645 24715 14724 24749
rect 14539 24681 14724 24715
rect 14539 24647 14611 24681
rect 14645 24647 14724 24681
rect 14539 24613 14724 24647
rect 14539 24579 14611 24613
rect 14645 24579 14724 24613
rect 14539 24545 14724 24579
rect 14539 24511 14611 24545
rect 14645 24511 14724 24545
rect 14539 24477 14724 24511
rect 14539 24443 14611 24477
rect 14645 24443 14724 24477
rect 14539 24409 14724 24443
rect 14539 24375 14611 24409
rect 14645 24375 14724 24409
rect 14539 24341 14724 24375
rect 14539 24307 14611 24341
rect 14645 24307 14724 24341
rect 14539 24273 14724 24307
rect 14539 24239 14611 24273
rect 14645 24239 14724 24273
rect 14539 24205 14724 24239
rect 14539 24171 14611 24205
rect 14645 24171 14724 24205
rect 14539 24137 14724 24171
rect 14539 24103 14611 24137
rect 14645 24103 14724 24137
rect 14539 24069 14724 24103
rect 14539 24035 14611 24069
rect 14645 24035 14724 24069
rect 14539 24001 14724 24035
rect 14539 23967 14611 24001
rect 14645 23967 14724 24001
rect 14539 23933 14724 23967
rect 14539 23899 14611 23933
rect 14645 23899 14724 23933
rect 14539 23865 14724 23899
rect 14539 23831 14611 23865
rect 14645 23831 14724 23865
rect 14539 23797 14724 23831
rect 14539 23763 14611 23797
rect 14645 23763 14724 23797
rect 14539 23729 14724 23763
rect 14539 23695 14611 23729
rect 14645 23695 14724 23729
rect 14539 23661 14724 23695
rect 14539 23627 14611 23661
rect 14645 23627 14724 23661
rect 14539 23593 14724 23627
rect 14539 23559 14611 23593
rect 14645 23559 14724 23593
rect 14539 23525 14724 23559
rect 14539 23491 14611 23525
rect 14645 23491 14724 23525
rect 14539 23457 14724 23491
rect 14539 23423 14611 23457
rect 14645 23423 14724 23457
rect 14539 23389 14724 23423
rect 14539 23355 14611 23389
rect 14645 23355 14724 23389
rect 14539 23321 14724 23355
rect 14539 23287 14611 23321
rect 14645 23287 14724 23321
rect 14539 23253 14724 23287
rect 14539 23219 14611 23253
rect 14645 23219 14724 23253
rect 14539 23185 14724 23219
rect 14539 23151 14611 23185
rect 14645 23151 14724 23185
rect 14539 23117 14724 23151
rect 14539 23083 14611 23117
rect 14645 23083 14724 23117
rect 14539 23049 14724 23083
rect 14539 23015 14611 23049
rect 14645 23015 14724 23049
rect 14539 22981 14724 23015
rect 14539 22947 14611 22981
rect 14645 22947 14724 22981
rect 14539 22913 14724 22947
rect 14539 22879 14611 22913
rect 14645 22879 14724 22913
rect 14539 22845 14724 22879
rect 14539 22811 14611 22845
rect 14645 22811 14724 22845
rect 14539 22777 14724 22811
rect 14539 22743 14611 22777
rect 14645 22743 14724 22777
rect 14539 22709 14724 22743
rect 14539 22675 14611 22709
rect 14645 22675 14724 22709
rect 14539 22641 14724 22675
rect 14539 22607 14611 22641
rect 14645 22607 14724 22641
rect 14539 22573 14724 22607
rect 14539 22539 14611 22573
rect 14645 22539 14724 22573
rect 14539 22505 14724 22539
rect 14539 22471 14611 22505
rect 14645 22471 14724 22505
rect 14539 22437 14724 22471
rect 14539 22403 14611 22437
rect 14645 22403 14724 22437
rect 14539 22369 14724 22403
rect 14539 22335 14611 22369
rect 14645 22335 14724 22369
rect 14539 22301 14724 22335
rect 14539 22267 14611 22301
rect 14645 22267 14724 22301
rect 14539 22233 14724 22267
rect 14539 22199 14611 22233
rect 14645 22199 14724 22233
rect 14539 22165 14724 22199
rect 14539 22131 14611 22165
rect 14645 22131 14724 22165
rect 14539 22097 14724 22131
rect 14539 22063 14611 22097
rect 14645 22063 14724 22097
rect 14539 22029 14724 22063
rect 14539 21995 14611 22029
rect 14645 21995 14724 22029
rect 14539 21961 14724 21995
rect 14539 21927 14611 21961
rect 14645 21927 14724 21961
rect 14539 21893 14724 21927
rect 14539 21859 14611 21893
rect 14645 21859 14724 21893
rect 14539 21825 14724 21859
rect 14539 21791 14611 21825
rect 14645 21791 14724 21825
rect 14539 21757 14724 21791
rect 14539 21723 14611 21757
rect 14645 21723 14724 21757
rect 14539 21689 14724 21723
rect 14539 21655 14611 21689
rect 14645 21655 14724 21689
rect 14539 21621 14724 21655
rect 14539 21587 14611 21621
rect 14645 21587 14724 21621
rect 14539 21553 14724 21587
rect 14539 21519 14611 21553
rect 14645 21519 14724 21553
rect 14539 21485 14724 21519
rect 14539 21451 14611 21485
rect 14645 21451 14724 21485
rect 14539 21417 14724 21451
rect 14539 21383 14611 21417
rect 14645 21383 14724 21417
rect 14539 21349 14724 21383
rect 14539 21315 14611 21349
rect 14645 21315 14724 21349
rect 14539 21281 14724 21315
rect 14539 21247 14611 21281
rect 14645 21247 14724 21281
rect 14539 21213 14724 21247
rect 14539 21179 14611 21213
rect 14645 21179 14724 21213
rect 14539 21145 14724 21179
rect 14539 21111 14611 21145
rect 14645 21111 14724 21145
rect 14539 21077 14724 21111
rect 14539 21043 14611 21077
rect 14645 21043 14724 21077
rect 14539 21009 14724 21043
rect 14539 20975 14611 21009
rect 14645 20975 14724 21009
rect 14539 20941 14724 20975
rect 14539 20907 14611 20941
rect 14645 20907 14724 20941
rect 14539 20873 14724 20907
rect 14539 20839 14611 20873
rect 14645 20839 14724 20873
rect 14539 20805 14724 20839
rect 14539 20771 14611 20805
rect 14645 20771 14724 20805
rect 14539 20737 14724 20771
rect 14539 20703 14611 20737
rect 14645 20703 14724 20737
rect 14539 20669 14724 20703
rect 14539 20635 14611 20669
rect 14645 20635 14724 20669
rect 14539 20601 14724 20635
rect 14539 20567 14611 20601
rect 14645 20567 14724 20601
rect 14539 20533 14724 20567
rect 14539 20499 14611 20533
rect 14645 20499 14724 20533
rect 14539 20465 14724 20499
rect 14539 20431 14611 20465
rect 14645 20431 14724 20465
rect 14539 20397 14724 20431
rect 14539 20363 14611 20397
rect 14645 20363 14724 20397
rect 14539 20329 14724 20363
rect 14539 20295 14611 20329
rect 14645 20295 14724 20329
rect 14539 20261 14724 20295
rect 14539 20227 14611 20261
rect 14645 20227 14724 20261
rect 14539 20193 14724 20227
rect 14539 20159 14611 20193
rect 14645 20159 14724 20193
rect 14539 20125 14724 20159
rect 14539 20091 14611 20125
rect 14645 20091 14724 20125
rect 14539 20057 14724 20091
rect 14539 20023 14611 20057
rect 14645 20023 14724 20057
rect 14539 19989 14724 20023
rect 14539 19955 14611 19989
rect 14645 19955 14724 19989
rect 14539 19921 14724 19955
rect 14539 19887 14611 19921
rect 14645 19887 14724 19921
rect 14539 19853 14724 19887
rect 14539 19819 14611 19853
rect 14645 19819 14724 19853
rect 14539 19785 14724 19819
rect 14539 19751 14611 19785
rect 14645 19751 14724 19785
rect 14539 19717 14724 19751
rect 14539 19683 14611 19717
rect 14645 19683 14724 19717
rect 14539 19649 14724 19683
rect 14539 19615 14611 19649
rect 14645 19615 14724 19649
rect 14539 19581 14724 19615
rect 14539 19547 14611 19581
rect 14645 19547 14724 19581
rect 14539 19513 14724 19547
rect 14539 19479 14611 19513
rect 14645 19479 14724 19513
rect 14539 19445 14724 19479
rect 14539 19411 14611 19445
rect 14645 19411 14724 19445
rect 14539 19377 14724 19411
rect 14539 19343 14611 19377
rect 14645 19343 14724 19377
rect 14539 19309 14724 19343
rect 14539 19275 14611 19309
rect 14645 19275 14724 19309
rect 14539 19241 14724 19275
rect 14539 19207 14611 19241
rect 14645 19207 14724 19241
rect 14539 19173 14724 19207
rect 14539 19139 14611 19173
rect 14645 19139 14724 19173
rect 14539 19105 14724 19139
rect 14539 19071 14611 19105
rect 14645 19071 14724 19105
rect 14539 19037 14724 19071
rect 14539 19003 14611 19037
rect 14645 19003 14724 19037
rect 14539 18969 14724 19003
rect 14539 18935 14611 18969
rect 14645 18935 14724 18969
rect 14539 18901 14724 18935
rect 14539 18867 14611 18901
rect 14645 18867 14724 18901
rect 14539 18833 14724 18867
rect 14539 18799 14611 18833
rect 14645 18799 14724 18833
rect 14539 18765 14724 18799
rect 14539 18731 14611 18765
rect 14645 18731 14724 18765
rect 14539 18697 14724 18731
rect 14539 18663 14611 18697
rect 14645 18663 14724 18697
rect 14539 18629 14724 18663
rect 14539 18595 14611 18629
rect 14645 18595 14724 18629
rect 14539 18561 14724 18595
rect 14539 18527 14611 18561
rect 14645 18527 14724 18561
rect 14539 18493 14724 18527
rect 14539 18459 14611 18493
rect 14645 18459 14724 18493
rect 14539 18425 14724 18459
rect 14539 18391 14611 18425
rect 14645 18391 14724 18425
rect 14539 18357 14724 18391
rect 14539 18323 14611 18357
rect 14645 18323 14724 18357
rect 14539 18289 14724 18323
rect 14539 18255 14611 18289
rect 14645 18255 14724 18289
rect 14539 18221 14724 18255
rect 14539 18187 14611 18221
rect 14645 18187 14724 18221
rect 14539 18153 14724 18187
rect 14539 18119 14611 18153
rect 14645 18119 14724 18153
rect 14539 18085 14724 18119
rect 14539 18051 14611 18085
rect 14645 18051 14724 18085
rect 14539 18017 14724 18051
rect 14539 17983 14611 18017
rect 14645 17983 14724 18017
rect 14539 17949 14724 17983
rect 14539 17915 14611 17949
rect 14645 17915 14724 17949
rect 14539 17881 14724 17915
rect 14539 17847 14611 17881
rect 14645 17847 14724 17881
rect 14539 17813 14724 17847
rect 14539 17779 14611 17813
rect 14645 17779 14724 17813
rect 14539 17745 14724 17779
rect 14539 17711 14611 17745
rect 14645 17711 14724 17745
rect 14539 17677 14724 17711
rect 14539 17643 14611 17677
rect 14645 17643 14724 17677
rect 14539 17609 14724 17643
rect 14539 17575 14611 17609
rect 14645 17575 14724 17609
rect 14539 17541 14724 17575
rect 14539 17507 14611 17541
rect 14645 17507 14724 17541
rect 14539 17473 14724 17507
rect 14539 17439 14611 17473
rect 14645 17439 14724 17473
rect 14539 17405 14724 17439
rect 14539 17371 14611 17405
rect 14645 17371 14724 17405
rect 14539 17337 14724 17371
rect 14539 17303 14611 17337
rect 14645 17303 14724 17337
rect 14539 17269 14724 17303
rect 14539 17235 14611 17269
rect 14645 17235 14724 17269
rect 14539 17201 14724 17235
rect 14539 17167 14611 17201
rect 14645 17167 14724 17201
rect 14539 17133 14724 17167
rect 14539 17099 14611 17133
rect 14645 17099 14724 17133
rect 14539 17065 14724 17099
rect 14539 17031 14611 17065
rect 14645 17031 14724 17065
rect 14539 16997 14724 17031
rect 14539 16963 14611 16997
rect 14645 16963 14724 16997
rect 14539 16929 14724 16963
rect 14539 16895 14611 16929
rect 14645 16895 14724 16929
rect 14539 16861 14724 16895
rect 14539 16827 14611 16861
rect 14645 16827 14724 16861
rect 14539 16793 14724 16827
rect 14539 16759 14611 16793
rect 14645 16759 14724 16793
rect 14539 16725 14724 16759
rect 14539 16691 14611 16725
rect 14645 16691 14724 16725
rect 14539 16657 14724 16691
rect 14539 16623 14611 16657
rect 14645 16623 14724 16657
rect 14539 16589 14724 16623
rect 14539 16555 14611 16589
rect 14645 16555 14724 16589
rect 14539 16521 14724 16555
rect 14539 16487 14611 16521
rect 14645 16487 14724 16521
rect 14539 16453 14724 16487
rect 14539 16419 14611 16453
rect 14645 16419 14724 16453
rect 14539 16385 14724 16419
rect 14539 16351 14611 16385
rect 14645 16351 14724 16385
rect 14539 16317 14724 16351
rect 14539 16283 14611 16317
rect 14645 16283 14724 16317
rect 14539 16249 14724 16283
rect 14539 16215 14611 16249
rect 14645 16215 14724 16249
rect 14539 16181 14724 16215
rect 14539 16147 14611 16181
rect 14645 16147 14724 16181
rect 14539 16113 14724 16147
rect 14539 16079 14611 16113
rect 14645 16079 14724 16113
rect 14539 16045 14724 16079
rect 14539 16011 14611 16045
rect 14645 16011 14724 16045
rect 14539 15977 14724 16011
rect 14539 15943 14611 15977
rect 14645 15943 14724 15977
rect 14539 15909 14724 15943
rect 14539 15875 14611 15909
rect 14645 15875 14724 15909
rect 14539 15841 14724 15875
rect 14539 15807 14611 15841
rect 14645 15807 14724 15841
rect 14539 15773 14724 15807
rect 14539 15739 14611 15773
rect 14645 15739 14724 15773
rect 14539 15705 14724 15739
rect 14539 15671 14611 15705
rect 14645 15671 14724 15705
rect 14539 15637 14724 15671
rect 14539 15603 14611 15637
rect 14645 15603 14724 15637
rect 14539 15569 14724 15603
rect 14539 15535 14611 15569
rect 14645 15535 14724 15569
rect 14539 15501 14724 15535
rect 14539 15467 14611 15501
rect 14645 15467 14724 15501
rect 14539 15433 14724 15467
rect 14539 15399 14611 15433
rect 14645 15399 14724 15433
rect 14539 15365 14724 15399
rect 14539 15331 14611 15365
rect 14645 15331 14724 15365
rect 14539 15297 14724 15331
rect 14539 15263 14611 15297
rect 14645 15263 14724 15297
rect 14539 15229 14724 15263
rect 14539 15195 14611 15229
rect 14645 15195 14724 15229
rect 14539 15161 14724 15195
rect 14539 15127 14611 15161
rect 14645 15127 14724 15161
rect 14539 15093 14724 15127
rect 14539 15059 14611 15093
rect 14645 15059 14724 15093
rect 14539 15025 14724 15059
rect 14539 14991 14611 15025
rect 14645 14991 14724 15025
rect 14539 14957 14724 14991
rect 14539 14923 14611 14957
rect 14645 14923 14724 14957
rect 14539 14889 14724 14923
rect 14539 14855 14611 14889
rect 14645 14855 14724 14889
rect 14539 14821 14724 14855
rect 14539 14787 14611 14821
rect 14645 14787 14724 14821
rect 14539 14753 14724 14787
rect 14539 14719 14611 14753
rect 14645 14719 14724 14753
rect 14539 14685 14724 14719
rect 14539 14651 14611 14685
rect 14645 14651 14724 14685
rect 14539 14617 14724 14651
rect 14539 14583 14611 14617
rect 14645 14583 14724 14617
rect 14539 14549 14724 14583
rect 14539 14515 14611 14549
rect 14645 14515 14724 14549
rect 14539 14481 14724 14515
rect 14539 14447 14611 14481
rect 14645 14447 14724 14481
rect 14539 14413 14724 14447
rect 14539 14379 14611 14413
rect 14645 14379 14724 14413
rect 14539 14345 14724 14379
rect 14539 14311 14611 14345
rect 14645 14311 14724 14345
rect 14539 14277 14724 14311
rect 14539 14243 14611 14277
rect 14645 14243 14724 14277
rect 14539 14209 14724 14243
rect 14539 14175 14611 14209
rect 14645 14175 14724 14209
rect 14539 14141 14724 14175
rect 14539 14107 14611 14141
rect 14645 14107 14724 14141
rect 14539 14073 14724 14107
rect 14539 14039 14611 14073
rect 14645 14039 14724 14073
rect 14539 14005 14724 14039
rect 14539 13971 14611 14005
rect 14645 13971 14724 14005
rect 14539 13937 14724 13971
rect 14539 13903 14611 13937
rect 14645 13903 14724 13937
rect 14539 13869 14724 13903
rect 14539 13835 14611 13869
rect 14645 13835 14724 13869
rect 14539 13801 14724 13835
rect 14539 13767 14611 13801
rect 14645 13767 14724 13801
rect 14539 13733 14724 13767
rect 14539 13699 14611 13733
rect 14645 13699 14724 13733
rect 14539 13665 14724 13699
rect 14539 13631 14611 13665
rect 14645 13631 14724 13665
rect 14539 13597 14724 13631
rect 14539 13563 14611 13597
rect 14645 13563 14724 13597
rect 14539 13529 14724 13563
rect 14539 13495 14611 13529
rect 14645 13495 14724 13529
rect 14539 13461 14724 13495
rect 14539 13427 14611 13461
rect 14645 13427 14724 13461
rect 14539 13393 14724 13427
rect 14539 13359 14611 13393
rect 14645 13359 14724 13393
rect 14539 13325 14724 13359
rect 14539 13291 14611 13325
rect 14645 13291 14724 13325
rect 14539 13257 14724 13291
rect 14539 13223 14611 13257
rect 14645 13223 14724 13257
rect 14539 13189 14724 13223
rect 14539 13155 14611 13189
rect 14645 13155 14724 13189
rect 14539 13121 14724 13155
rect 14539 13087 14611 13121
rect 14645 13087 14724 13121
rect 14539 13053 14724 13087
rect 14539 13019 14611 13053
rect 14645 13019 14724 13053
rect 14539 12985 14724 13019
rect 14539 12951 14611 12985
rect 14645 12951 14724 12985
rect 14539 12917 14724 12951
rect 14539 12883 14611 12917
rect 14645 12883 14724 12917
rect 14539 12849 14724 12883
rect 14539 12815 14611 12849
rect 14645 12815 14724 12849
rect 14539 12781 14724 12815
rect 14539 12747 14611 12781
rect 14645 12747 14724 12781
rect 14539 12713 14724 12747
rect 14539 12679 14611 12713
rect 14645 12679 14724 12713
rect 14539 12645 14724 12679
rect 14539 12611 14611 12645
rect 14645 12611 14724 12645
rect 14539 12577 14724 12611
rect 14539 12543 14611 12577
rect 14645 12543 14724 12577
rect 14539 12509 14724 12543
rect 14539 12475 14611 12509
rect 14645 12475 14724 12509
rect 14539 12441 14724 12475
rect 14539 12407 14611 12441
rect 14645 12407 14724 12441
rect 14539 12373 14724 12407
rect 14539 12339 14611 12373
rect 14645 12339 14724 12373
rect 14539 12305 14724 12339
rect 14539 12271 14611 12305
rect 14645 12271 14724 12305
rect 14539 12237 14724 12271
rect 14539 12203 14611 12237
rect 14645 12203 14724 12237
rect 14539 12169 14724 12203
rect 14539 12135 14611 12169
rect 14645 12135 14724 12169
rect 14539 12101 14724 12135
rect 14539 12067 14611 12101
rect 14645 12067 14724 12101
rect 14539 12033 14724 12067
rect 14539 11999 14611 12033
rect 14645 11999 14724 12033
rect 14539 11965 14724 11999
rect 14539 11931 14611 11965
rect 14645 11931 14724 11965
rect 14539 11897 14724 11931
rect 14539 11863 14611 11897
rect 14645 11863 14724 11897
rect 14539 11829 14724 11863
rect 14539 11795 14611 11829
rect 14645 11795 14724 11829
rect 14539 11761 14724 11795
rect 14539 11727 14611 11761
rect 14645 11727 14724 11761
rect 14539 11693 14724 11727
rect 14539 11659 14611 11693
rect 14645 11659 14724 11693
rect 14539 11625 14724 11659
rect 14539 11591 14611 11625
rect 14645 11591 14724 11625
rect 14539 11557 14724 11591
rect 14539 11523 14611 11557
rect 14645 11523 14724 11557
rect 14539 11489 14724 11523
rect 14539 11455 14611 11489
rect 14645 11455 14724 11489
rect 14539 11421 14724 11455
rect 14539 11387 14611 11421
rect 14645 11387 14724 11421
rect 14539 11353 14724 11387
rect 14539 11319 14611 11353
rect 14645 11319 14724 11353
rect 14539 11285 14724 11319
rect 14539 11251 14611 11285
rect 14645 11251 14724 11285
rect 14539 11217 14724 11251
rect 14539 11183 14611 11217
rect 14645 11183 14724 11217
rect 14539 11149 14724 11183
rect 14539 11115 14611 11149
rect 14645 11115 14724 11149
rect 14539 11081 14724 11115
rect 14539 11047 14611 11081
rect 14645 11047 14724 11081
rect 14539 11013 14724 11047
rect 14539 10979 14611 11013
rect 14645 10979 14724 11013
rect 14539 10945 14724 10979
rect 14539 10911 14611 10945
rect 14645 10911 14724 10945
rect 14539 10877 14724 10911
rect 14539 10843 14611 10877
rect 14645 10843 14724 10877
rect 14539 10809 14724 10843
rect 14539 10775 14611 10809
rect 14645 10775 14724 10809
rect 14539 10741 14724 10775
rect 14539 10707 14611 10741
rect 14645 10707 14724 10741
rect 14539 10673 14724 10707
rect 14539 10639 14611 10673
rect 14645 10639 14724 10673
rect 14539 10605 14724 10639
rect 14539 10571 14611 10605
rect 14645 10571 14724 10605
rect 14539 10537 14724 10571
rect 14539 10503 14611 10537
rect 14645 10503 14724 10537
rect 14539 10469 14724 10503
rect 14539 10435 14611 10469
rect 14645 10435 14724 10469
rect 14539 10401 14724 10435
rect 14539 10367 14611 10401
rect 14645 10367 14724 10401
rect 14539 10333 14724 10367
rect 14539 10299 14611 10333
rect 14645 10299 14724 10333
rect 14539 10265 14724 10299
rect 14539 10231 14611 10265
rect 14645 10231 14724 10265
rect 14539 10197 14724 10231
rect 14539 10163 14611 10197
rect 14645 10163 14724 10197
rect 14539 10129 14724 10163
rect 14539 10095 14611 10129
rect 14645 10095 14724 10129
rect 14539 10061 14724 10095
rect 14539 10027 14611 10061
rect 14645 10027 14724 10061
rect 14539 9993 14724 10027
rect 14539 9959 14611 9993
rect 14645 9959 14724 9993
rect 14539 9925 14724 9959
rect 14539 9891 14611 9925
rect 14645 9891 14724 9925
rect 14539 9857 14724 9891
rect 14539 9823 14611 9857
rect 14645 9823 14724 9857
rect 14539 9789 14724 9823
rect 14539 9755 14611 9789
rect 14645 9755 14724 9789
rect 14539 9721 14724 9755
rect 245 9655 430 9689
rect 245 9621 317 9655
rect 351 9621 430 9655
rect 245 9528 430 9621
rect 14539 9687 14611 9721
rect 14645 9687 14724 9721
rect 14539 9653 14724 9687
rect 14539 9619 14611 9653
rect 14645 9619 14724 9653
rect 14539 9528 14724 9619
rect 245 9450 14724 9528
rect 245 9416 506 9450
rect 540 9416 574 9450
rect 608 9416 642 9450
rect 676 9416 710 9450
rect 744 9416 778 9450
rect 812 9416 846 9450
rect 880 9416 914 9450
rect 948 9416 982 9450
rect 1016 9416 1050 9450
rect 1084 9416 1118 9450
rect 1152 9416 1186 9450
rect 1220 9416 1254 9450
rect 1288 9416 1322 9450
rect 1356 9416 1390 9450
rect 1424 9416 1458 9450
rect 1492 9416 1526 9450
rect 1560 9416 1594 9450
rect 1628 9416 1662 9450
rect 1696 9416 1730 9450
rect 1764 9416 1798 9450
rect 1832 9416 1866 9450
rect 1900 9416 1934 9450
rect 1968 9416 2002 9450
rect 2036 9416 2070 9450
rect 2104 9416 2138 9450
rect 2172 9416 2206 9450
rect 2240 9416 2274 9450
rect 2308 9416 2342 9450
rect 2376 9416 2410 9450
rect 2444 9416 2478 9450
rect 2512 9416 2546 9450
rect 2580 9416 2614 9450
rect 2648 9416 2682 9450
rect 2716 9416 2750 9450
rect 2784 9416 2818 9450
rect 2852 9416 2886 9450
rect 2920 9416 2954 9450
rect 2988 9416 3022 9450
rect 3056 9416 3090 9450
rect 3124 9416 3158 9450
rect 3192 9416 3226 9450
rect 3260 9416 3294 9450
rect 3328 9416 3362 9450
rect 3396 9416 3430 9450
rect 3464 9416 3498 9450
rect 3532 9416 3566 9450
rect 3600 9416 3634 9450
rect 3668 9416 3702 9450
rect 3736 9416 3770 9450
rect 3804 9416 3838 9450
rect 3872 9416 3906 9450
rect 3940 9416 3974 9450
rect 4008 9416 4042 9450
rect 4076 9416 4110 9450
rect 4144 9416 4178 9450
rect 4212 9416 4246 9450
rect 4280 9416 4314 9450
rect 4348 9416 4382 9450
rect 4416 9416 4450 9450
rect 4484 9416 4518 9450
rect 4552 9416 4586 9450
rect 4620 9416 4654 9450
rect 4688 9416 4722 9450
rect 4756 9416 4790 9450
rect 4824 9416 4858 9450
rect 4892 9416 4926 9450
rect 4960 9416 4994 9450
rect 5028 9416 5062 9450
rect 5096 9416 5130 9450
rect 5164 9416 5198 9450
rect 5232 9416 5266 9450
rect 5300 9416 5334 9450
rect 5368 9416 5402 9450
rect 5436 9416 5470 9450
rect 5504 9416 5538 9450
rect 5572 9416 5606 9450
rect 5640 9416 5674 9450
rect 5708 9416 5742 9450
rect 5776 9416 5810 9450
rect 5844 9416 5878 9450
rect 5912 9416 5946 9450
rect 5980 9416 6014 9450
rect 6048 9416 6082 9450
rect 6116 9416 6150 9450
rect 6184 9416 6218 9450
rect 6252 9416 6286 9450
rect 6320 9416 6354 9450
rect 6388 9416 6422 9450
rect 6456 9416 6490 9450
rect 6524 9416 6558 9450
rect 6592 9416 6626 9450
rect 6660 9416 6694 9450
rect 6728 9416 6762 9450
rect 6796 9416 6830 9450
rect 6864 9416 6898 9450
rect 6932 9416 6966 9450
rect 7000 9416 7034 9450
rect 7068 9416 7102 9450
rect 7136 9416 7170 9450
rect 7204 9416 7238 9450
rect 7272 9416 7306 9450
rect 7340 9416 7374 9450
rect 7408 9416 7442 9450
rect 7476 9416 7510 9450
rect 7544 9416 7578 9450
rect 7612 9416 7646 9450
rect 7680 9416 7714 9450
rect 7748 9416 7782 9450
rect 7816 9416 7850 9450
rect 7884 9416 7918 9450
rect 7952 9416 7986 9450
rect 8020 9416 8054 9450
rect 8088 9416 8122 9450
rect 8156 9416 8190 9450
rect 8224 9416 8258 9450
rect 8292 9416 8326 9450
rect 8360 9416 8394 9450
rect 8428 9416 8462 9450
rect 8496 9416 8530 9450
rect 8564 9416 8598 9450
rect 8632 9416 8666 9450
rect 8700 9416 8734 9450
rect 8768 9416 8802 9450
rect 8836 9416 8870 9450
rect 8904 9416 8938 9450
rect 8972 9416 9006 9450
rect 9040 9416 9074 9450
rect 9108 9416 9142 9450
rect 9176 9416 9210 9450
rect 9244 9416 9278 9450
rect 9312 9416 9346 9450
rect 9380 9416 9414 9450
rect 9448 9416 9482 9450
rect 9516 9416 9550 9450
rect 9584 9416 9618 9450
rect 9652 9416 9686 9450
rect 9720 9416 9754 9450
rect 9788 9416 9822 9450
rect 9856 9416 9890 9450
rect 9924 9416 9958 9450
rect 9992 9416 10026 9450
rect 10060 9416 10094 9450
rect 10128 9416 10162 9450
rect 10196 9416 10230 9450
rect 10264 9416 10298 9450
rect 10332 9416 10366 9450
rect 10400 9416 10434 9450
rect 10468 9416 10502 9450
rect 10536 9416 10570 9450
rect 10604 9416 10638 9450
rect 10672 9416 10706 9450
rect 10740 9416 10774 9450
rect 10808 9416 10842 9450
rect 10876 9416 10910 9450
rect 10944 9416 10978 9450
rect 11012 9416 11046 9450
rect 11080 9416 11114 9450
rect 11148 9416 11182 9450
rect 11216 9416 11250 9450
rect 11284 9416 11318 9450
rect 11352 9416 11386 9450
rect 11420 9416 11454 9450
rect 11488 9416 11522 9450
rect 11556 9416 11590 9450
rect 11624 9416 11658 9450
rect 11692 9416 11726 9450
rect 11760 9416 11794 9450
rect 11828 9416 11862 9450
rect 11896 9416 11930 9450
rect 11964 9416 11998 9450
rect 12032 9416 12066 9450
rect 12100 9416 12134 9450
rect 12168 9416 12202 9450
rect 12236 9416 12270 9450
rect 12304 9416 12338 9450
rect 12372 9416 12406 9450
rect 12440 9416 12474 9450
rect 12508 9416 12542 9450
rect 12576 9416 12610 9450
rect 12644 9416 12678 9450
rect 12712 9416 12746 9450
rect 12780 9416 12814 9450
rect 12848 9416 12882 9450
rect 12916 9416 12950 9450
rect 12984 9416 13018 9450
rect 13052 9416 13086 9450
rect 13120 9416 13154 9450
rect 13188 9416 13222 9450
rect 13256 9416 13290 9450
rect 13324 9416 13358 9450
rect 13392 9416 13426 9450
rect 13460 9416 13494 9450
rect 13528 9416 13562 9450
rect 13596 9416 13630 9450
rect 13664 9416 13698 9450
rect 13732 9416 13766 9450
rect 13800 9416 13834 9450
rect 13868 9416 13902 9450
rect 13936 9416 13970 9450
rect 14004 9416 14038 9450
rect 14072 9416 14106 9450
rect 14140 9416 14174 9450
rect 14208 9416 14242 9450
rect 14276 9416 14310 9450
rect 14344 9416 14378 9450
rect 14412 9416 14446 9450
rect 14480 9416 14724 9450
rect 245 9343 14724 9416
<< mvnsubdiff >>
rect 583 36177 14381 36227
rect 583 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14381 36177
rect 583 36093 14381 36143
rect 583 36032 715 36093
rect 583 35998 632 36032
rect 666 35998 715 36032
rect 583 35964 715 35998
rect 583 35930 632 35964
rect 666 35930 715 35964
rect 583 35896 715 35930
rect 583 35862 632 35896
rect 666 35862 715 35896
rect 583 35828 715 35862
rect 583 35794 632 35828
rect 666 35794 715 35828
rect 583 35760 715 35794
rect 583 35726 632 35760
rect 666 35726 715 35760
rect 583 35692 715 35726
rect 583 35658 632 35692
rect 666 35658 715 35692
rect 583 35624 715 35658
rect 583 35590 632 35624
rect 666 35590 715 35624
rect 583 35556 715 35590
rect 583 35522 632 35556
rect 666 35522 715 35556
rect 583 35488 715 35522
rect 583 35454 632 35488
rect 666 35454 715 35488
rect 583 35420 715 35454
rect 583 35386 632 35420
rect 666 35386 715 35420
rect 583 35352 715 35386
rect 583 35318 632 35352
rect 666 35318 715 35352
rect 583 35284 715 35318
rect 583 35250 632 35284
rect 666 35250 715 35284
rect 583 35216 715 35250
rect 583 35182 632 35216
rect 666 35182 715 35216
rect 583 35148 715 35182
rect 583 35114 632 35148
rect 666 35114 715 35148
rect 583 35080 715 35114
rect 583 35046 632 35080
rect 666 35046 715 35080
rect 583 35012 715 35046
rect 583 34978 632 35012
rect 666 34978 715 35012
rect 583 34944 715 34978
rect 583 34910 632 34944
rect 666 34910 715 34944
rect 583 34876 715 34910
rect 583 34842 632 34876
rect 666 34842 715 34876
rect 583 34808 715 34842
rect 583 34774 632 34808
rect 666 34774 715 34808
rect 583 34740 715 34774
rect 583 34706 632 34740
rect 666 34706 715 34740
rect 583 34672 715 34706
rect 14247 36032 14381 36093
rect 14247 35998 14297 36032
rect 14331 35998 14381 36032
rect 14247 35964 14381 35998
rect 14247 35930 14297 35964
rect 14331 35930 14381 35964
rect 14247 35896 14381 35930
rect 14247 35862 14297 35896
rect 14331 35862 14381 35896
rect 14247 35828 14381 35862
rect 14247 35794 14297 35828
rect 14331 35794 14381 35828
rect 14247 35760 14381 35794
rect 14247 35726 14297 35760
rect 14331 35726 14381 35760
rect 14247 35692 14381 35726
rect 14247 35658 14297 35692
rect 14331 35658 14381 35692
rect 14247 35624 14381 35658
rect 14247 35590 14297 35624
rect 14331 35590 14381 35624
rect 14247 35556 14381 35590
rect 14247 35522 14297 35556
rect 14331 35522 14381 35556
rect 14247 35488 14381 35522
rect 14247 35454 14297 35488
rect 14331 35454 14381 35488
rect 14247 35420 14381 35454
rect 14247 35386 14297 35420
rect 14331 35386 14381 35420
rect 14247 35352 14381 35386
rect 14247 35318 14297 35352
rect 14331 35318 14381 35352
rect 14247 35284 14381 35318
rect 14247 35250 14297 35284
rect 14331 35250 14381 35284
rect 14247 35216 14381 35250
rect 14247 35182 14297 35216
rect 14331 35182 14381 35216
rect 14247 35148 14381 35182
rect 14247 35114 14297 35148
rect 14331 35114 14381 35148
rect 14247 35080 14381 35114
rect 14247 35046 14297 35080
rect 14331 35046 14381 35080
rect 14247 35012 14381 35046
rect 14247 34978 14297 35012
rect 14331 34978 14381 35012
rect 14247 34944 14381 34978
rect 14247 34910 14297 34944
rect 14331 34910 14381 34944
rect 14247 34876 14381 34910
rect 14247 34842 14297 34876
rect 14331 34842 14381 34876
rect 14247 34808 14381 34842
rect 14247 34774 14297 34808
rect 14331 34774 14381 34808
rect 14247 34740 14381 34774
rect 14247 34706 14297 34740
rect 14331 34706 14381 34740
rect 583 34638 632 34672
rect 666 34638 715 34672
rect 583 34604 715 34638
rect 583 34570 632 34604
rect 666 34570 715 34604
rect 583 34536 715 34570
rect 583 34502 632 34536
rect 666 34502 715 34536
rect 583 34468 715 34502
rect 583 34434 632 34468
rect 666 34434 715 34468
rect 583 34400 715 34434
rect 583 34366 632 34400
rect 666 34366 715 34400
rect 583 34332 715 34366
rect 583 34298 632 34332
rect 666 34298 715 34332
rect 583 34264 715 34298
rect 583 34230 632 34264
rect 666 34230 715 34264
rect 583 34196 715 34230
rect 583 34162 632 34196
rect 666 34162 715 34196
rect 583 34128 715 34162
rect 583 34094 632 34128
rect 666 34094 715 34128
rect 583 34060 715 34094
rect 583 34026 632 34060
rect 666 34026 715 34060
rect 583 33992 715 34026
rect 583 33958 632 33992
rect 666 33958 715 33992
rect 583 33924 715 33958
rect 583 33890 632 33924
rect 666 33890 715 33924
rect 583 33856 715 33890
rect 583 33822 632 33856
rect 666 33822 715 33856
rect 583 33788 715 33822
rect 583 33754 632 33788
rect 666 33754 715 33788
rect 583 33720 715 33754
rect 583 33686 632 33720
rect 666 33686 715 33720
rect 583 33652 715 33686
rect 583 33618 632 33652
rect 666 33618 715 33652
rect 583 33584 715 33618
rect 583 33550 632 33584
rect 666 33550 715 33584
rect 583 33516 715 33550
rect 583 33482 632 33516
rect 666 33482 715 33516
rect 583 33448 715 33482
rect 583 33414 632 33448
rect 666 33414 715 33448
rect 583 33380 715 33414
rect 583 33346 632 33380
rect 666 33346 715 33380
rect 583 33312 715 33346
rect 583 33278 632 33312
rect 666 33278 715 33312
rect 583 33244 715 33278
rect 583 33210 632 33244
rect 666 33210 715 33244
rect 583 33176 715 33210
rect 583 33142 632 33176
rect 666 33142 715 33176
rect 583 33108 715 33142
rect 583 33074 632 33108
rect 666 33074 715 33108
rect 583 33040 715 33074
rect 583 33006 632 33040
rect 666 33006 715 33040
rect 583 32972 715 33006
rect 583 32938 632 32972
rect 666 32938 715 32972
rect 583 32904 715 32938
rect 583 32870 632 32904
rect 666 32870 715 32904
rect 583 32836 715 32870
rect 583 32802 632 32836
rect 666 32802 715 32836
rect 583 32768 715 32802
rect 583 32734 632 32768
rect 666 32734 715 32768
rect 583 32700 715 32734
rect 583 32666 632 32700
rect 666 32666 715 32700
rect 583 32632 715 32666
rect 583 32598 632 32632
rect 666 32598 715 32632
rect 583 32564 715 32598
rect 583 32530 632 32564
rect 666 32530 715 32564
rect 583 32496 715 32530
rect 583 32462 632 32496
rect 666 32462 715 32496
rect 583 32428 715 32462
rect 583 32394 632 32428
rect 666 32394 715 32428
rect 583 32360 715 32394
rect 583 32326 632 32360
rect 666 32326 715 32360
rect 583 32292 715 32326
rect 583 32258 632 32292
rect 666 32258 715 32292
rect 583 32224 715 32258
rect 583 32190 632 32224
rect 666 32190 715 32224
rect 583 32156 715 32190
rect 583 32122 632 32156
rect 666 32122 715 32156
rect 583 32088 715 32122
rect 583 32054 632 32088
rect 666 32054 715 32088
rect 583 32020 715 32054
rect 583 31986 632 32020
rect 666 31986 715 32020
rect 583 31952 715 31986
rect 583 31918 632 31952
rect 666 31918 715 31952
rect 583 31884 715 31918
rect 583 31850 632 31884
rect 666 31850 715 31884
rect 583 31816 715 31850
rect 583 31782 632 31816
rect 666 31782 715 31816
rect 583 31748 715 31782
rect 583 31714 632 31748
rect 666 31714 715 31748
rect 583 31680 715 31714
rect 583 31646 632 31680
rect 666 31646 715 31680
rect 583 31612 715 31646
rect 583 31578 632 31612
rect 666 31578 715 31612
rect 583 31544 715 31578
rect 583 31510 632 31544
rect 666 31510 715 31544
rect 583 31476 715 31510
rect 583 31442 632 31476
rect 666 31442 715 31476
rect 583 31408 715 31442
rect 583 31374 632 31408
rect 666 31374 715 31408
rect 583 31340 715 31374
rect 583 31306 632 31340
rect 666 31306 715 31340
rect 583 31272 715 31306
rect 583 31238 632 31272
rect 666 31238 715 31272
rect 583 31204 715 31238
rect 583 31170 632 31204
rect 666 31170 715 31204
rect 583 31136 715 31170
rect 583 31102 632 31136
rect 666 31102 715 31136
rect 583 31068 715 31102
rect 583 31034 632 31068
rect 666 31034 715 31068
rect 583 31000 715 31034
rect 583 30966 632 31000
rect 666 30966 715 31000
rect 583 30932 715 30966
rect 583 30898 632 30932
rect 666 30898 715 30932
rect 583 30864 715 30898
rect 583 30830 632 30864
rect 666 30830 715 30864
rect 583 30796 715 30830
rect 583 30762 632 30796
rect 666 30762 715 30796
rect 583 30728 715 30762
rect 583 30694 632 30728
rect 666 30694 715 30728
rect 583 30660 715 30694
rect 583 30626 632 30660
rect 666 30626 715 30660
rect 583 30592 715 30626
rect 583 30558 632 30592
rect 666 30558 715 30592
rect 583 30524 715 30558
rect 583 30490 632 30524
rect 666 30490 715 30524
rect 583 30456 715 30490
rect 583 30422 632 30456
rect 666 30422 715 30456
rect 583 30388 715 30422
rect 583 30354 632 30388
rect 666 30354 715 30388
rect 583 30320 715 30354
rect 583 30286 632 30320
rect 666 30286 715 30320
rect 583 30252 715 30286
rect 583 30218 632 30252
rect 666 30218 715 30252
rect 583 30184 715 30218
rect 583 30150 632 30184
rect 666 30150 715 30184
rect 583 30116 715 30150
rect 583 30082 632 30116
rect 666 30082 715 30116
rect 583 30048 715 30082
rect 583 30014 632 30048
rect 666 30014 715 30048
rect 583 29980 715 30014
rect 583 29946 632 29980
rect 666 29946 715 29980
rect 583 29912 715 29946
rect 583 29878 632 29912
rect 666 29878 715 29912
rect 583 29844 715 29878
rect 583 29810 632 29844
rect 666 29810 715 29844
rect 583 29776 715 29810
rect 583 29742 632 29776
rect 666 29742 715 29776
rect 583 29708 715 29742
rect 583 29674 632 29708
rect 666 29674 715 29708
rect 583 29640 715 29674
rect 583 29606 632 29640
rect 666 29606 715 29640
rect 583 29572 715 29606
rect 583 29538 632 29572
rect 666 29538 715 29572
rect 583 29504 715 29538
rect 583 29470 632 29504
rect 666 29470 715 29504
rect 583 29436 715 29470
rect 583 29402 632 29436
rect 666 29402 715 29436
rect 583 29368 715 29402
rect 583 29334 632 29368
rect 666 29334 715 29368
rect 583 29300 715 29334
rect 583 29266 632 29300
rect 666 29266 715 29300
rect 583 29232 715 29266
rect 583 29198 632 29232
rect 666 29198 715 29232
rect 583 29164 715 29198
rect 583 29130 632 29164
rect 666 29130 715 29164
rect 583 29096 715 29130
rect 583 29062 632 29096
rect 666 29062 715 29096
rect 583 29028 715 29062
rect 583 28994 632 29028
rect 666 28994 715 29028
rect 583 28960 715 28994
rect 583 28926 632 28960
rect 666 28926 715 28960
rect 583 28892 715 28926
rect 583 28858 632 28892
rect 666 28858 715 28892
rect 583 28824 715 28858
rect 583 28790 632 28824
rect 666 28790 715 28824
rect 583 28756 715 28790
rect 583 28722 632 28756
rect 666 28722 715 28756
rect 583 28688 715 28722
rect 583 28654 632 28688
rect 666 28654 715 28688
rect 583 28620 715 28654
rect 583 28586 632 28620
rect 666 28586 715 28620
rect 583 28552 715 28586
rect 583 28518 632 28552
rect 666 28518 715 28552
rect 583 28484 715 28518
rect 583 28450 632 28484
rect 666 28450 715 28484
rect 583 28416 715 28450
rect 583 28382 632 28416
rect 666 28382 715 28416
rect 583 28348 715 28382
rect 583 28314 632 28348
rect 666 28314 715 28348
rect 583 28280 715 28314
rect 583 28246 632 28280
rect 666 28246 715 28280
rect 583 28212 715 28246
rect 583 28178 632 28212
rect 666 28178 715 28212
rect 583 28144 715 28178
rect 583 28110 632 28144
rect 666 28110 715 28144
rect 583 28076 715 28110
rect 583 28042 632 28076
rect 666 28042 715 28076
rect 583 28008 715 28042
rect 583 27974 632 28008
rect 666 27974 715 28008
rect 583 27940 715 27974
rect 583 27906 632 27940
rect 666 27906 715 27940
rect 583 27872 715 27906
rect 583 27838 632 27872
rect 666 27838 715 27872
rect 583 27804 715 27838
rect 583 27770 632 27804
rect 666 27770 715 27804
rect 583 27736 715 27770
rect 583 27702 632 27736
rect 666 27702 715 27736
rect 583 27668 715 27702
rect 583 27634 632 27668
rect 666 27634 715 27668
rect 583 27600 715 27634
rect 583 27566 632 27600
rect 666 27566 715 27600
rect 583 27532 715 27566
rect 583 27498 632 27532
rect 666 27498 715 27532
rect 583 27464 715 27498
rect 583 27430 632 27464
rect 666 27430 715 27464
rect 583 27396 715 27430
rect 583 27362 632 27396
rect 666 27362 715 27396
rect 583 27328 715 27362
rect 583 27294 632 27328
rect 666 27294 715 27328
rect 583 27260 715 27294
rect 583 27226 632 27260
rect 666 27226 715 27260
rect 583 27192 715 27226
rect 583 27158 632 27192
rect 666 27158 715 27192
rect 583 27124 715 27158
rect 583 27090 632 27124
rect 666 27090 715 27124
rect 583 27056 715 27090
rect 583 27022 632 27056
rect 666 27022 715 27056
rect 583 26988 715 27022
rect 583 26954 632 26988
rect 666 26954 715 26988
rect 583 26920 715 26954
rect 583 26886 632 26920
rect 666 26886 715 26920
rect 583 26852 715 26886
rect 583 26818 632 26852
rect 666 26818 715 26852
rect 583 26784 715 26818
rect 583 26750 632 26784
rect 666 26750 715 26784
rect 583 26716 715 26750
rect 583 26682 632 26716
rect 666 26682 715 26716
rect 583 26648 715 26682
rect 583 26614 632 26648
rect 666 26614 715 26648
rect 583 26580 715 26614
rect 583 26546 632 26580
rect 666 26546 715 26580
rect 583 26512 715 26546
rect 583 26478 632 26512
rect 666 26478 715 26512
rect 583 26444 715 26478
rect 583 26410 632 26444
rect 666 26410 715 26444
rect 583 26376 715 26410
rect 583 26342 632 26376
rect 666 26342 715 26376
rect 583 26308 715 26342
rect 583 26274 632 26308
rect 666 26274 715 26308
rect 583 26240 715 26274
rect 583 26206 632 26240
rect 666 26206 715 26240
rect 583 26172 715 26206
rect 583 26138 632 26172
rect 666 26138 715 26172
rect 583 26104 715 26138
rect 583 26070 632 26104
rect 666 26070 715 26104
rect 583 26036 715 26070
rect 583 26002 632 26036
rect 666 26002 715 26036
rect 583 25968 715 26002
rect 583 25934 632 25968
rect 666 25934 715 25968
rect 583 25900 715 25934
rect 583 25866 632 25900
rect 666 25866 715 25900
rect 583 25832 715 25866
rect 583 25798 632 25832
rect 666 25798 715 25832
rect 583 25764 715 25798
rect 583 25730 632 25764
rect 666 25730 715 25764
rect 583 25696 715 25730
rect 583 25662 632 25696
rect 666 25662 715 25696
rect 583 25628 715 25662
rect 583 25594 632 25628
rect 666 25594 715 25628
rect 583 25560 715 25594
rect 583 25526 632 25560
rect 666 25526 715 25560
rect 583 25492 715 25526
rect 583 25458 632 25492
rect 666 25458 715 25492
rect 583 25424 715 25458
rect 583 25390 632 25424
rect 666 25390 715 25424
rect 583 25356 715 25390
rect 583 25322 632 25356
rect 666 25322 715 25356
rect 583 25288 715 25322
rect 583 25254 632 25288
rect 666 25254 715 25288
rect 583 25220 715 25254
rect 583 25186 632 25220
rect 666 25186 715 25220
rect 583 25152 715 25186
rect 583 25118 632 25152
rect 666 25118 715 25152
rect 583 25084 715 25118
rect 583 25050 632 25084
rect 666 25050 715 25084
rect 583 25016 715 25050
rect 583 24982 632 25016
rect 666 24982 715 25016
rect 583 24948 715 24982
rect 583 24914 632 24948
rect 666 24914 715 24948
rect 583 24880 715 24914
rect 583 24846 632 24880
rect 666 24846 715 24880
rect 583 24812 715 24846
rect 583 24778 632 24812
rect 666 24778 715 24812
rect 583 24744 715 24778
rect 583 24710 632 24744
rect 666 24710 715 24744
rect 583 24676 715 24710
rect 583 24642 632 24676
rect 666 24642 715 24676
rect 583 24608 715 24642
rect 583 24574 632 24608
rect 666 24574 715 24608
rect 583 24540 715 24574
rect 583 24506 632 24540
rect 666 24506 715 24540
rect 583 24472 715 24506
rect 583 24438 632 24472
rect 666 24438 715 24472
rect 583 24404 715 24438
rect 583 24370 632 24404
rect 666 24370 715 24404
rect 583 24336 715 24370
rect 583 24302 632 24336
rect 666 24302 715 24336
rect 583 24268 715 24302
rect 583 24234 632 24268
rect 666 24234 715 24268
rect 583 24200 715 24234
rect 583 24166 632 24200
rect 666 24166 715 24200
rect 583 24132 715 24166
rect 583 24098 632 24132
rect 666 24098 715 24132
rect 583 24064 715 24098
rect 583 24030 632 24064
rect 666 24030 715 24064
rect 583 23996 715 24030
rect 583 23962 632 23996
rect 666 23962 715 23996
rect 583 23928 715 23962
rect 583 23894 632 23928
rect 666 23894 715 23928
rect 583 23860 715 23894
rect 583 23826 632 23860
rect 666 23826 715 23860
rect 583 23792 715 23826
rect 583 23758 632 23792
rect 666 23758 715 23792
rect 583 23724 715 23758
rect 583 23690 632 23724
rect 666 23690 715 23724
rect 583 23656 715 23690
rect 583 23622 632 23656
rect 666 23622 715 23656
rect 583 23588 715 23622
rect 583 23554 632 23588
rect 666 23554 715 23588
rect 583 23520 715 23554
rect 583 23486 632 23520
rect 666 23486 715 23520
rect 583 23452 715 23486
rect 583 23418 632 23452
rect 666 23418 715 23452
rect 583 23384 715 23418
rect 583 23350 632 23384
rect 666 23350 715 23384
rect 583 23316 715 23350
rect 583 23282 632 23316
rect 666 23282 715 23316
rect 583 23248 715 23282
rect 583 23214 632 23248
rect 666 23214 715 23248
rect 583 23180 715 23214
rect 583 23146 632 23180
rect 666 23146 715 23180
rect 583 23112 715 23146
rect 583 23078 632 23112
rect 666 23078 715 23112
rect 583 23044 715 23078
rect 583 23010 632 23044
rect 666 23010 715 23044
rect 583 22976 715 23010
rect 583 22942 632 22976
rect 666 22942 715 22976
rect 583 22908 715 22942
rect 583 22874 632 22908
rect 666 22874 715 22908
rect 583 22840 715 22874
rect 583 22806 632 22840
rect 666 22806 715 22840
rect 583 22772 715 22806
rect 583 22738 632 22772
rect 666 22738 715 22772
rect 583 22704 715 22738
rect 583 22670 632 22704
rect 666 22670 715 22704
rect 583 22636 715 22670
rect 583 22602 632 22636
rect 666 22602 715 22636
rect 583 22568 715 22602
rect 583 22534 632 22568
rect 666 22534 715 22568
rect 583 22500 715 22534
rect 583 22466 632 22500
rect 666 22466 715 22500
rect 583 22432 715 22466
rect 583 22398 632 22432
rect 666 22398 715 22432
rect 583 22364 715 22398
rect 583 22330 632 22364
rect 666 22330 715 22364
rect 583 22296 715 22330
rect 583 22262 632 22296
rect 666 22262 715 22296
rect 583 22228 715 22262
rect 583 22194 632 22228
rect 666 22194 715 22228
rect 583 22160 715 22194
rect 583 22126 632 22160
rect 666 22126 715 22160
rect 583 22092 715 22126
rect 583 22058 632 22092
rect 666 22058 715 22092
rect 583 22024 715 22058
rect 583 21990 632 22024
rect 666 21990 715 22024
rect 583 21956 715 21990
rect 583 21922 632 21956
rect 666 21922 715 21956
rect 583 21888 715 21922
rect 583 21854 632 21888
rect 666 21854 715 21888
rect 583 21820 715 21854
rect 583 21786 632 21820
rect 666 21786 715 21820
rect 583 21752 715 21786
rect 583 21718 632 21752
rect 666 21718 715 21752
rect 583 21684 715 21718
rect 583 21650 632 21684
rect 666 21650 715 21684
rect 583 21616 715 21650
rect 583 21582 632 21616
rect 666 21582 715 21616
rect 583 21548 715 21582
rect 583 21514 632 21548
rect 666 21514 715 21548
rect 583 21480 715 21514
rect 583 21446 632 21480
rect 666 21446 715 21480
rect 583 21412 715 21446
rect 583 21378 632 21412
rect 666 21378 715 21412
rect 583 21344 715 21378
rect 583 21310 632 21344
rect 666 21310 715 21344
rect 583 21276 715 21310
rect 583 21242 632 21276
rect 666 21242 715 21276
rect 583 21208 715 21242
rect 583 21174 632 21208
rect 666 21174 715 21208
rect 583 21140 715 21174
rect 583 21106 632 21140
rect 666 21106 715 21140
rect 583 21072 715 21106
rect 583 21038 632 21072
rect 666 21038 715 21072
rect 583 21004 715 21038
rect 583 20970 632 21004
rect 666 20970 715 21004
rect 583 20936 715 20970
rect 583 20902 632 20936
rect 666 20902 715 20936
rect 583 20868 715 20902
rect 583 20834 632 20868
rect 666 20834 715 20868
rect 583 20800 715 20834
rect 583 20766 632 20800
rect 666 20766 715 20800
rect 583 20732 715 20766
rect 583 20698 632 20732
rect 666 20698 715 20732
rect 583 20664 715 20698
rect 583 20630 632 20664
rect 666 20630 715 20664
rect 583 20596 715 20630
rect 583 20562 632 20596
rect 666 20562 715 20596
rect 583 20528 715 20562
rect 583 20494 632 20528
rect 666 20494 715 20528
rect 583 20460 715 20494
rect 583 20426 632 20460
rect 666 20426 715 20460
rect 583 20392 715 20426
rect 583 20358 632 20392
rect 666 20358 715 20392
rect 583 20324 715 20358
rect 583 20290 632 20324
rect 666 20290 715 20324
rect 583 20256 715 20290
rect 583 20222 632 20256
rect 666 20222 715 20256
rect 583 20188 715 20222
rect 583 20154 632 20188
rect 666 20154 715 20188
rect 583 20120 715 20154
rect 583 20086 632 20120
rect 666 20086 715 20120
rect 583 20052 715 20086
rect 583 20018 632 20052
rect 666 20018 715 20052
rect 583 19984 715 20018
rect 583 19950 632 19984
rect 666 19950 715 19984
rect 583 19916 715 19950
rect 583 19882 632 19916
rect 666 19882 715 19916
rect 583 19848 715 19882
rect 583 19814 632 19848
rect 666 19814 715 19848
rect 583 19780 715 19814
rect 583 19746 632 19780
rect 666 19746 715 19780
rect 583 19712 715 19746
rect 583 19678 632 19712
rect 666 19678 715 19712
rect 583 19644 715 19678
rect 583 19610 632 19644
rect 666 19610 715 19644
rect 583 19576 715 19610
rect 583 19542 632 19576
rect 666 19542 715 19576
rect 583 19508 715 19542
rect 583 19474 632 19508
rect 666 19474 715 19508
rect 583 19440 715 19474
rect 583 19406 632 19440
rect 666 19406 715 19440
rect 583 19372 715 19406
rect 583 19338 632 19372
rect 666 19338 715 19372
rect 583 19304 715 19338
rect 583 19270 632 19304
rect 666 19270 715 19304
rect 583 19236 715 19270
rect 583 19202 632 19236
rect 666 19202 715 19236
rect 583 19168 715 19202
rect 583 19134 632 19168
rect 666 19134 715 19168
rect 583 19100 715 19134
rect 583 19066 632 19100
rect 666 19066 715 19100
rect 583 19032 715 19066
rect 583 18998 632 19032
rect 666 18998 715 19032
rect 583 18964 715 18998
rect 583 18930 632 18964
rect 666 18930 715 18964
rect 583 18896 715 18930
rect 583 18862 632 18896
rect 666 18862 715 18896
rect 583 18828 715 18862
rect 583 18794 632 18828
rect 666 18794 715 18828
rect 583 18760 715 18794
rect 583 18726 632 18760
rect 666 18726 715 18760
rect 583 18692 715 18726
rect 583 18658 632 18692
rect 666 18658 715 18692
rect 583 18624 715 18658
rect 583 18590 632 18624
rect 666 18590 715 18624
rect 583 18556 715 18590
rect 583 18522 632 18556
rect 666 18522 715 18556
rect 583 18488 715 18522
rect 583 18454 632 18488
rect 666 18454 715 18488
rect 583 18420 715 18454
rect 583 18386 632 18420
rect 666 18386 715 18420
rect 583 18352 715 18386
rect 583 18318 632 18352
rect 666 18318 715 18352
rect 583 18284 715 18318
rect 583 18250 632 18284
rect 666 18250 715 18284
rect 583 18216 715 18250
rect 583 18182 632 18216
rect 666 18182 715 18216
rect 583 18148 715 18182
rect 583 18114 632 18148
rect 666 18114 715 18148
rect 583 18080 715 18114
rect 583 18046 632 18080
rect 666 18046 715 18080
rect 583 18012 715 18046
rect 583 17978 632 18012
rect 666 17978 715 18012
rect 583 17944 715 17978
rect 583 17910 632 17944
rect 666 17910 715 17944
rect 583 17876 715 17910
rect 583 17842 632 17876
rect 666 17842 715 17876
rect 583 17808 715 17842
rect 583 17774 632 17808
rect 666 17774 715 17808
rect 583 17740 715 17774
rect 583 17706 632 17740
rect 666 17706 715 17740
rect 583 17672 715 17706
rect 583 17638 632 17672
rect 666 17638 715 17672
rect 583 17604 715 17638
rect 583 17570 632 17604
rect 666 17570 715 17604
rect 583 17536 715 17570
rect 583 17502 632 17536
rect 666 17502 715 17536
rect 583 17468 715 17502
rect 583 17434 632 17468
rect 666 17434 715 17468
rect 583 17400 715 17434
rect 583 17366 632 17400
rect 666 17366 715 17400
rect 583 17332 715 17366
rect 583 17298 632 17332
rect 666 17298 715 17332
rect 583 17264 715 17298
rect 583 17230 632 17264
rect 666 17230 715 17264
rect 583 17196 715 17230
rect 583 17162 632 17196
rect 666 17162 715 17196
rect 583 17128 715 17162
rect 583 17094 632 17128
rect 666 17094 715 17128
rect 583 17060 715 17094
rect 583 17026 632 17060
rect 666 17026 715 17060
rect 583 16992 715 17026
rect 583 16958 632 16992
rect 666 16958 715 16992
rect 583 16924 715 16958
rect 583 16890 632 16924
rect 666 16890 715 16924
rect 583 16856 715 16890
rect 583 16822 632 16856
rect 666 16822 715 16856
rect 583 16788 715 16822
rect 583 16754 632 16788
rect 666 16754 715 16788
rect 583 16720 715 16754
rect 583 16686 632 16720
rect 666 16686 715 16720
rect 583 16652 715 16686
rect 583 16618 632 16652
rect 666 16618 715 16652
rect 583 16584 715 16618
rect 583 16550 632 16584
rect 666 16550 715 16584
rect 583 16516 715 16550
rect 583 16482 632 16516
rect 666 16482 715 16516
rect 583 16448 715 16482
rect 583 16414 632 16448
rect 666 16414 715 16448
rect 583 16380 715 16414
rect 583 16346 632 16380
rect 666 16346 715 16380
rect 583 16312 715 16346
rect 583 16278 632 16312
rect 666 16278 715 16312
rect 583 16244 715 16278
rect 583 16210 632 16244
rect 666 16210 715 16244
rect 583 16176 715 16210
rect 583 16142 632 16176
rect 666 16142 715 16176
rect 583 16108 715 16142
rect 583 16074 632 16108
rect 666 16074 715 16108
rect 583 16040 715 16074
rect 583 16006 632 16040
rect 666 16006 715 16040
rect 583 15972 715 16006
rect 583 15938 632 15972
rect 666 15938 715 15972
rect 583 15904 715 15938
rect 583 15870 632 15904
rect 666 15870 715 15904
rect 583 15836 715 15870
rect 583 15802 632 15836
rect 666 15802 715 15836
rect 583 15768 715 15802
rect 583 15734 632 15768
rect 666 15734 715 15768
rect 583 15700 715 15734
rect 583 15666 632 15700
rect 666 15666 715 15700
rect 583 15632 715 15666
rect 583 15598 632 15632
rect 666 15598 715 15632
rect 583 15564 715 15598
rect 583 15530 632 15564
rect 666 15530 715 15564
rect 583 15496 715 15530
rect 583 15462 632 15496
rect 666 15462 715 15496
rect 583 15428 715 15462
rect 583 15394 632 15428
rect 666 15394 715 15428
rect 583 15360 715 15394
rect 583 15326 632 15360
rect 666 15326 715 15360
rect 583 15292 715 15326
rect 583 15258 632 15292
rect 666 15258 715 15292
rect 583 15224 715 15258
rect 583 15190 632 15224
rect 666 15190 715 15224
rect 583 15156 715 15190
rect 583 15122 632 15156
rect 666 15122 715 15156
rect 583 15088 715 15122
rect 583 15054 632 15088
rect 666 15054 715 15088
rect 583 15020 715 15054
rect 583 14986 632 15020
rect 666 14986 715 15020
rect 583 14952 715 14986
rect 583 14918 632 14952
rect 666 14918 715 14952
rect 583 14884 715 14918
rect 583 14850 632 14884
rect 666 14850 715 14884
rect 583 14816 715 14850
rect 583 14782 632 14816
rect 666 14782 715 14816
rect 583 14748 715 14782
rect 583 14714 632 14748
rect 666 14714 715 14748
rect 583 14680 715 14714
rect 583 14646 632 14680
rect 666 14646 715 14680
rect 583 14612 715 14646
rect 583 14578 632 14612
rect 666 14578 715 14612
rect 583 14544 715 14578
rect 583 14510 632 14544
rect 666 14510 715 14544
rect 583 14476 715 14510
rect 583 14442 632 14476
rect 666 14442 715 14476
rect 583 14408 715 14442
rect 583 14374 632 14408
rect 666 14374 715 14408
rect 583 14340 715 14374
rect 583 14306 632 14340
rect 666 14306 715 14340
rect 583 14272 715 14306
rect 583 14238 632 14272
rect 666 14238 715 14272
rect 583 14204 715 14238
rect 583 14170 632 14204
rect 666 14170 715 14204
rect 583 14136 715 14170
rect 583 14102 632 14136
rect 666 14102 715 14136
rect 583 14068 715 14102
rect 583 14034 632 14068
rect 666 14034 715 14068
rect 583 14000 715 14034
rect 583 13966 632 14000
rect 666 13966 715 14000
rect 583 13932 715 13966
rect 583 13898 632 13932
rect 666 13898 715 13932
rect 583 13864 715 13898
rect 583 13830 632 13864
rect 666 13830 715 13864
rect 583 13796 715 13830
rect 583 13762 632 13796
rect 666 13762 715 13796
rect 583 13728 715 13762
rect 583 13694 632 13728
rect 666 13694 715 13728
rect 583 13660 715 13694
rect 583 13626 632 13660
rect 666 13626 715 13660
rect 583 13592 715 13626
rect 583 13558 632 13592
rect 666 13558 715 13592
rect 583 13524 715 13558
rect 583 13490 632 13524
rect 666 13490 715 13524
rect 583 13456 715 13490
rect 583 13422 632 13456
rect 666 13422 715 13456
rect 583 13388 715 13422
rect 583 13354 632 13388
rect 666 13354 715 13388
rect 583 13320 715 13354
rect 583 13286 632 13320
rect 666 13286 715 13320
rect 583 13252 715 13286
rect 583 13218 632 13252
rect 666 13218 715 13252
rect 583 13184 715 13218
rect 583 13150 632 13184
rect 666 13150 715 13184
rect 583 13116 715 13150
rect 583 13082 632 13116
rect 666 13082 715 13116
rect 583 13048 715 13082
rect 583 13014 632 13048
rect 666 13014 715 13048
rect 583 12980 715 13014
rect 583 12946 632 12980
rect 666 12946 715 12980
rect 583 12912 715 12946
rect 583 12878 632 12912
rect 666 12878 715 12912
rect 583 12844 715 12878
rect 583 12810 632 12844
rect 666 12810 715 12844
rect 583 12776 715 12810
rect 583 12742 632 12776
rect 666 12742 715 12776
rect 583 12708 715 12742
rect 583 12674 632 12708
rect 666 12674 715 12708
rect 583 12640 715 12674
rect 583 12606 632 12640
rect 666 12606 715 12640
rect 583 12572 715 12606
rect 583 12538 632 12572
rect 666 12538 715 12572
rect 583 12504 715 12538
rect 583 12470 632 12504
rect 666 12470 715 12504
rect 583 12436 715 12470
rect 583 12402 632 12436
rect 666 12402 715 12436
rect 583 12368 715 12402
rect 583 12334 632 12368
rect 666 12334 715 12368
rect 583 12300 715 12334
rect 583 12266 632 12300
rect 666 12266 715 12300
rect 583 12232 715 12266
rect 583 12198 632 12232
rect 666 12198 715 12232
rect 583 12164 715 12198
rect 583 12130 632 12164
rect 666 12130 715 12164
rect 583 12096 715 12130
rect 583 12062 632 12096
rect 666 12062 715 12096
rect 583 12028 715 12062
rect 583 11994 632 12028
rect 666 11994 715 12028
rect 583 11960 715 11994
rect 583 11926 632 11960
rect 666 11926 715 11960
rect 583 11892 715 11926
rect 583 11858 632 11892
rect 666 11858 715 11892
rect 583 11824 715 11858
rect 583 11790 632 11824
rect 666 11790 715 11824
rect 583 11756 715 11790
rect 583 11722 632 11756
rect 666 11722 715 11756
rect 583 11688 715 11722
rect 583 11654 632 11688
rect 666 11654 715 11688
rect 583 11620 715 11654
rect 583 11586 632 11620
rect 666 11586 715 11620
rect 583 11552 715 11586
rect 583 11518 632 11552
rect 666 11518 715 11552
rect 583 11484 715 11518
rect 583 11450 632 11484
rect 666 11450 715 11484
rect 583 11416 715 11450
rect 583 11382 632 11416
rect 666 11382 715 11416
rect 583 11348 715 11382
rect 583 11314 632 11348
rect 666 11314 715 11348
rect 583 11280 715 11314
rect 583 11246 632 11280
rect 666 11246 715 11280
rect 583 11212 715 11246
rect 583 11178 632 11212
rect 666 11178 715 11212
rect 583 11144 715 11178
rect 583 11110 632 11144
rect 666 11110 715 11144
rect 583 11076 715 11110
rect 583 11042 632 11076
rect 666 11042 715 11076
rect 583 11008 715 11042
rect 583 10974 632 11008
rect 666 10974 715 11008
rect 583 10940 715 10974
rect 583 10906 632 10940
rect 666 10906 715 10940
rect 583 10872 715 10906
rect 583 10838 632 10872
rect 666 10838 715 10872
rect 583 10804 715 10838
rect 583 10770 632 10804
rect 666 10770 715 10804
rect 583 10736 715 10770
rect 583 10702 632 10736
rect 666 10702 715 10736
rect 583 10668 715 10702
rect 583 10634 632 10668
rect 666 10634 715 10668
rect 583 10600 715 10634
rect 583 10566 632 10600
rect 666 10566 715 10600
rect 583 10532 715 10566
rect 583 10498 632 10532
rect 666 10498 715 10532
rect 583 10464 715 10498
rect 583 10430 632 10464
rect 666 10430 715 10464
rect 583 10396 715 10430
rect 583 10362 632 10396
rect 666 10362 715 10396
rect 583 10328 715 10362
rect 583 10294 632 10328
rect 666 10294 715 10328
rect 583 10260 715 10294
rect 583 10226 632 10260
rect 666 10226 715 10260
rect 1659 31349 13357 31379
rect 1659 30975 2119 31349
rect 12897 30975 13357 31349
rect 1659 30945 13357 30975
rect 1659 30915 2093 30945
rect 1659 27481 1689 30915
rect 2063 27481 2093 30915
rect 1659 27451 2093 27481
rect 12923 30915 13357 30945
rect 12923 27481 12953 30915
rect 13327 27481 13357 30915
rect 12923 27451 13357 27481
rect 1659 27421 13357 27451
rect 1659 27047 2119 27421
rect 12897 27047 13357 27421
rect 1659 27017 13357 27047
rect 14247 34672 14381 34706
rect 14247 34638 14297 34672
rect 14331 34638 14381 34672
rect 14247 34604 14381 34638
rect 14247 34570 14297 34604
rect 14331 34570 14381 34604
rect 14247 34536 14381 34570
rect 14247 34502 14297 34536
rect 14331 34502 14381 34536
rect 14247 34468 14381 34502
rect 14247 34434 14297 34468
rect 14331 34434 14381 34468
rect 14247 34400 14381 34434
rect 14247 34366 14297 34400
rect 14331 34366 14381 34400
rect 14247 34332 14381 34366
rect 14247 34298 14297 34332
rect 14331 34298 14381 34332
rect 14247 34264 14381 34298
rect 14247 34230 14297 34264
rect 14331 34230 14381 34264
rect 14247 34196 14381 34230
rect 14247 34162 14297 34196
rect 14331 34162 14381 34196
rect 14247 34128 14381 34162
rect 14247 34094 14297 34128
rect 14331 34094 14381 34128
rect 14247 34060 14381 34094
rect 14247 34026 14297 34060
rect 14331 34026 14381 34060
rect 14247 33992 14381 34026
rect 14247 33958 14297 33992
rect 14331 33958 14381 33992
rect 14247 33924 14381 33958
rect 14247 33890 14297 33924
rect 14331 33890 14381 33924
rect 14247 33856 14381 33890
rect 14247 33822 14297 33856
rect 14331 33822 14381 33856
rect 14247 33788 14381 33822
rect 14247 33754 14297 33788
rect 14331 33754 14381 33788
rect 14247 33720 14381 33754
rect 14247 33686 14297 33720
rect 14331 33686 14381 33720
rect 14247 33652 14381 33686
rect 14247 33618 14297 33652
rect 14331 33618 14381 33652
rect 14247 33584 14381 33618
rect 14247 33550 14297 33584
rect 14331 33550 14381 33584
rect 14247 33516 14381 33550
rect 14247 33482 14297 33516
rect 14331 33482 14381 33516
rect 14247 33448 14381 33482
rect 14247 33414 14297 33448
rect 14331 33414 14381 33448
rect 14247 33380 14381 33414
rect 14247 33346 14297 33380
rect 14331 33346 14381 33380
rect 14247 33312 14381 33346
rect 14247 33278 14297 33312
rect 14331 33278 14381 33312
rect 14247 33244 14381 33278
rect 14247 33210 14297 33244
rect 14331 33210 14381 33244
rect 14247 33176 14381 33210
rect 14247 33142 14297 33176
rect 14331 33142 14381 33176
rect 14247 33108 14381 33142
rect 14247 33074 14297 33108
rect 14331 33074 14381 33108
rect 14247 33040 14381 33074
rect 14247 33006 14297 33040
rect 14331 33006 14381 33040
rect 14247 32972 14381 33006
rect 14247 32938 14297 32972
rect 14331 32938 14381 32972
rect 14247 32904 14381 32938
rect 14247 32870 14297 32904
rect 14331 32870 14381 32904
rect 14247 32836 14381 32870
rect 14247 32802 14297 32836
rect 14331 32802 14381 32836
rect 14247 32768 14381 32802
rect 14247 32734 14297 32768
rect 14331 32734 14381 32768
rect 14247 32700 14381 32734
rect 14247 32666 14297 32700
rect 14331 32666 14381 32700
rect 14247 32632 14381 32666
rect 14247 32598 14297 32632
rect 14331 32598 14381 32632
rect 14247 32564 14381 32598
rect 14247 32530 14297 32564
rect 14331 32530 14381 32564
rect 14247 32496 14381 32530
rect 14247 32462 14297 32496
rect 14331 32462 14381 32496
rect 14247 32428 14381 32462
rect 14247 32394 14297 32428
rect 14331 32394 14381 32428
rect 14247 32360 14381 32394
rect 14247 32326 14297 32360
rect 14331 32326 14381 32360
rect 14247 32292 14381 32326
rect 14247 32258 14297 32292
rect 14331 32258 14381 32292
rect 14247 32224 14381 32258
rect 14247 32190 14297 32224
rect 14331 32190 14381 32224
rect 14247 32156 14381 32190
rect 14247 32122 14297 32156
rect 14331 32122 14381 32156
rect 14247 32088 14381 32122
rect 14247 32054 14297 32088
rect 14331 32054 14381 32088
rect 14247 32020 14381 32054
rect 14247 31986 14297 32020
rect 14331 31986 14381 32020
rect 14247 31952 14381 31986
rect 14247 31918 14297 31952
rect 14331 31918 14381 31952
rect 14247 31884 14381 31918
rect 14247 31850 14297 31884
rect 14331 31850 14381 31884
rect 14247 31816 14381 31850
rect 14247 31782 14297 31816
rect 14331 31782 14381 31816
rect 14247 31748 14381 31782
rect 14247 31714 14297 31748
rect 14331 31714 14381 31748
rect 14247 31680 14381 31714
rect 14247 31646 14297 31680
rect 14331 31646 14381 31680
rect 14247 31612 14381 31646
rect 14247 31578 14297 31612
rect 14331 31578 14381 31612
rect 14247 31544 14381 31578
rect 14247 31510 14297 31544
rect 14331 31510 14381 31544
rect 14247 31476 14381 31510
rect 14247 31442 14297 31476
rect 14331 31442 14381 31476
rect 14247 31408 14381 31442
rect 14247 31374 14297 31408
rect 14331 31374 14381 31408
rect 14247 31340 14381 31374
rect 14247 31306 14297 31340
rect 14331 31306 14381 31340
rect 14247 31272 14381 31306
rect 14247 31238 14297 31272
rect 14331 31238 14381 31272
rect 14247 31204 14381 31238
rect 14247 31170 14297 31204
rect 14331 31170 14381 31204
rect 14247 31136 14381 31170
rect 14247 31102 14297 31136
rect 14331 31102 14381 31136
rect 14247 31068 14381 31102
rect 14247 31034 14297 31068
rect 14331 31034 14381 31068
rect 14247 31000 14381 31034
rect 14247 30966 14297 31000
rect 14331 30966 14381 31000
rect 14247 30932 14381 30966
rect 14247 30898 14297 30932
rect 14331 30898 14381 30932
rect 14247 30864 14381 30898
rect 14247 30830 14297 30864
rect 14331 30830 14381 30864
rect 14247 30796 14381 30830
rect 14247 30762 14297 30796
rect 14331 30762 14381 30796
rect 14247 30728 14381 30762
rect 14247 30694 14297 30728
rect 14331 30694 14381 30728
rect 14247 30660 14381 30694
rect 14247 30626 14297 30660
rect 14331 30626 14381 30660
rect 14247 30592 14381 30626
rect 14247 30558 14297 30592
rect 14331 30558 14381 30592
rect 14247 30524 14381 30558
rect 14247 30490 14297 30524
rect 14331 30490 14381 30524
rect 14247 30456 14381 30490
rect 14247 30422 14297 30456
rect 14331 30422 14381 30456
rect 14247 30388 14381 30422
rect 14247 30354 14297 30388
rect 14331 30354 14381 30388
rect 14247 30320 14381 30354
rect 14247 30286 14297 30320
rect 14331 30286 14381 30320
rect 14247 30252 14381 30286
rect 14247 30218 14297 30252
rect 14331 30218 14381 30252
rect 14247 30184 14381 30218
rect 14247 30150 14297 30184
rect 14331 30150 14381 30184
rect 14247 30116 14381 30150
rect 14247 30082 14297 30116
rect 14331 30082 14381 30116
rect 14247 30048 14381 30082
rect 14247 30014 14297 30048
rect 14331 30014 14381 30048
rect 14247 29980 14381 30014
rect 14247 29946 14297 29980
rect 14331 29946 14381 29980
rect 14247 29912 14381 29946
rect 14247 29878 14297 29912
rect 14331 29878 14381 29912
rect 14247 29844 14381 29878
rect 14247 29810 14297 29844
rect 14331 29810 14381 29844
rect 14247 29776 14381 29810
rect 14247 29742 14297 29776
rect 14331 29742 14381 29776
rect 14247 29708 14381 29742
rect 14247 29674 14297 29708
rect 14331 29674 14381 29708
rect 14247 29640 14381 29674
rect 14247 29606 14297 29640
rect 14331 29606 14381 29640
rect 14247 29572 14381 29606
rect 14247 29538 14297 29572
rect 14331 29538 14381 29572
rect 14247 29504 14381 29538
rect 14247 29470 14297 29504
rect 14331 29470 14381 29504
rect 14247 29436 14381 29470
rect 14247 29402 14297 29436
rect 14331 29402 14381 29436
rect 14247 29368 14381 29402
rect 14247 29334 14297 29368
rect 14331 29334 14381 29368
rect 14247 29300 14381 29334
rect 14247 29266 14297 29300
rect 14331 29266 14381 29300
rect 14247 29232 14381 29266
rect 14247 29198 14297 29232
rect 14331 29198 14381 29232
rect 14247 29164 14381 29198
rect 14247 29130 14297 29164
rect 14331 29130 14381 29164
rect 14247 29096 14381 29130
rect 14247 29062 14297 29096
rect 14331 29062 14381 29096
rect 14247 29028 14381 29062
rect 14247 28994 14297 29028
rect 14331 28994 14381 29028
rect 14247 28960 14381 28994
rect 14247 28926 14297 28960
rect 14331 28926 14381 28960
rect 14247 28892 14381 28926
rect 14247 28858 14297 28892
rect 14331 28858 14381 28892
rect 14247 28824 14381 28858
rect 14247 28790 14297 28824
rect 14331 28790 14381 28824
rect 14247 28756 14381 28790
rect 14247 28722 14297 28756
rect 14331 28722 14381 28756
rect 14247 28688 14381 28722
rect 14247 28654 14297 28688
rect 14331 28654 14381 28688
rect 14247 28620 14381 28654
rect 14247 28586 14297 28620
rect 14331 28586 14381 28620
rect 14247 28552 14381 28586
rect 14247 28518 14297 28552
rect 14331 28518 14381 28552
rect 14247 28484 14381 28518
rect 14247 28450 14297 28484
rect 14331 28450 14381 28484
rect 14247 28416 14381 28450
rect 14247 28382 14297 28416
rect 14331 28382 14381 28416
rect 14247 28348 14381 28382
rect 14247 28314 14297 28348
rect 14331 28314 14381 28348
rect 14247 28280 14381 28314
rect 14247 28246 14297 28280
rect 14331 28246 14381 28280
rect 14247 28212 14381 28246
rect 14247 28178 14297 28212
rect 14331 28178 14381 28212
rect 14247 28144 14381 28178
rect 14247 28110 14297 28144
rect 14331 28110 14381 28144
rect 14247 28076 14381 28110
rect 14247 28042 14297 28076
rect 14331 28042 14381 28076
rect 14247 28008 14381 28042
rect 14247 27974 14297 28008
rect 14331 27974 14381 28008
rect 14247 27940 14381 27974
rect 14247 27906 14297 27940
rect 14331 27906 14381 27940
rect 14247 27872 14381 27906
rect 14247 27838 14297 27872
rect 14331 27838 14381 27872
rect 14247 27804 14381 27838
rect 14247 27770 14297 27804
rect 14331 27770 14381 27804
rect 14247 27736 14381 27770
rect 14247 27702 14297 27736
rect 14331 27702 14381 27736
rect 14247 27668 14381 27702
rect 14247 27634 14297 27668
rect 14331 27634 14381 27668
rect 14247 27600 14381 27634
rect 14247 27566 14297 27600
rect 14331 27566 14381 27600
rect 14247 27532 14381 27566
rect 14247 27498 14297 27532
rect 14331 27498 14381 27532
rect 14247 27464 14381 27498
rect 14247 27430 14297 27464
rect 14331 27430 14381 27464
rect 14247 27396 14381 27430
rect 14247 27362 14297 27396
rect 14331 27362 14381 27396
rect 14247 27328 14381 27362
rect 14247 27294 14297 27328
rect 14331 27294 14381 27328
rect 14247 27260 14381 27294
rect 14247 27226 14297 27260
rect 14331 27226 14381 27260
rect 14247 27192 14381 27226
rect 14247 27158 14297 27192
rect 14331 27158 14381 27192
rect 14247 27124 14381 27158
rect 14247 27090 14297 27124
rect 14331 27090 14381 27124
rect 14247 27056 14381 27090
rect 14247 27022 14297 27056
rect 14331 27022 14381 27056
rect 14247 26988 14381 27022
rect 14247 26954 14297 26988
rect 14331 26954 14381 26988
rect 14247 26920 14381 26954
rect 14247 26886 14297 26920
rect 14331 26886 14381 26920
rect 14247 26852 14381 26886
rect 14247 26818 14297 26852
rect 14331 26818 14381 26852
rect 14247 26784 14381 26818
rect 14247 26750 14297 26784
rect 14331 26750 14381 26784
rect 14247 26716 14381 26750
rect 14247 26682 14297 26716
rect 14331 26682 14381 26716
rect 14247 26648 14381 26682
rect 14247 26614 14297 26648
rect 14331 26614 14381 26648
rect 14247 26580 14381 26614
rect 14247 26546 14297 26580
rect 14331 26546 14381 26580
rect 14247 26512 14381 26546
rect 14247 26478 14297 26512
rect 14331 26478 14381 26512
rect 14247 26444 14381 26478
rect 14247 26410 14297 26444
rect 14331 26410 14381 26444
rect 14247 26376 14381 26410
rect 14247 26342 14297 26376
rect 14331 26342 14381 26376
rect 14247 26308 14381 26342
rect 14247 26274 14297 26308
rect 14331 26274 14381 26308
rect 14247 26240 14381 26274
rect 14247 26206 14297 26240
rect 14331 26206 14381 26240
rect 14247 26172 14381 26206
rect 14247 26138 14297 26172
rect 14331 26138 14381 26172
rect 14247 26104 14381 26138
rect 14247 26070 14297 26104
rect 14331 26070 14381 26104
rect 14247 26036 14381 26070
rect 14247 26002 14297 26036
rect 14331 26002 14381 26036
rect 14247 25968 14381 26002
rect 14247 25934 14297 25968
rect 14331 25934 14381 25968
rect 14247 25900 14381 25934
rect 14247 25866 14297 25900
rect 14331 25866 14381 25900
rect 14247 25832 14381 25866
rect 14247 25798 14297 25832
rect 14331 25798 14381 25832
rect 14247 25764 14381 25798
rect 14247 25730 14297 25764
rect 14331 25730 14381 25764
rect 14247 25696 14381 25730
rect 14247 25662 14297 25696
rect 14331 25662 14381 25696
rect 14247 25628 14381 25662
rect 14247 25594 14297 25628
rect 14331 25594 14381 25628
rect 14247 25560 14381 25594
rect 14247 25526 14297 25560
rect 14331 25526 14381 25560
rect 14247 25492 14381 25526
rect 14247 25458 14297 25492
rect 14331 25458 14381 25492
rect 14247 25424 14381 25458
rect 14247 25390 14297 25424
rect 14331 25390 14381 25424
rect 14247 25356 14381 25390
rect 14247 25322 14297 25356
rect 14331 25322 14381 25356
rect 14247 25288 14381 25322
rect 14247 25254 14297 25288
rect 14331 25254 14381 25288
rect 14247 25220 14381 25254
rect 14247 25186 14297 25220
rect 14331 25186 14381 25220
rect 14247 25152 14381 25186
rect 14247 25118 14297 25152
rect 14331 25118 14381 25152
rect 14247 25084 14381 25118
rect 14247 25050 14297 25084
rect 14331 25050 14381 25084
rect 14247 25016 14381 25050
rect 14247 24982 14297 25016
rect 14331 24982 14381 25016
rect 14247 24948 14381 24982
rect 14247 24914 14297 24948
rect 14331 24914 14381 24948
rect 14247 24880 14381 24914
rect 14247 24846 14297 24880
rect 14331 24846 14381 24880
rect 14247 24812 14381 24846
rect 14247 24778 14297 24812
rect 14331 24778 14381 24812
rect 14247 24744 14381 24778
rect 14247 24710 14297 24744
rect 14331 24710 14381 24744
rect 14247 24676 14381 24710
rect 14247 24642 14297 24676
rect 14331 24642 14381 24676
rect 14247 24608 14381 24642
rect 14247 24574 14297 24608
rect 14331 24574 14381 24608
rect 14247 24540 14381 24574
rect 14247 24506 14297 24540
rect 14331 24506 14381 24540
rect 14247 24472 14381 24506
rect 14247 24438 14297 24472
rect 14331 24438 14381 24472
rect 14247 24404 14381 24438
rect 14247 24370 14297 24404
rect 14331 24370 14381 24404
rect 14247 24336 14381 24370
rect 14247 24302 14297 24336
rect 14331 24302 14381 24336
rect 14247 24268 14381 24302
rect 14247 24234 14297 24268
rect 14331 24234 14381 24268
rect 14247 24200 14381 24234
rect 14247 24166 14297 24200
rect 14331 24166 14381 24200
rect 14247 24132 14381 24166
rect 14247 24098 14297 24132
rect 14331 24098 14381 24132
rect 14247 24064 14381 24098
rect 14247 24030 14297 24064
rect 14331 24030 14381 24064
rect 14247 23996 14381 24030
rect 14247 23962 14297 23996
rect 14331 23962 14381 23996
rect 14247 23928 14381 23962
rect 14247 23894 14297 23928
rect 14331 23894 14381 23928
rect 14247 23860 14381 23894
rect 14247 23826 14297 23860
rect 14331 23826 14381 23860
rect 14247 23792 14381 23826
rect 14247 23758 14297 23792
rect 14331 23758 14381 23792
rect 14247 23724 14381 23758
rect 14247 23690 14297 23724
rect 14331 23690 14381 23724
rect 14247 23656 14381 23690
rect 14247 23622 14297 23656
rect 14331 23622 14381 23656
rect 14247 23588 14381 23622
rect 14247 23554 14297 23588
rect 14331 23554 14381 23588
rect 14247 23520 14381 23554
rect 14247 23486 14297 23520
rect 14331 23486 14381 23520
rect 14247 23452 14381 23486
rect 14247 23418 14297 23452
rect 14331 23418 14381 23452
rect 14247 23384 14381 23418
rect 14247 23350 14297 23384
rect 14331 23350 14381 23384
rect 14247 23316 14381 23350
rect 14247 23282 14297 23316
rect 14331 23282 14381 23316
rect 14247 23248 14381 23282
rect 14247 23214 14297 23248
rect 14331 23214 14381 23248
rect 14247 23180 14381 23214
rect 14247 23146 14297 23180
rect 14331 23146 14381 23180
rect 14247 23112 14381 23146
rect 14247 23078 14297 23112
rect 14331 23078 14381 23112
rect 14247 23044 14381 23078
rect 14247 23010 14297 23044
rect 14331 23010 14381 23044
rect 14247 22976 14381 23010
rect 14247 22942 14297 22976
rect 14331 22942 14381 22976
rect 14247 22908 14381 22942
rect 14247 22874 14297 22908
rect 14331 22874 14381 22908
rect 14247 22840 14381 22874
rect 14247 22806 14297 22840
rect 14331 22806 14381 22840
rect 14247 22772 14381 22806
rect 14247 22738 14297 22772
rect 14331 22738 14381 22772
rect 14247 22704 14381 22738
rect 14247 22670 14297 22704
rect 14331 22670 14381 22704
rect 14247 22636 14381 22670
rect 14247 22602 14297 22636
rect 14331 22602 14381 22636
rect 14247 22568 14381 22602
rect 14247 22534 14297 22568
rect 14331 22534 14381 22568
rect 14247 22500 14381 22534
rect 14247 22466 14297 22500
rect 14331 22466 14381 22500
rect 14247 22432 14381 22466
rect 14247 22398 14297 22432
rect 14331 22398 14381 22432
rect 14247 22364 14381 22398
rect 14247 22330 14297 22364
rect 14331 22330 14381 22364
rect 14247 22296 14381 22330
rect 14247 22262 14297 22296
rect 14331 22262 14381 22296
rect 14247 22228 14381 22262
rect 14247 22194 14297 22228
rect 14331 22194 14381 22228
rect 14247 22160 14381 22194
rect 14247 22126 14297 22160
rect 14331 22126 14381 22160
rect 14247 22092 14381 22126
rect 14247 22058 14297 22092
rect 14331 22058 14381 22092
rect 14247 22024 14381 22058
rect 14247 21990 14297 22024
rect 14331 21990 14381 22024
rect 14247 21956 14381 21990
rect 14247 21922 14297 21956
rect 14331 21922 14381 21956
rect 14247 21888 14381 21922
rect 14247 21854 14297 21888
rect 14331 21854 14381 21888
rect 14247 21820 14381 21854
rect 14247 21786 14297 21820
rect 14331 21786 14381 21820
rect 14247 21752 14381 21786
rect 14247 21718 14297 21752
rect 14331 21718 14381 21752
rect 14247 21684 14381 21718
rect 14247 21650 14297 21684
rect 14331 21650 14381 21684
rect 14247 21616 14381 21650
rect 14247 21582 14297 21616
rect 14331 21582 14381 21616
rect 14247 21548 14381 21582
rect 14247 21514 14297 21548
rect 14331 21514 14381 21548
rect 14247 21480 14381 21514
rect 14247 21446 14297 21480
rect 14331 21446 14381 21480
rect 14247 21412 14381 21446
rect 14247 21378 14297 21412
rect 14331 21378 14381 21412
rect 14247 21344 14381 21378
rect 14247 21310 14297 21344
rect 14331 21310 14381 21344
rect 14247 21276 14381 21310
rect 14247 21242 14297 21276
rect 14331 21242 14381 21276
rect 14247 21208 14381 21242
rect 14247 21174 14297 21208
rect 14331 21174 14381 21208
rect 14247 21140 14381 21174
rect 14247 21106 14297 21140
rect 14331 21106 14381 21140
rect 14247 21072 14381 21106
rect 14247 21038 14297 21072
rect 14331 21038 14381 21072
rect 14247 21004 14381 21038
rect 14247 20970 14297 21004
rect 14331 20970 14381 21004
rect 14247 20936 14381 20970
rect 14247 20902 14297 20936
rect 14331 20902 14381 20936
rect 14247 20868 14381 20902
rect 14247 20834 14297 20868
rect 14331 20834 14381 20868
rect 14247 20800 14381 20834
rect 14247 20766 14297 20800
rect 14331 20766 14381 20800
rect 14247 20732 14381 20766
rect 14247 20698 14297 20732
rect 14331 20698 14381 20732
rect 14247 20664 14381 20698
rect 14247 20630 14297 20664
rect 14331 20630 14381 20664
rect 14247 20596 14381 20630
rect 14247 20562 14297 20596
rect 14331 20562 14381 20596
rect 14247 20528 14381 20562
rect 14247 20494 14297 20528
rect 14331 20494 14381 20528
rect 14247 20460 14381 20494
rect 14247 20426 14297 20460
rect 14331 20426 14381 20460
rect 14247 20392 14381 20426
rect 14247 20358 14297 20392
rect 14331 20358 14381 20392
rect 14247 20324 14381 20358
rect 14247 20290 14297 20324
rect 14331 20290 14381 20324
rect 14247 20256 14381 20290
rect 14247 20222 14297 20256
rect 14331 20222 14381 20256
rect 14247 20188 14381 20222
rect 14247 20154 14297 20188
rect 14331 20154 14381 20188
rect 14247 20120 14381 20154
rect 14247 20086 14297 20120
rect 14331 20086 14381 20120
rect 14247 20052 14381 20086
rect 14247 20018 14297 20052
rect 14331 20018 14381 20052
rect 14247 19984 14381 20018
rect 14247 19950 14297 19984
rect 14331 19950 14381 19984
rect 14247 19916 14381 19950
rect 14247 19882 14297 19916
rect 14331 19882 14381 19916
rect 14247 19848 14381 19882
rect 14247 19814 14297 19848
rect 14331 19814 14381 19848
rect 14247 19780 14381 19814
rect 14247 19746 14297 19780
rect 14331 19746 14381 19780
rect 14247 19712 14381 19746
rect 14247 19678 14297 19712
rect 14331 19678 14381 19712
rect 14247 19644 14381 19678
rect 14247 19610 14297 19644
rect 14331 19610 14381 19644
rect 14247 19576 14381 19610
rect 14247 19542 14297 19576
rect 14331 19542 14381 19576
rect 14247 19508 14381 19542
rect 14247 19474 14297 19508
rect 14331 19474 14381 19508
rect 14247 19440 14381 19474
rect 14247 19406 14297 19440
rect 14331 19406 14381 19440
rect 14247 19372 14381 19406
rect 14247 19338 14297 19372
rect 14331 19338 14381 19372
rect 14247 19304 14381 19338
rect 14247 19270 14297 19304
rect 14331 19270 14381 19304
rect 14247 19236 14381 19270
rect 14247 19202 14297 19236
rect 14331 19202 14381 19236
rect 14247 19168 14381 19202
rect 14247 19134 14297 19168
rect 14331 19134 14381 19168
rect 14247 19100 14381 19134
rect 14247 19066 14297 19100
rect 14331 19066 14381 19100
rect 14247 19032 14381 19066
rect 14247 18998 14297 19032
rect 14331 18998 14381 19032
rect 14247 18964 14381 18998
rect 14247 18930 14297 18964
rect 14331 18930 14381 18964
rect 14247 18896 14381 18930
rect 14247 18862 14297 18896
rect 14331 18862 14381 18896
rect 14247 18828 14381 18862
rect 14247 18794 14297 18828
rect 14331 18794 14381 18828
rect 14247 18760 14381 18794
rect 14247 18726 14297 18760
rect 14331 18726 14381 18760
rect 14247 18692 14381 18726
rect 14247 18658 14297 18692
rect 14331 18658 14381 18692
rect 14247 18624 14381 18658
rect 14247 18590 14297 18624
rect 14331 18590 14381 18624
rect 14247 18556 14381 18590
rect 14247 18522 14297 18556
rect 14331 18522 14381 18556
rect 14247 18488 14381 18522
rect 14247 18454 14297 18488
rect 14331 18454 14381 18488
rect 14247 18420 14381 18454
rect 14247 18386 14297 18420
rect 14331 18386 14381 18420
rect 14247 18352 14381 18386
rect 14247 18318 14297 18352
rect 14331 18318 14381 18352
rect 14247 18284 14381 18318
rect 14247 18250 14297 18284
rect 14331 18250 14381 18284
rect 14247 18216 14381 18250
rect 14247 18182 14297 18216
rect 14331 18182 14381 18216
rect 14247 18148 14381 18182
rect 14247 18114 14297 18148
rect 14331 18114 14381 18148
rect 14247 18080 14381 18114
rect 14247 18046 14297 18080
rect 14331 18046 14381 18080
rect 14247 18012 14381 18046
rect 14247 17978 14297 18012
rect 14331 17978 14381 18012
rect 14247 17944 14381 17978
rect 14247 17910 14297 17944
rect 14331 17910 14381 17944
rect 14247 17876 14381 17910
rect 14247 17842 14297 17876
rect 14331 17842 14381 17876
rect 14247 17808 14381 17842
rect 14247 17774 14297 17808
rect 14331 17774 14381 17808
rect 14247 17740 14381 17774
rect 14247 17706 14297 17740
rect 14331 17706 14381 17740
rect 14247 17672 14381 17706
rect 14247 17638 14297 17672
rect 14331 17638 14381 17672
rect 14247 17604 14381 17638
rect 14247 17570 14297 17604
rect 14331 17570 14381 17604
rect 14247 17536 14381 17570
rect 14247 17502 14297 17536
rect 14331 17502 14381 17536
rect 14247 17468 14381 17502
rect 14247 17434 14297 17468
rect 14331 17434 14381 17468
rect 14247 17400 14381 17434
rect 14247 17366 14297 17400
rect 14331 17366 14381 17400
rect 14247 17332 14381 17366
rect 14247 17298 14297 17332
rect 14331 17298 14381 17332
rect 14247 17264 14381 17298
rect 14247 17230 14297 17264
rect 14331 17230 14381 17264
rect 14247 17196 14381 17230
rect 14247 17162 14297 17196
rect 14331 17162 14381 17196
rect 14247 17128 14381 17162
rect 14247 17094 14297 17128
rect 14331 17094 14381 17128
rect 14247 17060 14381 17094
rect 14247 17026 14297 17060
rect 14331 17026 14381 17060
rect 14247 16992 14381 17026
rect 14247 16958 14297 16992
rect 14331 16958 14381 16992
rect 14247 16924 14381 16958
rect 14247 16890 14297 16924
rect 14331 16890 14381 16924
rect 14247 16856 14381 16890
rect 14247 16822 14297 16856
rect 14331 16822 14381 16856
rect 14247 16788 14381 16822
rect 14247 16754 14297 16788
rect 14331 16754 14381 16788
rect 14247 16720 14381 16754
rect 14247 16686 14297 16720
rect 14331 16686 14381 16720
rect 14247 16652 14381 16686
rect 14247 16618 14297 16652
rect 14331 16618 14381 16652
rect 14247 16584 14381 16618
rect 14247 16550 14297 16584
rect 14331 16550 14381 16584
rect 14247 16516 14381 16550
rect 14247 16482 14297 16516
rect 14331 16482 14381 16516
rect 14247 16448 14381 16482
rect 14247 16414 14297 16448
rect 14331 16414 14381 16448
rect 14247 16380 14381 16414
rect 14247 16346 14297 16380
rect 14331 16346 14381 16380
rect 14247 16312 14381 16346
rect 14247 16278 14297 16312
rect 14331 16278 14381 16312
rect 14247 16244 14381 16278
rect 14247 16210 14297 16244
rect 14331 16210 14381 16244
rect 14247 16176 14381 16210
rect 14247 16142 14297 16176
rect 14331 16142 14381 16176
rect 14247 16108 14381 16142
rect 14247 16074 14297 16108
rect 14331 16074 14381 16108
rect 14247 16040 14381 16074
rect 14247 16006 14297 16040
rect 14331 16006 14381 16040
rect 14247 15972 14381 16006
rect 14247 15938 14297 15972
rect 14331 15938 14381 15972
rect 14247 15904 14381 15938
rect 14247 15870 14297 15904
rect 14331 15870 14381 15904
rect 14247 15836 14381 15870
rect 14247 15802 14297 15836
rect 14331 15802 14381 15836
rect 14247 15768 14381 15802
rect 14247 15734 14297 15768
rect 14331 15734 14381 15768
rect 14247 15700 14381 15734
rect 14247 15666 14297 15700
rect 14331 15666 14381 15700
rect 14247 15632 14381 15666
rect 14247 15598 14297 15632
rect 14331 15598 14381 15632
rect 14247 15564 14381 15598
rect 14247 15530 14297 15564
rect 14331 15530 14381 15564
rect 14247 15496 14381 15530
rect 14247 15462 14297 15496
rect 14331 15462 14381 15496
rect 14247 15428 14381 15462
rect 14247 15394 14297 15428
rect 14331 15394 14381 15428
rect 14247 15360 14381 15394
rect 14247 15326 14297 15360
rect 14331 15326 14381 15360
rect 14247 15292 14381 15326
rect 14247 15258 14297 15292
rect 14331 15258 14381 15292
rect 14247 15224 14381 15258
rect 14247 15190 14297 15224
rect 14331 15190 14381 15224
rect 14247 15156 14381 15190
rect 14247 15122 14297 15156
rect 14331 15122 14381 15156
rect 14247 15088 14381 15122
rect 14247 15054 14297 15088
rect 14331 15054 14381 15088
rect 14247 15020 14381 15054
rect 14247 14986 14297 15020
rect 14331 14986 14381 15020
rect 14247 14952 14381 14986
rect 14247 14918 14297 14952
rect 14331 14918 14381 14952
rect 14247 14884 14381 14918
rect 14247 14850 14297 14884
rect 14331 14850 14381 14884
rect 14247 14816 14381 14850
rect 14247 14782 14297 14816
rect 14331 14782 14381 14816
rect 14247 14748 14381 14782
rect 14247 14714 14297 14748
rect 14331 14714 14381 14748
rect 14247 14680 14381 14714
rect 14247 14646 14297 14680
rect 14331 14646 14381 14680
rect 14247 14612 14381 14646
rect 14247 14578 14297 14612
rect 14331 14578 14381 14612
rect 14247 14544 14381 14578
rect 14247 14510 14297 14544
rect 14331 14510 14381 14544
rect 14247 14476 14381 14510
rect 14247 14442 14297 14476
rect 14331 14442 14381 14476
rect 14247 14408 14381 14442
rect 14247 14374 14297 14408
rect 14331 14374 14381 14408
rect 14247 14340 14381 14374
rect 14247 14306 14297 14340
rect 14331 14306 14381 14340
rect 14247 14272 14381 14306
rect 14247 14238 14297 14272
rect 14331 14238 14381 14272
rect 14247 14204 14381 14238
rect 14247 14170 14297 14204
rect 14331 14170 14381 14204
rect 14247 14136 14381 14170
rect 14247 14102 14297 14136
rect 14331 14102 14381 14136
rect 14247 14068 14381 14102
rect 14247 14034 14297 14068
rect 14331 14034 14381 14068
rect 14247 14000 14381 14034
rect 14247 13966 14297 14000
rect 14331 13966 14381 14000
rect 14247 13932 14381 13966
rect 14247 13898 14297 13932
rect 14331 13898 14381 13932
rect 14247 13864 14381 13898
rect 14247 13830 14297 13864
rect 14331 13830 14381 13864
rect 14247 13796 14381 13830
rect 14247 13762 14297 13796
rect 14331 13762 14381 13796
rect 14247 13728 14381 13762
rect 14247 13694 14297 13728
rect 14331 13694 14381 13728
rect 14247 13660 14381 13694
rect 14247 13626 14297 13660
rect 14331 13626 14381 13660
rect 14247 13592 14381 13626
rect 14247 13558 14297 13592
rect 14331 13558 14381 13592
rect 14247 13524 14381 13558
rect 14247 13490 14297 13524
rect 14331 13490 14381 13524
rect 14247 13456 14381 13490
rect 14247 13422 14297 13456
rect 14331 13422 14381 13456
rect 14247 13388 14381 13422
rect 14247 13354 14297 13388
rect 14331 13354 14381 13388
rect 14247 13320 14381 13354
rect 14247 13286 14297 13320
rect 14331 13286 14381 13320
rect 14247 13252 14381 13286
rect 14247 13218 14297 13252
rect 14331 13218 14381 13252
rect 14247 13184 14381 13218
rect 14247 13150 14297 13184
rect 14331 13150 14381 13184
rect 14247 13116 14381 13150
rect 14247 13082 14297 13116
rect 14331 13082 14381 13116
rect 14247 13048 14381 13082
rect 14247 13014 14297 13048
rect 14331 13014 14381 13048
rect 14247 12980 14381 13014
rect 14247 12946 14297 12980
rect 14331 12946 14381 12980
rect 14247 12912 14381 12946
rect 14247 12878 14297 12912
rect 14331 12878 14381 12912
rect 14247 12844 14381 12878
rect 14247 12810 14297 12844
rect 14331 12810 14381 12844
rect 14247 12776 14381 12810
rect 14247 12742 14297 12776
rect 14331 12742 14381 12776
rect 14247 12708 14381 12742
rect 14247 12674 14297 12708
rect 14331 12674 14381 12708
rect 14247 12640 14381 12674
rect 14247 12606 14297 12640
rect 14331 12606 14381 12640
rect 14247 12572 14381 12606
rect 14247 12538 14297 12572
rect 14331 12538 14381 12572
rect 14247 12504 14381 12538
rect 14247 12470 14297 12504
rect 14331 12470 14381 12504
rect 14247 12436 14381 12470
rect 14247 12402 14297 12436
rect 14331 12402 14381 12436
rect 14247 12368 14381 12402
rect 14247 12334 14297 12368
rect 14331 12334 14381 12368
rect 14247 12300 14381 12334
rect 14247 12266 14297 12300
rect 14331 12266 14381 12300
rect 14247 12232 14381 12266
rect 14247 12198 14297 12232
rect 14331 12198 14381 12232
rect 14247 12164 14381 12198
rect 14247 12130 14297 12164
rect 14331 12130 14381 12164
rect 14247 12096 14381 12130
rect 14247 12062 14297 12096
rect 14331 12062 14381 12096
rect 14247 12028 14381 12062
rect 14247 11994 14297 12028
rect 14331 11994 14381 12028
rect 14247 11960 14381 11994
rect 14247 11926 14297 11960
rect 14331 11926 14381 11960
rect 14247 11892 14381 11926
rect 14247 11858 14297 11892
rect 14331 11858 14381 11892
rect 14247 11824 14381 11858
rect 14247 11790 14297 11824
rect 14331 11790 14381 11824
rect 14247 11756 14381 11790
rect 14247 11722 14297 11756
rect 14331 11722 14381 11756
rect 14247 11688 14381 11722
rect 14247 11654 14297 11688
rect 14331 11654 14381 11688
rect 14247 11620 14381 11654
rect 14247 11586 14297 11620
rect 14331 11586 14381 11620
rect 14247 11552 14381 11586
rect 14247 11518 14297 11552
rect 14331 11518 14381 11552
rect 14247 11484 14381 11518
rect 14247 11450 14297 11484
rect 14331 11450 14381 11484
rect 14247 11416 14381 11450
rect 14247 11382 14297 11416
rect 14331 11382 14381 11416
rect 14247 11348 14381 11382
rect 14247 11314 14297 11348
rect 14331 11314 14381 11348
rect 14247 11280 14381 11314
rect 14247 11246 14297 11280
rect 14331 11246 14381 11280
rect 14247 11212 14381 11246
rect 14247 11178 14297 11212
rect 14331 11178 14381 11212
rect 14247 11144 14381 11178
rect 14247 11110 14297 11144
rect 14331 11110 14381 11144
rect 14247 11076 14381 11110
rect 14247 11042 14297 11076
rect 14331 11042 14381 11076
rect 14247 11008 14381 11042
rect 14247 10974 14297 11008
rect 14331 10974 14381 11008
rect 14247 10940 14381 10974
rect 14247 10906 14297 10940
rect 14331 10906 14381 10940
rect 14247 10872 14381 10906
rect 14247 10838 14297 10872
rect 14331 10838 14381 10872
rect 14247 10804 14381 10838
rect 14247 10770 14297 10804
rect 14331 10770 14381 10804
rect 14247 10736 14381 10770
rect 14247 10702 14297 10736
rect 14331 10702 14381 10736
rect 14247 10668 14381 10702
rect 14247 10634 14297 10668
rect 14331 10634 14381 10668
rect 14247 10600 14381 10634
rect 14247 10566 14297 10600
rect 14331 10566 14381 10600
rect 14247 10532 14381 10566
rect 14247 10498 14297 10532
rect 14331 10498 14381 10532
rect 14247 10464 14381 10498
rect 14247 10430 14297 10464
rect 14331 10430 14381 10464
rect 14247 10396 14381 10430
rect 14247 10362 14297 10396
rect 14331 10362 14381 10396
rect 14247 10328 14381 10362
rect 14247 10294 14297 10328
rect 14331 10294 14381 10328
rect 14247 10260 14381 10294
rect 583 10192 715 10226
rect 583 10158 632 10192
rect 666 10158 715 10192
rect 583 10124 715 10158
rect 583 10090 632 10124
rect 666 10090 715 10124
rect 583 10056 715 10090
rect 583 10022 632 10056
rect 666 10022 715 10056
rect 583 9988 715 10022
rect 583 9954 632 9988
rect 666 9954 715 9988
rect 583 9920 715 9954
rect 583 9886 632 9920
rect 666 9886 715 9920
rect 583 9825 715 9886
rect 14247 10226 14297 10260
rect 14331 10226 14381 10260
rect 14247 10192 14381 10226
rect 14247 10158 14297 10192
rect 14331 10158 14381 10192
rect 14247 10124 14381 10158
rect 14247 10090 14297 10124
rect 14331 10090 14381 10124
rect 14247 10056 14381 10090
rect 14247 10022 14297 10056
rect 14331 10022 14381 10056
rect 14247 9988 14381 10022
rect 14247 9954 14297 9988
rect 14331 9954 14381 9988
rect 14247 9920 14381 9954
rect 14247 9886 14297 9920
rect 14331 9886 14381 9920
rect 14247 9825 14381 9886
rect 583 9775 14381 9825
rect 583 9741 740 9775
rect 774 9741 808 9775
rect 842 9741 915 9775
rect 949 9741 983 9775
rect 1017 9741 1051 9775
rect 1085 9741 1119 9775
rect 1153 9741 1187 9775
rect 1221 9741 1255 9775
rect 1289 9741 1323 9775
rect 1357 9741 1391 9775
rect 1425 9741 1459 9775
rect 1493 9741 1527 9775
rect 1561 9741 1595 9775
rect 1629 9741 1663 9775
rect 1697 9741 1731 9775
rect 1765 9741 1799 9775
rect 1833 9741 1867 9775
rect 1901 9741 1935 9775
rect 1969 9741 2003 9775
rect 2037 9741 2121 9775
rect 2155 9741 2189 9775
rect 2223 9741 2257 9775
rect 2291 9741 2325 9775
rect 2359 9741 2393 9775
rect 2427 9741 2461 9775
rect 2495 9741 2529 9775
rect 2563 9741 2597 9775
rect 2631 9741 2665 9775
rect 2699 9741 2733 9775
rect 2767 9741 2801 9775
rect 2835 9741 2869 9775
rect 2903 9741 2937 9775
rect 2971 9741 3005 9775
rect 3039 9741 3073 9775
rect 3107 9741 3141 9775
rect 3175 9741 3209 9775
rect 3243 9741 3277 9775
rect 3311 9741 3345 9775
rect 3379 9741 3413 9775
rect 3447 9741 3481 9775
rect 3515 9741 3549 9775
rect 3583 9741 3617 9775
rect 3651 9741 3685 9775
rect 3719 9741 3753 9775
rect 3787 9741 3821 9775
rect 3855 9741 3889 9775
rect 3923 9741 3957 9775
rect 3991 9741 4025 9775
rect 4059 9741 4093 9775
rect 4127 9741 4161 9775
rect 4195 9741 4229 9775
rect 4263 9741 4297 9775
rect 4331 9741 4365 9775
rect 4399 9741 4433 9775
rect 4467 9741 4501 9775
rect 4535 9741 4569 9775
rect 4603 9741 4637 9775
rect 4671 9741 4705 9775
rect 4739 9741 4773 9775
rect 4807 9741 4841 9775
rect 4875 9741 4909 9775
rect 4943 9741 4977 9775
rect 5011 9741 5045 9775
rect 5079 9741 5113 9775
rect 5147 9741 5181 9775
rect 5215 9741 5249 9775
rect 5283 9741 5317 9775
rect 5351 9741 5385 9775
rect 5419 9741 5453 9775
rect 5487 9741 5521 9775
rect 5555 9741 5589 9775
rect 5623 9741 5657 9775
rect 5691 9741 5725 9775
rect 5759 9741 5793 9775
rect 5827 9741 5861 9775
rect 5895 9741 5929 9775
rect 5963 9741 5997 9775
rect 6031 9741 6065 9775
rect 6099 9741 6133 9775
rect 6167 9741 6201 9775
rect 6235 9741 6269 9775
rect 6303 9741 6337 9775
rect 6371 9741 6405 9775
rect 6439 9741 6473 9775
rect 6507 9741 6541 9775
rect 6575 9741 6609 9775
rect 6643 9741 6677 9775
rect 6711 9741 6745 9775
rect 6779 9741 6813 9775
rect 6847 9741 6881 9775
rect 6915 9741 6949 9775
rect 6983 9741 7017 9775
rect 7051 9741 7085 9775
rect 7119 9741 7153 9775
rect 7187 9741 7221 9775
rect 7255 9741 7289 9775
rect 7323 9741 7357 9775
rect 7391 9741 7425 9775
rect 7459 9741 7493 9775
rect 7527 9741 7561 9775
rect 7595 9741 7629 9775
rect 7663 9741 7697 9775
rect 7731 9741 7765 9775
rect 7799 9741 7833 9775
rect 7867 9741 7901 9775
rect 7935 9741 7969 9775
rect 8003 9741 8037 9775
rect 8071 9741 8105 9775
rect 8139 9741 8173 9775
rect 8207 9741 8241 9775
rect 8275 9741 8309 9775
rect 8343 9741 8377 9775
rect 8411 9741 8445 9775
rect 8479 9741 8513 9775
rect 8547 9741 8581 9775
rect 8615 9741 8649 9775
rect 8683 9741 8717 9775
rect 8751 9741 8785 9775
rect 8819 9741 8853 9775
rect 8887 9741 8921 9775
rect 8955 9741 8989 9775
rect 9023 9741 9057 9775
rect 9091 9741 9125 9775
rect 9159 9741 9193 9775
rect 9227 9741 9261 9775
rect 9295 9741 9329 9775
rect 9363 9741 9397 9775
rect 9431 9741 9465 9775
rect 9499 9741 9533 9775
rect 9567 9741 9601 9775
rect 9635 9741 9669 9775
rect 9703 9741 9737 9775
rect 9771 9741 9805 9775
rect 9839 9741 9873 9775
rect 9907 9741 9941 9775
rect 9975 9741 10009 9775
rect 10043 9741 10077 9775
rect 10111 9741 10145 9775
rect 10179 9741 10213 9775
rect 10247 9741 10281 9775
rect 10315 9741 10349 9775
rect 10383 9741 10417 9775
rect 10451 9741 10485 9775
rect 10519 9741 10553 9775
rect 10587 9741 10621 9775
rect 10655 9741 10689 9775
rect 10723 9741 10757 9775
rect 10791 9741 10825 9775
rect 10859 9741 10893 9775
rect 10927 9741 10961 9775
rect 10995 9741 11029 9775
rect 11063 9741 11097 9775
rect 11131 9741 11165 9775
rect 11199 9741 11233 9775
rect 11267 9741 11301 9775
rect 11335 9741 11369 9775
rect 11403 9741 11437 9775
rect 11471 9741 11505 9775
rect 11539 9741 11573 9775
rect 11607 9741 11641 9775
rect 11675 9741 11709 9775
rect 11743 9741 11777 9775
rect 11811 9741 11845 9775
rect 11879 9741 11913 9775
rect 11947 9741 11981 9775
rect 12015 9741 12049 9775
rect 12083 9741 12117 9775
rect 12151 9741 12185 9775
rect 12219 9741 12253 9775
rect 12287 9741 12321 9775
rect 12355 9741 12389 9775
rect 12423 9741 12457 9775
rect 12491 9741 12525 9775
rect 12559 9741 12593 9775
rect 12627 9741 12661 9775
rect 12695 9741 12729 9775
rect 12763 9741 12797 9775
rect 12831 9774 14115 9775
rect 12831 9741 12915 9774
rect 583 9740 12915 9741
rect 12949 9740 12983 9774
rect 13017 9740 13051 9774
rect 13085 9740 13119 9774
rect 13153 9740 13187 9774
rect 13221 9740 13255 9774
rect 13289 9740 13323 9774
rect 13357 9740 13391 9774
rect 13425 9740 13459 9774
rect 13493 9740 13527 9774
rect 13561 9740 13595 9774
rect 13629 9740 13663 9774
rect 13697 9740 13731 9774
rect 13765 9740 13799 9774
rect 13833 9740 13867 9774
rect 13901 9740 13935 9774
rect 13969 9740 14003 9774
rect 14037 9741 14115 9774
rect 14149 9741 14183 9775
rect 14217 9741 14381 9775
rect 14037 9740 14381 9741
rect 583 9691 14381 9740
<< mvpsubdiffcont >>
rect 532 36464 566 36498
rect 600 36464 634 36498
rect 668 36464 702 36498
rect 736 36464 770 36498
rect 804 36464 838 36498
rect 872 36464 906 36498
rect 940 36464 974 36498
rect 1008 36464 1042 36498
rect 1076 36464 1110 36498
rect 1144 36464 1178 36498
rect 1212 36464 1246 36498
rect 1280 36464 1314 36498
rect 1348 36464 1382 36498
rect 1416 36464 1450 36498
rect 1484 36464 1518 36498
rect 1552 36464 1586 36498
rect 1620 36464 1654 36498
rect 1688 36464 1722 36498
rect 1756 36464 1790 36498
rect 1824 36464 1858 36498
rect 1892 36464 1926 36498
rect 1960 36464 1994 36498
rect 2028 36464 2062 36498
rect 2096 36464 2130 36498
rect 2164 36464 2198 36498
rect 2232 36464 2266 36498
rect 2300 36464 2334 36498
rect 2368 36464 2402 36498
rect 2436 36464 2470 36498
rect 2504 36464 2538 36498
rect 2572 36464 2606 36498
rect 2640 36464 2674 36498
rect 2708 36464 2742 36498
rect 2776 36464 2810 36498
rect 2844 36464 2878 36498
rect 2912 36464 2946 36498
rect 2980 36464 3014 36498
rect 3048 36464 3082 36498
rect 3116 36464 3150 36498
rect 3184 36464 3218 36498
rect 3252 36464 3286 36498
rect 3320 36464 3354 36498
rect 3388 36464 3422 36498
rect 3456 36464 3490 36498
rect 3524 36464 3558 36498
rect 3592 36464 3626 36498
rect 3660 36464 3694 36498
rect 3728 36464 3762 36498
rect 3796 36464 3830 36498
rect 3864 36464 3898 36498
rect 3932 36464 3966 36498
rect 4000 36464 4034 36498
rect 4068 36464 4102 36498
rect 4136 36464 4170 36498
rect 4204 36464 4238 36498
rect 4272 36464 4306 36498
rect 4340 36464 4374 36498
rect 4408 36464 4442 36498
rect 4476 36464 4510 36498
rect 4544 36464 4578 36498
rect 4612 36464 4646 36498
rect 4680 36464 4714 36498
rect 4748 36464 4782 36498
rect 4816 36464 4850 36498
rect 4884 36464 4918 36498
rect 4952 36464 4986 36498
rect 5020 36464 5054 36498
rect 5088 36464 5122 36498
rect 5156 36464 5190 36498
rect 5224 36464 5258 36498
rect 5292 36464 5326 36498
rect 5360 36464 5394 36498
rect 5428 36464 5462 36498
rect 5496 36464 5530 36498
rect 5564 36464 5598 36498
rect 5632 36464 5666 36498
rect 5700 36464 5734 36498
rect 5768 36464 5802 36498
rect 5836 36464 5870 36498
rect 5904 36464 5938 36498
rect 5972 36464 6006 36498
rect 6040 36464 6074 36498
rect 6108 36464 6142 36498
rect 6176 36464 6210 36498
rect 6244 36464 6278 36498
rect 6312 36464 6346 36498
rect 6380 36464 6414 36498
rect 6448 36464 6482 36498
rect 6516 36464 6550 36498
rect 6584 36464 6618 36498
rect 6652 36464 6686 36498
rect 6720 36464 6754 36498
rect 6788 36464 6822 36498
rect 6856 36464 6890 36498
rect 6924 36464 6958 36498
rect 6992 36464 7026 36498
rect 7060 36464 7094 36498
rect 7128 36464 7162 36498
rect 7196 36464 7230 36498
rect 7264 36464 7298 36498
rect 7332 36464 7366 36498
rect 7400 36464 7434 36498
rect 7468 36464 7502 36498
rect 7536 36464 7570 36498
rect 7604 36464 7638 36498
rect 7672 36464 7706 36498
rect 7740 36464 7774 36498
rect 7808 36464 7842 36498
rect 7876 36464 7910 36498
rect 7944 36464 7978 36498
rect 8012 36464 8046 36498
rect 8080 36464 8114 36498
rect 8148 36464 8182 36498
rect 8216 36464 8250 36498
rect 8284 36464 8318 36498
rect 8352 36464 8386 36498
rect 8420 36464 8454 36498
rect 8488 36464 8522 36498
rect 8556 36464 8590 36498
rect 8624 36464 8658 36498
rect 8692 36464 8726 36498
rect 8760 36464 8794 36498
rect 8828 36464 8862 36498
rect 8896 36464 8930 36498
rect 8964 36464 8998 36498
rect 9032 36464 9066 36498
rect 9100 36464 9134 36498
rect 9168 36464 9202 36498
rect 9236 36464 9270 36498
rect 9304 36464 9338 36498
rect 9372 36464 9406 36498
rect 9440 36464 9474 36498
rect 9508 36464 9542 36498
rect 9576 36464 9610 36498
rect 9644 36464 9678 36498
rect 9712 36464 9746 36498
rect 9780 36464 9814 36498
rect 9848 36464 9882 36498
rect 9916 36464 9950 36498
rect 9984 36464 10018 36498
rect 10052 36464 10086 36498
rect 10120 36464 10154 36498
rect 10188 36464 10222 36498
rect 10256 36464 10290 36498
rect 10324 36464 10358 36498
rect 10392 36464 10426 36498
rect 10460 36464 10494 36498
rect 10528 36464 10562 36498
rect 10596 36464 10630 36498
rect 10664 36464 10698 36498
rect 10732 36464 10766 36498
rect 10800 36464 10834 36498
rect 10868 36464 10902 36498
rect 10936 36464 10970 36498
rect 11004 36464 11038 36498
rect 11072 36464 11106 36498
rect 11140 36464 11174 36498
rect 11208 36464 11242 36498
rect 11276 36464 11310 36498
rect 11344 36464 11378 36498
rect 11412 36464 11446 36498
rect 11480 36464 11514 36498
rect 11548 36464 11582 36498
rect 11616 36464 11650 36498
rect 11684 36464 11718 36498
rect 11752 36464 11786 36498
rect 11820 36464 11854 36498
rect 11888 36464 11922 36498
rect 11956 36464 11990 36498
rect 12024 36464 12058 36498
rect 12092 36464 12126 36498
rect 12160 36464 12194 36498
rect 12228 36464 12262 36498
rect 12296 36464 12330 36498
rect 12364 36464 12398 36498
rect 12432 36464 12466 36498
rect 12500 36464 12534 36498
rect 12568 36464 12602 36498
rect 12636 36464 12670 36498
rect 12704 36464 12738 36498
rect 12772 36464 12806 36498
rect 12840 36464 12874 36498
rect 12908 36464 12942 36498
rect 12976 36464 13010 36498
rect 13044 36464 13078 36498
rect 13112 36464 13146 36498
rect 13180 36464 13214 36498
rect 13248 36464 13282 36498
rect 13316 36464 13350 36498
rect 13384 36464 13418 36498
rect 13452 36464 13486 36498
rect 13520 36464 13554 36498
rect 13588 36464 13622 36498
rect 13656 36464 13690 36498
rect 13724 36464 13758 36498
rect 13792 36464 13826 36498
rect 13860 36464 13894 36498
rect 13928 36464 13962 36498
rect 13996 36464 14030 36498
rect 14064 36464 14098 36498
rect 14132 36464 14166 36498
rect 14200 36464 14234 36498
rect 14268 36464 14302 36498
rect 14336 36464 14370 36498
rect 14404 36464 14438 36498
rect 14472 36464 14506 36498
rect 317 36277 351 36311
rect 317 36209 351 36243
rect 14611 36275 14645 36309
rect 317 36141 351 36175
rect 317 36073 351 36107
rect 317 36005 351 36039
rect 317 35937 351 35971
rect 317 35869 351 35903
rect 317 35801 351 35835
rect 317 35733 351 35767
rect 317 35665 351 35699
rect 317 35597 351 35631
rect 317 35529 351 35563
rect 317 35461 351 35495
rect 317 35393 351 35427
rect 317 35325 351 35359
rect 317 35257 351 35291
rect 317 35189 351 35223
rect 317 35121 351 35155
rect 317 35053 351 35087
rect 317 34985 351 35019
rect 317 34917 351 34951
rect 317 34849 351 34883
rect 317 34781 351 34815
rect 317 34713 351 34747
rect 317 34645 351 34679
rect 317 34577 351 34611
rect 317 34509 351 34543
rect 317 34441 351 34475
rect 317 34373 351 34407
rect 317 34305 351 34339
rect 317 34237 351 34271
rect 317 34169 351 34203
rect 317 34101 351 34135
rect 317 34033 351 34067
rect 317 33965 351 33999
rect 317 33897 351 33931
rect 317 33829 351 33863
rect 317 33761 351 33795
rect 317 33693 351 33727
rect 317 33625 351 33659
rect 317 33557 351 33591
rect 317 33489 351 33523
rect 317 33421 351 33455
rect 317 33353 351 33387
rect 317 33285 351 33319
rect 317 33217 351 33251
rect 317 33149 351 33183
rect 317 33081 351 33115
rect 317 33013 351 33047
rect 317 32945 351 32979
rect 317 32877 351 32911
rect 317 32809 351 32843
rect 317 32741 351 32775
rect 317 32673 351 32707
rect 317 32605 351 32639
rect 317 32537 351 32571
rect 317 32469 351 32503
rect 317 32401 351 32435
rect 317 32333 351 32367
rect 317 32265 351 32299
rect 317 32197 351 32231
rect 317 32129 351 32163
rect 317 32061 351 32095
rect 317 31993 351 32027
rect 317 31925 351 31959
rect 317 31857 351 31891
rect 317 31789 351 31823
rect 317 31721 351 31755
rect 317 31653 351 31687
rect 317 31585 351 31619
rect 317 31517 351 31551
rect 317 31449 351 31483
rect 317 31381 351 31415
rect 317 31313 351 31347
rect 317 31245 351 31279
rect 317 31177 351 31211
rect 317 31109 351 31143
rect 317 31041 351 31075
rect 317 30973 351 31007
rect 317 30905 351 30939
rect 317 30837 351 30871
rect 317 30769 351 30803
rect 317 30701 351 30735
rect 317 30633 351 30667
rect 317 30565 351 30599
rect 317 30497 351 30531
rect 317 30429 351 30463
rect 317 30361 351 30395
rect 317 30293 351 30327
rect 317 30225 351 30259
rect 317 30157 351 30191
rect 317 30089 351 30123
rect 317 30021 351 30055
rect 317 29953 351 29987
rect 317 29885 351 29919
rect 317 29817 351 29851
rect 317 29749 351 29783
rect 317 29681 351 29715
rect 317 29613 351 29647
rect 317 29545 351 29579
rect 317 29477 351 29511
rect 317 29409 351 29443
rect 317 29341 351 29375
rect 317 29273 351 29307
rect 317 29205 351 29239
rect 317 29137 351 29171
rect 317 29069 351 29103
rect 317 29001 351 29035
rect 317 28933 351 28967
rect 317 28865 351 28899
rect 317 28797 351 28831
rect 317 28729 351 28763
rect 317 28661 351 28695
rect 317 28593 351 28627
rect 317 28525 351 28559
rect 317 28457 351 28491
rect 317 28389 351 28423
rect 317 28321 351 28355
rect 317 28253 351 28287
rect 317 28185 351 28219
rect 317 28117 351 28151
rect 317 28049 351 28083
rect 317 27981 351 28015
rect 317 27913 351 27947
rect 317 27845 351 27879
rect 317 27777 351 27811
rect 317 27709 351 27743
rect 317 27641 351 27675
rect 317 27573 351 27607
rect 317 27505 351 27539
rect 317 27437 351 27471
rect 317 27369 351 27403
rect 317 27301 351 27335
rect 317 27233 351 27267
rect 317 27165 351 27199
rect 317 27097 351 27131
rect 317 27029 351 27063
rect 317 26961 351 26995
rect 317 26893 351 26927
rect 317 26825 351 26859
rect 317 26757 351 26791
rect 317 26689 351 26723
rect 317 26621 351 26655
rect 317 26553 351 26587
rect 317 26485 351 26519
rect 317 26417 351 26451
rect 317 26349 351 26383
rect 317 26281 351 26315
rect 317 26213 351 26247
rect 317 26145 351 26179
rect 317 26077 351 26111
rect 317 26009 351 26043
rect 317 25941 351 25975
rect 317 25873 351 25907
rect 317 25805 351 25839
rect 317 25737 351 25771
rect 317 25669 351 25703
rect 317 25601 351 25635
rect 317 25533 351 25567
rect 317 25465 351 25499
rect 317 25397 351 25431
rect 317 25329 351 25363
rect 317 25261 351 25295
rect 317 25193 351 25227
rect 317 25125 351 25159
rect 317 25057 351 25091
rect 317 24989 351 25023
rect 317 24921 351 24955
rect 317 24853 351 24887
rect 317 24785 351 24819
rect 317 24717 351 24751
rect 317 24649 351 24683
rect 317 24581 351 24615
rect 317 24513 351 24547
rect 317 24445 351 24479
rect 317 24377 351 24411
rect 317 24309 351 24343
rect 317 24241 351 24275
rect 317 24173 351 24207
rect 317 24105 351 24139
rect 317 24037 351 24071
rect 317 23969 351 24003
rect 317 23901 351 23935
rect 317 23833 351 23867
rect 317 23765 351 23799
rect 317 23697 351 23731
rect 317 23629 351 23663
rect 317 23561 351 23595
rect 317 23493 351 23527
rect 317 23425 351 23459
rect 317 23357 351 23391
rect 317 23289 351 23323
rect 317 23221 351 23255
rect 317 23153 351 23187
rect 317 23085 351 23119
rect 317 23017 351 23051
rect 317 22949 351 22983
rect 317 22881 351 22915
rect 317 22813 351 22847
rect 317 22745 351 22779
rect 317 22677 351 22711
rect 317 22609 351 22643
rect 317 22541 351 22575
rect 317 22473 351 22507
rect 317 22405 351 22439
rect 317 22337 351 22371
rect 317 22269 351 22303
rect 317 22201 351 22235
rect 317 22133 351 22167
rect 317 22065 351 22099
rect 317 21997 351 22031
rect 317 21929 351 21963
rect 317 21861 351 21895
rect 317 21793 351 21827
rect 317 21725 351 21759
rect 317 21657 351 21691
rect 317 21589 351 21623
rect 317 21521 351 21555
rect 317 21453 351 21487
rect 317 21385 351 21419
rect 317 21317 351 21351
rect 317 21249 351 21283
rect 317 21181 351 21215
rect 317 21113 351 21147
rect 317 21045 351 21079
rect 317 20977 351 21011
rect 317 20909 351 20943
rect 317 20841 351 20875
rect 317 20773 351 20807
rect 317 20705 351 20739
rect 317 20637 351 20671
rect 317 20569 351 20603
rect 317 20501 351 20535
rect 317 20433 351 20467
rect 317 20365 351 20399
rect 317 20297 351 20331
rect 317 20229 351 20263
rect 317 20161 351 20195
rect 317 20093 351 20127
rect 317 20025 351 20059
rect 317 19957 351 19991
rect 317 19889 351 19923
rect 317 19821 351 19855
rect 317 19753 351 19787
rect 317 19685 351 19719
rect 317 19617 351 19651
rect 317 19549 351 19583
rect 317 19481 351 19515
rect 317 19413 351 19447
rect 317 19345 351 19379
rect 317 19277 351 19311
rect 317 19209 351 19243
rect 317 19141 351 19175
rect 317 19073 351 19107
rect 317 19005 351 19039
rect 317 18937 351 18971
rect 317 18869 351 18903
rect 317 18801 351 18835
rect 317 18733 351 18767
rect 317 18665 351 18699
rect 317 18597 351 18631
rect 317 18529 351 18563
rect 317 18461 351 18495
rect 317 18393 351 18427
rect 317 18325 351 18359
rect 317 18257 351 18291
rect 317 18189 351 18223
rect 317 18121 351 18155
rect 317 18053 351 18087
rect 317 17985 351 18019
rect 317 17917 351 17951
rect 317 17849 351 17883
rect 317 17781 351 17815
rect 317 17713 351 17747
rect 317 17645 351 17679
rect 317 17577 351 17611
rect 317 17509 351 17543
rect 317 17441 351 17475
rect 317 17373 351 17407
rect 317 17305 351 17339
rect 317 17237 351 17271
rect 317 17169 351 17203
rect 317 17101 351 17135
rect 317 17033 351 17067
rect 317 16965 351 16999
rect 317 16897 351 16931
rect 317 16829 351 16863
rect 317 16761 351 16795
rect 317 16693 351 16727
rect 317 16625 351 16659
rect 317 16557 351 16591
rect 317 16489 351 16523
rect 317 16421 351 16455
rect 317 16353 351 16387
rect 317 16285 351 16319
rect 317 16217 351 16251
rect 317 16149 351 16183
rect 317 16081 351 16115
rect 317 16013 351 16047
rect 317 15945 351 15979
rect 317 15877 351 15911
rect 317 15809 351 15843
rect 317 15741 351 15775
rect 317 15673 351 15707
rect 317 15605 351 15639
rect 317 15537 351 15571
rect 317 15469 351 15503
rect 317 15401 351 15435
rect 317 15333 351 15367
rect 317 15265 351 15299
rect 317 15197 351 15231
rect 317 15129 351 15163
rect 317 15061 351 15095
rect 317 14993 351 15027
rect 317 14925 351 14959
rect 317 14857 351 14891
rect 317 14789 351 14823
rect 317 14721 351 14755
rect 317 14653 351 14687
rect 317 14585 351 14619
rect 317 14517 351 14551
rect 317 14449 351 14483
rect 317 14381 351 14415
rect 317 14313 351 14347
rect 317 14245 351 14279
rect 317 14177 351 14211
rect 317 14109 351 14143
rect 317 14041 351 14075
rect 317 13973 351 14007
rect 317 13905 351 13939
rect 317 13837 351 13871
rect 317 13769 351 13803
rect 317 13701 351 13735
rect 317 13633 351 13667
rect 317 13565 351 13599
rect 317 13497 351 13531
rect 317 13429 351 13463
rect 317 13361 351 13395
rect 317 13293 351 13327
rect 317 13225 351 13259
rect 317 13157 351 13191
rect 317 13089 351 13123
rect 317 13021 351 13055
rect 317 12953 351 12987
rect 317 12885 351 12919
rect 317 12817 351 12851
rect 317 12749 351 12783
rect 317 12681 351 12715
rect 317 12613 351 12647
rect 317 12545 351 12579
rect 317 12477 351 12511
rect 317 12409 351 12443
rect 317 12341 351 12375
rect 317 12273 351 12307
rect 317 12205 351 12239
rect 317 12137 351 12171
rect 317 12069 351 12103
rect 317 12001 351 12035
rect 317 11933 351 11967
rect 317 11865 351 11899
rect 317 11797 351 11831
rect 317 11729 351 11763
rect 317 11661 351 11695
rect 317 11593 351 11627
rect 317 11525 351 11559
rect 317 11457 351 11491
rect 317 11389 351 11423
rect 317 11321 351 11355
rect 317 11253 351 11287
rect 317 11185 351 11219
rect 317 11117 351 11151
rect 317 11049 351 11083
rect 317 10981 351 11015
rect 317 10913 351 10947
rect 317 10845 351 10879
rect 317 10777 351 10811
rect 317 10709 351 10743
rect 317 10641 351 10675
rect 317 10573 351 10607
rect 317 10505 351 10539
rect 317 10437 351 10471
rect 317 10369 351 10403
rect 317 10301 351 10335
rect 317 10233 351 10267
rect 317 10165 351 10199
rect 317 10097 351 10131
rect 317 10029 351 10063
rect 317 9961 351 9995
rect 317 9893 351 9927
rect 317 9825 351 9859
rect 317 9757 351 9791
rect 317 9689 351 9723
rect 1327 34616 1361 34650
rect 1395 34616 1429 34650
rect 1463 34616 1497 34650
rect 1531 34616 1565 34650
rect 1599 34616 1633 34650
rect 1667 34616 1701 34650
rect 1735 34616 1769 34650
rect 1803 34616 1837 34650
rect 1871 34616 1905 34650
rect 1939 34616 1973 34650
rect 2007 34616 2041 34650
rect 2075 34616 2109 34650
rect 2143 34616 2177 34650
rect 2211 34616 2245 34650
rect 2279 34616 2313 34650
rect 2347 34616 2381 34650
rect 2415 34616 2449 34650
rect 2483 34616 2517 34650
rect 2551 34616 2585 34650
rect 2619 34616 2653 34650
rect 2687 34616 2721 34650
rect 2755 34616 2789 34650
rect 2823 34616 2857 34650
rect 2891 34616 2925 34650
rect 2959 34616 2993 34650
rect 3027 34616 3061 34650
rect 3095 34616 3129 34650
rect 3163 34616 3197 34650
rect 3231 34616 3265 34650
rect 3299 34616 3333 34650
rect 3367 34616 3401 34650
rect 3435 34616 3469 34650
rect 3503 34616 3537 34650
rect 3571 34616 3605 34650
rect 3639 34616 3673 34650
rect 3707 34616 3741 34650
rect 3775 34616 3809 34650
rect 3843 34616 3877 34650
rect 3911 34616 3945 34650
rect 3979 34616 4013 34650
rect 4047 34616 4081 34650
rect 4115 34616 4149 34650
rect 4183 34616 4217 34650
rect 4251 34616 4285 34650
rect 4319 34616 4353 34650
rect 4387 34616 4421 34650
rect 4455 34616 4489 34650
rect 4523 34616 4557 34650
rect 4591 34616 4625 34650
rect 4659 34616 4693 34650
rect 4727 34616 4761 34650
rect 4795 34616 4829 34650
rect 4863 34616 4897 34650
rect 4931 34616 4965 34650
rect 4999 34616 5033 34650
rect 5067 34616 5101 34650
rect 5135 34616 5169 34650
rect 5203 34616 5237 34650
rect 5271 34616 5305 34650
rect 5339 34616 5373 34650
rect 5407 34616 5441 34650
rect 5475 34616 5509 34650
rect 5543 34616 5577 34650
rect 5611 34616 5645 34650
rect 5679 34616 5713 34650
rect 5747 34616 5781 34650
rect 5815 34616 5849 34650
rect 5883 34616 5917 34650
rect 5951 34616 5985 34650
rect 6019 34616 6053 34650
rect 6087 34616 6121 34650
rect 6155 34616 6189 34650
rect 6223 34616 6257 34650
rect 6291 34616 6325 34650
rect 6359 34616 6393 34650
rect 6427 34616 6461 34650
rect 6495 34616 6529 34650
rect 6563 34616 6597 34650
rect 6631 34616 6665 34650
rect 6699 34616 6733 34650
rect 6767 34616 6801 34650
rect 6835 34616 6869 34650
rect 6903 34616 6937 34650
rect 6971 34616 7005 34650
rect 7039 34616 7073 34650
rect 7107 34616 7141 34650
rect 7175 34616 7209 34650
rect 7243 34616 7277 34650
rect 7311 34616 7345 34650
rect 7379 34616 7413 34650
rect 7447 34616 7481 34650
rect 7515 34616 7549 34650
rect 7583 34616 7617 34650
rect 7651 34616 7685 34650
rect 7719 34616 7753 34650
rect 7787 34616 7821 34650
rect 7855 34616 7889 34650
rect 7923 34616 7957 34650
rect 7991 34616 8025 34650
rect 8059 34616 8093 34650
rect 8127 34616 8161 34650
rect 8195 34616 8229 34650
rect 8263 34616 8297 34650
rect 8331 34616 8365 34650
rect 8399 34616 8433 34650
rect 8467 34616 8501 34650
rect 8535 34616 8569 34650
rect 8603 34616 8637 34650
rect 8671 34616 8705 34650
rect 8739 34616 8773 34650
rect 8807 34616 8841 34650
rect 8875 34616 8909 34650
rect 8943 34616 8977 34650
rect 9011 34616 9045 34650
rect 9079 34616 9113 34650
rect 9147 34616 9181 34650
rect 9215 34616 9249 34650
rect 9283 34616 9317 34650
rect 9351 34616 9385 34650
rect 9419 34616 9453 34650
rect 9487 34616 9521 34650
rect 9555 34616 9589 34650
rect 9623 34616 9657 34650
rect 9691 34616 9725 34650
rect 9759 34616 9793 34650
rect 9827 34616 9861 34650
rect 9895 34616 9929 34650
rect 9963 34616 9997 34650
rect 10031 34616 10065 34650
rect 10099 34616 10133 34650
rect 10167 34616 10201 34650
rect 10235 34616 10269 34650
rect 10303 34616 10337 34650
rect 10371 34616 10405 34650
rect 10439 34616 10473 34650
rect 10507 34616 10541 34650
rect 10575 34616 10609 34650
rect 10643 34616 10677 34650
rect 10711 34616 10745 34650
rect 10779 34616 10813 34650
rect 10847 34616 10881 34650
rect 10915 34616 10949 34650
rect 10983 34616 11017 34650
rect 11051 34616 11085 34650
rect 11119 34616 11153 34650
rect 11187 34616 11221 34650
rect 11255 34616 11289 34650
rect 11323 34616 11357 34650
rect 11391 34616 11425 34650
rect 11459 34616 11493 34650
rect 11527 34616 11561 34650
rect 11595 34616 11629 34650
rect 11663 34616 11697 34650
rect 11731 34616 11765 34650
rect 11799 34616 11833 34650
rect 11867 34616 11901 34650
rect 11935 34616 11969 34650
rect 12003 34616 12037 34650
rect 12071 34616 12105 34650
rect 12139 34616 12173 34650
rect 12207 34616 12241 34650
rect 12275 34616 12309 34650
rect 12343 34616 12377 34650
rect 12411 34616 12445 34650
rect 12479 34616 12513 34650
rect 12547 34616 12581 34650
rect 12615 34616 12649 34650
rect 12683 34616 12717 34650
rect 12751 34616 12785 34650
rect 12819 34616 12853 34650
rect 12887 34616 12921 34650
rect 12955 34616 12989 34650
rect 13023 34616 13057 34650
rect 13091 34616 13125 34650
rect 13159 34616 13193 34650
rect 13227 34616 13261 34650
rect 13295 34616 13329 34650
rect 13363 34616 13397 34650
rect 13431 34616 13465 34650
rect 13499 34616 13533 34650
rect 13567 34616 13601 34650
rect 13635 34616 13669 34650
rect 1192 34487 1226 34521
rect 1192 34419 1226 34453
rect 1192 34351 1226 34385
rect 1192 34283 1226 34317
rect 1192 34215 1226 34249
rect 1192 34147 1226 34181
rect 1192 34079 1226 34113
rect 1192 34011 1226 34045
rect 1192 33943 1226 33977
rect 1192 33875 1226 33909
rect 1192 33807 1226 33841
rect 1192 33739 1226 33773
rect 1192 33671 1226 33705
rect 1192 33603 1226 33637
rect 1192 33535 1226 33569
rect 1192 33467 1226 33501
rect 1192 33399 1226 33433
rect 1192 33331 1226 33365
rect 1192 33263 1226 33297
rect 1192 33195 1226 33229
rect 1192 33127 1226 33161
rect 1192 33059 1226 33093
rect 1192 32991 1226 33025
rect 1192 32923 1226 32957
rect 1192 32855 1226 32889
rect 1192 32787 1226 32821
rect 1192 32719 1226 32753
rect 1192 32651 1226 32685
rect 1192 32583 1226 32617
rect 1192 32515 1226 32549
rect 1192 32447 1226 32481
rect 1192 32379 1226 32413
rect 1192 32311 1226 32345
rect 1192 32243 1226 32277
rect 1192 32175 1226 32209
rect 1192 32107 1226 32141
rect 1192 32039 1226 32073
rect 1192 31971 1226 32005
rect 1192 31903 1226 31937
rect 1192 31835 1226 31869
rect 1192 31767 1226 31801
rect 1192 31699 1226 31733
rect 1192 31631 1226 31665
rect 1192 31563 1226 31597
rect 1192 31495 1226 31529
rect 1192 31427 1226 31461
rect 1192 31359 1226 31393
rect 13768 34500 13802 34534
rect 13768 34432 13802 34466
rect 13768 34364 13802 34398
rect 13768 34296 13802 34330
rect 13768 34228 13802 34262
rect 13768 34160 13802 34194
rect 13768 34092 13802 34126
rect 13768 34024 13802 34058
rect 13768 33956 13802 33990
rect 13768 33888 13802 33922
rect 13768 33820 13802 33854
rect 13768 33752 13802 33786
rect 13768 33684 13802 33718
rect 13768 33616 13802 33650
rect 13768 33548 13802 33582
rect 13768 33480 13802 33514
rect 13768 33412 13802 33446
rect 13768 33344 13802 33378
rect 13768 33276 13802 33310
rect 13768 33208 13802 33242
rect 13768 33140 13802 33174
rect 13768 33072 13802 33106
rect 13768 33004 13802 33038
rect 13768 32936 13802 32970
rect 13768 32868 13802 32902
rect 13768 32800 13802 32834
rect 13768 32732 13802 32766
rect 13768 32664 13802 32698
rect 13768 32596 13802 32630
rect 13768 32528 13802 32562
rect 13768 32460 13802 32494
rect 13768 32392 13802 32426
rect 13768 32324 13802 32358
rect 13768 32256 13802 32290
rect 13768 32188 13802 32222
rect 13768 32120 13802 32154
rect 13768 32052 13802 32086
rect 13768 31984 13802 32018
rect 13768 31916 13802 31950
rect 13768 31848 13802 31882
rect 13768 31780 13802 31814
rect 13768 31712 13802 31746
rect 13768 31644 13802 31678
rect 13768 31576 13802 31610
rect 13768 31508 13802 31542
rect 13768 31440 13802 31474
rect 1192 31291 1226 31325
rect 1192 31223 1226 31257
rect 1192 31155 1226 31189
rect 1192 31087 1226 31121
rect 1192 31019 1226 31053
rect 1192 30951 1226 30985
rect 1192 30883 1226 30917
rect 1192 30815 1226 30849
rect 1192 30747 1226 30781
rect 1192 30679 1226 30713
rect 1192 30611 1226 30645
rect 1192 30543 1226 30577
rect 1192 30475 1226 30509
rect 1192 30407 1226 30441
rect 1192 30339 1226 30373
rect 1192 30271 1226 30305
rect 1192 30203 1226 30237
rect 1192 30135 1226 30169
rect 1192 30067 1226 30101
rect 1192 29999 1226 30033
rect 1192 29931 1226 29965
rect 1192 29863 1226 29897
rect 1192 29795 1226 29829
rect 1192 29727 1226 29761
rect 1192 29659 1226 29693
rect 1192 29591 1226 29625
rect 1192 29523 1226 29557
rect 1192 29455 1226 29489
rect 1192 29387 1226 29421
rect 1192 29319 1226 29353
rect 1192 29251 1226 29285
rect 1192 29183 1226 29217
rect 1192 29115 1226 29149
rect 1192 29047 1226 29081
rect 1192 28979 1226 29013
rect 1192 28911 1226 28945
rect 1192 28843 1226 28877
rect 1192 28775 1226 28809
rect 1192 28707 1226 28741
rect 1192 28639 1226 28673
rect 1192 28571 1226 28605
rect 1192 28503 1226 28537
rect 1192 28435 1226 28469
rect 1192 28367 1226 28401
rect 1192 28299 1226 28333
rect 1192 28231 1226 28265
rect 1192 28163 1226 28197
rect 1192 28095 1226 28129
rect 1192 28027 1226 28061
rect 1192 27959 1226 27993
rect 1192 27891 1226 27925
rect 1192 27823 1226 27857
rect 1192 27755 1226 27789
rect 1192 27687 1226 27721
rect 1192 27619 1226 27653
rect 1192 27551 1226 27585
rect 1192 27483 1226 27517
rect 1192 27415 1226 27449
rect 1192 27347 1226 27381
rect 1192 27279 1226 27313
rect 1192 27211 1226 27245
rect 1192 27143 1226 27177
rect 1192 27075 1226 27109
rect 1192 27007 1226 27041
rect 13768 31372 13802 31406
rect 13768 31304 13802 31338
rect 13768 31236 13802 31270
rect 13768 31168 13802 31202
rect 13768 31100 13802 31134
rect 13768 31032 13802 31066
rect 13768 30964 13802 30998
rect 13768 30896 13802 30930
rect 13768 30828 13802 30862
rect 13768 30760 13802 30794
rect 13768 30692 13802 30726
rect 13768 30624 13802 30658
rect 13768 30556 13802 30590
rect 13768 30488 13802 30522
rect 13768 30420 13802 30454
rect 13768 30352 13802 30386
rect 13768 30284 13802 30318
rect 13768 30216 13802 30250
rect 13768 30148 13802 30182
rect 13768 30080 13802 30114
rect 13768 30012 13802 30046
rect 13768 29944 13802 29978
rect 13768 29876 13802 29910
rect 13768 29808 13802 29842
rect 13768 29740 13802 29774
rect 13768 29672 13802 29706
rect 13768 29604 13802 29638
rect 13768 29536 13802 29570
rect 13768 29468 13802 29502
rect 13768 29400 13802 29434
rect 13768 29332 13802 29366
rect 13768 29264 13802 29298
rect 13768 29196 13802 29230
rect 13768 29128 13802 29162
rect 13768 29060 13802 29094
rect 13768 28992 13802 29026
rect 13768 28924 13802 28958
rect 13768 28856 13802 28890
rect 13768 28788 13802 28822
rect 13768 28720 13802 28754
rect 13768 28652 13802 28686
rect 13768 28584 13802 28618
rect 13768 28516 13802 28550
rect 13768 28448 13802 28482
rect 13768 28380 13802 28414
rect 13768 28312 13802 28346
rect 13768 28244 13802 28278
rect 13768 28176 13802 28210
rect 13768 28108 13802 28142
rect 13768 28040 13802 28074
rect 13768 27972 13802 28006
rect 13768 27904 13802 27938
rect 13768 27836 13802 27870
rect 13768 27768 13802 27802
rect 13768 27700 13802 27734
rect 13768 27632 13802 27666
rect 13768 27564 13802 27598
rect 13768 27496 13802 27530
rect 13768 27428 13802 27462
rect 13768 27360 13802 27394
rect 13768 27292 13802 27326
rect 13768 27224 13802 27258
rect 13768 27156 13802 27190
rect 13768 27088 13802 27122
rect 13768 27020 13802 27054
rect 1192 26939 1226 26973
rect 1192 26871 1226 26905
rect 1192 26803 1226 26837
rect 1192 26735 1226 26769
rect 1192 26667 1226 26701
rect 1192 26599 1226 26633
rect 1192 26531 1226 26565
rect 1192 26463 1226 26497
rect 1192 26395 1226 26429
rect 1192 26327 1226 26361
rect 1192 26259 1226 26293
rect 1192 26191 1226 26225
rect 1192 26123 1226 26157
rect 1192 26055 1226 26089
rect 1192 25987 1226 26021
rect 1192 25919 1226 25953
rect 1192 25851 1226 25885
rect 1192 25783 1226 25817
rect 1192 25715 1226 25749
rect 1192 25647 1226 25681
rect 1192 25579 1226 25613
rect 1192 25511 1226 25545
rect 1192 25443 1226 25477
rect 1192 25375 1226 25409
rect 1192 25307 1226 25341
rect 1192 25239 1226 25273
rect 1192 25171 1226 25205
rect 1192 25103 1226 25137
rect 1192 25035 1226 25069
rect 1192 24967 1226 25001
rect 1192 24899 1226 24933
rect 1192 24831 1226 24865
rect 1192 24763 1226 24797
rect 1192 24695 1226 24729
rect 1192 24627 1226 24661
rect 1192 24559 1226 24593
rect 1192 24491 1226 24525
rect 1192 24423 1226 24457
rect 1192 24355 1226 24389
rect 1192 24287 1226 24321
rect 1192 24219 1226 24253
rect 1192 24151 1226 24185
rect 1192 24083 1226 24117
rect 1192 24015 1226 24049
rect 1192 23947 1226 23981
rect 1192 23879 1226 23913
rect 1192 23811 1226 23845
rect 1192 23743 1226 23777
rect 1192 23675 1226 23709
rect 1192 23607 1226 23641
rect 1192 23539 1226 23573
rect 1192 23471 1226 23505
rect 1192 23403 1226 23437
rect 1192 23335 1226 23369
rect 1192 23267 1226 23301
rect 1192 23199 1226 23233
rect 1192 23131 1226 23165
rect 1192 23063 1226 23097
rect 1192 22995 1226 23029
rect 1192 22927 1226 22961
rect 1192 22859 1226 22893
rect 1192 22791 1226 22825
rect 1192 22723 1226 22757
rect 1192 22655 1226 22689
rect 1192 22587 1226 22621
rect 1192 22519 1226 22553
rect 1192 22451 1226 22485
rect 1192 22383 1226 22417
rect 1192 22315 1226 22349
rect 1192 22247 1226 22281
rect 1192 22179 1226 22213
rect 1192 22111 1226 22145
rect 1192 22043 1226 22077
rect 1192 21975 1226 22009
rect 1192 21907 1226 21941
rect 1192 21839 1226 21873
rect 1192 21771 1226 21805
rect 1192 21703 1226 21737
rect 1192 21635 1226 21669
rect 1192 21567 1226 21601
rect 1192 21499 1226 21533
rect 1192 21431 1226 21465
rect 1192 21363 1226 21397
rect 1192 21295 1226 21329
rect 1192 21227 1226 21261
rect 1192 21159 1226 21193
rect 1192 21091 1226 21125
rect 1192 21023 1226 21057
rect 1192 20955 1226 20989
rect 1192 20887 1226 20921
rect 1192 20819 1226 20853
rect 1192 20751 1226 20785
rect 1192 20683 1226 20717
rect 1192 20615 1226 20649
rect 1192 20547 1226 20581
rect 1192 20479 1226 20513
rect 1192 20411 1226 20445
rect 1192 20343 1226 20377
rect 1192 20275 1226 20309
rect 1192 20207 1226 20241
rect 1192 20139 1226 20173
rect 1192 20071 1226 20105
rect 1192 20003 1226 20037
rect 1192 19935 1226 19969
rect 1192 19867 1226 19901
rect 1192 19799 1226 19833
rect 1192 19731 1226 19765
rect 1192 19663 1226 19697
rect 1192 19595 1226 19629
rect 1192 19527 1226 19561
rect 1192 19459 1226 19493
rect 1192 19391 1226 19425
rect 1192 19323 1226 19357
rect 1192 19255 1226 19289
rect 1192 19187 1226 19221
rect 1192 19119 1226 19153
rect 1192 19051 1226 19085
rect 1192 18983 1226 19017
rect 1192 18915 1226 18949
rect 1192 18847 1226 18881
rect 1192 18779 1226 18813
rect 1192 18711 1226 18745
rect 1192 18643 1226 18677
rect 1192 18575 1226 18609
rect 1192 18507 1226 18541
rect 1192 18439 1226 18473
rect 1192 18371 1226 18405
rect 1192 18303 1226 18337
rect 1192 18235 1226 18269
rect 1192 18167 1226 18201
rect 1192 18099 1226 18133
rect 1192 18031 1226 18065
rect 1192 17963 1226 17997
rect 1192 17895 1226 17929
rect 1192 17827 1226 17861
rect 1192 17759 1226 17793
rect 1192 17691 1226 17725
rect 1192 17623 1226 17657
rect 1192 17555 1226 17589
rect 1192 17487 1226 17521
rect 1192 17419 1226 17453
rect 1192 17351 1226 17385
rect 1192 17283 1226 17317
rect 1192 17215 1226 17249
rect 1192 17147 1226 17181
rect 1192 17079 1226 17113
rect 1192 17011 1226 17045
rect 1192 16943 1226 16977
rect 1192 16875 1226 16909
rect 1192 16807 1226 16841
rect 1192 16739 1226 16773
rect 1192 16671 1226 16705
rect 1192 16603 1226 16637
rect 1192 16535 1226 16569
rect 1192 16467 1226 16501
rect 1192 16399 1226 16433
rect 1192 16331 1226 16365
rect 1192 16263 1226 16297
rect 1192 16195 1226 16229
rect 1192 16127 1226 16161
rect 1192 16059 1226 16093
rect 1192 15991 1226 16025
rect 1192 15923 1226 15957
rect 1192 15855 1226 15889
rect 1192 15787 1226 15821
rect 1192 15719 1226 15753
rect 1192 15651 1226 15685
rect 1192 15583 1226 15617
rect 1192 15515 1226 15549
rect 1192 15447 1226 15481
rect 1192 15379 1226 15413
rect 1192 15311 1226 15345
rect 1192 15243 1226 15277
rect 1192 15175 1226 15209
rect 1192 15107 1226 15141
rect 1192 15039 1226 15073
rect 1192 14971 1226 15005
rect 1192 14903 1226 14937
rect 1192 14835 1226 14869
rect 1192 14767 1226 14801
rect 1192 14699 1226 14733
rect 1192 14631 1226 14665
rect 1192 14563 1226 14597
rect 1192 14495 1226 14529
rect 1192 14427 1226 14461
rect 1192 14359 1226 14393
rect 1192 14291 1226 14325
rect 1192 14223 1226 14257
rect 1192 14155 1226 14189
rect 1192 14087 1226 14121
rect 1192 14019 1226 14053
rect 1192 13951 1226 13985
rect 1192 13883 1226 13917
rect 1192 13815 1226 13849
rect 1192 13747 1226 13781
rect 1192 13679 1226 13713
rect 1192 13611 1226 13645
rect 1192 13543 1226 13577
rect 1192 13475 1226 13509
rect 1192 13407 1226 13441
rect 1192 13339 1226 13373
rect 1192 13271 1226 13305
rect 1192 13203 1226 13237
rect 1192 13135 1226 13169
rect 1192 13067 1226 13101
rect 1192 12999 1226 13033
rect 1192 12931 1226 12965
rect 1192 12863 1226 12897
rect 1192 12795 1226 12829
rect 1192 12727 1226 12761
rect 1192 12659 1226 12693
rect 1192 12591 1226 12625
rect 1192 12523 1226 12557
rect 1192 12455 1226 12489
rect 1192 12387 1226 12421
rect 1192 12319 1226 12353
rect 1192 12251 1226 12285
rect 1192 12183 1226 12217
rect 1192 12115 1226 12149
rect 1192 12047 1226 12081
rect 1192 11979 1226 12013
rect 1192 11911 1226 11945
rect 1192 11843 1226 11877
rect 1192 11775 1226 11809
rect 1192 11707 1226 11741
rect 1192 11639 1226 11673
rect 1192 11571 1226 11605
rect 1192 11503 1226 11537
rect 1192 11435 1226 11469
rect 1192 11367 1226 11401
rect 1192 11299 1226 11333
rect 1192 11231 1226 11265
rect 1192 11163 1226 11197
rect 1192 11095 1226 11129
rect 1192 11027 1226 11061
rect 1192 10959 1226 10993
rect 1192 10891 1226 10925
rect 1192 10823 1226 10857
rect 1192 10755 1226 10789
rect 1192 10687 1226 10721
rect 1192 10619 1226 10653
rect 1192 10551 1226 10585
rect 1192 10483 1226 10517
rect 1192 10415 1226 10449
rect 13768 26952 13802 26986
rect 13768 26884 13802 26918
rect 13768 26816 13802 26850
rect 13768 26748 13802 26782
rect 13768 26680 13802 26714
rect 13768 26612 13802 26646
rect 13768 26544 13802 26578
rect 13768 26476 13802 26510
rect 13768 26408 13802 26442
rect 13768 26340 13802 26374
rect 13768 26272 13802 26306
rect 13768 26204 13802 26238
rect 13768 26136 13802 26170
rect 13768 26068 13802 26102
rect 13768 26000 13802 26034
rect 13768 25932 13802 25966
rect 13768 25864 13802 25898
rect 13768 25796 13802 25830
rect 13768 25728 13802 25762
rect 13768 25660 13802 25694
rect 13768 25592 13802 25626
rect 13768 25524 13802 25558
rect 13768 25456 13802 25490
rect 13768 25388 13802 25422
rect 13768 25320 13802 25354
rect 13768 25252 13802 25286
rect 13768 25184 13802 25218
rect 13768 25116 13802 25150
rect 13768 25048 13802 25082
rect 13768 24980 13802 25014
rect 13768 24912 13802 24946
rect 13768 24844 13802 24878
rect 13768 24776 13802 24810
rect 13768 24708 13802 24742
rect 13768 24640 13802 24674
rect 13768 24572 13802 24606
rect 13768 24504 13802 24538
rect 13768 24436 13802 24470
rect 13768 24368 13802 24402
rect 13768 24300 13802 24334
rect 13768 24232 13802 24266
rect 13768 24164 13802 24198
rect 13768 24096 13802 24130
rect 13768 24028 13802 24062
rect 13768 23960 13802 23994
rect 13768 23892 13802 23926
rect 13768 23824 13802 23858
rect 13768 23756 13802 23790
rect 13768 23688 13802 23722
rect 13768 23620 13802 23654
rect 13768 23552 13802 23586
rect 13768 23484 13802 23518
rect 13768 23416 13802 23450
rect 13768 23348 13802 23382
rect 13768 23280 13802 23314
rect 13768 23212 13802 23246
rect 13768 23144 13802 23178
rect 13768 23076 13802 23110
rect 13768 23008 13802 23042
rect 13768 22940 13802 22974
rect 13768 22872 13802 22906
rect 13768 22804 13802 22838
rect 13768 22736 13802 22770
rect 13768 22668 13802 22702
rect 13768 22600 13802 22634
rect 13768 22532 13802 22566
rect 13768 22464 13802 22498
rect 13768 22396 13802 22430
rect 13768 22328 13802 22362
rect 13768 22260 13802 22294
rect 13768 22192 13802 22226
rect 13768 22124 13802 22158
rect 13768 22056 13802 22090
rect 13768 21988 13802 22022
rect 13768 21920 13802 21954
rect 13768 21852 13802 21886
rect 13768 21784 13802 21818
rect 13768 21716 13802 21750
rect 13768 21648 13802 21682
rect 13768 21580 13802 21614
rect 13768 21512 13802 21546
rect 13768 21444 13802 21478
rect 13768 21376 13802 21410
rect 13768 21308 13802 21342
rect 13768 21240 13802 21274
rect 13768 21172 13802 21206
rect 13768 21104 13802 21138
rect 13768 21036 13802 21070
rect 13768 20968 13802 21002
rect 13768 20900 13802 20934
rect 13768 20832 13802 20866
rect 13768 20764 13802 20798
rect 13768 20696 13802 20730
rect 13768 20628 13802 20662
rect 13768 20560 13802 20594
rect 13768 20492 13802 20526
rect 13768 20424 13802 20458
rect 13768 20356 13802 20390
rect 13768 20288 13802 20322
rect 13768 20220 13802 20254
rect 13768 20152 13802 20186
rect 13768 20084 13802 20118
rect 13768 20016 13802 20050
rect 13768 19948 13802 19982
rect 13768 19880 13802 19914
rect 13768 19812 13802 19846
rect 13768 19744 13802 19778
rect 13768 19676 13802 19710
rect 13768 19608 13802 19642
rect 13768 19540 13802 19574
rect 13768 19472 13802 19506
rect 13768 19404 13802 19438
rect 13768 19336 13802 19370
rect 13768 19268 13802 19302
rect 13768 19200 13802 19234
rect 13768 19132 13802 19166
rect 13768 19064 13802 19098
rect 13768 18996 13802 19030
rect 13768 18928 13802 18962
rect 13768 18860 13802 18894
rect 13768 18792 13802 18826
rect 13768 18724 13802 18758
rect 13768 18656 13802 18690
rect 13768 18588 13802 18622
rect 13768 18520 13802 18554
rect 13768 18452 13802 18486
rect 13768 18384 13802 18418
rect 13768 18316 13802 18350
rect 13768 18248 13802 18282
rect 13768 18180 13802 18214
rect 13768 18112 13802 18146
rect 13768 18044 13802 18078
rect 13768 17976 13802 18010
rect 13768 17908 13802 17942
rect 13768 17840 13802 17874
rect 13768 17772 13802 17806
rect 13768 17704 13802 17738
rect 13768 17636 13802 17670
rect 13768 17568 13802 17602
rect 13768 17500 13802 17534
rect 13768 17432 13802 17466
rect 13768 17364 13802 17398
rect 13768 17296 13802 17330
rect 13768 17228 13802 17262
rect 13768 17160 13802 17194
rect 13768 17092 13802 17126
rect 13768 17024 13802 17058
rect 13768 16956 13802 16990
rect 13768 16888 13802 16922
rect 13768 16820 13802 16854
rect 13768 16752 13802 16786
rect 13768 16684 13802 16718
rect 13768 16616 13802 16650
rect 13768 16548 13802 16582
rect 13768 16480 13802 16514
rect 13768 16412 13802 16446
rect 13768 16344 13802 16378
rect 13768 16276 13802 16310
rect 13768 16208 13802 16242
rect 13768 16140 13802 16174
rect 13768 16072 13802 16106
rect 13768 16004 13802 16038
rect 13768 15936 13802 15970
rect 13768 15868 13802 15902
rect 13768 15800 13802 15834
rect 13768 15732 13802 15766
rect 13768 15664 13802 15698
rect 13768 15596 13802 15630
rect 13768 15528 13802 15562
rect 13768 15460 13802 15494
rect 13768 15392 13802 15426
rect 13768 15324 13802 15358
rect 13768 15256 13802 15290
rect 13768 15188 13802 15222
rect 13768 15120 13802 15154
rect 13768 15052 13802 15086
rect 13768 14984 13802 15018
rect 13768 14916 13802 14950
rect 13768 14848 13802 14882
rect 13768 14780 13802 14814
rect 13768 14712 13802 14746
rect 13768 14644 13802 14678
rect 13768 14576 13802 14610
rect 13768 14508 13802 14542
rect 13768 14440 13802 14474
rect 13768 14372 13802 14406
rect 13768 14304 13802 14338
rect 13768 14236 13802 14270
rect 13768 14168 13802 14202
rect 13768 14100 13802 14134
rect 13768 14032 13802 14066
rect 13768 13964 13802 13998
rect 13768 13896 13802 13930
rect 13768 13828 13802 13862
rect 13768 13760 13802 13794
rect 13768 13692 13802 13726
rect 13768 13624 13802 13658
rect 13768 13556 13802 13590
rect 13768 13488 13802 13522
rect 13768 13420 13802 13454
rect 13768 13352 13802 13386
rect 13768 13284 13802 13318
rect 13768 13216 13802 13250
rect 13768 13148 13802 13182
rect 13768 13080 13802 13114
rect 13768 13012 13802 13046
rect 13768 12944 13802 12978
rect 13768 12876 13802 12910
rect 13768 12808 13802 12842
rect 13768 12740 13802 12774
rect 13768 12672 13802 12706
rect 13768 12604 13802 12638
rect 13768 12536 13802 12570
rect 13768 12468 13802 12502
rect 13768 12400 13802 12434
rect 13768 12332 13802 12366
rect 13768 12264 13802 12298
rect 13768 12196 13802 12230
rect 13768 12128 13802 12162
rect 13768 12060 13802 12094
rect 13768 11992 13802 12026
rect 13768 11924 13802 11958
rect 13768 11856 13802 11890
rect 13768 11788 13802 11822
rect 13768 11720 13802 11754
rect 13768 11652 13802 11686
rect 13768 11584 13802 11618
rect 13768 11516 13802 11550
rect 13768 11448 13802 11482
rect 13768 11380 13802 11414
rect 13768 11312 13802 11346
rect 13768 11244 13802 11278
rect 13768 11176 13802 11210
rect 13768 11108 13802 11142
rect 13768 11040 13802 11074
rect 13768 10972 13802 11006
rect 13768 10904 13802 10938
rect 13768 10836 13802 10870
rect 13768 10768 13802 10802
rect 13768 10700 13802 10734
rect 13768 10632 13802 10666
rect 13768 10564 13802 10598
rect 13768 10496 13802 10530
rect 13768 10428 13802 10462
rect 13768 10360 13802 10394
rect 1329 10284 1363 10318
rect 1397 10284 1431 10318
rect 1465 10284 1499 10318
rect 1533 10284 1567 10318
rect 1601 10284 1635 10318
rect 1669 10284 1703 10318
rect 1737 10284 1771 10318
rect 1805 10284 1839 10318
rect 1873 10284 1907 10318
rect 1941 10284 1975 10318
rect 2009 10284 2043 10318
rect 2077 10284 2111 10318
rect 2145 10284 2179 10318
rect 2213 10284 2247 10318
rect 2281 10284 2315 10318
rect 2349 10284 2383 10318
rect 2417 10284 2451 10318
rect 2485 10284 2519 10318
rect 2553 10284 2587 10318
rect 2621 10284 2655 10318
rect 2689 10284 2723 10318
rect 2757 10284 2791 10318
rect 2825 10284 2859 10318
rect 2893 10284 2927 10318
rect 2961 10284 2995 10318
rect 3029 10284 3063 10318
rect 3097 10284 3131 10318
rect 3165 10284 3199 10318
rect 3233 10284 3267 10318
rect 3301 10284 3335 10318
rect 3369 10284 3403 10318
rect 3437 10284 3471 10318
rect 3505 10284 3539 10318
rect 3573 10284 3607 10318
rect 3641 10284 3675 10318
rect 3709 10284 3743 10318
rect 3777 10284 3811 10318
rect 3845 10284 3879 10318
rect 3913 10284 3947 10318
rect 3981 10284 4015 10318
rect 4049 10284 4083 10318
rect 4117 10284 4151 10318
rect 4185 10284 4219 10318
rect 4253 10284 4287 10318
rect 4321 10284 4355 10318
rect 4389 10284 4423 10318
rect 4457 10284 4491 10318
rect 4525 10284 4559 10318
rect 4593 10284 4627 10318
rect 4661 10284 4695 10318
rect 4729 10284 4763 10318
rect 4797 10284 4831 10318
rect 4865 10284 4899 10318
rect 4933 10284 4967 10318
rect 5001 10284 5035 10318
rect 5069 10284 5103 10318
rect 5137 10284 5171 10318
rect 5205 10284 5239 10318
rect 5273 10284 5307 10318
rect 5341 10284 5375 10318
rect 5409 10284 5443 10318
rect 5477 10284 5511 10318
rect 5545 10284 5579 10318
rect 5613 10284 5647 10318
rect 5681 10284 5715 10318
rect 5749 10284 5783 10318
rect 5817 10284 5851 10318
rect 5885 10284 5919 10318
rect 5953 10284 5987 10318
rect 6021 10284 6055 10318
rect 6089 10284 6123 10318
rect 6157 10284 6191 10318
rect 6225 10284 6259 10318
rect 6293 10284 6327 10318
rect 6361 10284 6395 10318
rect 6429 10284 6463 10318
rect 6497 10284 6531 10318
rect 6565 10284 6599 10318
rect 6633 10284 6667 10318
rect 6701 10284 6735 10318
rect 6769 10284 6803 10318
rect 6837 10284 6871 10318
rect 6905 10284 6939 10318
rect 6973 10284 7007 10318
rect 7041 10284 7075 10318
rect 7109 10284 7143 10318
rect 7177 10284 7211 10318
rect 7245 10284 7279 10318
rect 7313 10284 7347 10318
rect 7381 10284 7415 10318
rect 7449 10284 7483 10318
rect 7517 10284 7551 10318
rect 7585 10284 7619 10318
rect 7653 10284 7687 10318
rect 7721 10284 7755 10318
rect 7789 10284 7823 10318
rect 7857 10284 7891 10318
rect 7925 10284 7959 10318
rect 7993 10284 8027 10318
rect 8061 10284 8095 10318
rect 8129 10284 8163 10318
rect 8197 10284 8231 10318
rect 8265 10284 8299 10318
rect 8333 10284 8367 10318
rect 8401 10284 8435 10318
rect 8469 10284 8503 10318
rect 8537 10284 8571 10318
rect 8605 10284 8639 10318
rect 8673 10284 8707 10318
rect 8741 10284 8775 10318
rect 8809 10284 8843 10318
rect 8877 10284 8911 10318
rect 8945 10284 8979 10318
rect 9013 10284 9047 10318
rect 9081 10284 9115 10318
rect 9149 10284 9183 10318
rect 9217 10284 9251 10318
rect 9285 10284 9319 10318
rect 9353 10284 9387 10318
rect 9421 10284 9455 10318
rect 9489 10284 9523 10318
rect 9557 10284 9591 10318
rect 9625 10284 9659 10318
rect 9693 10284 9727 10318
rect 9761 10284 9795 10318
rect 9829 10284 9863 10318
rect 9897 10284 9931 10318
rect 9965 10284 9999 10318
rect 10033 10284 10067 10318
rect 10101 10284 10135 10318
rect 10169 10284 10203 10318
rect 10237 10284 10271 10318
rect 10305 10284 10339 10318
rect 10373 10284 10407 10318
rect 10441 10284 10475 10318
rect 10509 10284 10543 10318
rect 10577 10284 10611 10318
rect 10645 10284 10679 10318
rect 10713 10284 10747 10318
rect 10781 10284 10815 10318
rect 10849 10284 10883 10318
rect 10917 10284 10951 10318
rect 10985 10284 11019 10318
rect 11053 10284 11087 10318
rect 11121 10284 11155 10318
rect 11189 10284 11223 10318
rect 11257 10284 11291 10318
rect 11325 10284 11359 10318
rect 11393 10284 11427 10318
rect 11461 10284 11495 10318
rect 11529 10284 11563 10318
rect 11597 10284 11631 10318
rect 11665 10284 11699 10318
rect 11733 10284 11767 10318
rect 11801 10284 11835 10318
rect 11869 10284 11903 10318
rect 11937 10284 11971 10318
rect 12005 10284 12039 10318
rect 12073 10284 12107 10318
rect 12141 10284 12175 10318
rect 12209 10284 12243 10318
rect 12277 10284 12311 10318
rect 12345 10284 12379 10318
rect 12413 10284 12447 10318
rect 12481 10284 12515 10318
rect 12549 10284 12583 10318
rect 12617 10284 12651 10318
rect 12685 10284 12719 10318
rect 12753 10284 12787 10318
rect 12821 10284 12855 10318
rect 12889 10284 12923 10318
rect 12957 10284 12991 10318
rect 13025 10284 13059 10318
rect 13093 10284 13127 10318
rect 13161 10284 13195 10318
rect 13229 10284 13263 10318
rect 13297 10284 13331 10318
rect 13365 10284 13399 10318
rect 13433 10284 13467 10318
rect 13501 10284 13535 10318
rect 13569 10284 13603 10318
rect 13637 10284 13671 10318
rect 14611 36207 14645 36241
rect 14611 36139 14645 36173
rect 14611 36071 14645 36105
rect 14611 36003 14645 36037
rect 14611 35935 14645 35969
rect 14611 35867 14645 35901
rect 14611 35799 14645 35833
rect 14611 35731 14645 35765
rect 14611 35663 14645 35697
rect 14611 35595 14645 35629
rect 14611 35527 14645 35561
rect 14611 35459 14645 35493
rect 14611 35391 14645 35425
rect 14611 35323 14645 35357
rect 14611 35255 14645 35289
rect 14611 35187 14645 35221
rect 14611 35119 14645 35153
rect 14611 35051 14645 35085
rect 14611 34983 14645 35017
rect 14611 34915 14645 34949
rect 14611 34847 14645 34881
rect 14611 34779 14645 34813
rect 14611 34711 14645 34745
rect 14611 34643 14645 34677
rect 14611 34575 14645 34609
rect 14611 34507 14645 34541
rect 14611 34439 14645 34473
rect 14611 34371 14645 34405
rect 14611 34303 14645 34337
rect 14611 34235 14645 34269
rect 14611 34167 14645 34201
rect 14611 34099 14645 34133
rect 14611 34031 14645 34065
rect 14611 33963 14645 33997
rect 14611 33895 14645 33929
rect 14611 33827 14645 33861
rect 14611 33759 14645 33793
rect 14611 33691 14645 33725
rect 14611 33623 14645 33657
rect 14611 33555 14645 33589
rect 14611 33487 14645 33521
rect 14611 33419 14645 33453
rect 14611 33351 14645 33385
rect 14611 33283 14645 33317
rect 14611 33215 14645 33249
rect 14611 33147 14645 33181
rect 14611 33079 14645 33113
rect 14611 33011 14645 33045
rect 14611 32943 14645 32977
rect 14611 32875 14645 32909
rect 14611 32807 14645 32841
rect 14611 32739 14645 32773
rect 14611 32671 14645 32705
rect 14611 32603 14645 32637
rect 14611 32535 14645 32569
rect 14611 32467 14645 32501
rect 14611 32399 14645 32433
rect 14611 32331 14645 32365
rect 14611 32263 14645 32297
rect 14611 32195 14645 32229
rect 14611 32127 14645 32161
rect 14611 32059 14645 32093
rect 14611 31991 14645 32025
rect 14611 31923 14645 31957
rect 14611 31855 14645 31889
rect 14611 31787 14645 31821
rect 14611 31719 14645 31753
rect 14611 31651 14645 31685
rect 14611 31583 14645 31617
rect 14611 31515 14645 31549
rect 14611 31447 14645 31481
rect 14611 31379 14645 31413
rect 14611 31311 14645 31345
rect 14611 31243 14645 31277
rect 14611 31175 14645 31209
rect 14611 31107 14645 31141
rect 14611 31039 14645 31073
rect 14611 30971 14645 31005
rect 14611 30903 14645 30937
rect 14611 30835 14645 30869
rect 14611 30767 14645 30801
rect 14611 30699 14645 30733
rect 14611 30631 14645 30665
rect 14611 30563 14645 30597
rect 14611 30495 14645 30529
rect 14611 30427 14645 30461
rect 14611 30359 14645 30393
rect 14611 30291 14645 30325
rect 14611 30223 14645 30257
rect 14611 30155 14645 30189
rect 14611 30087 14645 30121
rect 14611 30019 14645 30053
rect 14611 29951 14645 29985
rect 14611 29883 14645 29917
rect 14611 29815 14645 29849
rect 14611 29747 14645 29781
rect 14611 29679 14645 29713
rect 14611 29611 14645 29645
rect 14611 29543 14645 29577
rect 14611 29475 14645 29509
rect 14611 29407 14645 29441
rect 14611 29339 14645 29373
rect 14611 29271 14645 29305
rect 14611 29203 14645 29237
rect 14611 29135 14645 29169
rect 14611 29067 14645 29101
rect 14611 28999 14645 29033
rect 14611 28931 14645 28965
rect 14611 28863 14645 28897
rect 14611 28795 14645 28829
rect 14611 28727 14645 28761
rect 14611 28659 14645 28693
rect 14611 28591 14645 28625
rect 14611 28523 14645 28557
rect 14611 28455 14645 28489
rect 14611 28387 14645 28421
rect 14611 28319 14645 28353
rect 14611 28251 14645 28285
rect 14611 28183 14645 28217
rect 14611 28115 14645 28149
rect 14611 28047 14645 28081
rect 14611 27979 14645 28013
rect 14611 27911 14645 27945
rect 14611 27843 14645 27877
rect 14611 27775 14645 27809
rect 14611 27707 14645 27741
rect 14611 27639 14645 27673
rect 14611 27571 14645 27605
rect 14611 27503 14645 27537
rect 14611 27435 14645 27469
rect 14611 27367 14645 27401
rect 14611 27299 14645 27333
rect 14611 27231 14645 27265
rect 14611 27163 14645 27197
rect 14611 27095 14645 27129
rect 14611 27027 14645 27061
rect 14611 26959 14645 26993
rect 14611 26891 14645 26925
rect 14611 26823 14645 26857
rect 14611 26755 14645 26789
rect 14611 26687 14645 26721
rect 14611 26619 14645 26653
rect 14611 26551 14645 26585
rect 14611 26483 14645 26517
rect 14611 26415 14645 26449
rect 14611 26347 14645 26381
rect 14611 26279 14645 26313
rect 14611 26211 14645 26245
rect 14611 26143 14645 26177
rect 14611 26075 14645 26109
rect 14611 26007 14645 26041
rect 14611 25939 14645 25973
rect 14611 25871 14645 25905
rect 14611 25803 14645 25837
rect 14611 25735 14645 25769
rect 14611 25667 14645 25701
rect 14611 25599 14645 25633
rect 14611 25531 14645 25565
rect 14611 25463 14645 25497
rect 14611 25395 14645 25429
rect 14611 25327 14645 25361
rect 14611 25259 14645 25293
rect 14611 25191 14645 25225
rect 14611 25123 14645 25157
rect 14611 25055 14645 25089
rect 14611 24987 14645 25021
rect 14611 24919 14645 24953
rect 14611 24851 14645 24885
rect 14611 24783 14645 24817
rect 14611 24715 14645 24749
rect 14611 24647 14645 24681
rect 14611 24579 14645 24613
rect 14611 24511 14645 24545
rect 14611 24443 14645 24477
rect 14611 24375 14645 24409
rect 14611 24307 14645 24341
rect 14611 24239 14645 24273
rect 14611 24171 14645 24205
rect 14611 24103 14645 24137
rect 14611 24035 14645 24069
rect 14611 23967 14645 24001
rect 14611 23899 14645 23933
rect 14611 23831 14645 23865
rect 14611 23763 14645 23797
rect 14611 23695 14645 23729
rect 14611 23627 14645 23661
rect 14611 23559 14645 23593
rect 14611 23491 14645 23525
rect 14611 23423 14645 23457
rect 14611 23355 14645 23389
rect 14611 23287 14645 23321
rect 14611 23219 14645 23253
rect 14611 23151 14645 23185
rect 14611 23083 14645 23117
rect 14611 23015 14645 23049
rect 14611 22947 14645 22981
rect 14611 22879 14645 22913
rect 14611 22811 14645 22845
rect 14611 22743 14645 22777
rect 14611 22675 14645 22709
rect 14611 22607 14645 22641
rect 14611 22539 14645 22573
rect 14611 22471 14645 22505
rect 14611 22403 14645 22437
rect 14611 22335 14645 22369
rect 14611 22267 14645 22301
rect 14611 22199 14645 22233
rect 14611 22131 14645 22165
rect 14611 22063 14645 22097
rect 14611 21995 14645 22029
rect 14611 21927 14645 21961
rect 14611 21859 14645 21893
rect 14611 21791 14645 21825
rect 14611 21723 14645 21757
rect 14611 21655 14645 21689
rect 14611 21587 14645 21621
rect 14611 21519 14645 21553
rect 14611 21451 14645 21485
rect 14611 21383 14645 21417
rect 14611 21315 14645 21349
rect 14611 21247 14645 21281
rect 14611 21179 14645 21213
rect 14611 21111 14645 21145
rect 14611 21043 14645 21077
rect 14611 20975 14645 21009
rect 14611 20907 14645 20941
rect 14611 20839 14645 20873
rect 14611 20771 14645 20805
rect 14611 20703 14645 20737
rect 14611 20635 14645 20669
rect 14611 20567 14645 20601
rect 14611 20499 14645 20533
rect 14611 20431 14645 20465
rect 14611 20363 14645 20397
rect 14611 20295 14645 20329
rect 14611 20227 14645 20261
rect 14611 20159 14645 20193
rect 14611 20091 14645 20125
rect 14611 20023 14645 20057
rect 14611 19955 14645 19989
rect 14611 19887 14645 19921
rect 14611 19819 14645 19853
rect 14611 19751 14645 19785
rect 14611 19683 14645 19717
rect 14611 19615 14645 19649
rect 14611 19547 14645 19581
rect 14611 19479 14645 19513
rect 14611 19411 14645 19445
rect 14611 19343 14645 19377
rect 14611 19275 14645 19309
rect 14611 19207 14645 19241
rect 14611 19139 14645 19173
rect 14611 19071 14645 19105
rect 14611 19003 14645 19037
rect 14611 18935 14645 18969
rect 14611 18867 14645 18901
rect 14611 18799 14645 18833
rect 14611 18731 14645 18765
rect 14611 18663 14645 18697
rect 14611 18595 14645 18629
rect 14611 18527 14645 18561
rect 14611 18459 14645 18493
rect 14611 18391 14645 18425
rect 14611 18323 14645 18357
rect 14611 18255 14645 18289
rect 14611 18187 14645 18221
rect 14611 18119 14645 18153
rect 14611 18051 14645 18085
rect 14611 17983 14645 18017
rect 14611 17915 14645 17949
rect 14611 17847 14645 17881
rect 14611 17779 14645 17813
rect 14611 17711 14645 17745
rect 14611 17643 14645 17677
rect 14611 17575 14645 17609
rect 14611 17507 14645 17541
rect 14611 17439 14645 17473
rect 14611 17371 14645 17405
rect 14611 17303 14645 17337
rect 14611 17235 14645 17269
rect 14611 17167 14645 17201
rect 14611 17099 14645 17133
rect 14611 17031 14645 17065
rect 14611 16963 14645 16997
rect 14611 16895 14645 16929
rect 14611 16827 14645 16861
rect 14611 16759 14645 16793
rect 14611 16691 14645 16725
rect 14611 16623 14645 16657
rect 14611 16555 14645 16589
rect 14611 16487 14645 16521
rect 14611 16419 14645 16453
rect 14611 16351 14645 16385
rect 14611 16283 14645 16317
rect 14611 16215 14645 16249
rect 14611 16147 14645 16181
rect 14611 16079 14645 16113
rect 14611 16011 14645 16045
rect 14611 15943 14645 15977
rect 14611 15875 14645 15909
rect 14611 15807 14645 15841
rect 14611 15739 14645 15773
rect 14611 15671 14645 15705
rect 14611 15603 14645 15637
rect 14611 15535 14645 15569
rect 14611 15467 14645 15501
rect 14611 15399 14645 15433
rect 14611 15331 14645 15365
rect 14611 15263 14645 15297
rect 14611 15195 14645 15229
rect 14611 15127 14645 15161
rect 14611 15059 14645 15093
rect 14611 14991 14645 15025
rect 14611 14923 14645 14957
rect 14611 14855 14645 14889
rect 14611 14787 14645 14821
rect 14611 14719 14645 14753
rect 14611 14651 14645 14685
rect 14611 14583 14645 14617
rect 14611 14515 14645 14549
rect 14611 14447 14645 14481
rect 14611 14379 14645 14413
rect 14611 14311 14645 14345
rect 14611 14243 14645 14277
rect 14611 14175 14645 14209
rect 14611 14107 14645 14141
rect 14611 14039 14645 14073
rect 14611 13971 14645 14005
rect 14611 13903 14645 13937
rect 14611 13835 14645 13869
rect 14611 13767 14645 13801
rect 14611 13699 14645 13733
rect 14611 13631 14645 13665
rect 14611 13563 14645 13597
rect 14611 13495 14645 13529
rect 14611 13427 14645 13461
rect 14611 13359 14645 13393
rect 14611 13291 14645 13325
rect 14611 13223 14645 13257
rect 14611 13155 14645 13189
rect 14611 13087 14645 13121
rect 14611 13019 14645 13053
rect 14611 12951 14645 12985
rect 14611 12883 14645 12917
rect 14611 12815 14645 12849
rect 14611 12747 14645 12781
rect 14611 12679 14645 12713
rect 14611 12611 14645 12645
rect 14611 12543 14645 12577
rect 14611 12475 14645 12509
rect 14611 12407 14645 12441
rect 14611 12339 14645 12373
rect 14611 12271 14645 12305
rect 14611 12203 14645 12237
rect 14611 12135 14645 12169
rect 14611 12067 14645 12101
rect 14611 11999 14645 12033
rect 14611 11931 14645 11965
rect 14611 11863 14645 11897
rect 14611 11795 14645 11829
rect 14611 11727 14645 11761
rect 14611 11659 14645 11693
rect 14611 11591 14645 11625
rect 14611 11523 14645 11557
rect 14611 11455 14645 11489
rect 14611 11387 14645 11421
rect 14611 11319 14645 11353
rect 14611 11251 14645 11285
rect 14611 11183 14645 11217
rect 14611 11115 14645 11149
rect 14611 11047 14645 11081
rect 14611 10979 14645 11013
rect 14611 10911 14645 10945
rect 14611 10843 14645 10877
rect 14611 10775 14645 10809
rect 14611 10707 14645 10741
rect 14611 10639 14645 10673
rect 14611 10571 14645 10605
rect 14611 10503 14645 10537
rect 14611 10435 14645 10469
rect 14611 10367 14645 10401
rect 14611 10299 14645 10333
rect 14611 10231 14645 10265
rect 14611 10163 14645 10197
rect 14611 10095 14645 10129
rect 14611 10027 14645 10061
rect 14611 9959 14645 9993
rect 14611 9891 14645 9925
rect 14611 9823 14645 9857
rect 14611 9755 14645 9789
rect 317 9621 351 9655
rect 14611 9687 14645 9721
rect 14611 9619 14645 9653
rect 506 9416 540 9450
rect 574 9416 608 9450
rect 642 9416 676 9450
rect 710 9416 744 9450
rect 778 9416 812 9450
rect 846 9416 880 9450
rect 914 9416 948 9450
rect 982 9416 1016 9450
rect 1050 9416 1084 9450
rect 1118 9416 1152 9450
rect 1186 9416 1220 9450
rect 1254 9416 1288 9450
rect 1322 9416 1356 9450
rect 1390 9416 1424 9450
rect 1458 9416 1492 9450
rect 1526 9416 1560 9450
rect 1594 9416 1628 9450
rect 1662 9416 1696 9450
rect 1730 9416 1764 9450
rect 1798 9416 1832 9450
rect 1866 9416 1900 9450
rect 1934 9416 1968 9450
rect 2002 9416 2036 9450
rect 2070 9416 2104 9450
rect 2138 9416 2172 9450
rect 2206 9416 2240 9450
rect 2274 9416 2308 9450
rect 2342 9416 2376 9450
rect 2410 9416 2444 9450
rect 2478 9416 2512 9450
rect 2546 9416 2580 9450
rect 2614 9416 2648 9450
rect 2682 9416 2716 9450
rect 2750 9416 2784 9450
rect 2818 9416 2852 9450
rect 2886 9416 2920 9450
rect 2954 9416 2988 9450
rect 3022 9416 3056 9450
rect 3090 9416 3124 9450
rect 3158 9416 3192 9450
rect 3226 9416 3260 9450
rect 3294 9416 3328 9450
rect 3362 9416 3396 9450
rect 3430 9416 3464 9450
rect 3498 9416 3532 9450
rect 3566 9416 3600 9450
rect 3634 9416 3668 9450
rect 3702 9416 3736 9450
rect 3770 9416 3804 9450
rect 3838 9416 3872 9450
rect 3906 9416 3940 9450
rect 3974 9416 4008 9450
rect 4042 9416 4076 9450
rect 4110 9416 4144 9450
rect 4178 9416 4212 9450
rect 4246 9416 4280 9450
rect 4314 9416 4348 9450
rect 4382 9416 4416 9450
rect 4450 9416 4484 9450
rect 4518 9416 4552 9450
rect 4586 9416 4620 9450
rect 4654 9416 4688 9450
rect 4722 9416 4756 9450
rect 4790 9416 4824 9450
rect 4858 9416 4892 9450
rect 4926 9416 4960 9450
rect 4994 9416 5028 9450
rect 5062 9416 5096 9450
rect 5130 9416 5164 9450
rect 5198 9416 5232 9450
rect 5266 9416 5300 9450
rect 5334 9416 5368 9450
rect 5402 9416 5436 9450
rect 5470 9416 5504 9450
rect 5538 9416 5572 9450
rect 5606 9416 5640 9450
rect 5674 9416 5708 9450
rect 5742 9416 5776 9450
rect 5810 9416 5844 9450
rect 5878 9416 5912 9450
rect 5946 9416 5980 9450
rect 6014 9416 6048 9450
rect 6082 9416 6116 9450
rect 6150 9416 6184 9450
rect 6218 9416 6252 9450
rect 6286 9416 6320 9450
rect 6354 9416 6388 9450
rect 6422 9416 6456 9450
rect 6490 9416 6524 9450
rect 6558 9416 6592 9450
rect 6626 9416 6660 9450
rect 6694 9416 6728 9450
rect 6762 9416 6796 9450
rect 6830 9416 6864 9450
rect 6898 9416 6932 9450
rect 6966 9416 7000 9450
rect 7034 9416 7068 9450
rect 7102 9416 7136 9450
rect 7170 9416 7204 9450
rect 7238 9416 7272 9450
rect 7306 9416 7340 9450
rect 7374 9416 7408 9450
rect 7442 9416 7476 9450
rect 7510 9416 7544 9450
rect 7578 9416 7612 9450
rect 7646 9416 7680 9450
rect 7714 9416 7748 9450
rect 7782 9416 7816 9450
rect 7850 9416 7884 9450
rect 7918 9416 7952 9450
rect 7986 9416 8020 9450
rect 8054 9416 8088 9450
rect 8122 9416 8156 9450
rect 8190 9416 8224 9450
rect 8258 9416 8292 9450
rect 8326 9416 8360 9450
rect 8394 9416 8428 9450
rect 8462 9416 8496 9450
rect 8530 9416 8564 9450
rect 8598 9416 8632 9450
rect 8666 9416 8700 9450
rect 8734 9416 8768 9450
rect 8802 9416 8836 9450
rect 8870 9416 8904 9450
rect 8938 9416 8972 9450
rect 9006 9416 9040 9450
rect 9074 9416 9108 9450
rect 9142 9416 9176 9450
rect 9210 9416 9244 9450
rect 9278 9416 9312 9450
rect 9346 9416 9380 9450
rect 9414 9416 9448 9450
rect 9482 9416 9516 9450
rect 9550 9416 9584 9450
rect 9618 9416 9652 9450
rect 9686 9416 9720 9450
rect 9754 9416 9788 9450
rect 9822 9416 9856 9450
rect 9890 9416 9924 9450
rect 9958 9416 9992 9450
rect 10026 9416 10060 9450
rect 10094 9416 10128 9450
rect 10162 9416 10196 9450
rect 10230 9416 10264 9450
rect 10298 9416 10332 9450
rect 10366 9416 10400 9450
rect 10434 9416 10468 9450
rect 10502 9416 10536 9450
rect 10570 9416 10604 9450
rect 10638 9416 10672 9450
rect 10706 9416 10740 9450
rect 10774 9416 10808 9450
rect 10842 9416 10876 9450
rect 10910 9416 10944 9450
rect 10978 9416 11012 9450
rect 11046 9416 11080 9450
rect 11114 9416 11148 9450
rect 11182 9416 11216 9450
rect 11250 9416 11284 9450
rect 11318 9416 11352 9450
rect 11386 9416 11420 9450
rect 11454 9416 11488 9450
rect 11522 9416 11556 9450
rect 11590 9416 11624 9450
rect 11658 9416 11692 9450
rect 11726 9416 11760 9450
rect 11794 9416 11828 9450
rect 11862 9416 11896 9450
rect 11930 9416 11964 9450
rect 11998 9416 12032 9450
rect 12066 9416 12100 9450
rect 12134 9416 12168 9450
rect 12202 9416 12236 9450
rect 12270 9416 12304 9450
rect 12338 9416 12372 9450
rect 12406 9416 12440 9450
rect 12474 9416 12508 9450
rect 12542 9416 12576 9450
rect 12610 9416 12644 9450
rect 12678 9416 12712 9450
rect 12746 9416 12780 9450
rect 12814 9416 12848 9450
rect 12882 9416 12916 9450
rect 12950 9416 12984 9450
rect 13018 9416 13052 9450
rect 13086 9416 13120 9450
rect 13154 9416 13188 9450
rect 13222 9416 13256 9450
rect 13290 9416 13324 9450
rect 13358 9416 13392 9450
rect 13426 9416 13460 9450
rect 13494 9416 13528 9450
rect 13562 9416 13596 9450
rect 13630 9416 13664 9450
rect 13698 9416 13732 9450
rect 13766 9416 13800 9450
rect 13834 9416 13868 9450
rect 13902 9416 13936 9450
rect 13970 9416 14004 9450
rect 14038 9416 14072 9450
rect 14106 9416 14140 9450
rect 14174 9416 14208 9450
rect 14242 9416 14276 9450
rect 14310 9416 14344 9450
rect 14378 9416 14412 9450
rect 14446 9416 14480 9450
<< mvnsubdiffcont >>
rect 766 36143 800 36177
rect 834 36143 868 36177
rect 902 36143 936 36177
rect 970 36143 1004 36177
rect 1038 36143 1072 36177
rect 1106 36143 1140 36177
rect 1174 36143 1208 36177
rect 1242 36143 1276 36177
rect 1310 36143 1344 36177
rect 1378 36143 1412 36177
rect 1446 36143 1480 36177
rect 1514 36143 1548 36177
rect 1582 36143 1616 36177
rect 1650 36143 1684 36177
rect 1718 36143 1752 36177
rect 1786 36143 1820 36177
rect 1854 36143 1888 36177
rect 1922 36143 1956 36177
rect 1990 36143 2024 36177
rect 2058 36143 2092 36177
rect 2126 36143 2160 36177
rect 2194 36143 2228 36177
rect 2262 36143 2296 36177
rect 2330 36143 2364 36177
rect 2398 36143 2432 36177
rect 2466 36143 2500 36177
rect 2534 36143 2568 36177
rect 2602 36143 2636 36177
rect 2670 36143 2704 36177
rect 2738 36143 2772 36177
rect 2806 36143 2840 36177
rect 2874 36143 2908 36177
rect 2942 36143 2976 36177
rect 3010 36143 3044 36177
rect 3078 36143 3112 36177
rect 3146 36143 3180 36177
rect 3214 36143 3248 36177
rect 3282 36143 3316 36177
rect 3350 36143 3384 36177
rect 3418 36143 3452 36177
rect 3486 36143 3520 36177
rect 3554 36143 3588 36177
rect 3622 36143 3656 36177
rect 3690 36143 3724 36177
rect 3758 36143 3792 36177
rect 3826 36143 3860 36177
rect 3894 36143 3928 36177
rect 3962 36143 3996 36177
rect 4030 36143 4064 36177
rect 4098 36143 4132 36177
rect 4166 36143 4200 36177
rect 4234 36143 4268 36177
rect 4302 36143 4336 36177
rect 4370 36143 4404 36177
rect 4438 36143 4472 36177
rect 4506 36143 4540 36177
rect 4574 36143 4608 36177
rect 4642 36143 4676 36177
rect 4710 36143 4744 36177
rect 4778 36143 4812 36177
rect 4846 36143 4880 36177
rect 4914 36143 4948 36177
rect 4982 36143 5016 36177
rect 5050 36143 5084 36177
rect 5118 36143 5152 36177
rect 5186 36143 5220 36177
rect 5254 36143 5288 36177
rect 5322 36143 5356 36177
rect 5390 36143 5424 36177
rect 5458 36143 5492 36177
rect 5526 36143 5560 36177
rect 5594 36143 5628 36177
rect 5662 36143 5696 36177
rect 5730 36143 5764 36177
rect 5798 36143 5832 36177
rect 5866 36143 5900 36177
rect 5934 36143 5968 36177
rect 6002 36143 6036 36177
rect 6070 36143 6104 36177
rect 6138 36143 6172 36177
rect 6206 36143 6240 36177
rect 6274 36143 6308 36177
rect 6342 36143 6376 36177
rect 6410 36143 6444 36177
rect 6478 36143 6512 36177
rect 6546 36143 6580 36177
rect 6614 36143 6648 36177
rect 6682 36143 6716 36177
rect 6750 36143 6784 36177
rect 6818 36143 6852 36177
rect 6886 36143 6920 36177
rect 6954 36143 6988 36177
rect 7022 36143 7056 36177
rect 7090 36143 7124 36177
rect 7158 36143 7192 36177
rect 7226 36143 7260 36177
rect 7294 36143 7328 36177
rect 7362 36143 7396 36177
rect 7430 36143 7464 36177
rect 7498 36143 7532 36177
rect 7566 36143 7600 36177
rect 7634 36143 7668 36177
rect 7702 36143 7736 36177
rect 7770 36143 7804 36177
rect 7838 36143 7872 36177
rect 7906 36143 7940 36177
rect 7974 36143 8008 36177
rect 8042 36143 8076 36177
rect 8110 36143 8144 36177
rect 8178 36143 8212 36177
rect 8246 36143 8280 36177
rect 8314 36143 8348 36177
rect 8382 36143 8416 36177
rect 8450 36143 8484 36177
rect 8518 36143 8552 36177
rect 8586 36143 8620 36177
rect 8654 36143 8688 36177
rect 8722 36143 8756 36177
rect 8790 36143 8824 36177
rect 8858 36143 8892 36177
rect 8926 36143 8960 36177
rect 8994 36143 9028 36177
rect 9062 36143 9096 36177
rect 9130 36143 9164 36177
rect 9198 36143 9232 36177
rect 9266 36143 9300 36177
rect 9334 36143 9368 36177
rect 9402 36143 9436 36177
rect 9470 36143 9504 36177
rect 9538 36143 9572 36177
rect 9606 36143 9640 36177
rect 9674 36143 9708 36177
rect 9742 36143 9776 36177
rect 9810 36143 9844 36177
rect 9878 36143 9912 36177
rect 9946 36143 9980 36177
rect 10014 36143 10048 36177
rect 10082 36143 10116 36177
rect 10150 36143 10184 36177
rect 10218 36143 10252 36177
rect 10286 36143 10320 36177
rect 10354 36143 10388 36177
rect 10422 36143 10456 36177
rect 10490 36143 10524 36177
rect 10558 36143 10592 36177
rect 10626 36143 10660 36177
rect 10694 36143 10728 36177
rect 10762 36143 10796 36177
rect 10830 36143 10864 36177
rect 10898 36143 10932 36177
rect 10966 36143 11000 36177
rect 11034 36143 11068 36177
rect 11102 36143 11136 36177
rect 11170 36143 11204 36177
rect 11238 36143 11272 36177
rect 11306 36143 11340 36177
rect 11374 36143 11408 36177
rect 11442 36143 11476 36177
rect 11510 36143 11544 36177
rect 11578 36143 11612 36177
rect 11646 36143 11680 36177
rect 11714 36143 11748 36177
rect 11782 36143 11816 36177
rect 11850 36143 11884 36177
rect 11918 36143 11952 36177
rect 11986 36143 12020 36177
rect 12054 36143 12088 36177
rect 12122 36143 12156 36177
rect 12190 36143 12224 36177
rect 12258 36143 12292 36177
rect 12326 36143 12360 36177
rect 12394 36143 12428 36177
rect 12462 36143 12496 36177
rect 12530 36143 12564 36177
rect 12598 36143 12632 36177
rect 12666 36143 12700 36177
rect 12734 36143 12768 36177
rect 12802 36143 12836 36177
rect 12870 36143 12904 36177
rect 12938 36143 12972 36177
rect 13006 36143 13040 36177
rect 13074 36143 13108 36177
rect 13142 36143 13176 36177
rect 13210 36143 13244 36177
rect 13278 36143 13312 36177
rect 13346 36143 13380 36177
rect 13414 36143 13448 36177
rect 13482 36143 13516 36177
rect 13550 36143 13584 36177
rect 13618 36143 13652 36177
rect 13686 36143 13720 36177
rect 13754 36143 13788 36177
rect 13822 36143 13856 36177
rect 13890 36143 13924 36177
rect 13958 36143 13992 36177
rect 14026 36143 14060 36177
rect 14094 36143 14128 36177
rect 14162 36143 14196 36177
rect 632 35998 666 36032
rect 632 35930 666 35964
rect 632 35862 666 35896
rect 632 35794 666 35828
rect 632 35726 666 35760
rect 632 35658 666 35692
rect 632 35590 666 35624
rect 632 35522 666 35556
rect 632 35454 666 35488
rect 632 35386 666 35420
rect 632 35318 666 35352
rect 632 35250 666 35284
rect 632 35182 666 35216
rect 632 35114 666 35148
rect 632 35046 666 35080
rect 632 34978 666 35012
rect 632 34910 666 34944
rect 632 34842 666 34876
rect 632 34774 666 34808
rect 632 34706 666 34740
rect 14297 35998 14331 36032
rect 14297 35930 14331 35964
rect 14297 35862 14331 35896
rect 14297 35794 14331 35828
rect 14297 35726 14331 35760
rect 14297 35658 14331 35692
rect 14297 35590 14331 35624
rect 14297 35522 14331 35556
rect 14297 35454 14331 35488
rect 14297 35386 14331 35420
rect 14297 35318 14331 35352
rect 14297 35250 14331 35284
rect 14297 35182 14331 35216
rect 14297 35114 14331 35148
rect 14297 35046 14331 35080
rect 14297 34978 14331 35012
rect 14297 34910 14331 34944
rect 14297 34842 14331 34876
rect 14297 34774 14331 34808
rect 14297 34706 14331 34740
rect 632 34638 666 34672
rect 632 34570 666 34604
rect 632 34502 666 34536
rect 632 34434 666 34468
rect 632 34366 666 34400
rect 632 34298 666 34332
rect 632 34230 666 34264
rect 632 34162 666 34196
rect 632 34094 666 34128
rect 632 34026 666 34060
rect 632 33958 666 33992
rect 632 33890 666 33924
rect 632 33822 666 33856
rect 632 33754 666 33788
rect 632 33686 666 33720
rect 632 33618 666 33652
rect 632 33550 666 33584
rect 632 33482 666 33516
rect 632 33414 666 33448
rect 632 33346 666 33380
rect 632 33278 666 33312
rect 632 33210 666 33244
rect 632 33142 666 33176
rect 632 33074 666 33108
rect 632 33006 666 33040
rect 632 32938 666 32972
rect 632 32870 666 32904
rect 632 32802 666 32836
rect 632 32734 666 32768
rect 632 32666 666 32700
rect 632 32598 666 32632
rect 632 32530 666 32564
rect 632 32462 666 32496
rect 632 32394 666 32428
rect 632 32326 666 32360
rect 632 32258 666 32292
rect 632 32190 666 32224
rect 632 32122 666 32156
rect 632 32054 666 32088
rect 632 31986 666 32020
rect 632 31918 666 31952
rect 632 31850 666 31884
rect 632 31782 666 31816
rect 632 31714 666 31748
rect 632 31646 666 31680
rect 632 31578 666 31612
rect 632 31510 666 31544
rect 632 31442 666 31476
rect 632 31374 666 31408
rect 632 31306 666 31340
rect 632 31238 666 31272
rect 632 31170 666 31204
rect 632 31102 666 31136
rect 632 31034 666 31068
rect 632 30966 666 31000
rect 632 30898 666 30932
rect 632 30830 666 30864
rect 632 30762 666 30796
rect 632 30694 666 30728
rect 632 30626 666 30660
rect 632 30558 666 30592
rect 632 30490 666 30524
rect 632 30422 666 30456
rect 632 30354 666 30388
rect 632 30286 666 30320
rect 632 30218 666 30252
rect 632 30150 666 30184
rect 632 30082 666 30116
rect 632 30014 666 30048
rect 632 29946 666 29980
rect 632 29878 666 29912
rect 632 29810 666 29844
rect 632 29742 666 29776
rect 632 29674 666 29708
rect 632 29606 666 29640
rect 632 29538 666 29572
rect 632 29470 666 29504
rect 632 29402 666 29436
rect 632 29334 666 29368
rect 632 29266 666 29300
rect 632 29198 666 29232
rect 632 29130 666 29164
rect 632 29062 666 29096
rect 632 28994 666 29028
rect 632 28926 666 28960
rect 632 28858 666 28892
rect 632 28790 666 28824
rect 632 28722 666 28756
rect 632 28654 666 28688
rect 632 28586 666 28620
rect 632 28518 666 28552
rect 632 28450 666 28484
rect 632 28382 666 28416
rect 632 28314 666 28348
rect 632 28246 666 28280
rect 632 28178 666 28212
rect 632 28110 666 28144
rect 632 28042 666 28076
rect 632 27974 666 28008
rect 632 27906 666 27940
rect 632 27838 666 27872
rect 632 27770 666 27804
rect 632 27702 666 27736
rect 632 27634 666 27668
rect 632 27566 666 27600
rect 632 27498 666 27532
rect 632 27430 666 27464
rect 632 27362 666 27396
rect 632 27294 666 27328
rect 632 27226 666 27260
rect 632 27158 666 27192
rect 632 27090 666 27124
rect 632 27022 666 27056
rect 632 26954 666 26988
rect 632 26886 666 26920
rect 632 26818 666 26852
rect 632 26750 666 26784
rect 632 26682 666 26716
rect 632 26614 666 26648
rect 632 26546 666 26580
rect 632 26478 666 26512
rect 632 26410 666 26444
rect 632 26342 666 26376
rect 632 26274 666 26308
rect 632 26206 666 26240
rect 632 26138 666 26172
rect 632 26070 666 26104
rect 632 26002 666 26036
rect 632 25934 666 25968
rect 632 25866 666 25900
rect 632 25798 666 25832
rect 632 25730 666 25764
rect 632 25662 666 25696
rect 632 25594 666 25628
rect 632 25526 666 25560
rect 632 25458 666 25492
rect 632 25390 666 25424
rect 632 25322 666 25356
rect 632 25254 666 25288
rect 632 25186 666 25220
rect 632 25118 666 25152
rect 632 25050 666 25084
rect 632 24982 666 25016
rect 632 24914 666 24948
rect 632 24846 666 24880
rect 632 24778 666 24812
rect 632 24710 666 24744
rect 632 24642 666 24676
rect 632 24574 666 24608
rect 632 24506 666 24540
rect 632 24438 666 24472
rect 632 24370 666 24404
rect 632 24302 666 24336
rect 632 24234 666 24268
rect 632 24166 666 24200
rect 632 24098 666 24132
rect 632 24030 666 24064
rect 632 23962 666 23996
rect 632 23894 666 23928
rect 632 23826 666 23860
rect 632 23758 666 23792
rect 632 23690 666 23724
rect 632 23622 666 23656
rect 632 23554 666 23588
rect 632 23486 666 23520
rect 632 23418 666 23452
rect 632 23350 666 23384
rect 632 23282 666 23316
rect 632 23214 666 23248
rect 632 23146 666 23180
rect 632 23078 666 23112
rect 632 23010 666 23044
rect 632 22942 666 22976
rect 632 22874 666 22908
rect 632 22806 666 22840
rect 632 22738 666 22772
rect 632 22670 666 22704
rect 632 22602 666 22636
rect 632 22534 666 22568
rect 632 22466 666 22500
rect 632 22398 666 22432
rect 632 22330 666 22364
rect 632 22262 666 22296
rect 632 22194 666 22228
rect 632 22126 666 22160
rect 632 22058 666 22092
rect 632 21990 666 22024
rect 632 21922 666 21956
rect 632 21854 666 21888
rect 632 21786 666 21820
rect 632 21718 666 21752
rect 632 21650 666 21684
rect 632 21582 666 21616
rect 632 21514 666 21548
rect 632 21446 666 21480
rect 632 21378 666 21412
rect 632 21310 666 21344
rect 632 21242 666 21276
rect 632 21174 666 21208
rect 632 21106 666 21140
rect 632 21038 666 21072
rect 632 20970 666 21004
rect 632 20902 666 20936
rect 632 20834 666 20868
rect 632 20766 666 20800
rect 632 20698 666 20732
rect 632 20630 666 20664
rect 632 20562 666 20596
rect 632 20494 666 20528
rect 632 20426 666 20460
rect 632 20358 666 20392
rect 632 20290 666 20324
rect 632 20222 666 20256
rect 632 20154 666 20188
rect 632 20086 666 20120
rect 632 20018 666 20052
rect 632 19950 666 19984
rect 632 19882 666 19916
rect 632 19814 666 19848
rect 632 19746 666 19780
rect 632 19678 666 19712
rect 632 19610 666 19644
rect 632 19542 666 19576
rect 632 19474 666 19508
rect 632 19406 666 19440
rect 632 19338 666 19372
rect 632 19270 666 19304
rect 632 19202 666 19236
rect 632 19134 666 19168
rect 632 19066 666 19100
rect 632 18998 666 19032
rect 632 18930 666 18964
rect 632 18862 666 18896
rect 632 18794 666 18828
rect 632 18726 666 18760
rect 632 18658 666 18692
rect 632 18590 666 18624
rect 632 18522 666 18556
rect 632 18454 666 18488
rect 632 18386 666 18420
rect 632 18318 666 18352
rect 632 18250 666 18284
rect 632 18182 666 18216
rect 632 18114 666 18148
rect 632 18046 666 18080
rect 632 17978 666 18012
rect 632 17910 666 17944
rect 632 17842 666 17876
rect 632 17774 666 17808
rect 632 17706 666 17740
rect 632 17638 666 17672
rect 632 17570 666 17604
rect 632 17502 666 17536
rect 632 17434 666 17468
rect 632 17366 666 17400
rect 632 17298 666 17332
rect 632 17230 666 17264
rect 632 17162 666 17196
rect 632 17094 666 17128
rect 632 17026 666 17060
rect 632 16958 666 16992
rect 632 16890 666 16924
rect 632 16822 666 16856
rect 632 16754 666 16788
rect 632 16686 666 16720
rect 632 16618 666 16652
rect 632 16550 666 16584
rect 632 16482 666 16516
rect 632 16414 666 16448
rect 632 16346 666 16380
rect 632 16278 666 16312
rect 632 16210 666 16244
rect 632 16142 666 16176
rect 632 16074 666 16108
rect 632 16006 666 16040
rect 632 15938 666 15972
rect 632 15870 666 15904
rect 632 15802 666 15836
rect 632 15734 666 15768
rect 632 15666 666 15700
rect 632 15598 666 15632
rect 632 15530 666 15564
rect 632 15462 666 15496
rect 632 15394 666 15428
rect 632 15326 666 15360
rect 632 15258 666 15292
rect 632 15190 666 15224
rect 632 15122 666 15156
rect 632 15054 666 15088
rect 632 14986 666 15020
rect 632 14918 666 14952
rect 632 14850 666 14884
rect 632 14782 666 14816
rect 632 14714 666 14748
rect 632 14646 666 14680
rect 632 14578 666 14612
rect 632 14510 666 14544
rect 632 14442 666 14476
rect 632 14374 666 14408
rect 632 14306 666 14340
rect 632 14238 666 14272
rect 632 14170 666 14204
rect 632 14102 666 14136
rect 632 14034 666 14068
rect 632 13966 666 14000
rect 632 13898 666 13932
rect 632 13830 666 13864
rect 632 13762 666 13796
rect 632 13694 666 13728
rect 632 13626 666 13660
rect 632 13558 666 13592
rect 632 13490 666 13524
rect 632 13422 666 13456
rect 632 13354 666 13388
rect 632 13286 666 13320
rect 632 13218 666 13252
rect 632 13150 666 13184
rect 632 13082 666 13116
rect 632 13014 666 13048
rect 632 12946 666 12980
rect 632 12878 666 12912
rect 632 12810 666 12844
rect 632 12742 666 12776
rect 632 12674 666 12708
rect 632 12606 666 12640
rect 632 12538 666 12572
rect 632 12470 666 12504
rect 632 12402 666 12436
rect 632 12334 666 12368
rect 632 12266 666 12300
rect 632 12198 666 12232
rect 632 12130 666 12164
rect 632 12062 666 12096
rect 632 11994 666 12028
rect 632 11926 666 11960
rect 632 11858 666 11892
rect 632 11790 666 11824
rect 632 11722 666 11756
rect 632 11654 666 11688
rect 632 11586 666 11620
rect 632 11518 666 11552
rect 632 11450 666 11484
rect 632 11382 666 11416
rect 632 11314 666 11348
rect 632 11246 666 11280
rect 632 11178 666 11212
rect 632 11110 666 11144
rect 632 11042 666 11076
rect 632 10974 666 11008
rect 632 10906 666 10940
rect 632 10838 666 10872
rect 632 10770 666 10804
rect 632 10702 666 10736
rect 632 10634 666 10668
rect 632 10566 666 10600
rect 632 10498 666 10532
rect 632 10430 666 10464
rect 632 10362 666 10396
rect 632 10294 666 10328
rect 632 10226 666 10260
rect 2119 30975 12897 31349
rect 1689 27481 2063 30915
rect 12953 27481 13327 30915
rect 2119 27047 12897 27421
rect 14297 34638 14331 34672
rect 14297 34570 14331 34604
rect 14297 34502 14331 34536
rect 14297 34434 14331 34468
rect 14297 34366 14331 34400
rect 14297 34298 14331 34332
rect 14297 34230 14331 34264
rect 14297 34162 14331 34196
rect 14297 34094 14331 34128
rect 14297 34026 14331 34060
rect 14297 33958 14331 33992
rect 14297 33890 14331 33924
rect 14297 33822 14331 33856
rect 14297 33754 14331 33788
rect 14297 33686 14331 33720
rect 14297 33618 14331 33652
rect 14297 33550 14331 33584
rect 14297 33482 14331 33516
rect 14297 33414 14331 33448
rect 14297 33346 14331 33380
rect 14297 33278 14331 33312
rect 14297 33210 14331 33244
rect 14297 33142 14331 33176
rect 14297 33074 14331 33108
rect 14297 33006 14331 33040
rect 14297 32938 14331 32972
rect 14297 32870 14331 32904
rect 14297 32802 14331 32836
rect 14297 32734 14331 32768
rect 14297 32666 14331 32700
rect 14297 32598 14331 32632
rect 14297 32530 14331 32564
rect 14297 32462 14331 32496
rect 14297 32394 14331 32428
rect 14297 32326 14331 32360
rect 14297 32258 14331 32292
rect 14297 32190 14331 32224
rect 14297 32122 14331 32156
rect 14297 32054 14331 32088
rect 14297 31986 14331 32020
rect 14297 31918 14331 31952
rect 14297 31850 14331 31884
rect 14297 31782 14331 31816
rect 14297 31714 14331 31748
rect 14297 31646 14331 31680
rect 14297 31578 14331 31612
rect 14297 31510 14331 31544
rect 14297 31442 14331 31476
rect 14297 31374 14331 31408
rect 14297 31306 14331 31340
rect 14297 31238 14331 31272
rect 14297 31170 14331 31204
rect 14297 31102 14331 31136
rect 14297 31034 14331 31068
rect 14297 30966 14331 31000
rect 14297 30898 14331 30932
rect 14297 30830 14331 30864
rect 14297 30762 14331 30796
rect 14297 30694 14331 30728
rect 14297 30626 14331 30660
rect 14297 30558 14331 30592
rect 14297 30490 14331 30524
rect 14297 30422 14331 30456
rect 14297 30354 14331 30388
rect 14297 30286 14331 30320
rect 14297 30218 14331 30252
rect 14297 30150 14331 30184
rect 14297 30082 14331 30116
rect 14297 30014 14331 30048
rect 14297 29946 14331 29980
rect 14297 29878 14331 29912
rect 14297 29810 14331 29844
rect 14297 29742 14331 29776
rect 14297 29674 14331 29708
rect 14297 29606 14331 29640
rect 14297 29538 14331 29572
rect 14297 29470 14331 29504
rect 14297 29402 14331 29436
rect 14297 29334 14331 29368
rect 14297 29266 14331 29300
rect 14297 29198 14331 29232
rect 14297 29130 14331 29164
rect 14297 29062 14331 29096
rect 14297 28994 14331 29028
rect 14297 28926 14331 28960
rect 14297 28858 14331 28892
rect 14297 28790 14331 28824
rect 14297 28722 14331 28756
rect 14297 28654 14331 28688
rect 14297 28586 14331 28620
rect 14297 28518 14331 28552
rect 14297 28450 14331 28484
rect 14297 28382 14331 28416
rect 14297 28314 14331 28348
rect 14297 28246 14331 28280
rect 14297 28178 14331 28212
rect 14297 28110 14331 28144
rect 14297 28042 14331 28076
rect 14297 27974 14331 28008
rect 14297 27906 14331 27940
rect 14297 27838 14331 27872
rect 14297 27770 14331 27804
rect 14297 27702 14331 27736
rect 14297 27634 14331 27668
rect 14297 27566 14331 27600
rect 14297 27498 14331 27532
rect 14297 27430 14331 27464
rect 14297 27362 14331 27396
rect 14297 27294 14331 27328
rect 14297 27226 14331 27260
rect 14297 27158 14331 27192
rect 14297 27090 14331 27124
rect 14297 27022 14331 27056
rect 14297 26954 14331 26988
rect 14297 26886 14331 26920
rect 14297 26818 14331 26852
rect 14297 26750 14331 26784
rect 14297 26682 14331 26716
rect 14297 26614 14331 26648
rect 14297 26546 14331 26580
rect 14297 26478 14331 26512
rect 14297 26410 14331 26444
rect 14297 26342 14331 26376
rect 14297 26274 14331 26308
rect 14297 26206 14331 26240
rect 14297 26138 14331 26172
rect 14297 26070 14331 26104
rect 14297 26002 14331 26036
rect 14297 25934 14331 25968
rect 14297 25866 14331 25900
rect 14297 25798 14331 25832
rect 14297 25730 14331 25764
rect 14297 25662 14331 25696
rect 14297 25594 14331 25628
rect 14297 25526 14331 25560
rect 14297 25458 14331 25492
rect 14297 25390 14331 25424
rect 14297 25322 14331 25356
rect 14297 25254 14331 25288
rect 14297 25186 14331 25220
rect 14297 25118 14331 25152
rect 14297 25050 14331 25084
rect 14297 24982 14331 25016
rect 14297 24914 14331 24948
rect 14297 24846 14331 24880
rect 14297 24778 14331 24812
rect 14297 24710 14331 24744
rect 14297 24642 14331 24676
rect 14297 24574 14331 24608
rect 14297 24506 14331 24540
rect 14297 24438 14331 24472
rect 14297 24370 14331 24404
rect 14297 24302 14331 24336
rect 14297 24234 14331 24268
rect 14297 24166 14331 24200
rect 14297 24098 14331 24132
rect 14297 24030 14331 24064
rect 14297 23962 14331 23996
rect 14297 23894 14331 23928
rect 14297 23826 14331 23860
rect 14297 23758 14331 23792
rect 14297 23690 14331 23724
rect 14297 23622 14331 23656
rect 14297 23554 14331 23588
rect 14297 23486 14331 23520
rect 14297 23418 14331 23452
rect 14297 23350 14331 23384
rect 14297 23282 14331 23316
rect 14297 23214 14331 23248
rect 14297 23146 14331 23180
rect 14297 23078 14331 23112
rect 14297 23010 14331 23044
rect 14297 22942 14331 22976
rect 14297 22874 14331 22908
rect 14297 22806 14331 22840
rect 14297 22738 14331 22772
rect 14297 22670 14331 22704
rect 14297 22602 14331 22636
rect 14297 22534 14331 22568
rect 14297 22466 14331 22500
rect 14297 22398 14331 22432
rect 14297 22330 14331 22364
rect 14297 22262 14331 22296
rect 14297 22194 14331 22228
rect 14297 22126 14331 22160
rect 14297 22058 14331 22092
rect 14297 21990 14331 22024
rect 14297 21922 14331 21956
rect 14297 21854 14331 21888
rect 14297 21786 14331 21820
rect 14297 21718 14331 21752
rect 14297 21650 14331 21684
rect 14297 21582 14331 21616
rect 14297 21514 14331 21548
rect 14297 21446 14331 21480
rect 14297 21378 14331 21412
rect 14297 21310 14331 21344
rect 14297 21242 14331 21276
rect 14297 21174 14331 21208
rect 14297 21106 14331 21140
rect 14297 21038 14331 21072
rect 14297 20970 14331 21004
rect 14297 20902 14331 20936
rect 14297 20834 14331 20868
rect 14297 20766 14331 20800
rect 14297 20698 14331 20732
rect 14297 20630 14331 20664
rect 14297 20562 14331 20596
rect 14297 20494 14331 20528
rect 14297 20426 14331 20460
rect 14297 20358 14331 20392
rect 14297 20290 14331 20324
rect 14297 20222 14331 20256
rect 14297 20154 14331 20188
rect 14297 20086 14331 20120
rect 14297 20018 14331 20052
rect 14297 19950 14331 19984
rect 14297 19882 14331 19916
rect 14297 19814 14331 19848
rect 14297 19746 14331 19780
rect 14297 19678 14331 19712
rect 14297 19610 14331 19644
rect 14297 19542 14331 19576
rect 14297 19474 14331 19508
rect 14297 19406 14331 19440
rect 14297 19338 14331 19372
rect 14297 19270 14331 19304
rect 14297 19202 14331 19236
rect 14297 19134 14331 19168
rect 14297 19066 14331 19100
rect 14297 18998 14331 19032
rect 14297 18930 14331 18964
rect 14297 18862 14331 18896
rect 14297 18794 14331 18828
rect 14297 18726 14331 18760
rect 14297 18658 14331 18692
rect 14297 18590 14331 18624
rect 14297 18522 14331 18556
rect 14297 18454 14331 18488
rect 14297 18386 14331 18420
rect 14297 18318 14331 18352
rect 14297 18250 14331 18284
rect 14297 18182 14331 18216
rect 14297 18114 14331 18148
rect 14297 18046 14331 18080
rect 14297 17978 14331 18012
rect 14297 17910 14331 17944
rect 14297 17842 14331 17876
rect 14297 17774 14331 17808
rect 14297 17706 14331 17740
rect 14297 17638 14331 17672
rect 14297 17570 14331 17604
rect 14297 17502 14331 17536
rect 14297 17434 14331 17468
rect 14297 17366 14331 17400
rect 14297 17298 14331 17332
rect 14297 17230 14331 17264
rect 14297 17162 14331 17196
rect 14297 17094 14331 17128
rect 14297 17026 14331 17060
rect 14297 16958 14331 16992
rect 14297 16890 14331 16924
rect 14297 16822 14331 16856
rect 14297 16754 14331 16788
rect 14297 16686 14331 16720
rect 14297 16618 14331 16652
rect 14297 16550 14331 16584
rect 14297 16482 14331 16516
rect 14297 16414 14331 16448
rect 14297 16346 14331 16380
rect 14297 16278 14331 16312
rect 14297 16210 14331 16244
rect 14297 16142 14331 16176
rect 14297 16074 14331 16108
rect 14297 16006 14331 16040
rect 14297 15938 14331 15972
rect 14297 15870 14331 15904
rect 14297 15802 14331 15836
rect 14297 15734 14331 15768
rect 14297 15666 14331 15700
rect 14297 15598 14331 15632
rect 14297 15530 14331 15564
rect 14297 15462 14331 15496
rect 14297 15394 14331 15428
rect 14297 15326 14331 15360
rect 14297 15258 14331 15292
rect 14297 15190 14331 15224
rect 14297 15122 14331 15156
rect 14297 15054 14331 15088
rect 14297 14986 14331 15020
rect 14297 14918 14331 14952
rect 14297 14850 14331 14884
rect 14297 14782 14331 14816
rect 14297 14714 14331 14748
rect 14297 14646 14331 14680
rect 14297 14578 14331 14612
rect 14297 14510 14331 14544
rect 14297 14442 14331 14476
rect 14297 14374 14331 14408
rect 14297 14306 14331 14340
rect 14297 14238 14331 14272
rect 14297 14170 14331 14204
rect 14297 14102 14331 14136
rect 14297 14034 14331 14068
rect 14297 13966 14331 14000
rect 14297 13898 14331 13932
rect 14297 13830 14331 13864
rect 14297 13762 14331 13796
rect 14297 13694 14331 13728
rect 14297 13626 14331 13660
rect 14297 13558 14331 13592
rect 14297 13490 14331 13524
rect 14297 13422 14331 13456
rect 14297 13354 14331 13388
rect 14297 13286 14331 13320
rect 14297 13218 14331 13252
rect 14297 13150 14331 13184
rect 14297 13082 14331 13116
rect 14297 13014 14331 13048
rect 14297 12946 14331 12980
rect 14297 12878 14331 12912
rect 14297 12810 14331 12844
rect 14297 12742 14331 12776
rect 14297 12674 14331 12708
rect 14297 12606 14331 12640
rect 14297 12538 14331 12572
rect 14297 12470 14331 12504
rect 14297 12402 14331 12436
rect 14297 12334 14331 12368
rect 14297 12266 14331 12300
rect 14297 12198 14331 12232
rect 14297 12130 14331 12164
rect 14297 12062 14331 12096
rect 14297 11994 14331 12028
rect 14297 11926 14331 11960
rect 14297 11858 14331 11892
rect 14297 11790 14331 11824
rect 14297 11722 14331 11756
rect 14297 11654 14331 11688
rect 14297 11586 14331 11620
rect 14297 11518 14331 11552
rect 14297 11450 14331 11484
rect 14297 11382 14331 11416
rect 14297 11314 14331 11348
rect 14297 11246 14331 11280
rect 14297 11178 14331 11212
rect 14297 11110 14331 11144
rect 14297 11042 14331 11076
rect 14297 10974 14331 11008
rect 14297 10906 14331 10940
rect 14297 10838 14331 10872
rect 14297 10770 14331 10804
rect 14297 10702 14331 10736
rect 14297 10634 14331 10668
rect 14297 10566 14331 10600
rect 14297 10498 14331 10532
rect 14297 10430 14331 10464
rect 14297 10362 14331 10396
rect 14297 10294 14331 10328
rect 632 10158 666 10192
rect 632 10090 666 10124
rect 632 10022 666 10056
rect 632 9954 666 9988
rect 632 9886 666 9920
rect 14297 10226 14331 10260
rect 14297 10158 14331 10192
rect 14297 10090 14331 10124
rect 14297 10022 14331 10056
rect 14297 9954 14331 9988
rect 14297 9886 14331 9920
rect 740 9741 774 9775
rect 808 9741 842 9775
rect 915 9741 949 9775
rect 983 9741 1017 9775
rect 1051 9741 1085 9775
rect 1119 9741 1153 9775
rect 1187 9741 1221 9775
rect 1255 9741 1289 9775
rect 1323 9741 1357 9775
rect 1391 9741 1425 9775
rect 1459 9741 1493 9775
rect 1527 9741 1561 9775
rect 1595 9741 1629 9775
rect 1663 9741 1697 9775
rect 1731 9741 1765 9775
rect 1799 9741 1833 9775
rect 1867 9741 1901 9775
rect 1935 9741 1969 9775
rect 2003 9741 2037 9775
rect 2121 9741 2155 9775
rect 2189 9741 2223 9775
rect 2257 9741 2291 9775
rect 2325 9741 2359 9775
rect 2393 9741 2427 9775
rect 2461 9741 2495 9775
rect 2529 9741 2563 9775
rect 2597 9741 2631 9775
rect 2665 9741 2699 9775
rect 2733 9741 2767 9775
rect 2801 9741 2835 9775
rect 2869 9741 2903 9775
rect 2937 9741 2971 9775
rect 3005 9741 3039 9775
rect 3073 9741 3107 9775
rect 3141 9741 3175 9775
rect 3209 9741 3243 9775
rect 3277 9741 3311 9775
rect 3345 9741 3379 9775
rect 3413 9741 3447 9775
rect 3481 9741 3515 9775
rect 3549 9741 3583 9775
rect 3617 9741 3651 9775
rect 3685 9741 3719 9775
rect 3753 9741 3787 9775
rect 3821 9741 3855 9775
rect 3889 9741 3923 9775
rect 3957 9741 3991 9775
rect 4025 9741 4059 9775
rect 4093 9741 4127 9775
rect 4161 9741 4195 9775
rect 4229 9741 4263 9775
rect 4297 9741 4331 9775
rect 4365 9741 4399 9775
rect 4433 9741 4467 9775
rect 4501 9741 4535 9775
rect 4569 9741 4603 9775
rect 4637 9741 4671 9775
rect 4705 9741 4739 9775
rect 4773 9741 4807 9775
rect 4841 9741 4875 9775
rect 4909 9741 4943 9775
rect 4977 9741 5011 9775
rect 5045 9741 5079 9775
rect 5113 9741 5147 9775
rect 5181 9741 5215 9775
rect 5249 9741 5283 9775
rect 5317 9741 5351 9775
rect 5385 9741 5419 9775
rect 5453 9741 5487 9775
rect 5521 9741 5555 9775
rect 5589 9741 5623 9775
rect 5657 9741 5691 9775
rect 5725 9741 5759 9775
rect 5793 9741 5827 9775
rect 5861 9741 5895 9775
rect 5929 9741 5963 9775
rect 5997 9741 6031 9775
rect 6065 9741 6099 9775
rect 6133 9741 6167 9775
rect 6201 9741 6235 9775
rect 6269 9741 6303 9775
rect 6337 9741 6371 9775
rect 6405 9741 6439 9775
rect 6473 9741 6507 9775
rect 6541 9741 6575 9775
rect 6609 9741 6643 9775
rect 6677 9741 6711 9775
rect 6745 9741 6779 9775
rect 6813 9741 6847 9775
rect 6881 9741 6915 9775
rect 6949 9741 6983 9775
rect 7017 9741 7051 9775
rect 7085 9741 7119 9775
rect 7153 9741 7187 9775
rect 7221 9741 7255 9775
rect 7289 9741 7323 9775
rect 7357 9741 7391 9775
rect 7425 9741 7459 9775
rect 7493 9741 7527 9775
rect 7561 9741 7595 9775
rect 7629 9741 7663 9775
rect 7697 9741 7731 9775
rect 7765 9741 7799 9775
rect 7833 9741 7867 9775
rect 7901 9741 7935 9775
rect 7969 9741 8003 9775
rect 8037 9741 8071 9775
rect 8105 9741 8139 9775
rect 8173 9741 8207 9775
rect 8241 9741 8275 9775
rect 8309 9741 8343 9775
rect 8377 9741 8411 9775
rect 8445 9741 8479 9775
rect 8513 9741 8547 9775
rect 8581 9741 8615 9775
rect 8649 9741 8683 9775
rect 8717 9741 8751 9775
rect 8785 9741 8819 9775
rect 8853 9741 8887 9775
rect 8921 9741 8955 9775
rect 8989 9741 9023 9775
rect 9057 9741 9091 9775
rect 9125 9741 9159 9775
rect 9193 9741 9227 9775
rect 9261 9741 9295 9775
rect 9329 9741 9363 9775
rect 9397 9741 9431 9775
rect 9465 9741 9499 9775
rect 9533 9741 9567 9775
rect 9601 9741 9635 9775
rect 9669 9741 9703 9775
rect 9737 9741 9771 9775
rect 9805 9741 9839 9775
rect 9873 9741 9907 9775
rect 9941 9741 9975 9775
rect 10009 9741 10043 9775
rect 10077 9741 10111 9775
rect 10145 9741 10179 9775
rect 10213 9741 10247 9775
rect 10281 9741 10315 9775
rect 10349 9741 10383 9775
rect 10417 9741 10451 9775
rect 10485 9741 10519 9775
rect 10553 9741 10587 9775
rect 10621 9741 10655 9775
rect 10689 9741 10723 9775
rect 10757 9741 10791 9775
rect 10825 9741 10859 9775
rect 10893 9741 10927 9775
rect 10961 9741 10995 9775
rect 11029 9741 11063 9775
rect 11097 9741 11131 9775
rect 11165 9741 11199 9775
rect 11233 9741 11267 9775
rect 11301 9741 11335 9775
rect 11369 9741 11403 9775
rect 11437 9741 11471 9775
rect 11505 9741 11539 9775
rect 11573 9741 11607 9775
rect 11641 9741 11675 9775
rect 11709 9741 11743 9775
rect 11777 9741 11811 9775
rect 11845 9741 11879 9775
rect 11913 9741 11947 9775
rect 11981 9741 12015 9775
rect 12049 9741 12083 9775
rect 12117 9741 12151 9775
rect 12185 9741 12219 9775
rect 12253 9741 12287 9775
rect 12321 9741 12355 9775
rect 12389 9741 12423 9775
rect 12457 9741 12491 9775
rect 12525 9741 12559 9775
rect 12593 9741 12627 9775
rect 12661 9741 12695 9775
rect 12729 9741 12763 9775
rect 12797 9741 12831 9775
rect 12915 9740 12949 9774
rect 12983 9740 13017 9774
rect 13051 9740 13085 9774
rect 13119 9740 13153 9774
rect 13187 9740 13221 9774
rect 13255 9740 13289 9774
rect 13323 9740 13357 9774
rect 13391 9740 13425 9774
rect 13459 9740 13493 9774
rect 13527 9740 13561 9774
rect 13595 9740 13629 9774
rect 13663 9740 13697 9774
rect 13731 9740 13765 9774
rect 13799 9740 13833 9774
rect 13867 9740 13901 9774
rect 13935 9740 13969 9774
rect 14003 9740 14037 9774
rect 14115 9741 14149 9775
rect 14183 9741 14217 9775
<< locali >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36464 532 36498
rect 590 36464 600 36498
rect 662 36464 668 36498
rect 734 36464 736 36498
rect 770 36464 772 36498
rect 838 36464 844 36498
rect 906 36464 916 36498
rect 974 36464 988 36498
rect 1042 36464 1060 36498
rect 1110 36464 1132 36498
rect 1178 36464 1204 36498
rect 1246 36464 1276 36498
rect 1314 36464 1348 36498
rect 1382 36464 1416 36498
rect 1454 36464 1484 36498
rect 1526 36464 1552 36498
rect 1598 36464 1620 36498
rect 1670 36464 1688 36498
rect 1742 36464 1756 36498
rect 1814 36464 1824 36498
rect 1886 36464 1892 36498
rect 1958 36464 1960 36498
rect 1994 36464 1996 36498
rect 2062 36464 2068 36498
rect 2130 36464 2140 36498
rect 2198 36464 2212 36498
rect 2266 36464 2284 36498
rect 2334 36464 2356 36498
rect 2402 36464 2428 36498
rect 2470 36464 2500 36498
rect 2538 36464 2572 36498
rect 2606 36464 2640 36498
rect 2678 36464 2708 36498
rect 2750 36464 2776 36498
rect 2822 36464 2844 36498
rect 2894 36464 2912 36498
rect 2966 36464 2980 36498
rect 3038 36464 3048 36498
rect 3110 36464 3116 36498
rect 3182 36464 3184 36498
rect 3218 36464 3220 36498
rect 3286 36464 3292 36498
rect 3354 36464 3364 36498
rect 3422 36464 3436 36498
rect 3490 36464 3508 36498
rect 3558 36464 3580 36498
rect 3626 36464 3652 36498
rect 3694 36464 3724 36498
rect 3762 36464 3796 36498
rect 3830 36464 3864 36498
rect 3902 36464 3932 36498
rect 3974 36464 4000 36498
rect 4046 36464 4068 36498
rect 4118 36464 4136 36498
rect 4190 36464 4204 36498
rect 4262 36464 4272 36498
rect 4334 36464 4340 36498
rect 4406 36464 4408 36498
rect 4442 36464 4444 36498
rect 4510 36464 4516 36498
rect 4578 36464 4588 36498
rect 4646 36464 4660 36498
rect 4714 36464 4732 36498
rect 4782 36464 4804 36498
rect 4850 36464 4876 36498
rect 4918 36464 4948 36498
rect 4986 36464 5020 36498
rect 5054 36464 5088 36498
rect 5126 36464 5156 36498
rect 5198 36464 5224 36498
rect 5270 36464 5292 36498
rect 5342 36464 5360 36498
rect 5414 36464 5428 36498
rect 5486 36464 5496 36498
rect 5558 36464 5564 36498
rect 5630 36464 5632 36498
rect 5666 36464 5668 36498
rect 5734 36464 5740 36498
rect 5802 36464 5812 36498
rect 5870 36464 5884 36498
rect 5938 36464 5956 36498
rect 6006 36464 6028 36498
rect 6074 36464 6100 36498
rect 6142 36464 6172 36498
rect 6210 36464 6244 36498
rect 6278 36464 6312 36498
rect 6350 36464 6380 36498
rect 6422 36464 6448 36498
rect 6494 36464 6516 36498
rect 6566 36464 6584 36498
rect 6638 36464 6652 36498
rect 6710 36464 6720 36498
rect 6782 36464 6788 36498
rect 6854 36464 6856 36498
rect 6890 36464 6892 36498
rect 6958 36464 6964 36498
rect 7026 36464 7036 36498
rect 7094 36464 7108 36498
rect 7162 36464 7180 36498
rect 7230 36464 7252 36498
rect 7298 36464 7324 36498
rect 7366 36464 7396 36498
rect 7434 36464 7468 36498
rect 7502 36464 7536 36498
rect 7574 36464 7604 36498
rect 7646 36464 7672 36498
rect 7718 36464 7740 36498
rect 7790 36464 7808 36498
rect 7862 36464 7876 36498
rect 7934 36464 7944 36498
rect 8006 36464 8012 36498
rect 8078 36464 8080 36498
rect 8114 36464 8116 36498
rect 8182 36464 8188 36498
rect 8250 36464 8260 36498
rect 8318 36464 8332 36498
rect 8386 36464 8404 36498
rect 8454 36464 8476 36498
rect 8522 36464 8548 36498
rect 8590 36464 8620 36498
rect 8658 36464 8692 36498
rect 8726 36464 8760 36498
rect 8798 36464 8828 36498
rect 8870 36464 8896 36498
rect 8942 36464 8964 36498
rect 9014 36464 9032 36498
rect 9086 36464 9100 36498
rect 9158 36464 9168 36498
rect 9230 36464 9236 36498
rect 9302 36464 9304 36498
rect 9338 36464 9340 36498
rect 9406 36464 9412 36498
rect 9474 36464 9484 36498
rect 9542 36464 9556 36498
rect 9610 36464 9628 36498
rect 9678 36464 9700 36498
rect 9746 36464 9772 36498
rect 9814 36464 9844 36498
rect 9882 36464 9916 36498
rect 9950 36464 9984 36498
rect 10022 36464 10052 36498
rect 10094 36464 10120 36498
rect 10166 36464 10188 36498
rect 10238 36464 10256 36498
rect 10310 36464 10324 36498
rect 10382 36464 10392 36498
rect 10454 36464 10460 36498
rect 10526 36464 10528 36498
rect 10562 36464 10564 36498
rect 10630 36464 10636 36498
rect 10698 36464 10708 36498
rect 10766 36464 10780 36498
rect 10834 36464 10852 36498
rect 10902 36464 10924 36498
rect 10970 36464 10996 36498
rect 11038 36464 11068 36498
rect 11106 36464 11140 36498
rect 11174 36464 11208 36498
rect 11246 36464 11276 36498
rect 11318 36464 11344 36498
rect 11390 36464 11412 36498
rect 11462 36464 11480 36498
rect 11534 36464 11548 36498
rect 11606 36464 11616 36498
rect 11678 36464 11684 36498
rect 11750 36464 11752 36498
rect 11786 36464 11788 36498
rect 11854 36464 11860 36498
rect 11922 36464 11932 36498
rect 11990 36464 12004 36498
rect 12058 36464 12076 36498
rect 12126 36464 12148 36498
rect 12194 36464 12220 36498
rect 12262 36464 12292 36498
rect 12330 36464 12364 36498
rect 12398 36464 12432 36498
rect 12470 36464 12500 36498
rect 12542 36464 12568 36498
rect 12614 36464 12636 36498
rect 12686 36464 12704 36498
rect 12758 36464 12772 36498
rect 12830 36464 12840 36498
rect 12902 36464 12908 36498
rect 12974 36464 12976 36498
rect 13010 36464 13012 36498
rect 13078 36464 13084 36498
rect 13146 36464 13156 36498
rect 13214 36464 13228 36498
rect 13282 36464 13300 36498
rect 13350 36464 13372 36498
rect 13418 36464 13444 36498
rect 13486 36464 13516 36498
rect 13554 36464 13588 36498
rect 13622 36464 13656 36498
rect 13694 36464 13724 36498
rect 13766 36464 13792 36498
rect 13838 36464 13860 36498
rect 13910 36464 13928 36498
rect 13982 36464 13996 36498
rect 14054 36464 14064 36498
rect 14126 36464 14132 36498
rect 14198 36464 14200 36498
rect 14234 36464 14236 36498
rect 14302 36464 14308 36498
rect 14370 36464 14380 36498
rect 14438 36464 14472 36498
rect 14506 36464 14724 36498
rect 245 36462 14724 36464
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36311 430 36389
rect 245 36277 317 36311
rect 351 36277 430 36311
rect 245 36265 430 36277
rect 245 36243 320 36265
rect 245 36209 317 36243
rect 354 36231 430 36265
rect 351 36209 430 36231
rect 245 36193 430 36209
rect 14539 36309 14724 36389
rect 14539 36275 14611 36309
rect 14645 36275 14724 36309
rect 14539 36262 14724 36275
rect 14539 36241 14614 36262
rect 14539 36207 14611 36241
rect 14648 36228 14724 36262
rect 14645 36207 14724 36228
rect 245 36175 320 36193
rect 245 36141 317 36175
rect 354 36159 430 36193
rect 351 36141 430 36159
rect 245 36121 430 36141
rect 245 36107 320 36121
rect 245 36073 317 36107
rect 354 36087 430 36121
rect 351 36073 430 36087
rect 245 36049 430 36073
rect 245 36039 320 36049
rect 245 36005 317 36039
rect 354 36015 430 36049
rect 351 36005 430 36015
rect 245 35977 430 36005
rect 245 35971 320 35977
rect 245 35937 317 35971
rect 354 35943 430 35977
rect 351 35937 430 35943
rect 245 35905 430 35937
rect 245 35903 320 35905
rect 245 35869 317 35903
rect 354 35871 430 35905
rect 351 35869 430 35871
rect 245 35835 430 35869
rect 245 35801 317 35835
rect 351 35833 430 35835
rect 245 35799 320 35801
rect 354 35799 430 35833
rect 245 35767 430 35799
rect 245 35733 317 35767
rect 351 35761 430 35767
rect 245 35727 320 35733
rect 354 35727 430 35761
rect 245 35699 430 35727
rect 245 35665 317 35699
rect 351 35689 430 35699
rect 245 35655 320 35665
rect 354 35655 430 35689
rect 245 35631 430 35655
rect 245 35597 317 35631
rect 351 35617 430 35631
rect 245 35583 320 35597
rect 354 35583 430 35617
rect 245 35563 430 35583
rect 245 35529 317 35563
rect 351 35545 430 35563
rect 245 35511 320 35529
rect 354 35511 430 35545
rect 245 35495 430 35511
rect 245 35461 317 35495
rect 351 35473 430 35495
rect 245 35439 320 35461
rect 354 35439 430 35473
rect 245 35427 430 35439
rect 245 35393 317 35427
rect 351 35401 430 35427
rect 245 35367 320 35393
rect 354 35367 430 35401
rect 245 35359 430 35367
rect 245 35325 317 35359
rect 351 35329 430 35359
rect 245 35295 320 35325
rect 354 35295 430 35329
rect 245 35291 430 35295
rect 245 35257 317 35291
rect 351 35257 430 35291
rect 245 35223 320 35257
rect 354 35223 430 35257
rect 245 35189 317 35223
rect 351 35189 430 35223
rect 245 35185 430 35189
rect 245 35155 320 35185
rect 245 35121 317 35155
rect 354 35151 430 35185
rect 351 35121 430 35151
rect 245 35113 430 35121
rect 245 35087 320 35113
rect 245 35053 317 35087
rect 354 35079 430 35113
rect 351 35053 430 35079
rect 245 35041 430 35053
rect 245 35019 320 35041
rect 245 34985 317 35019
rect 354 35007 430 35041
rect 351 34985 430 35007
rect 245 34969 430 34985
rect 245 34951 320 34969
rect 245 34917 317 34951
rect 354 34935 430 34969
rect 351 34917 430 34935
rect 245 34897 430 34917
rect 245 34883 320 34897
rect 245 34849 317 34883
rect 354 34863 430 34897
rect 351 34849 430 34863
rect 245 34825 430 34849
rect 245 34815 320 34825
rect 245 34781 317 34815
rect 354 34791 430 34825
rect 351 34781 430 34791
rect 245 34753 430 34781
rect 245 34747 320 34753
rect 245 34713 317 34747
rect 354 34719 430 34753
rect 351 34713 430 34719
rect 245 34681 430 34713
rect 245 34679 320 34681
rect 245 34645 317 34679
rect 354 34647 430 34681
rect 351 34645 430 34647
rect 245 34611 430 34645
rect 245 34577 317 34611
rect 351 34609 430 34611
rect 245 34575 320 34577
rect 354 34575 430 34609
rect 245 34543 430 34575
rect 245 34509 317 34543
rect 351 34537 430 34543
rect 245 34503 320 34509
rect 354 34503 430 34537
rect 245 34475 430 34503
rect 245 34441 317 34475
rect 351 34465 430 34475
rect 245 34431 320 34441
rect 354 34431 430 34465
rect 245 34407 430 34431
rect 245 34373 317 34407
rect 351 34393 430 34407
rect 245 34359 320 34373
rect 354 34359 430 34393
rect 245 34339 430 34359
rect 245 34305 317 34339
rect 351 34321 430 34339
rect 245 34287 320 34305
rect 354 34287 430 34321
rect 245 34271 430 34287
rect 245 34237 317 34271
rect 351 34249 430 34271
rect 245 34215 320 34237
rect 354 34215 430 34249
rect 245 34203 430 34215
rect 245 34169 317 34203
rect 351 34177 430 34203
rect 245 34143 320 34169
rect 354 34143 430 34177
rect 245 34135 430 34143
rect 245 34101 317 34135
rect 351 34105 430 34135
rect 245 34071 320 34101
rect 354 34071 430 34105
rect 245 34067 430 34071
rect 245 34033 317 34067
rect 351 34033 430 34067
rect 245 33999 320 34033
rect 354 33999 430 34033
rect 245 33965 317 33999
rect 351 33965 430 33999
rect 245 33961 430 33965
rect 245 33931 320 33961
rect 245 33897 317 33931
rect 354 33927 430 33961
rect 351 33897 430 33927
rect 245 33889 430 33897
rect 245 33863 320 33889
rect 245 33829 317 33863
rect 354 33855 430 33889
rect 351 33829 430 33855
rect 245 33817 430 33829
rect 245 33795 320 33817
rect 245 33761 317 33795
rect 354 33783 430 33817
rect 351 33761 430 33783
rect 245 33745 430 33761
rect 245 33727 320 33745
rect 245 33693 317 33727
rect 354 33711 430 33745
rect 351 33693 430 33711
rect 245 33673 430 33693
rect 245 33659 320 33673
rect 245 33625 317 33659
rect 354 33639 430 33673
rect 351 33625 430 33639
rect 245 33601 430 33625
rect 245 33591 320 33601
rect 245 33557 317 33591
rect 354 33567 430 33601
rect 351 33557 430 33567
rect 245 33529 430 33557
rect 245 33523 320 33529
rect 245 33489 317 33523
rect 354 33495 430 33529
rect 351 33489 430 33495
rect 245 33457 430 33489
rect 245 33455 320 33457
rect 245 33421 317 33455
rect 354 33423 430 33457
rect 351 33421 430 33423
rect 245 33387 430 33421
rect 245 33353 317 33387
rect 351 33385 430 33387
rect 245 33351 320 33353
rect 354 33351 430 33385
rect 245 33319 430 33351
rect 245 33285 317 33319
rect 351 33313 430 33319
rect 245 33279 320 33285
rect 354 33279 430 33313
rect 245 33251 430 33279
rect 245 33217 317 33251
rect 351 33241 430 33251
rect 245 33207 320 33217
rect 354 33207 430 33241
rect 245 33183 430 33207
rect 245 33149 317 33183
rect 351 33169 430 33183
rect 245 33135 320 33149
rect 354 33135 430 33169
rect 245 33115 430 33135
rect 245 33081 317 33115
rect 351 33097 430 33115
rect 245 33063 320 33081
rect 354 33063 430 33097
rect 245 33047 430 33063
rect 245 33013 317 33047
rect 351 33025 430 33047
rect 245 32991 320 33013
rect 354 32991 430 33025
rect 245 32979 430 32991
rect 245 32945 317 32979
rect 351 32953 430 32979
rect 245 32919 320 32945
rect 354 32919 430 32953
rect 245 32911 430 32919
rect 245 32877 317 32911
rect 351 32881 430 32911
rect 245 32847 320 32877
rect 354 32847 430 32881
rect 245 32843 430 32847
rect 245 32809 317 32843
rect 351 32809 430 32843
rect 245 32775 320 32809
rect 354 32775 430 32809
rect 245 32741 317 32775
rect 351 32741 430 32775
rect 245 32737 430 32741
rect 245 32707 320 32737
rect 245 32673 317 32707
rect 354 32703 430 32737
rect 351 32673 430 32703
rect 245 32665 430 32673
rect 245 32639 320 32665
rect 245 32605 317 32639
rect 354 32631 430 32665
rect 351 32605 430 32631
rect 245 32593 430 32605
rect 245 32571 320 32593
rect 245 32537 317 32571
rect 354 32559 430 32593
rect 351 32537 430 32559
rect 245 32521 430 32537
rect 245 32503 320 32521
rect 245 32469 317 32503
rect 354 32487 430 32521
rect 351 32469 430 32487
rect 245 32449 430 32469
rect 245 32435 320 32449
rect 245 32401 317 32435
rect 354 32415 430 32449
rect 351 32401 430 32415
rect 245 32377 430 32401
rect 245 32367 320 32377
rect 245 32333 317 32367
rect 354 32343 430 32377
rect 351 32333 430 32343
rect 245 32305 430 32333
rect 245 32299 320 32305
rect 245 32265 317 32299
rect 354 32271 430 32305
rect 351 32265 430 32271
rect 245 32233 430 32265
rect 245 32231 320 32233
rect 245 32197 317 32231
rect 354 32199 430 32233
rect 351 32197 430 32199
rect 245 32163 430 32197
rect 245 32129 317 32163
rect 351 32161 430 32163
rect 245 32127 320 32129
rect 354 32127 430 32161
rect 245 32095 430 32127
rect 245 32061 317 32095
rect 351 32089 430 32095
rect 245 32055 320 32061
rect 354 32055 430 32089
rect 245 32027 430 32055
rect 245 31993 317 32027
rect 351 32017 430 32027
rect 245 31983 320 31993
rect 354 31983 430 32017
rect 245 31959 430 31983
rect 245 31925 317 31959
rect 351 31945 430 31959
rect 245 31911 320 31925
rect 354 31911 430 31945
rect 245 31891 430 31911
rect 245 31857 317 31891
rect 351 31873 430 31891
rect 245 31839 320 31857
rect 354 31839 430 31873
rect 245 31823 430 31839
rect 245 31789 317 31823
rect 351 31801 430 31823
rect 245 31767 320 31789
rect 354 31767 430 31801
rect 245 31755 430 31767
rect 245 31721 317 31755
rect 351 31729 430 31755
rect 245 31695 320 31721
rect 354 31695 430 31729
rect 245 31687 430 31695
rect 245 31653 317 31687
rect 351 31657 430 31687
rect 245 31623 320 31653
rect 354 31623 430 31657
rect 245 31619 430 31623
rect 245 31585 317 31619
rect 351 31585 430 31619
rect 245 31551 320 31585
rect 354 31551 430 31585
rect 245 31517 317 31551
rect 351 31517 430 31551
rect 245 31513 430 31517
rect 245 31483 320 31513
rect 245 31449 317 31483
rect 354 31479 430 31513
rect 351 31449 430 31479
rect 245 31441 430 31449
rect 245 31415 320 31441
rect 245 31381 317 31415
rect 354 31407 430 31441
rect 351 31381 430 31407
rect 245 31369 430 31381
rect 245 31347 320 31369
rect 245 31313 317 31347
rect 354 31335 430 31369
rect 351 31313 430 31335
rect 245 31297 430 31313
rect 245 31279 320 31297
rect 245 31245 317 31279
rect 354 31263 430 31297
rect 351 31245 430 31263
rect 245 31225 430 31245
rect 245 31211 320 31225
rect 245 31177 317 31211
rect 354 31191 430 31225
rect 351 31177 430 31191
rect 245 31153 430 31177
rect 245 31143 320 31153
rect 245 31109 317 31143
rect 354 31119 430 31153
rect 351 31109 430 31119
rect 245 31081 430 31109
rect 245 31075 320 31081
rect 245 31041 317 31075
rect 354 31047 430 31081
rect 351 31041 430 31047
rect 245 31009 430 31041
rect 245 31007 320 31009
rect 245 30973 317 31007
rect 354 30975 430 31009
rect 351 30973 430 30975
rect 245 30939 430 30973
rect 245 30905 317 30939
rect 351 30937 430 30939
rect 245 30903 320 30905
rect 354 30903 430 30937
rect 245 30871 430 30903
rect 245 30837 317 30871
rect 351 30865 430 30871
rect 245 30831 320 30837
rect 354 30831 430 30865
rect 245 30803 430 30831
rect 245 30769 317 30803
rect 351 30793 430 30803
rect 245 30759 320 30769
rect 354 30759 430 30793
rect 245 30735 430 30759
rect 245 30701 317 30735
rect 351 30721 430 30735
rect 245 30687 320 30701
rect 354 30687 430 30721
rect 245 30667 430 30687
rect 245 30633 317 30667
rect 351 30649 430 30667
rect 245 30615 320 30633
rect 354 30615 430 30649
rect 245 30599 430 30615
rect 245 30565 317 30599
rect 351 30577 430 30599
rect 245 30543 320 30565
rect 354 30543 430 30577
rect 245 30531 430 30543
rect 245 30497 317 30531
rect 351 30505 430 30531
rect 245 30471 320 30497
rect 354 30471 430 30505
rect 245 30463 430 30471
rect 245 30429 317 30463
rect 351 30433 430 30463
rect 245 30399 320 30429
rect 354 30399 430 30433
rect 245 30395 430 30399
rect 245 30361 317 30395
rect 351 30361 430 30395
rect 245 30327 320 30361
rect 354 30327 430 30361
rect 245 30293 317 30327
rect 351 30293 430 30327
rect 245 30289 430 30293
rect 245 30259 320 30289
rect 245 30225 317 30259
rect 354 30255 430 30289
rect 351 30225 430 30255
rect 245 30217 430 30225
rect 245 30191 320 30217
rect 245 30157 317 30191
rect 354 30183 430 30217
rect 351 30157 430 30183
rect 245 30145 430 30157
rect 245 30123 320 30145
rect 245 30089 317 30123
rect 354 30111 430 30145
rect 351 30089 430 30111
rect 245 30073 430 30089
rect 245 30055 320 30073
rect 245 30021 317 30055
rect 354 30039 430 30073
rect 351 30021 430 30039
rect 245 30001 430 30021
rect 245 29987 320 30001
rect 245 29953 317 29987
rect 354 29967 430 30001
rect 351 29953 430 29967
rect 245 29929 430 29953
rect 245 29919 320 29929
rect 245 29885 317 29919
rect 354 29895 430 29929
rect 351 29885 430 29895
rect 245 29857 430 29885
rect 245 29851 320 29857
rect 245 29817 317 29851
rect 354 29823 430 29857
rect 351 29817 430 29823
rect 245 29785 430 29817
rect 245 29783 320 29785
rect 245 29749 317 29783
rect 354 29751 430 29785
rect 351 29749 430 29751
rect 245 29715 430 29749
rect 245 29681 317 29715
rect 351 29713 430 29715
rect 245 29679 320 29681
rect 354 29679 430 29713
rect 245 29647 430 29679
rect 245 29613 317 29647
rect 351 29641 430 29647
rect 245 29607 320 29613
rect 354 29607 430 29641
rect 245 29579 430 29607
rect 245 29545 317 29579
rect 351 29569 430 29579
rect 245 29535 320 29545
rect 354 29535 430 29569
rect 245 29511 430 29535
rect 245 29477 317 29511
rect 351 29497 430 29511
rect 245 29463 320 29477
rect 354 29463 430 29497
rect 245 29443 430 29463
rect 245 29409 317 29443
rect 351 29425 430 29443
rect 245 29391 320 29409
rect 354 29391 430 29425
rect 245 29375 430 29391
rect 245 29341 317 29375
rect 351 29353 430 29375
rect 245 29319 320 29341
rect 354 29319 430 29353
rect 245 29307 430 29319
rect 245 29273 317 29307
rect 351 29281 430 29307
rect 245 29247 320 29273
rect 354 29247 430 29281
rect 245 29239 430 29247
rect 245 29205 317 29239
rect 351 29209 430 29239
rect 245 29175 320 29205
rect 354 29175 430 29209
rect 245 29171 430 29175
rect 245 29137 317 29171
rect 351 29137 430 29171
rect 245 29103 320 29137
rect 354 29103 430 29137
rect 245 29069 317 29103
rect 351 29069 430 29103
rect 245 29065 430 29069
rect 245 29035 320 29065
rect 245 29001 317 29035
rect 354 29031 430 29065
rect 351 29001 430 29031
rect 245 28993 430 29001
rect 245 28967 320 28993
rect 245 28933 317 28967
rect 354 28959 430 28993
rect 351 28933 430 28959
rect 245 28921 430 28933
rect 245 28899 320 28921
rect 245 28865 317 28899
rect 354 28887 430 28921
rect 351 28865 430 28887
rect 245 28849 430 28865
rect 245 28831 320 28849
rect 245 28797 317 28831
rect 354 28815 430 28849
rect 351 28797 430 28815
rect 245 28777 430 28797
rect 245 28763 320 28777
rect 245 28729 317 28763
rect 354 28743 430 28777
rect 351 28729 430 28743
rect 245 28705 430 28729
rect 245 28695 320 28705
rect 245 28661 317 28695
rect 354 28671 430 28705
rect 351 28661 430 28671
rect 245 28633 430 28661
rect 245 28627 320 28633
rect 245 28593 317 28627
rect 354 28599 430 28633
rect 351 28593 430 28599
rect 245 28561 430 28593
rect 245 28559 320 28561
rect 245 28525 317 28559
rect 354 28527 430 28561
rect 351 28525 430 28527
rect 245 28491 430 28525
rect 245 28457 317 28491
rect 351 28489 430 28491
rect 245 28455 320 28457
rect 354 28455 430 28489
rect 245 28423 430 28455
rect 245 28389 317 28423
rect 351 28417 430 28423
rect 245 28383 320 28389
rect 354 28383 430 28417
rect 245 28355 430 28383
rect 245 28321 317 28355
rect 351 28345 430 28355
rect 245 28311 320 28321
rect 354 28311 430 28345
rect 245 28287 430 28311
rect 245 28253 317 28287
rect 351 28273 430 28287
rect 245 28239 320 28253
rect 354 28239 430 28273
rect 245 28219 430 28239
rect 245 28185 317 28219
rect 351 28201 430 28219
rect 245 28167 320 28185
rect 354 28167 430 28201
rect 245 28151 430 28167
rect 245 28117 317 28151
rect 351 28129 430 28151
rect 245 28095 320 28117
rect 354 28095 430 28129
rect 245 28083 430 28095
rect 245 28049 317 28083
rect 351 28057 430 28083
rect 245 28023 320 28049
rect 354 28023 430 28057
rect 245 28015 430 28023
rect 245 27981 317 28015
rect 351 27985 430 28015
rect 245 27951 320 27981
rect 354 27951 430 27985
rect 245 27947 430 27951
rect 245 27913 317 27947
rect 351 27913 430 27947
rect 245 27879 320 27913
rect 354 27879 430 27913
rect 245 27845 317 27879
rect 351 27845 430 27879
rect 245 27841 430 27845
rect 245 27811 320 27841
rect 245 27777 317 27811
rect 354 27807 430 27841
rect 351 27777 430 27807
rect 245 27769 430 27777
rect 245 27743 320 27769
rect 245 27709 317 27743
rect 354 27735 430 27769
rect 351 27709 430 27735
rect 245 27697 430 27709
rect 245 27675 320 27697
rect 245 27641 317 27675
rect 354 27663 430 27697
rect 351 27641 430 27663
rect 245 27625 430 27641
rect 245 27607 320 27625
rect 245 27573 317 27607
rect 354 27591 430 27625
rect 351 27573 430 27591
rect 245 27553 430 27573
rect 245 27539 320 27553
rect 245 27505 317 27539
rect 354 27519 430 27553
rect 351 27505 430 27519
rect 245 27481 430 27505
rect 245 27471 320 27481
rect 245 27437 317 27471
rect 354 27447 430 27481
rect 351 27437 430 27447
rect 245 27409 430 27437
rect 245 27403 320 27409
rect 245 27369 317 27403
rect 354 27375 430 27409
rect 351 27369 430 27375
rect 245 27337 430 27369
rect 245 27335 320 27337
rect 245 27301 317 27335
rect 354 27303 430 27337
rect 351 27301 430 27303
rect 245 27267 430 27301
rect 245 27233 317 27267
rect 351 27265 430 27267
rect 245 27231 320 27233
rect 354 27231 430 27265
rect 245 27199 430 27231
rect 245 27165 317 27199
rect 351 27193 430 27199
rect 245 27159 320 27165
rect 354 27159 430 27193
rect 245 27131 430 27159
rect 245 27097 317 27131
rect 351 27121 430 27131
rect 245 27087 320 27097
rect 354 27087 430 27121
rect 245 27063 430 27087
rect 245 27029 317 27063
rect 351 27049 430 27063
rect 245 27015 320 27029
rect 354 27015 430 27049
rect 245 26995 430 27015
rect 245 26961 317 26995
rect 351 26977 430 26995
rect 245 26943 320 26961
rect 354 26943 430 26977
rect 245 26927 430 26943
rect 245 26893 317 26927
rect 351 26905 430 26927
rect 245 26871 320 26893
rect 354 26871 430 26905
rect 245 26859 430 26871
rect 245 26825 317 26859
rect 351 26833 430 26859
rect 245 26799 320 26825
rect 354 26799 430 26833
rect 245 26791 430 26799
rect 245 26757 317 26791
rect 351 26761 430 26791
rect 245 26727 320 26757
rect 354 26727 430 26761
rect 245 26723 430 26727
rect 245 26689 317 26723
rect 351 26689 430 26723
rect 245 26655 320 26689
rect 354 26655 430 26689
rect 245 26621 317 26655
rect 351 26621 430 26655
rect 245 26617 430 26621
rect 245 26587 320 26617
rect 245 26553 317 26587
rect 354 26583 430 26617
rect 351 26553 430 26583
rect 245 26545 430 26553
rect 245 26519 320 26545
rect 245 26485 317 26519
rect 354 26511 430 26545
rect 351 26485 430 26511
rect 245 26473 430 26485
rect 245 26451 320 26473
rect 245 26417 317 26451
rect 354 26439 430 26473
rect 351 26417 430 26439
rect 245 26401 430 26417
rect 245 26383 320 26401
rect 245 26349 317 26383
rect 354 26367 430 26401
rect 351 26349 430 26367
rect 245 26329 430 26349
rect 245 26315 320 26329
rect 245 26281 317 26315
rect 354 26295 430 26329
rect 351 26281 430 26295
rect 245 26257 430 26281
rect 245 26247 320 26257
rect 245 26213 317 26247
rect 354 26223 430 26257
rect 351 26213 430 26223
rect 245 26185 430 26213
rect 245 26179 320 26185
rect 245 26145 317 26179
rect 354 26151 430 26185
rect 351 26145 430 26151
rect 245 26113 430 26145
rect 245 26111 320 26113
rect 245 26077 317 26111
rect 354 26079 430 26113
rect 351 26077 430 26079
rect 245 26043 430 26077
rect 245 26009 317 26043
rect 351 26041 430 26043
rect 245 26007 320 26009
rect 354 26007 430 26041
rect 245 25975 430 26007
rect 245 25941 317 25975
rect 351 25969 430 25975
rect 245 25935 320 25941
rect 354 25935 430 25969
rect 245 25907 430 25935
rect 245 25873 317 25907
rect 351 25897 430 25907
rect 245 25863 320 25873
rect 354 25863 430 25897
rect 245 25839 430 25863
rect 245 25805 317 25839
rect 351 25825 430 25839
rect 245 25791 320 25805
rect 354 25791 430 25825
rect 245 25771 430 25791
rect 245 25737 317 25771
rect 351 25753 430 25771
rect 245 25719 320 25737
rect 354 25719 430 25753
rect 245 25703 430 25719
rect 245 25669 317 25703
rect 351 25681 430 25703
rect 245 25647 320 25669
rect 354 25647 430 25681
rect 245 25635 430 25647
rect 245 25601 317 25635
rect 351 25609 430 25635
rect 245 25575 320 25601
rect 354 25575 430 25609
rect 245 25567 430 25575
rect 245 25533 317 25567
rect 351 25537 430 25567
rect 245 25503 320 25533
rect 354 25503 430 25537
rect 245 25499 430 25503
rect 245 25465 317 25499
rect 351 25465 430 25499
rect 245 25431 320 25465
rect 354 25431 430 25465
rect 245 25397 317 25431
rect 351 25397 430 25431
rect 245 25393 430 25397
rect 245 25363 320 25393
rect 245 25329 317 25363
rect 354 25359 430 25393
rect 351 25329 430 25359
rect 245 25321 430 25329
rect 245 25295 320 25321
rect 245 25261 317 25295
rect 354 25287 430 25321
rect 351 25261 430 25287
rect 245 25249 430 25261
rect 245 25227 320 25249
rect 245 25193 317 25227
rect 354 25215 430 25249
rect 351 25193 430 25215
rect 245 25177 430 25193
rect 245 25159 320 25177
rect 245 25125 317 25159
rect 354 25143 430 25177
rect 351 25125 430 25143
rect 245 25105 430 25125
rect 245 25091 320 25105
rect 245 25057 317 25091
rect 354 25071 430 25105
rect 351 25057 430 25071
rect 245 25033 430 25057
rect 245 25023 320 25033
rect 245 24989 317 25023
rect 354 24999 430 25033
rect 351 24989 430 24999
rect 245 24961 430 24989
rect 245 24955 320 24961
rect 245 24921 317 24955
rect 354 24927 430 24961
rect 351 24921 430 24927
rect 245 24889 430 24921
rect 245 24887 320 24889
rect 245 24853 317 24887
rect 354 24855 430 24889
rect 351 24853 430 24855
rect 245 24819 430 24853
rect 245 24785 317 24819
rect 351 24817 430 24819
rect 245 24783 320 24785
rect 354 24783 430 24817
rect 245 24751 430 24783
rect 245 24717 317 24751
rect 351 24745 430 24751
rect 245 24711 320 24717
rect 354 24711 430 24745
rect 245 24683 430 24711
rect 245 24649 317 24683
rect 351 24673 430 24683
rect 245 24639 320 24649
rect 354 24639 430 24673
rect 245 24615 430 24639
rect 245 24581 317 24615
rect 351 24601 430 24615
rect 245 24567 320 24581
rect 354 24567 430 24601
rect 245 24547 430 24567
rect 245 24513 317 24547
rect 351 24529 430 24547
rect 245 24495 320 24513
rect 354 24495 430 24529
rect 245 24479 430 24495
rect 245 24445 317 24479
rect 351 24457 430 24479
rect 245 24423 320 24445
rect 354 24423 430 24457
rect 245 24411 430 24423
rect 245 24377 317 24411
rect 351 24385 430 24411
rect 245 24351 320 24377
rect 354 24351 430 24385
rect 245 24343 430 24351
rect 245 24309 317 24343
rect 351 24313 430 24343
rect 245 24279 320 24309
rect 354 24279 430 24313
rect 245 24275 430 24279
rect 245 24241 317 24275
rect 351 24241 430 24275
rect 245 24207 320 24241
rect 354 24207 430 24241
rect 245 24173 317 24207
rect 351 24173 430 24207
rect 245 24169 430 24173
rect 245 24139 320 24169
rect 245 24105 317 24139
rect 354 24135 430 24169
rect 351 24105 430 24135
rect 245 24097 430 24105
rect 245 24071 320 24097
rect 245 24037 317 24071
rect 354 24063 430 24097
rect 351 24037 430 24063
rect 245 24025 430 24037
rect 245 24003 320 24025
rect 245 23969 317 24003
rect 354 23991 430 24025
rect 351 23969 430 23991
rect 245 23953 430 23969
rect 245 23935 320 23953
rect 245 23901 317 23935
rect 354 23919 430 23953
rect 351 23901 430 23919
rect 245 23881 430 23901
rect 245 23867 320 23881
rect 245 23833 317 23867
rect 354 23847 430 23881
rect 351 23833 430 23847
rect 245 23809 430 23833
rect 245 23799 320 23809
rect 245 23765 317 23799
rect 354 23775 430 23809
rect 351 23765 430 23775
rect 245 23737 430 23765
rect 245 23731 320 23737
rect 245 23697 317 23731
rect 354 23703 430 23737
rect 351 23697 430 23703
rect 245 23665 430 23697
rect 245 23663 320 23665
rect 245 23629 317 23663
rect 354 23631 430 23665
rect 351 23629 430 23631
rect 245 23595 430 23629
rect 245 23561 317 23595
rect 351 23593 430 23595
rect 245 23559 320 23561
rect 354 23559 430 23593
rect 245 23527 430 23559
rect 245 23493 317 23527
rect 351 23521 430 23527
rect 245 23487 320 23493
rect 354 23487 430 23521
rect 245 23459 430 23487
rect 245 23425 317 23459
rect 351 23449 430 23459
rect 245 23415 320 23425
rect 354 23415 430 23449
rect 245 23391 430 23415
rect 245 23357 317 23391
rect 351 23377 430 23391
rect 245 23343 320 23357
rect 354 23343 430 23377
rect 245 23323 430 23343
rect 245 23289 317 23323
rect 351 23305 430 23323
rect 245 23271 320 23289
rect 354 23271 430 23305
rect 245 23255 430 23271
rect 245 23221 317 23255
rect 351 23233 430 23255
rect 245 23199 320 23221
rect 354 23199 430 23233
rect 245 23187 430 23199
rect 245 23153 317 23187
rect 351 23161 430 23187
rect 245 23127 320 23153
rect 354 23127 430 23161
rect 245 23119 430 23127
rect 245 23085 317 23119
rect 351 23089 430 23119
rect 245 23055 320 23085
rect 354 23055 430 23089
rect 245 23051 430 23055
rect 245 23017 317 23051
rect 351 23017 430 23051
rect 245 22983 320 23017
rect 354 22983 430 23017
rect 245 22949 317 22983
rect 351 22949 430 22983
rect 245 22945 430 22949
rect 245 22915 320 22945
rect 245 22881 317 22915
rect 354 22911 430 22945
rect 351 22881 430 22911
rect 245 22873 430 22881
rect 245 22847 320 22873
rect 245 22813 317 22847
rect 354 22839 430 22873
rect 351 22813 430 22839
rect 245 22801 430 22813
rect 245 22779 320 22801
rect 245 22745 317 22779
rect 354 22767 430 22801
rect 351 22745 430 22767
rect 245 22729 430 22745
rect 245 22711 320 22729
rect 245 22677 317 22711
rect 354 22695 430 22729
rect 351 22677 430 22695
rect 245 22657 430 22677
rect 245 22643 320 22657
rect 245 22609 317 22643
rect 354 22623 430 22657
rect 351 22609 430 22623
rect 245 22585 430 22609
rect 245 22575 320 22585
rect 245 22541 317 22575
rect 354 22551 430 22585
rect 351 22541 430 22551
rect 245 22513 430 22541
rect 245 22507 320 22513
rect 245 22473 317 22507
rect 354 22479 430 22513
rect 351 22473 430 22479
rect 245 22441 430 22473
rect 245 22439 320 22441
rect 245 22405 317 22439
rect 354 22407 430 22441
rect 351 22405 430 22407
rect 245 22371 430 22405
rect 245 22337 317 22371
rect 351 22369 430 22371
rect 245 22335 320 22337
rect 354 22335 430 22369
rect 245 22303 430 22335
rect 245 22269 317 22303
rect 351 22297 430 22303
rect 245 22263 320 22269
rect 354 22263 430 22297
rect 245 22235 430 22263
rect 245 22201 317 22235
rect 351 22225 430 22235
rect 245 22191 320 22201
rect 354 22191 430 22225
rect 245 22167 430 22191
rect 245 22133 317 22167
rect 351 22153 430 22167
rect 245 22119 320 22133
rect 354 22119 430 22153
rect 245 22099 430 22119
rect 245 22065 317 22099
rect 351 22081 430 22099
rect 245 22047 320 22065
rect 354 22047 430 22081
rect 245 22031 430 22047
rect 245 21997 317 22031
rect 351 22009 430 22031
rect 245 21975 320 21997
rect 354 21975 430 22009
rect 245 21963 430 21975
rect 245 21929 317 21963
rect 351 21937 430 21963
rect 245 21903 320 21929
rect 354 21903 430 21937
rect 245 21895 430 21903
rect 245 21861 317 21895
rect 351 21865 430 21895
rect 245 21831 320 21861
rect 354 21831 430 21865
rect 245 21827 430 21831
rect 245 21793 317 21827
rect 351 21793 430 21827
rect 245 21759 320 21793
rect 354 21759 430 21793
rect 245 21725 317 21759
rect 351 21725 430 21759
rect 245 21721 430 21725
rect 245 21691 320 21721
rect 245 21657 317 21691
rect 354 21687 430 21721
rect 351 21657 430 21687
rect 245 21649 430 21657
rect 245 21623 320 21649
rect 245 21589 317 21623
rect 354 21615 430 21649
rect 351 21589 430 21615
rect 245 21577 430 21589
rect 245 21555 320 21577
rect 245 21521 317 21555
rect 354 21543 430 21577
rect 351 21521 430 21543
rect 245 21505 430 21521
rect 245 21487 320 21505
rect 245 21453 317 21487
rect 354 21471 430 21505
rect 351 21453 430 21471
rect 245 21433 430 21453
rect 245 21419 320 21433
rect 245 21385 317 21419
rect 354 21399 430 21433
rect 351 21385 430 21399
rect 245 21361 430 21385
rect 245 21351 320 21361
rect 245 21317 317 21351
rect 354 21327 430 21361
rect 351 21317 430 21327
rect 245 21289 430 21317
rect 245 21283 320 21289
rect 245 21249 317 21283
rect 354 21255 430 21289
rect 351 21249 430 21255
rect 245 21217 430 21249
rect 245 21215 320 21217
rect 245 21181 317 21215
rect 354 21183 430 21217
rect 351 21181 430 21183
rect 245 21147 430 21181
rect 245 21113 317 21147
rect 351 21145 430 21147
rect 245 21111 320 21113
rect 354 21111 430 21145
rect 245 21079 430 21111
rect 245 21045 317 21079
rect 351 21073 430 21079
rect 245 21039 320 21045
rect 354 21039 430 21073
rect 245 21011 430 21039
rect 245 20977 317 21011
rect 351 21001 430 21011
rect 245 20967 320 20977
rect 354 20967 430 21001
rect 245 20943 430 20967
rect 245 20909 317 20943
rect 351 20929 430 20943
rect 245 20895 320 20909
rect 354 20895 430 20929
rect 245 20875 430 20895
rect 245 20841 317 20875
rect 351 20857 430 20875
rect 245 20823 320 20841
rect 354 20823 430 20857
rect 245 20807 430 20823
rect 245 20773 317 20807
rect 351 20785 430 20807
rect 245 20751 320 20773
rect 354 20751 430 20785
rect 245 20739 430 20751
rect 245 20705 317 20739
rect 351 20713 430 20739
rect 245 20679 320 20705
rect 354 20679 430 20713
rect 245 20671 430 20679
rect 245 20637 317 20671
rect 351 20641 430 20671
rect 245 20607 320 20637
rect 354 20607 430 20641
rect 245 20603 430 20607
rect 245 20569 317 20603
rect 351 20569 430 20603
rect 245 20535 320 20569
rect 354 20535 430 20569
rect 245 20501 317 20535
rect 351 20501 430 20535
rect 245 20497 430 20501
rect 245 20467 320 20497
rect 245 20433 317 20467
rect 354 20463 430 20497
rect 351 20433 430 20463
rect 245 20425 430 20433
rect 245 20399 320 20425
rect 245 20365 317 20399
rect 354 20391 430 20425
rect 351 20365 430 20391
rect 245 20353 430 20365
rect 245 20331 320 20353
rect 245 20297 317 20331
rect 354 20319 430 20353
rect 351 20297 430 20319
rect 245 20281 430 20297
rect 245 20263 320 20281
rect 245 20229 317 20263
rect 354 20247 430 20281
rect 351 20229 430 20247
rect 245 20209 430 20229
rect 245 20195 320 20209
rect 245 20161 317 20195
rect 354 20175 430 20209
rect 351 20161 430 20175
rect 245 20137 430 20161
rect 245 20127 320 20137
rect 245 20093 317 20127
rect 354 20103 430 20137
rect 351 20093 430 20103
rect 245 20065 430 20093
rect 245 20059 320 20065
rect 245 20025 317 20059
rect 354 20031 430 20065
rect 351 20025 430 20031
rect 245 19993 430 20025
rect 245 19991 320 19993
rect 245 19957 317 19991
rect 354 19959 430 19993
rect 351 19957 430 19959
rect 245 19923 430 19957
rect 245 19889 317 19923
rect 351 19921 430 19923
rect 245 19887 320 19889
rect 354 19887 430 19921
rect 245 19855 430 19887
rect 245 19821 317 19855
rect 351 19849 430 19855
rect 245 19815 320 19821
rect 354 19815 430 19849
rect 245 19787 430 19815
rect 245 19753 317 19787
rect 351 19777 430 19787
rect 245 19743 320 19753
rect 354 19743 430 19777
rect 245 19719 430 19743
rect 245 19685 317 19719
rect 351 19705 430 19719
rect 245 19671 320 19685
rect 354 19671 430 19705
rect 245 19651 430 19671
rect 245 19617 317 19651
rect 351 19633 430 19651
rect 245 19599 320 19617
rect 354 19599 430 19633
rect 245 19583 430 19599
rect 245 19549 317 19583
rect 351 19561 430 19583
rect 245 19527 320 19549
rect 354 19527 430 19561
rect 245 19515 430 19527
rect 245 19481 317 19515
rect 351 19489 430 19515
rect 245 19455 320 19481
rect 354 19455 430 19489
rect 245 19447 430 19455
rect 245 19413 317 19447
rect 351 19417 430 19447
rect 245 19383 320 19413
rect 354 19383 430 19417
rect 245 19379 430 19383
rect 245 19345 317 19379
rect 351 19345 430 19379
rect 245 19311 320 19345
rect 354 19311 430 19345
rect 245 19277 317 19311
rect 351 19277 430 19311
rect 245 19273 430 19277
rect 245 19243 320 19273
rect 245 19209 317 19243
rect 354 19239 430 19273
rect 351 19209 430 19239
rect 245 19201 430 19209
rect 245 19175 320 19201
rect 245 19141 317 19175
rect 354 19167 430 19201
rect 351 19141 430 19167
rect 245 19129 430 19141
rect 245 19107 320 19129
rect 245 19073 317 19107
rect 354 19095 430 19129
rect 351 19073 430 19095
rect 245 19057 430 19073
rect 245 19039 320 19057
rect 245 19005 317 19039
rect 354 19023 430 19057
rect 351 19005 430 19023
rect 245 18985 430 19005
rect 245 18971 320 18985
rect 245 18937 317 18971
rect 354 18951 430 18985
rect 351 18937 430 18951
rect 245 18913 430 18937
rect 245 18903 320 18913
rect 245 18869 317 18903
rect 354 18879 430 18913
rect 351 18869 430 18879
rect 245 18841 430 18869
rect 245 18835 320 18841
rect 245 18801 317 18835
rect 354 18807 430 18841
rect 351 18801 430 18807
rect 245 18769 430 18801
rect 245 18767 320 18769
rect 245 18733 317 18767
rect 354 18735 430 18769
rect 351 18733 430 18735
rect 245 18699 430 18733
rect 245 18665 317 18699
rect 351 18697 430 18699
rect 245 18663 320 18665
rect 354 18663 430 18697
rect 245 18631 430 18663
rect 245 18597 317 18631
rect 351 18625 430 18631
rect 245 18591 320 18597
rect 354 18591 430 18625
rect 245 18563 430 18591
rect 245 18529 317 18563
rect 351 18553 430 18563
rect 245 18519 320 18529
rect 354 18519 430 18553
rect 245 18495 430 18519
rect 245 18461 317 18495
rect 351 18481 430 18495
rect 245 18447 320 18461
rect 354 18447 430 18481
rect 245 18427 430 18447
rect 245 18393 317 18427
rect 351 18409 430 18427
rect 245 18375 320 18393
rect 354 18375 430 18409
rect 245 18359 430 18375
rect 245 18325 317 18359
rect 351 18337 430 18359
rect 245 18303 320 18325
rect 354 18303 430 18337
rect 245 18291 430 18303
rect 245 18257 317 18291
rect 351 18265 430 18291
rect 245 18231 320 18257
rect 354 18231 430 18265
rect 245 18223 430 18231
rect 245 18189 317 18223
rect 351 18193 430 18223
rect 245 18159 320 18189
rect 354 18159 430 18193
rect 245 18155 430 18159
rect 245 18121 317 18155
rect 351 18121 430 18155
rect 245 18087 320 18121
rect 354 18087 430 18121
rect 245 18053 317 18087
rect 351 18053 430 18087
rect 245 18049 430 18053
rect 245 18019 320 18049
rect 245 17985 317 18019
rect 354 18015 430 18049
rect 351 17985 430 18015
rect 245 17977 430 17985
rect 245 17951 320 17977
rect 245 17917 317 17951
rect 354 17943 430 17977
rect 351 17917 430 17943
rect 245 17905 430 17917
rect 245 17883 320 17905
rect 245 17849 317 17883
rect 354 17871 430 17905
rect 351 17849 430 17871
rect 245 17833 430 17849
rect 245 17815 320 17833
rect 245 17781 317 17815
rect 354 17799 430 17833
rect 351 17781 430 17799
rect 245 17761 430 17781
rect 245 17747 320 17761
rect 245 17713 317 17747
rect 354 17727 430 17761
rect 351 17713 430 17727
rect 245 17689 430 17713
rect 245 17679 320 17689
rect 245 17645 317 17679
rect 354 17655 430 17689
rect 351 17645 430 17655
rect 245 17617 430 17645
rect 245 17611 320 17617
rect 245 17577 317 17611
rect 354 17583 430 17617
rect 351 17577 430 17583
rect 245 17545 430 17577
rect 245 17543 320 17545
rect 245 17509 317 17543
rect 354 17511 430 17545
rect 351 17509 430 17511
rect 245 17475 430 17509
rect 245 17441 317 17475
rect 351 17473 430 17475
rect 245 17439 320 17441
rect 354 17439 430 17473
rect 245 17407 430 17439
rect 245 17373 317 17407
rect 351 17401 430 17407
rect 245 17367 320 17373
rect 354 17367 430 17401
rect 245 17339 430 17367
rect 245 17305 317 17339
rect 351 17329 430 17339
rect 245 17295 320 17305
rect 354 17295 430 17329
rect 245 17271 430 17295
rect 245 17237 317 17271
rect 351 17257 430 17271
rect 245 17223 320 17237
rect 354 17223 430 17257
rect 245 17203 430 17223
rect 245 17169 317 17203
rect 351 17185 430 17203
rect 245 17151 320 17169
rect 354 17151 430 17185
rect 245 17135 430 17151
rect 245 17101 317 17135
rect 351 17113 430 17135
rect 245 17079 320 17101
rect 354 17079 430 17113
rect 245 17067 430 17079
rect 245 17033 317 17067
rect 351 17041 430 17067
rect 245 17007 320 17033
rect 354 17007 430 17041
rect 245 16999 430 17007
rect 245 16965 317 16999
rect 351 16969 430 16999
rect 245 16935 320 16965
rect 354 16935 430 16969
rect 245 16931 430 16935
rect 245 16897 317 16931
rect 351 16897 430 16931
rect 245 16863 320 16897
rect 354 16863 430 16897
rect 245 16829 317 16863
rect 351 16829 430 16863
rect 245 16825 430 16829
rect 245 16795 320 16825
rect 245 16761 317 16795
rect 354 16791 430 16825
rect 351 16761 430 16791
rect 245 16753 430 16761
rect 245 16727 320 16753
rect 245 16693 317 16727
rect 354 16719 430 16753
rect 351 16693 430 16719
rect 245 16681 430 16693
rect 245 16659 320 16681
rect 245 16625 317 16659
rect 354 16647 430 16681
rect 351 16625 430 16647
rect 245 16609 430 16625
rect 245 16591 320 16609
rect 245 16557 317 16591
rect 354 16575 430 16609
rect 351 16557 430 16575
rect 245 16537 430 16557
rect 245 16523 320 16537
rect 245 16489 317 16523
rect 354 16503 430 16537
rect 351 16489 430 16503
rect 245 16465 430 16489
rect 245 16455 320 16465
rect 245 16421 317 16455
rect 354 16431 430 16465
rect 351 16421 430 16431
rect 245 16393 430 16421
rect 245 16387 320 16393
rect 245 16353 317 16387
rect 354 16359 430 16393
rect 351 16353 430 16359
rect 245 16321 430 16353
rect 245 16319 320 16321
rect 245 16285 317 16319
rect 354 16287 430 16321
rect 351 16285 430 16287
rect 245 16251 430 16285
rect 245 16217 317 16251
rect 351 16249 430 16251
rect 245 16215 320 16217
rect 354 16215 430 16249
rect 245 16183 430 16215
rect 245 16149 317 16183
rect 351 16177 430 16183
rect 245 16143 320 16149
rect 354 16143 430 16177
rect 245 16115 430 16143
rect 245 16081 317 16115
rect 351 16105 430 16115
rect 245 16071 320 16081
rect 354 16071 430 16105
rect 245 16047 430 16071
rect 245 16013 317 16047
rect 351 16033 430 16047
rect 245 15999 320 16013
rect 354 15999 430 16033
rect 245 15979 430 15999
rect 245 15945 317 15979
rect 351 15961 430 15979
rect 245 15927 320 15945
rect 354 15927 430 15961
rect 245 15911 430 15927
rect 245 15877 317 15911
rect 351 15889 430 15911
rect 245 15855 320 15877
rect 354 15855 430 15889
rect 245 15843 430 15855
rect 245 15809 317 15843
rect 351 15817 430 15843
rect 245 15783 320 15809
rect 354 15783 430 15817
rect 245 15775 430 15783
rect 245 15741 317 15775
rect 351 15745 430 15775
rect 245 15711 320 15741
rect 354 15711 430 15745
rect 245 15707 430 15711
rect 245 15673 317 15707
rect 351 15673 430 15707
rect 245 15639 320 15673
rect 354 15639 430 15673
rect 245 15605 317 15639
rect 351 15605 430 15639
rect 245 15601 430 15605
rect 245 15571 320 15601
rect 245 15537 317 15571
rect 354 15567 430 15601
rect 351 15537 430 15567
rect 245 15529 430 15537
rect 245 15503 320 15529
rect 245 15469 317 15503
rect 354 15495 430 15529
rect 351 15469 430 15495
rect 245 15457 430 15469
rect 245 15435 320 15457
rect 245 15401 317 15435
rect 354 15423 430 15457
rect 351 15401 430 15423
rect 245 15385 430 15401
rect 245 15367 320 15385
rect 245 15333 317 15367
rect 354 15351 430 15385
rect 351 15333 430 15351
rect 245 15313 430 15333
rect 245 15299 320 15313
rect 245 15265 317 15299
rect 354 15279 430 15313
rect 351 15265 430 15279
rect 245 15241 430 15265
rect 245 15231 320 15241
rect 245 15197 317 15231
rect 354 15207 430 15241
rect 351 15197 430 15207
rect 245 15169 430 15197
rect 245 15163 320 15169
rect 245 15129 317 15163
rect 354 15135 430 15169
rect 351 15129 430 15135
rect 245 15097 430 15129
rect 245 15095 320 15097
rect 245 15061 317 15095
rect 354 15063 430 15097
rect 351 15061 430 15063
rect 245 15027 430 15061
rect 245 14993 317 15027
rect 351 15025 430 15027
rect 245 14991 320 14993
rect 354 14991 430 15025
rect 245 14959 430 14991
rect 245 14925 317 14959
rect 351 14953 430 14959
rect 245 14919 320 14925
rect 354 14919 430 14953
rect 245 14891 430 14919
rect 245 14857 317 14891
rect 351 14881 430 14891
rect 245 14847 320 14857
rect 354 14847 430 14881
rect 245 14823 430 14847
rect 245 14789 317 14823
rect 351 14809 430 14823
rect 245 14775 320 14789
rect 354 14775 430 14809
rect 245 14755 430 14775
rect 245 14721 317 14755
rect 351 14737 430 14755
rect 245 14703 320 14721
rect 354 14703 430 14737
rect 245 14687 430 14703
rect 245 14653 317 14687
rect 351 14665 430 14687
rect 245 14631 320 14653
rect 354 14631 430 14665
rect 245 14619 430 14631
rect 245 14585 317 14619
rect 351 14593 430 14619
rect 245 14559 320 14585
rect 354 14559 430 14593
rect 245 14551 430 14559
rect 245 14517 317 14551
rect 351 14521 430 14551
rect 245 14487 320 14517
rect 354 14487 430 14521
rect 245 14483 430 14487
rect 245 14449 317 14483
rect 351 14449 430 14483
rect 245 14415 320 14449
rect 354 14415 430 14449
rect 245 14381 317 14415
rect 351 14381 430 14415
rect 245 14377 430 14381
rect 245 14347 320 14377
rect 245 14313 317 14347
rect 354 14343 430 14377
rect 351 14313 430 14343
rect 245 14305 430 14313
rect 245 14279 320 14305
rect 245 14245 317 14279
rect 354 14271 430 14305
rect 351 14245 430 14271
rect 245 14233 430 14245
rect 245 14211 320 14233
rect 245 14177 317 14211
rect 354 14199 430 14233
rect 351 14177 430 14199
rect 245 14161 430 14177
rect 245 14143 320 14161
rect 245 14109 317 14143
rect 354 14127 430 14161
rect 351 14109 430 14127
rect 245 14089 430 14109
rect 245 14075 320 14089
rect 245 14041 317 14075
rect 354 14055 430 14089
rect 351 14041 430 14055
rect 245 14017 430 14041
rect 245 14007 320 14017
rect 245 13973 317 14007
rect 354 13983 430 14017
rect 351 13973 430 13983
rect 245 13945 430 13973
rect 245 13939 320 13945
rect 245 13905 317 13939
rect 354 13911 430 13945
rect 351 13905 430 13911
rect 245 13873 430 13905
rect 245 13871 320 13873
rect 245 13837 317 13871
rect 354 13839 430 13873
rect 351 13837 430 13839
rect 245 13803 430 13837
rect 245 13769 317 13803
rect 351 13801 430 13803
rect 245 13767 320 13769
rect 354 13767 430 13801
rect 245 13735 430 13767
rect 245 13701 317 13735
rect 351 13729 430 13735
rect 245 13695 320 13701
rect 354 13695 430 13729
rect 245 13667 430 13695
rect 245 13633 317 13667
rect 351 13657 430 13667
rect 245 13623 320 13633
rect 354 13623 430 13657
rect 245 13599 430 13623
rect 245 13565 317 13599
rect 351 13585 430 13599
rect 245 13551 320 13565
rect 354 13551 430 13585
rect 245 13531 430 13551
rect 245 13497 317 13531
rect 351 13513 430 13531
rect 245 13479 320 13497
rect 354 13479 430 13513
rect 245 13463 430 13479
rect 245 13429 317 13463
rect 351 13441 430 13463
rect 245 13407 320 13429
rect 354 13407 430 13441
rect 245 13395 430 13407
rect 245 13361 317 13395
rect 351 13369 430 13395
rect 245 13335 320 13361
rect 354 13335 430 13369
rect 245 13327 430 13335
rect 245 13293 317 13327
rect 351 13297 430 13327
rect 245 13263 320 13293
rect 354 13263 430 13297
rect 245 13259 430 13263
rect 245 13225 317 13259
rect 351 13225 430 13259
rect 245 13191 320 13225
rect 354 13191 430 13225
rect 245 13157 317 13191
rect 351 13157 430 13191
rect 245 13153 430 13157
rect 245 13123 320 13153
rect 245 13089 317 13123
rect 354 13119 430 13153
rect 351 13089 430 13119
rect 245 13081 430 13089
rect 245 13055 320 13081
rect 245 13021 317 13055
rect 354 13047 430 13081
rect 351 13021 430 13047
rect 245 13009 430 13021
rect 245 12987 320 13009
rect 245 12953 317 12987
rect 354 12975 430 13009
rect 351 12953 430 12975
rect 245 12937 430 12953
rect 245 12919 320 12937
rect 245 12885 317 12919
rect 354 12903 430 12937
rect 351 12885 430 12903
rect 245 12865 430 12885
rect 245 12851 320 12865
rect 245 12817 317 12851
rect 354 12831 430 12865
rect 351 12817 430 12831
rect 245 12793 430 12817
rect 245 12783 320 12793
rect 245 12749 317 12783
rect 354 12759 430 12793
rect 351 12749 430 12759
rect 245 12721 430 12749
rect 245 12715 320 12721
rect 245 12681 317 12715
rect 354 12687 430 12721
rect 351 12681 430 12687
rect 245 12649 430 12681
rect 245 12647 320 12649
rect 245 12613 317 12647
rect 354 12615 430 12649
rect 351 12613 430 12615
rect 245 12579 430 12613
rect 245 12545 317 12579
rect 351 12577 430 12579
rect 245 12543 320 12545
rect 354 12543 430 12577
rect 245 12511 430 12543
rect 245 12477 317 12511
rect 351 12505 430 12511
rect 245 12471 320 12477
rect 354 12471 430 12505
rect 245 12443 430 12471
rect 245 12409 317 12443
rect 351 12433 430 12443
rect 245 12399 320 12409
rect 354 12399 430 12433
rect 245 12375 430 12399
rect 245 12341 317 12375
rect 351 12361 430 12375
rect 245 12327 320 12341
rect 354 12327 430 12361
rect 245 12307 430 12327
rect 245 12273 317 12307
rect 351 12289 430 12307
rect 245 12255 320 12273
rect 354 12255 430 12289
rect 245 12239 430 12255
rect 245 12205 317 12239
rect 351 12217 430 12239
rect 245 12183 320 12205
rect 354 12183 430 12217
rect 245 12171 430 12183
rect 245 12137 317 12171
rect 351 12145 430 12171
rect 245 12111 320 12137
rect 354 12111 430 12145
rect 245 12103 430 12111
rect 245 12069 317 12103
rect 351 12073 430 12103
rect 245 12039 320 12069
rect 354 12039 430 12073
rect 245 12035 430 12039
rect 245 12001 317 12035
rect 351 12001 430 12035
rect 245 11967 320 12001
rect 354 11967 430 12001
rect 245 11933 317 11967
rect 351 11933 430 11967
rect 245 11929 430 11933
rect 245 11899 320 11929
rect 245 11865 317 11899
rect 354 11895 430 11929
rect 351 11865 430 11895
rect 245 11857 430 11865
rect 245 11831 320 11857
rect 245 11797 317 11831
rect 354 11823 430 11857
rect 351 11797 430 11823
rect 245 11785 430 11797
rect 245 11763 320 11785
rect 245 11729 317 11763
rect 354 11751 430 11785
rect 351 11729 430 11751
rect 245 11713 430 11729
rect 245 11695 320 11713
rect 245 11661 317 11695
rect 354 11679 430 11713
rect 351 11661 430 11679
rect 245 11641 430 11661
rect 245 11627 320 11641
rect 245 11593 317 11627
rect 354 11607 430 11641
rect 351 11593 430 11607
rect 245 11569 430 11593
rect 245 11559 320 11569
rect 245 11525 317 11559
rect 354 11535 430 11569
rect 351 11525 430 11535
rect 245 11497 430 11525
rect 245 11491 320 11497
rect 245 11457 317 11491
rect 354 11463 430 11497
rect 351 11457 430 11463
rect 245 11425 430 11457
rect 245 11423 320 11425
rect 245 11389 317 11423
rect 354 11391 430 11425
rect 351 11389 430 11391
rect 245 11355 430 11389
rect 245 11321 317 11355
rect 351 11353 430 11355
rect 245 11319 320 11321
rect 354 11319 430 11353
rect 245 11287 430 11319
rect 245 11253 317 11287
rect 351 11281 430 11287
rect 245 11247 320 11253
rect 354 11247 430 11281
rect 245 11219 430 11247
rect 245 11185 317 11219
rect 351 11209 430 11219
rect 245 11175 320 11185
rect 354 11175 430 11209
rect 245 11151 430 11175
rect 245 11117 317 11151
rect 351 11137 430 11151
rect 245 11103 320 11117
rect 354 11103 430 11137
rect 245 11083 430 11103
rect 245 11049 317 11083
rect 351 11065 430 11083
rect 245 11031 320 11049
rect 354 11031 430 11065
rect 245 11015 430 11031
rect 245 10981 317 11015
rect 351 10993 430 11015
rect 245 10959 320 10981
rect 354 10959 430 10993
rect 245 10947 430 10959
rect 245 10913 317 10947
rect 351 10921 430 10947
rect 245 10887 320 10913
rect 354 10887 430 10921
rect 245 10879 430 10887
rect 245 10845 317 10879
rect 351 10849 430 10879
rect 245 10815 320 10845
rect 354 10815 430 10849
rect 245 10811 430 10815
rect 245 10777 317 10811
rect 351 10777 430 10811
rect 245 10743 320 10777
rect 354 10743 430 10777
rect 245 10709 317 10743
rect 351 10709 430 10743
rect 245 10705 430 10709
rect 245 10675 320 10705
rect 245 10641 317 10675
rect 354 10671 430 10705
rect 351 10641 430 10671
rect 245 10633 430 10641
rect 245 10607 320 10633
rect 245 10573 317 10607
rect 354 10599 430 10633
rect 351 10573 430 10599
rect 245 10561 430 10573
rect 245 10539 320 10561
rect 245 10505 317 10539
rect 354 10527 430 10561
rect 351 10505 430 10527
rect 245 10489 430 10505
rect 245 10471 320 10489
rect 245 10437 317 10471
rect 354 10455 430 10489
rect 351 10437 430 10455
rect 245 10417 430 10437
rect 245 10403 320 10417
rect 245 10369 317 10403
rect 354 10383 430 10417
rect 351 10369 430 10383
rect 245 10345 430 10369
rect 245 10335 320 10345
rect 245 10301 317 10335
rect 354 10311 430 10345
rect 351 10301 430 10311
rect 245 10273 430 10301
rect 245 10267 320 10273
rect 245 10233 317 10267
rect 354 10239 430 10273
rect 351 10233 430 10239
rect 245 10201 430 10233
rect 245 10199 320 10201
rect 245 10165 317 10199
rect 354 10167 430 10201
rect 351 10165 430 10167
rect 245 10131 430 10165
rect 245 10097 317 10131
rect 351 10129 430 10131
rect 245 10095 320 10097
rect 354 10095 430 10129
rect 245 10063 430 10095
rect 245 10029 317 10063
rect 351 10057 430 10063
rect 245 10023 320 10029
rect 354 10023 430 10057
rect 245 9995 430 10023
rect 245 9961 317 9995
rect 351 9985 430 9995
rect 245 9951 320 9961
rect 354 9951 430 9985
rect 245 9927 430 9951
rect 245 9893 317 9927
rect 351 9913 430 9927
rect 245 9879 320 9893
rect 354 9879 430 9913
rect 245 9859 430 9879
rect 245 9825 317 9859
rect 351 9841 430 9859
rect 245 9807 320 9825
rect 354 9807 430 9841
rect 245 9791 430 9807
rect 245 9757 317 9791
rect 351 9769 430 9791
rect 245 9735 320 9757
rect 354 9735 430 9769
rect 245 9723 430 9735
rect 245 9689 317 9723
rect 351 9697 430 9723
rect 603 36177 14361 36207
rect 603 36143 766 36177
rect 800 36143 834 36177
rect 868 36143 902 36177
rect 936 36143 970 36177
rect 1004 36143 1038 36177
rect 1072 36143 1106 36177
rect 1140 36143 1174 36177
rect 1208 36143 1242 36177
rect 1276 36143 1310 36177
rect 1344 36143 1378 36177
rect 1412 36143 1446 36177
rect 1480 36143 1514 36177
rect 1548 36143 1582 36177
rect 1616 36143 1650 36177
rect 1684 36143 1718 36177
rect 1752 36143 1786 36177
rect 1820 36143 1854 36177
rect 1888 36143 1922 36177
rect 1956 36143 1990 36177
rect 2024 36143 2058 36177
rect 2092 36143 2126 36177
rect 2160 36143 2194 36177
rect 2228 36143 2262 36177
rect 2296 36143 2330 36177
rect 2364 36143 2398 36177
rect 2432 36143 2466 36177
rect 2500 36143 2534 36177
rect 2568 36143 2602 36177
rect 2636 36143 2670 36177
rect 2704 36143 2738 36177
rect 2772 36143 2806 36177
rect 2840 36143 2874 36177
rect 2908 36143 2942 36177
rect 2976 36143 3010 36177
rect 3044 36143 3078 36177
rect 3112 36143 3146 36177
rect 3180 36143 3214 36177
rect 3248 36143 3282 36177
rect 3316 36143 3350 36177
rect 3384 36143 3418 36177
rect 3452 36143 3486 36177
rect 3520 36143 3554 36177
rect 3588 36143 3622 36177
rect 3656 36143 3690 36177
rect 3724 36143 3758 36177
rect 3792 36143 3826 36177
rect 3860 36143 3894 36177
rect 3928 36143 3962 36177
rect 3996 36143 4030 36177
rect 4064 36143 4098 36177
rect 4132 36143 4166 36177
rect 4200 36143 4234 36177
rect 4268 36143 4302 36177
rect 4336 36143 4370 36177
rect 4404 36143 4438 36177
rect 4472 36143 4506 36177
rect 4540 36143 4574 36177
rect 4608 36143 4642 36177
rect 4676 36143 4710 36177
rect 4744 36143 4778 36177
rect 4812 36143 4846 36177
rect 4880 36143 4914 36177
rect 4948 36143 4982 36177
rect 5016 36143 5050 36177
rect 5084 36143 5118 36177
rect 5152 36143 5186 36177
rect 5220 36143 5254 36177
rect 5288 36143 5322 36177
rect 5356 36143 5390 36177
rect 5424 36143 5458 36177
rect 5492 36143 5526 36177
rect 5560 36143 5594 36177
rect 5628 36143 5662 36177
rect 5696 36143 5730 36177
rect 5764 36143 5798 36177
rect 5832 36143 5866 36177
rect 5900 36143 5934 36177
rect 5968 36143 6002 36177
rect 6036 36143 6070 36177
rect 6104 36143 6138 36177
rect 6172 36143 6206 36177
rect 6240 36143 6274 36177
rect 6308 36143 6342 36177
rect 6376 36143 6410 36177
rect 6444 36143 6478 36177
rect 6512 36143 6546 36177
rect 6580 36143 6614 36177
rect 6648 36143 6682 36177
rect 6716 36143 6750 36177
rect 6784 36143 6818 36177
rect 6852 36143 6886 36177
rect 6920 36143 6954 36177
rect 6988 36143 7022 36177
rect 7056 36143 7090 36177
rect 7124 36143 7158 36177
rect 7192 36143 7226 36177
rect 7260 36143 7294 36177
rect 7328 36143 7362 36177
rect 7396 36143 7430 36177
rect 7464 36143 7498 36177
rect 7532 36143 7566 36177
rect 7600 36143 7634 36177
rect 7668 36143 7702 36177
rect 7736 36143 7770 36177
rect 7804 36143 7838 36177
rect 7872 36143 7906 36177
rect 7940 36143 7974 36177
rect 8008 36143 8042 36177
rect 8076 36143 8110 36177
rect 8144 36143 8178 36177
rect 8212 36143 8246 36177
rect 8280 36143 8314 36177
rect 8348 36143 8382 36177
rect 8416 36143 8450 36177
rect 8484 36143 8518 36177
rect 8552 36143 8586 36177
rect 8620 36143 8654 36177
rect 8688 36143 8722 36177
rect 8756 36143 8790 36177
rect 8824 36143 8858 36177
rect 8892 36143 8926 36177
rect 8960 36143 8994 36177
rect 9028 36143 9062 36177
rect 9096 36143 9130 36177
rect 9164 36143 9198 36177
rect 9232 36143 9266 36177
rect 9300 36143 9334 36177
rect 9368 36143 9402 36177
rect 9436 36143 9470 36177
rect 9504 36143 9538 36177
rect 9572 36143 9606 36177
rect 9640 36143 9674 36177
rect 9708 36143 9742 36177
rect 9776 36143 9810 36177
rect 9844 36143 9878 36177
rect 9912 36143 9946 36177
rect 9980 36143 10014 36177
rect 10048 36143 10082 36177
rect 10116 36143 10150 36177
rect 10184 36143 10218 36177
rect 10252 36143 10286 36177
rect 10320 36143 10354 36177
rect 10388 36143 10422 36177
rect 10456 36143 10490 36177
rect 10524 36143 10558 36177
rect 10592 36143 10626 36177
rect 10660 36143 10694 36177
rect 10728 36143 10762 36177
rect 10796 36143 10830 36177
rect 10864 36143 10898 36177
rect 10932 36143 10966 36177
rect 11000 36143 11034 36177
rect 11068 36143 11102 36177
rect 11136 36143 11170 36177
rect 11204 36143 11238 36177
rect 11272 36143 11306 36177
rect 11340 36143 11374 36177
rect 11408 36143 11442 36177
rect 11476 36143 11510 36177
rect 11544 36143 11578 36177
rect 11612 36143 11646 36177
rect 11680 36143 11714 36177
rect 11748 36143 11782 36177
rect 11816 36143 11850 36177
rect 11884 36143 11918 36177
rect 11952 36143 11986 36177
rect 12020 36143 12054 36177
rect 12088 36143 12122 36177
rect 12156 36143 12190 36177
rect 12224 36143 12258 36177
rect 12292 36143 12326 36177
rect 12360 36143 12394 36177
rect 12428 36143 12462 36177
rect 12496 36143 12530 36177
rect 12564 36143 12598 36177
rect 12632 36143 12666 36177
rect 12700 36143 12734 36177
rect 12768 36143 12802 36177
rect 12836 36143 12870 36177
rect 12904 36143 12938 36177
rect 12972 36143 13006 36177
rect 13040 36143 13074 36177
rect 13108 36143 13142 36177
rect 13176 36143 13210 36177
rect 13244 36143 13278 36177
rect 13312 36143 13346 36177
rect 13380 36143 13414 36177
rect 13448 36143 13482 36177
rect 13516 36143 13550 36177
rect 13584 36143 13618 36177
rect 13652 36143 13686 36177
rect 13720 36143 13754 36177
rect 13788 36143 13822 36177
rect 13856 36143 13890 36177
rect 13924 36143 13958 36177
rect 13992 36143 14026 36177
rect 14060 36143 14094 36177
rect 14128 36143 14162 36177
rect 14196 36143 14361 36177
rect 603 36032 14361 36143
rect 603 35998 632 36032
rect 666 36003 14297 36032
rect 666 35998 1007 36003
rect 603 35969 1007 35998
rect 1041 35969 1079 36003
rect 1113 35969 1151 36003
rect 1185 35969 1223 36003
rect 1257 35969 1295 36003
rect 1329 35969 1367 36003
rect 1401 35969 1439 36003
rect 1473 35969 1511 36003
rect 1545 35969 1583 36003
rect 1617 35969 1655 36003
rect 1689 35969 1727 36003
rect 1761 35969 1799 36003
rect 1833 35969 1871 36003
rect 1905 35969 1943 36003
rect 1977 35969 2015 36003
rect 2049 35969 2087 36003
rect 2121 35969 2159 36003
rect 2193 35969 2231 36003
rect 2265 35969 2303 36003
rect 2337 35969 2375 36003
rect 2409 35969 2447 36003
rect 2481 35969 2519 36003
rect 2553 35969 2591 36003
rect 2625 35969 2663 36003
rect 2697 35969 2735 36003
rect 2769 35969 2807 36003
rect 2841 35969 2879 36003
rect 2913 35969 2951 36003
rect 2985 35969 3023 36003
rect 3057 35969 3095 36003
rect 3129 35969 3167 36003
rect 3201 35969 3239 36003
rect 3273 35969 3311 36003
rect 3345 35969 3383 36003
rect 3417 35969 3455 36003
rect 3489 35969 3527 36003
rect 3561 35969 3599 36003
rect 3633 35969 3671 36003
rect 3705 35969 3743 36003
rect 3777 35969 3815 36003
rect 3849 35969 3887 36003
rect 3921 35969 3959 36003
rect 3993 35969 4031 36003
rect 4065 35969 4103 36003
rect 4137 35969 4175 36003
rect 4209 35969 4247 36003
rect 4281 35969 4319 36003
rect 4353 35969 4391 36003
rect 4425 35969 4463 36003
rect 4497 35969 4535 36003
rect 4569 35969 4607 36003
rect 4641 35969 4679 36003
rect 4713 35969 4751 36003
rect 4785 35969 4823 36003
rect 4857 35969 4895 36003
rect 4929 35969 4967 36003
rect 5001 35969 5039 36003
rect 5073 35969 5111 36003
rect 5145 35969 5183 36003
rect 5217 35969 5255 36003
rect 5289 35969 5327 36003
rect 5361 35969 5399 36003
rect 5433 35969 5471 36003
rect 5505 35969 5543 36003
rect 5577 35969 5615 36003
rect 5649 35969 5687 36003
rect 5721 35969 5759 36003
rect 5793 35969 5831 36003
rect 5865 35969 5903 36003
rect 5937 35969 5975 36003
rect 6009 35969 6047 36003
rect 6081 35969 6119 36003
rect 6153 35969 6191 36003
rect 6225 35969 6263 36003
rect 6297 35969 6335 36003
rect 6369 35969 6407 36003
rect 6441 35969 6479 36003
rect 6513 35969 6551 36003
rect 6585 35969 6623 36003
rect 6657 35969 6695 36003
rect 6729 35969 6767 36003
rect 6801 35969 6839 36003
rect 6873 35969 6911 36003
rect 6945 35969 6983 36003
rect 7017 35969 7055 36003
rect 7089 35969 7127 36003
rect 7161 35969 7199 36003
rect 7233 35969 7271 36003
rect 7305 35969 7343 36003
rect 7377 35969 7415 36003
rect 7449 35969 7487 36003
rect 7521 35969 7559 36003
rect 7593 35969 7631 36003
rect 7665 35969 7703 36003
rect 7737 35969 7775 36003
rect 7809 35969 7847 36003
rect 7881 35969 7919 36003
rect 7953 35969 7991 36003
rect 8025 35969 8063 36003
rect 8097 35969 8135 36003
rect 8169 35969 8207 36003
rect 8241 35969 8279 36003
rect 8313 35969 8351 36003
rect 8385 35969 8423 36003
rect 8457 35969 8495 36003
rect 8529 35969 8567 36003
rect 8601 35969 8639 36003
rect 8673 35969 8711 36003
rect 8745 35969 8783 36003
rect 8817 35969 8855 36003
rect 8889 35969 8927 36003
rect 8961 35969 8999 36003
rect 9033 35969 9071 36003
rect 9105 35969 9143 36003
rect 9177 35969 9215 36003
rect 9249 35969 9287 36003
rect 9321 35969 9359 36003
rect 9393 35969 9431 36003
rect 9465 35969 9503 36003
rect 9537 35969 9575 36003
rect 9609 35969 9647 36003
rect 9681 35969 9719 36003
rect 9753 35969 9791 36003
rect 9825 35969 9863 36003
rect 9897 35969 9935 36003
rect 9969 35969 10007 36003
rect 10041 35969 10079 36003
rect 10113 35969 10151 36003
rect 10185 35969 10223 36003
rect 10257 35969 10295 36003
rect 10329 35969 10367 36003
rect 10401 35969 10439 36003
rect 10473 35969 10511 36003
rect 10545 35969 10583 36003
rect 10617 35969 10655 36003
rect 10689 35969 10727 36003
rect 10761 35969 10799 36003
rect 10833 35969 10871 36003
rect 10905 35969 10943 36003
rect 10977 35969 11015 36003
rect 11049 35969 11087 36003
rect 11121 35969 11159 36003
rect 11193 35969 11231 36003
rect 11265 35969 11303 36003
rect 11337 35969 11375 36003
rect 11409 35969 11447 36003
rect 11481 35969 11519 36003
rect 11553 35969 11591 36003
rect 11625 35969 11663 36003
rect 11697 35969 11735 36003
rect 11769 35969 11807 36003
rect 11841 35969 11879 36003
rect 11913 35969 11951 36003
rect 11985 35969 12023 36003
rect 12057 35969 12095 36003
rect 12129 35969 12167 36003
rect 12201 35969 12239 36003
rect 12273 35969 12311 36003
rect 12345 35969 12383 36003
rect 12417 35969 12455 36003
rect 12489 35969 12527 36003
rect 12561 35969 12599 36003
rect 12633 35969 12671 36003
rect 12705 35969 12743 36003
rect 12777 35969 12815 36003
rect 12849 35969 12887 36003
rect 12921 35969 12959 36003
rect 12993 35969 13031 36003
rect 13065 35969 13103 36003
rect 13137 35969 13175 36003
rect 13209 35969 13247 36003
rect 13281 35969 13319 36003
rect 13353 35969 13391 36003
rect 13425 35969 13463 36003
rect 13497 35969 13535 36003
rect 13569 35969 13607 36003
rect 13641 35969 13679 36003
rect 13713 35969 13751 36003
rect 13785 35969 13823 36003
rect 13857 35969 13895 36003
rect 13929 35969 13967 36003
rect 14001 35998 14297 36003
rect 14331 35998 14361 36032
rect 14001 35969 14361 35998
rect 603 35964 14361 35969
rect 603 35930 632 35964
rect 666 35930 14297 35964
rect 14331 35930 14361 35964
rect 603 35896 14361 35930
rect 603 35862 632 35896
rect 666 35884 14297 35896
rect 666 35862 807 35884
rect 603 35850 807 35862
rect 841 35862 14297 35884
rect 14331 35862 14361 35896
rect 841 35850 14361 35862
rect 603 35828 14361 35850
rect 603 35794 632 35828
rect 666 35812 14297 35828
rect 666 35794 807 35812
rect 603 35778 807 35794
rect 841 35805 14297 35812
rect 841 35778 14142 35805
rect 603 35771 14142 35778
rect 14176 35794 14297 35805
rect 14331 35794 14361 35828
rect 14176 35771 14361 35794
rect 603 35760 14361 35771
rect 603 35726 632 35760
rect 666 35740 14297 35760
rect 666 35726 807 35740
rect 603 35706 807 35726
rect 841 35733 14297 35740
rect 841 35706 14142 35733
rect 603 35699 14142 35706
rect 14176 35726 14297 35733
rect 14331 35726 14361 35760
rect 14176 35699 14361 35726
rect 603 35692 14361 35699
rect 603 35658 632 35692
rect 666 35668 14297 35692
rect 666 35658 807 35668
rect 603 35634 807 35658
rect 841 35661 14297 35668
rect 841 35634 14142 35661
rect 603 35627 14142 35634
rect 14176 35658 14297 35661
rect 14331 35658 14361 35692
rect 14176 35627 14361 35658
rect 603 35624 14361 35627
rect 603 35590 632 35624
rect 666 35596 14297 35624
rect 666 35590 807 35596
rect 603 35562 807 35590
rect 841 35590 14297 35596
rect 14331 35590 14361 35624
rect 841 35589 14361 35590
rect 841 35562 14142 35589
rect 603 35556 14142 35562
rect 603 35522 632 35556
rect 666 35555 14142 35556
rect 14176 35556 14361 35589
rect 14176 35555 14297 35556
rect 666 35524 14297 35555
rect 666 35522 807 35524
rect 603 35490 807 35522
rect 841 35522 14297 35524
rect 14331 35522 14361 35556
rect 841 35517 14361 35522
rect 841 35490 14142 35517
rect 603 35488 14142 35490
rect 603 35454 632 35488
rect 666 35483 14142 35488
rect 14176 35488 14361 35517
rect 14176 35483 14297 35488
rect 666 35454 14297 35483
rect 14331 35454 14361 35488
rect 603 35452 14361 35454
rect 603 35420 807 35452
rect 603 35386 632 35420
rect 666 35418 807 35420
rect 841 35445 14361 35452
rect 841 35418 14142 35445
rect 666 35411 14142 35418
rect 14176 35420 14361 35445
rect 14176 35411 14297 35420
rect 666 35386 14297 35411
rect 14331 35386 14361 35420
rect 603 35380 14361 35386
rect 603 35352 807 35380
rect 603 35318 632 35352
rect 666 35346 807 35352
rect 841 35373 14361 35380
rect 841 35346 14142 35373
rect 666 35339 14142 35346
rect 14176 35352 14361 35373
rect 14176 35339 14297 35352
rect 666 35318 14297 35339
rect 14331 35318 14361 35352
rect 603 35308 14361 35318
rect 603 35284 807 35308
rect 603 35250 632 35284
rect 666 35274 807 35284
rect 841 35301 14361 35308
rect 841 35274 14142 35301
rect 666 35267 14142 35274
rect 14176 35284 14361 35301
rect 14176 35267 14297 35284
rect 666 35250 14297 35267
rect 14331 35250 14361 35284
rect 603 35236 14361 35250
rect 603 35216 807 35236
rect 603 35182 632 35216
rect 666 35202 807 35216
rect 841 35229 14361 35236
rect 841 35202 14142 35229
rect 666 35195 14142 35202
rect 14176 35216 14361 35229
rect 14176 35195 14297 35216
rect 666 35182 14297 35195
rect 14331 35182 14361 35216
rect 603 35164 14361 35182
rect 603 35148 807 35164
rect 603 35114 632 35148
rect 666 35130 807 35148
rect 841 35157 14361 35164
rect 841 35130 14142 35157
rect 666 35123 14142 35130
rect 14176 35148 14361 35157
rect 14176 35123 14297 35148
rect 666 35114 14297 35123
rect 14331 35114 14361 35148
rect 603 35092 14361 35114
rect 603 35080 807 35092
rect 603 35046 632 35080
rect 666 35058 807 35080
rect 841 35085 14361 35092
rect 841 35058 14142 35085
rect 666 35051 14142 35058
rect 14176 35080 14361 35085
rect 14176 35051 14297 35080
rect 666 35046 14297 35051
rect 14331 35046 14361 35080
rect 603 35020 14361 35046
rect 603 35012 807 35020
rect 603 34978 632 35012
rect 666 34986 807 35012
rect 841 35013 14361 35020
rect 841 34986 14142 35013
rect 666 34979 14142 34986
rect 14176 35012 14361 35013
rect 14176 34979 14297 35012
rect 666 34978 14297 34979
rect 14331 34978 14361 35012
rect 603 34948 14361 34978
rect 603 34944 807 34948
rect 603 34910 632 34944
rect 666 34914 807 34944
rect 841 34944 14361 34948
rect 841 34941 14297 34944
rect 841 34914 14142 34941
rect 666 34910 14142 34914
rect 603 34907 14142 34910
rect 14176 34910 14297 34941
rect 14331 34910 14361 34944
rect 14176 34907 14361 34910
rect 603 34876 14361 34907
rect 603 34842 632 34876
rect 666 34842 807 34876
rect 841 34869 14297 34876
rect 841 34842 14142 34869
rect 603 34835 14142 34842
rect 14176 34842 14297 34869
rect 14331 34842 14361 34876
rect 14176 34835 14361 34842
rect 603 34831 14361 34835
rect 603 34808 1026 34831
rect 603 34774 632 34808
rect 666 34804 1026 34808
rect 666 34774 807 34804
rect 603 34770 807 34774
rect 841 34770 1026 34804
rect 603 34740 1026 34770
rect 603 34706 632 34740
rect 666 34732 1026 34740
rect 666 34706 807 34732
rect 603 34698 807 34706
rect 841 34698 1026 34732
rect 603 34672 1026 34698
rect 13968 34808 14361 34831
rect 13968 34797 14297 34808
rect 13968 34763 14142 34797
rect 14176 34774 14297 34797
rect 14331 34774 14361 34808
rect 14176 34763 14361 34774
rect 13968 34740 14361 34763
rect 13968 34725 14297 34740
rect 603 34638 632 34672
rect 666 34660 1026 34672
rect 666 34638 807 34660
rect 603 34626 807 34638
rect 841 34626 1026 34660
rect 603 34604 1026 34626
rect 603 34570 632 34604
rect 666 34588 1026 34604
rect 666 34570 807 34588
rect 603 34554 807 34570
rect 841 34554 1026 34588
rect 603 34536 1026 34554
rect 603 34502 632 34536
rect 666 34516 1026 34536
rect 666 34502 807 34516
rect 603 34482 807 34502
rect 841 34482 1026 34516
rect 603 34468 1026 34482
rect 603 34434 632 34468
rect 666 34444 1026 34468
rect 666 34434 807 34444
rect 603 34410 807 34434
rect 841 34410 1026 34444
rect 603 34400 1026 34410
rect 603 34366 632 34400
rect 666 34372 1026 34400
rect 666 34366 807 34372
rect 603 34338 807 34366
rect 841 34338 1026 34372
rect 603 34332 1026 34338
rect 603 34298 632 34332
rect 666 34300 1026 34332
rect 666 34298 807 34300
rect 603 34266 807 34298
rect 841 34266 1026 34300
rect 603 34264 1026 34266
rect 603 34230 632 34264
rect 666 34230 1026 34264
rect 603 34228 1026 34230
rect 603 34196 807 34228
rect 603 34162 632 34196
rect 666 34194 807 34196
rect 841 34194 1026 34228
rect 666 34162 1026 34194
rect 603 34156 1026 34162
rect 603 34128 807 34156
rect 603 34094 632 34128
rect 666 34122 807 34128
rect 841 34122 1026 34156
rect 666 34094 1026 34122
rect 603 34084 1026 34094
rect 603 34060 807 34084
rect 603 34026 632 34060
rect 666 34050 807 34060
rect 841 34050 1026 34084
rect 666 34026 1026 34050
rect 603 34012 1026 34026
rect 603 33992 807 34012
rect 603 33958 632 33992
rect 666 33978 807 33992
rect 841 33978 1026 34012
rect 666 33958 1026 33978
rect 603 33940 1026 33958
rect 603 33924 807 33940
rect 603 33890 632 33924
rect 666 33906 807 33924
rect 841 33906 1026 33940
rect 666 33890 1026 33906
rect 603 33868 1026 33890
rect 603 33856 807 33868
rect 603 33822 632 33856
rect 666 33834 807 33856
rect 841 33834 1026 33868
rect 666 33822 1026 33834
rect 603 33796 1026 33822
rect 603 33788 807 33796
rect 603 33754 632 33788
rect 666 33762 807 33788
rect 841 33762 1026 33796
rect 666 33754 1026 33762
rect 603 33724 1026 33754
rect 603 33720 807 33724
rect 603 33686 632 33720
rect 666 33690 807 33720
rect 841 33690 1026 33724
rect 666 33686 1026 33690
rect 603 33652 1026 33686
rect 603 33618 632 33652
rect 666 33618 807 33652
rect 841 33618 1026 33652
rect 603 33584 1026 33618
rect 603 33550 632 33584
rect 666 33580 1026 33584
rect 666 33550 807 33580
rect 603 33546 807 33550
rect 841 33546 1026 33580
rect 603 33516 1026 33546
rect 603 33482 632 33516
rect 666 33508 1026 33516
rect 666 33482 807 33508
rect 603 33474 807 33482
rect 841 33474 1026 33508
rect 603 33448 1026 33474
rect 603 33414 632 33448
rect 666 33436 1026 33448
rect 666 33414 807 33436
rect 603 33402 807 33414
rect 841 33402 1026 33436
rect 603 33380 1026 33402
rect 603 33346 632 33380
rect 666 33364 1026 33380
rect 666 33346 807 33364
rect 603 33330 807 33346
rect 841 33330 1026 33364
rect 603 33312 1026 33330
rect 603 33278 632 33312
rect 666 33292 1026 33312
rect 666 33278 807 33292
rect 603 33258 807 33278
rect 841 33258 1026 33292
rect 603 33244 1026 33258
rect 603 33210 632 33244
rect 666 33220 1026 33244
rect 666 33210 807 33220
rect 603 33186 807 33210
rect 841 33186 1026 33220
rect 603 33176 1026 33186
rect 603 33142 632 33176
rect 666 33148 1026 33176
rect 666 33142 807 33148
rect 603 33114 807 33142
rect 841 33114 1026 33148
rect 603 33108 1026 33114
rect 603 33074 632 33108
rect 666 33076 1026 33108
rect 666 33074 807 33076
rect 603 33042 807 33074
rect 841 33042 1026 33076
rect 603 33040 1026 33042
rect 603 33006 632 33040
rect 666 33006 1026 33040
rect 603 33004 1026 33006
rect 603 32972 807 33004
rect 603 32938 632 32972
rect 666 32970 807 32972
rect 841 32970 1026 33004
rect 666 32938 1026 32970
rect 603 32932 1026 32938
rect 603 32904 807 32932
rect 603 32870 632 32904
rect 666 32898 807 32904
rect 841 32898 1026 32932
rect 666 32870 1026 32898
rect 603 32860 1026 32870
rect 603 32836 807 32860
rect 603 32802 632 32836
rect 666 32826 807 32836
rect 841 32826 1026 32860
rect 666 32802 1026 32826
rect 603 32788 1026 32802
rect 603 32768 807 32788
rect 603 32734 632 32768
rect 666 32754 807 32768
rect 841 32754 1026 32788
rect 666 32734 1026 32754
rect 603 32716 1026 32734
rect 603 32700 807 32716
rect 603 32666 632 32700
rect 666 32682 807 32700
rect 841 32682 1026 32716
rect 666 32666 1026 32682
rect 603 32644 1026 32666
rect 603 32632 807 32644
rect 603 32598 632 32632
rect 666 32610 807 32632
rect 841 32610 1026 32644
rect 666 32598 1026 32610
rect 603 32572 1026 32598
rect 603 32564 807 32572
rect 603 32530 632 32564
rect 666 32538 807 32564
rect 841 32538 1026 32572
rect 666 32530 1026 32538
rect 603 32500 1026 32530
rect 603 32496 807 32500
rect 603 32462 632 32496
rect 666 32466 807 32496
rect 841 32466 1026 32500
rect 666 32462 1026 32466
rect 603 32428 1026 32462
rect 603 32394 632 32428
rect 666 32394 807 32428
rect 841 32394 1026 32428
rect 603 32360 1026 32394
rect 603 32326 632 32360
rect 666 32356 1026 32360
rect 666 32326 807 32356
rect 603 32322 807 32326
rect 841 32322 1026 32356
rect 603 32292 1026 32322
rect 603 32258 632 32292
rect 666 32284 1026 32292
rect 666 32258 807 32284
rect 603 32250 807 32258
rect 841 32250 1026 32284
rect 603 32224 1026 32250
rect 603 32190 632 32224
rect 666 32212 1026 32224
rect 666 32190 807 32212
rect 603 32178 807 32190
rect 841 32178 1026 32212
rect 603 32156 1026 32178
rect 603 32122 632 32156
rect 666 32140 1026 32156
rect 666 32122 807 32140
rect 603 32106 807 32122
rect 841 32106 1026 32140
rect 603 32088 1026 32106
rect 603 32054 632 32088
rect 666 32068 1026 32088
rect 666 32054 807 32068
rect 603 32034 807 32054
rect 841 32034 1026 32068
rect 603 32020 1026 32034
rect 603 31986 632 32020
rect 666 31996 1026 32020
rect 666 31986 807 31996
rect 603 31962 807 31986
rect 841 31962 1026 31996
rect 603 31952 1026 31962
rect 603 31918 632 31952
rect 666 31924 1026 31952
rect 666 31918 807 31924
rect 603 31890 807 31918
rect 841 31890 1026 31924
rect 603 31884 1026 31890
rect 603 31850 632 31884
rect 666 31852 1026 31884
rect 666 31850 807 31852
rect 603 31818 807 31850
rect 841 31818 1026 31852
rect 603 31816 1026 31818
rect 603 31782 632 31816
rect 666 31782 1026 31816
rect 603 31780 1026 31782
rect 603 31748 807 31780
rect 603 31714 632 31748
rect 666 31746 807 31748
rect 841 31746 1026 31780
rect 666 31714 1026 31746
rect 603 31708 1026 31714
rect 603 31680 807 31708
rect 603 31646 632 31680
rect 666 31674 807 31680
rect 841 31674 1026 31708
rect 666 31646 1026 31674
rect 603 31636 1026 31646
rect 603 31612 807 31636
rect 603 31578 632 31612
rect 666 31602 807 31612
rect 841 31602 1026 31636
rect 666 31578 1026 31602
rect 603 31564 1026 31578
rect 603 31544 807 31564
rect 603 31510 632 31544
rect 666 31530 807 31544
rect 841 31530 1026 31564
rect 666 31510 1026 31530
rect 603 31492 1026 31510
rect 603 31476 807 31492
rect 603 31442 632 31476
rect 666 31458 807 31476
rect 841 31458 1026 31492
rect 666 31442 1026 31458
rect 603 31420 1026 31442
rect 603 31408 807 31420
rect 603 31374 632 31408
rect 666 31386 807 31408
rect 841 31386 1026 31420
rect 666 31374 1026 31386
rect 603 31348 1026 31374
rect 603 31340 807 31348
rect 603 31306 632 31340
rect 666 31314 807 31340
rect 841 31314 1026 31348
rect 666 31306 1026 31314
rect 603 31276 1026 31306
rect 603 31272 807 31276
rect 603 31238 632 31272
rect 666 31242 807 31272
rect 841 31242 1026 31276
rect 666 31238 1026 31242
rect 603 31204 1026 31238
rect 603 31170 632 31204
rect 666 31170 807 31204
rect 841 31170 1026 31204
rect 603 31136 1026 31170
rect 603 31102 632 31136
rect 666 31132 1026 31136
rect 666 31102 807 31132
rect 603 31098 807 31102
rect 841 31098 1026 31132
rect 603 31068 1026 31098
rect 603 31034 632 31068
rect 666 31060 1026 31068
rect 666 31034 807 31060
rect 603 31026 807 31034
rect 841 31026 1026 31060
rect 603 31000 1026 31026
rect 603 30966 632 31000
rect 666 30988 1026 31000
rect 666 30966 807 30988
rect 603 30954 807 30966
rect 841 30954 1026 30988
rect 603 30932 1026 30954
rect 603 30898 632 30932
rect 666 30916 1026 30932
rect 666 30898 807 30916
rect 603 30882 807 30898
rect 841 30882 1026 30916
rect 603 30864 1026 30882
rect 603 30830 632 30864
rect 666 30844 1026 30864
rect 666 30830 807 30844
rect 603 30810 807 30830
rect 841 30810 1026 30844
rect 603 30796 1026 30810
rect 603 30762 632 30796
rect 666 30772 1026 30796
rect 666 30762 807 30772
rect 603 30738 807 30762
rect 841 30738 1026 30772
rect 603 30728 1026 30738
rect 603 30694 632 30728
rect 666 30700 1026 30728
rect 666 30694 807 30700
rect 603 30666 807 30694
rect 841 30666 1026 30700
rect 603 30660 1026 30666
rect 603 30626 632 30660
rect 666 30628 1026 30660
rect 666 30626 807 30628
rect 603 30594 807 30626
rect 841 30594 1026 30628
rect 603 30592 1026 30594
rect 603 30558 632 30592
rect 666 30558 1026 30592
rect 603 30556 1026 30558
rect 603 30524 807 30556
rect 603 30490 632 30524
rect 666 30522 807 30524
rect 841 30522 1026 30556
rect 666 30490 1026 30522
rect 603 30484 1026 30490
rect 603 30456 807 30484
rect 603 30422 632 30456
rect 666 30450 807 30456
rect 841 30450 1026 30484
rect 666 30422 1026 30450
rect 603 30412 1026 30422
rect 603 30388 807 30412
rect 603 30354 632 30388
rect 666 30378 807 30388
rect 841 30378 1026 30412
rect 666 30354 1026 30378
rect 603 30340 1026 30354
rect 603 30320 807 30340
rect 603 30286 632 30320
rect 666 30306 807 30320
rect 841 30306 1026 30340
rect 666 30286 1026 30306
rect 603 30268 1026 30286
rect 603 30252 807 30268
rect 603 30218 632 30252
rect 666 30234 807 30252
rect 841 30234 1026 30268
rect 666 30218 1026 30234
rect 603 30196 1026 30218
rect 603 30184 807 30196
rect 603 30150 632 30184
rect 666 30162 807 30184
rect 841 30162 1026 30196
rect 666 30150 1026 30162
rect 603 30124 1026 30150
rect 603 30116 807 30124
rect 603 30082 632 30116
rect 666 30090 807 30116
rect 841 30090 1026 30124
rect 666 30082 1026 30090
rect 603 30052 1026 30082
rect 603 30048 807 30052
rect 603 30014 632 30048
rect 666 30018 807 30048
rect 841 30018 1026 30052
rect 666 30014 1026 30018
rect 603 29980 1026 30014
rect 603 29946 632 29980
rect 666 29946 807 29980
rect 841 29946 1026 29980
rect 603 29912 1026 29946
rect 603 29878 632 29912
rect 666 29908 1026 29912
rect 666 29878 807 29908
rect 603 29874 807 29878
rect 841 29874 1026 29908
rect 603 29844 1026 29874
rect 603 29810 632 29844
rect 666 29836 1026 29844
rect 666 29810 807 29836
rect 603 29802 807 29810
rect 841 29802 1026 29836
rect 603 29776 1026 29802
rect 603 29742 632 29776
rect 666 29764 1026 29776
rect 666 29742 807 29764
rect 603 29730 807 29742
rect 841 29730 1026 29764
rect 603 29708 1026 29730
rect 603 29674 632 29708
rect 666 29692 1026 29708
rect 666 29674 807 29692
rect 603 29658 807 29674
rect 841 29658 1026 29692
rect 603 29640 1026 29658
rect 603 29606 632 29640
rect 666 29620 1026 29640
rect 666 29606 807 29620
rect 603 29586 807 29606
rect 841 29586 1026 29620
rect 603 29572 1026 29586
rect 603 29538 632 29572
rect 666 29548 1026 29572
rect 666 29538 807 29548
rect 603 29514 807 29538
rect 841 29514 1026 29548
rect 603 29504 1026 29514
rect 603 29470 632 29504
rect 666 29476 1026 29504
rect 666 29470 807 29476
rect 603 29442 807 29470
rect 841 29442 1026 29476
rect 603 29436 1026 29442
rect 603 29402 632 29436
rect 666 29404 1026 29436
rect 666 29402 807 29404
rect 603 29370 807 29402
rect 841 29370 1026 29404
rect 603 29368 1026 29370
rect 603 29334 632 29368
rect 666 29334 1026 29368
rect 603 29332 1026 29334
rect 603 29300 807 29332
rect 603 29266 632 29300
rect 666 29298 807 29300
rect 841 29298 1026 29332
rect 666 29266 1026 29298
rect 603 29260 1026 29266
rect 603 29232 807 29260
rect 603 29198 632 29232
rect 666 29226 807 29232
rect 841 29226 1026 29260
rect 666 29198 1026 29226
rect 603 29188 1026 29198
rect 603 29164 807 29188
rect 603 29130 632 29164
rect 666 29154 807 29164
rect 841 29154 1026 29188
rect 666 29130 1026 29154
rect 603 29116 1026 29130
rect 603 29096 807 29116
rect 603 29062 632 29096
rect 666 29082 807 29096
rect 841 29082 1026 29116
rect 666 29062 1026 29082
rect 603 29044 1026 29062
rect 603 29028 807 29044
rect 603 28994 632 29028
rect 666 29010 807 29028
rect 841 29010 1026 29044
rect 666 28994 1026 29010
rect 603 28972 1026 28994
rect 603 28960 807 28972
rect 603 28926 632 28960
rect 666 28938 807 28960
rect 841 28938 1026 28972
rect 666 28926 1026 28938
rect 603 28900 1026 28926
rect 603 28892 807 28900
rect 603 28858 632 28892
rect 666 28866 807 28892
rect 841 28866 1026 28900
rect 666 28858 1026 28866
rect 603 28828 1026 28858
rect 603 28824 807 28828
rect 603 28790 632 28824
rect 666 28794 807 28824
rect 841 28794 1026 28828
rect 666 28790 1026 28794
rect 603 28756 1026 28790
rect 603 28722 632 28756
rect 666 28722 807 28756
rect 841 28722 1026 28756
rect 603 28688 1026 28722
rect 603 28654 632 28688
rect 666 28684 1026 28688
rect 666 28654 807 28684
rect 603 28650 807 28654
rect 841 28650 1026 28684
rect 603 28620 1026 28650
rect 603 28586 632 28620
rect 666 28612 1026 28620
rect 666 28586 807 28612
rect 603 28578 807 28586
rect 841 28578 1026 28612
rect 603 28552 1026 28578
rect 603 28518 632 28552
rect 666 28540 1026 28552
rect 666 28518 807 28540
rect 603 28506 807 28518
rect 841 28506 1026 28540
rect 603 28484 1026 28506
rect 603 28450 632 28484
rect 666 28468 1026 28484
rect 666 28450 807 28468
rect 603 28434 807 28450
rect 841 28434 1026 28468
rect 603 28416 1026 28434
rect 603 28382 632 28416
rect 666 28396 1026 28416
rect 666 28382 807 28396
rect 603 28362 807 28382
rect 841 28362 1026 28396
rect 603 28348 1026 28362
rect 603 28314 632 28348
rect 666 28324 1026 28348
rect 666 28314 807 28324
rect 603 28290 807 28314
rect 841 28290 1026 28324
rect 603 28280 1026 28290
rect 603 28246 632 28280
rect 666 28252 1026 28280
rect 666 28246 807 28252
rect 603 28218 807 28246
rect 841 28218 1026 28252
rect 603 28212 1026 28218
rect 603 28178 632 28212
rect 666 28180 1026 28212
rect 666 28178 807 28180
rect 603 28146 807 28178
rect 841 28146 1026 28180
rect 603 28144 1026 28146
rect 603 28110 632 28144
rect 666 28110 1026 28144
rect 603 28108 1026 28110
rect 603 28076 807 28108
rect 603 28042 632 28076
rect 666 28074 807 28076
rect 841 28074 1026 28108
rect 666 28042 1026 28074
rect 603 28036 1026 28042
rect 603 28008 807 28036
rect 603 27974 632 28008
rect 666 28002 807 28008
rect 841 28002 1026 28036
rect 666 27974 1026 28002
rect 603 27964 1026 27974
rect 603 27940 807 27964
rect 603 27906 632 27940
rect 666 27930 807 27940
rect 841 27930 1026 27964
rect 666 27906 1026 27930
rect 603 27892 1026 27906
rect 603 27872 807 27892
rect 603 27838 632 27872
rect 666 27858 807 27872
rect 841 27858 1026 27892
rect 666 27838 1026 27858
rect 603 27820 1026 27838
rect 603 27804 807 27820
rect 603 27770 632 27804
rect 666 27786 807 27804
rect 841 27786 1026 27820
rect 666 27770 1026 27786
rect 603 27748 1026 27770
rect 603 27736 807 27748
rect 603 27702 632 27736
rect 666 27714 807 27736
rect 841 27714 1026 27748
rect 666 27702 1026 27714
rect 603 27676 1026 27702
rect 603 27668 807 27676
rect 603 27634 632 27668
rect 666 27642 807 27668
rect 841 27642 1026 27676
rect 666 27634 1026 27642
rect 603 27604 1026 27634
rect 603 27600 807 27604
rect 603 27566 632 27600
rect 666 27570 807 27600
rect 841 27570 1026 27604
rect 666 27566 1026 27570
rect 603 27532 1026 27566
rect 603 27498 632 27532
rect 666 27498 807 27532
rect 841 27498 1026 27532
rect 603 27464 1026 27498
rect 603 27430 632 27464
rect 666 27460 1026 27464
rect 666 27430 807 27460
rect 603 27426 807 27430
rect 841 27426 1026 27460
rect 603 27396 1026 27426
rect 603 27362 632 27396
rect 666 27388 1026 27396
rect 666 27362 807 27388
rect 603 27354 807 27362
rect 841 27354 1026 27388
rect 603 27328 1026 27354
rect 603 27294 632 27328
rect 666 27316 1026 27328
rect 666 27294 807 27316
rect 603 27282 807 27294
rect 841 27282 1026 27316
rect 603 27260 1026 27282
rect 603 27226 632 27260
rect 666 27244 1026 27260
rect 666 27226 807 27244
rect 603 27210 807 27226
rect 841 27210 1026 27244
rect 603 27192 1026 27210
rect 603 27158 632 27192
rect 666 27172 1026 27192
rect 666 27158 807 27172
rect 603 27138 807 27158
rect 841 27138 1026 27172
rect 603 27124 1026 27138
rect 603 27090 632 27124
rect 666 27100 1026 27124
rect 666 27090 807 27100
rect 603 27066 807 27090
rect 841 27066 1026 27100
rect 603 27056 1026 27066
rect 603 27022 632 27056
rect 666 27028 1026 27056
rect 666 27022 807 27028
rect 603 26994 807 27022
rect 841 26994 1026 27028
rect 603 26988 1026 26994
rect 603 26954 632 26988
rect 666 26956 1026 26988
rect 666 26954 807 26956
rect 603 26922 807 26954
rect 841 26922 1026 26956
rect 603 26920 1026 26922
rect 603 26886 632 26920
rect 666 26886 1026 26920
rect 603 26884 1026 26886
rect 603 26852 807 26884
rect 603 26818 632 26852
rect 666 26850 807 26852
rect 841 26850 1026 26884
rect 666 26818 1026 26850
rect 603 26812 1026 26818
rect 603 26784 807 26812
rect 603 26750 632 26784
rect 666 26778 807 26784
rect 841 26778 1026 26812
rect 666 26750 1026 26778
rect 603 26740 1026 26750
rect 603 26716 807 26740
rect 603 26682 632 26716
rect 666 26706 807 26716
rect 841 26706 1026 26740
rect 666 26682 1026 26706
rect 603 26668 1026 26682
rect 603 26648 807 26668
rect 603 26614 632 26648
rect 666 26634 807 26648
rect 841 26634 1026 26668
rect 666 26614 1026 26634
rect 603 26596 1026 26614
rect 603 26580 807 26596
rect 603 26546 632 26580
rect 666 26562 807 26580
rect 841 26562 1026 26596
rect 666 26546 1026 26562
rect 603 26524 1026 26546
rect 603 26512 807 26524
rect 603 26478 632 26512
rect 666 26490 807 26512
rect 841 26490 1026 26524
rect 666 26478 1026 26490
rect 603 26452 1026 26478
rect 603 26444 807 26452
rect 603 26410 632 26444
rect 666 26418 807 26444
rect 841 26418 1026 26452
rect 666 26410 1026 26418
rect 603 26380 1026 26410
rect 603 26376 807 26380
rect 603 26342 632 26376
rect 666 26346 807 26376
rect 841 26346 1026 26380
rect 666 26342 1026 26346
rect 603 26308 1026 26342
rect 603 26274 632 26308
rect 666 26274 807 26308
rect 841 26274 1026 26308
rect 603 26240 1026 26274
rect 603 26206 632 26240
rect 666 26236 1026 26240
rect 666 26206 807 26236
rect 603 26202 807 26206
rect 841 26202 1026 26236
rect 603 26172 1026 26202
rect 603 26138 632 26172
rect 666 26164 1026 26172
rect 666 26138 807 26164
rect 603 26130 807 26138
rect 841 26130 1026 26164
rect 603 26104 1026 26130
rect 603 26070 632 26104
rect 666 26092 1026 26104
rect 666 26070 807 26092
rect 603 26058 807 26070
rect 841 26058 1026 26092
rect 603 26036 1026 26058
rect 603 26002 632 26036
rect 666 26020 1026 26036
rect 666 26002 807 26020
rect 603 25986 807 26002
rect 841 25986 1026 26020
rect 603 25968 1026 25986
rect 603 25934 632 25968
rect 666 25948 1026 25968
rect 666 25934 807 25948
rect 603 25914 807 25934
rect 841 25914 1026 25948
rect 603 25900 1026 25914
rect 603 25866 632 25900
rect 666 25876 1026 25900
rect 666 25866 807 25876
rect 603 25842 807 25866
rect 841 25842 1026 25876
rect 603 25832 1026 25842
rect 603 25798 632 25832
rect 666 25804 1026 25832
rect 666 25798 807 25804
rect 603 25770 807 25798
rect 841 25770 1026 25804
rect 603 25764 1026 25770
rect 603 25730 632 25764
rect 666 25732 1026 25764
rect 666 25730 807 25732
rect 603 25698 807 25730
rect 841 25698 1026 25732
rect 603 25696 1026 25698
rect 603 25662 632 25696
rect 666 25662 1026 25696
rect 603 25660 1026 25662
rect 603 25628 807 25660
rect 603 25594 632 25628
rect 666 25626 807 25628
rect 841 25626 1026 25660
rect 666 25594 1026 25626
rect 603 25588 1026 25594
rect 603 25560 807 25588
rect 603 25526 632 25560
rect 666 25554 807 25560
rect 841 25554 1026 25588
rect 666 25526 1026 25554
rect 603 25516 1026 25526
rect 603 25492 807 25516
rect 603 25458 632 25492
rect 666 25482 807 25492
rect 841 25482 1026 25516
rect 666 25458 1026 25482
rect 603 25444 1026 25458
rect 603 25424 807 25444
rect 603 25390 632 25424
rect 666 25410 807 25424
rect 841 25410 1026 25444
rect 666 25390 1026 25410
rect 603 25372 1026 25390
rect 603 25356 807 25372
rect 603 25322 632 25356
rect 666 25338 807 25356
rect 841 25338 1026 25372
rect 666 25322 1026 25338
rect 603 25300 1026 25322
rect 603 25288 807 25300
rect 603 25254 632 25288
rect 666 25266 807 25288
rect 841 25266 1026 25300
rect 666 25254 1026 25266
rect 603 25228 1026 25254
rect 603 25220 807 25228
rect 603 25186 632 25220
rect 666 25194 807 25220
rect 841 25194 1026 25228
rect 666 25186 1026 25194
rect 603 25156 1026 25186
rect 603 25152 807 25156
rect 603 25118 632 25152
rect 666 25122 807 25152
rect 841 25122 1026 25156
rect 666 25118 1026 25122
rect 603 25084 1026 25118
rect 603 25050 632 25084
rect 666 25050 807 25084
rect 841 25050 1026 25084
rect 603 25016 1026 25050
rect 603 24982 632 25016
rect 666 25012 1026 25016
rect 666 24982 807 25012
rect 603 24978 807 24982
rect 841 24978 1026 25012
rect 603 24948 1026 24978
rect 603 24914 632 24948
rect 666 24940 1026 24948
rect 666 24914 807 24940
rect 603 24906 807 24914
rect 841 24906 1026 24940
rect 603 24880 1026 24906
rect 603 24846 632 24880
rect 666 24868 1026 24880
rect 666 24846 807 24868
rect 603 24834 807 24846
rect 841 24834 1026 24868
rect 603 24812 1026 24834
rect 603 24778 632 24812
rect 666 24796 1026 24812
rect 666 24778 807 24796
rect 603 24762 807 24778
rect 841 24762 1026 24796
rect 603 24744 1026 24762
rect 603 24710 632 24744
rect 666 24724 1026 24744
rect 666 24710 807 24724
rect 603 24690 807 24710
rect 841 24690 1026 24724
rect 603 24676 1026 24690
rect 603 24642 632 24676
rect 666 24652 1026 24676
rect 666 24642 807 24652
rect 603 24618 807 24642
rect 841 24618 1026 24652
rect 603 24608 1026 24618
rect 603 24574 632 24608
rect 666 24580 1026 24608
rect 666 24574 807 24580
rect 603 24546 807 24574
rect 841 24546 1026 24580
rect 603 24540 1026 24546
rect 603 24506 632 24540
rect 666 24508 1026 24540
rect 666 24506 807 24508
rect 603 24474 807 24506
rect 841 24474 1026 24508
rect 603 24472 1026 24474
rect 603 24438 632 24472
rect 666 24438 1026 24472
rect 603 24436 1026 24438
rect 603 24404 807 24436
rect 603 24370 632 24404
rect 666 24402 807 24404
rect 841 24402 1026 24436
rect 666 24370 1026 24402
rect 603 24364 1026 24370
rect 603 24336 807 24364
rect 603 24302 632 24336
rect 666 24330 807 24336
rect 841 24330 1026 24364
rect 666 24302 1026 24330
rect 603 24292 1026 24302
rect 603 24268 807 24292
rect 603 24234 632 24268
rect 666 24258 807 24268
rect 841 24258 1026 24292
rect 666 24234 1026 24258
rect 603 24220 1026 24234
rect 603 24200 807 24220
rect 603 24166 632 24200
rect 666 24186 807 24200
rect 841 24186 1026 24220
rect 666 24166 1026 24186
rect 603 24148 1026 24166
rect 603 24132 807 24148
rect 603 24098 632 24132
rect 666 24114 807 24132
rect 841 24114 1026 24148
rect 666 24098 1026 24114
rect 603 24076 1026 24098
rect 603 24064 807 24076
rect 603 24030 632 24064
rect 666 24042 807 24064
rect 841 24042 1026 24076
rect 666 24030 1026 24042
rect 603 24004 1026 24030
rect 603 23996 807 24004
rect 603 23962 632 23996
rect 666 23970 807 23996
rect 841 23970 1026 24004
rect 666 23962 1026 23970
rect 603 23932 1026 23962
rect 603 23928 807 23932
rect 603 23894 632 23928
rect 666 23898 807 23928
rect 841 23898 1026 23932
rect 666 23894 1026 23898
rect 603 23860 1026 23894
rect 603 23826 632 23860
rect 666 23826 807 23860
rect 841 23826 1026 23860
rect 603 23792 1026 23826
rect 603 23758 632 23792
rect 666 23788 1026 23792
rect 666 23758 807 23788
rect 603 23754 807 23758
rect 841 23754 1026 23788
rect 603 23724 1026 23754
rect 603 23690 632 23724
rect 666 23716 1026 23724
rect 666 23690 807 23716
rect 603 23682 807 23690
rect 841 23682 1026 23716
rect 603 23656 1026 23682
rect 603 23622 632 23656
rect 666 23644 1026 23656
rect 666 23622 807 23644
rect 603 23610 807 23622
rect 841 23610 1026 23644
rect 603 23588 1026 23610
rect 603 23554 632 23588
rect 666 23572 1026 23588
rect 666 23554 807 23572
rect 603 23538 807 23554
rect 841 23538 1026 23572
rect 603 23520 1026 23538
rect 603 23486 632 23520
rect 666 23500 1026 23520
rect 666 23486 807 23500
rect 603 23466 807 23486
rect 841 23466 1026 23500
rect 603 23452 1026 23466
rect 603 23418 632 23452
rect 666 23428 1026 23452
rect 666 23418 807 23428
rect 603 23394 807 23418
rect 841 23394 1026 23428
rect 603 23384 1026 23394
rect 603 23350 632 23384
rect 666 23356 1026 23384
rect 666 23350 807 23356
rect 603 23322 807 23350
rect 841 23322 1026 23356
rect 603 23316 1026 23322
rect 603 23282 632 23316
rect 666 23284 1026 23316
rect 666 23282 807 23284
rect 603 23250 807 23282
rect 841 23250 1026 23284
rect 603 23248 1026 23250
rect 603 23214 632 23248
rect 666 23214 1026 23248
rect 603 23212 1026 23214
rect 603 23180 807 23212
rect 603 23146 632 23180
rect 666 23178 807 23180
rect 841 23178 1026 23212
rect 666 23146 1026 23178
rect 603 23140 1026 23146
rect 603 23112 807 23140
rect 603 23078 632 23112
rect 666 23106 807 23112
rect 841 23106 1026 23140
rect 666 23078 1026 23106
rect 603 23068 1026 23078
rect 603 23044 807 23068
rect 603 23010 632 23044
rect 666 23034 807 23044
rect 841 23034 1026 23068
rect 666 23010 1026 23034
rect 603 22996 1026 23010
rect 603 22976 807 22996
rect 603 22942 632 22976
rect 666 22962 807 22976
rect 841 22962 1026 22996
rect 666 22942 1026 22962
rect 603 22924 1026 22942
rect 603 22908 807 22924
rect 603 22874 632 22908
rect 666 22890 807 22908
rect 841 22890 1026 22924
rect 666 22874 1026 22890
rect 603 22852 1026 22874
rect 603 22840 807 22852
rect 603 22806 632 22840
rect 666 22818 807 22840
rect 841 22818 1026 22852
rect 666 22806 1026 22818
rect 603 22780 1026 22806
rect 603 22772 807 22780
rect 603 22738 632 22772
rect 666 22746 807 22772
rect 841 22746 1026 22780
rect 666 22738 1026 22746
rect 603 22708 1026 22738
rect 603 22704 807 22708
rect 603 22670 632 22704
rect 666 22674 807 22704
rect 841 22674 1026 22708
rect 666 22670 1026 22674
rect 603 22636 1026 22670
rect 603 22602 632 22636
rect 666 22602 807 22636
rect 841 22602 1026 22636
rect 603 22568 1026 22602
rect 603 22534 632 22568
rect 666 22564 1026 22568
rect 666 22534 807 22564
rect 603 22530 807 22534
rect 841 22530 1026 22564
rect 603 22500 1026 22530
rect 603 22466 632 22500
rect 666 22492 1026 22500
rect 666 22466 807 22492
rect 603 22458 807 22466
rect 841 22458 1026 22492
rect 603 22432 1026 22458
rect 603 22398 632 22432
rect 666 22420 1026 22432
rect 666 22398 807 22420
rect 603 22386 807 22398
rect 841 22386 1026 22420
rect 603 22364 1026 22386
rect 603 22330 632 22364
rect 666 22348 1026 22364
rect 666 22330 807 22348
rect 603 22314 807 22330
rect 841 22314 1026 22348
rect 603 22296 1026 22314
rect 603 22262 632 22296
rect 666 22276 1026 22296
rect 666 22262 807 22276
rect 603 22242 807 22262
rect 841 22242 1026 22276
rect 603 22228 1026 22242
rect 603 22194 632 22228
rect 666 22204 1026 22228
rect 666 22194 807 22204
rect 603 22170 807 22194
rect 841 22170 1026 22204
rect 603 22160 1026 22170
rect 603 22126 632 22160
rect 666 22132 1026 22160
rect 666 22126 807 22132
rect 603 22098 807 22126
rect 841 22098 1026 22132
rect 603 22092 1026 22098
rect 603 22058 632 22092
rect 666 22060 1026 22092
rect 666 22058 807 22060
rect 603 22026 807 22058
rect 841 22026 1026 22060
rect 603 22024 1026 22026
rect 603 21990 632 22024
rect 666 21990 1026 22024
rect 603 21988 1026 21990
rect 603 21956 807 21988
rect 603 21922 632 21956
rect 666 21954 807 21956
rect 841 21954 1026 21988
rect 666 21922 1026 21954
rect 603 21916 1026 21922
rect 603 21888 807 21916
rect 603 21854 632 21888
rect 666 21882 807 21888
rect 841 21882 1026 21916
rect 666 21854 1026 21882
rect 603 21844 1026 21854
rect 603 21820 807 21844
rect 603 21786 632 21820
rect 666 21810 807 21820
rect 841 21810 1026 21844
rect 666 21786 1026 21810
rect 603 21772 1026 21786
rect 603 21752 807 21772
rect 603 21718 632 21752
rect 666 21738 807 21752
rect 841 21738 1026 21772
rect 666 21718 1026 21738
rect 603 21700 1026 21718
rect 603 21684 807 21700
rect 603 21650 632 21684
rect 666 21666 807 21684
rect 841 21666 1026 21700
rect 666 21650 1026 21666
rect 603 21628 1026 21650
rect 603 21616 807 21628
rect 603 21582 632 21616
rect 666 21594 807 21616
rect 841 21594 1026 21628
rect 666 21582 1026 21594
rect 603 21556 1026 21582
rect 603 21548 807 21556
rect 603 21514 632 21548
rect 666 21522 807 21548
rect 841 21522 1026 21556
rect 666 21514 1026 21522
rect 603 21484 1026 21514
rect 603 21480 807 21484
rect 603 21446 632 21480
rect 666 21450 807 21480
rect 841 21450 1026 21484
rect 666 21446 1026 21450
rect 603 21412 1026 21446
rect 603 21378 632 21412
rect 666 21378 807 21412
rect 841 21378 1026 21412
rect 603 21344 1026 21378
rect 603 21310 632 21344
rect 666 21340 1026 21344
rect 666 21310 807 21340
rect 603 21306 807 21310
rect 841 21306 1026 21340
rect 603 21276 1026 21306
rect 603 21242 632 21276
rect 666 21268 1026 21276
rect 666 21242 807 21268
rect 603 21234 807 21242
rect 841 21234 1026 21268
rect 603 21208 1026 21234
rect 603 21174 632 21208
rect 666 21196 1026 21208
rect 666 21174 807 21196
rect 603 21162 807 21174
rect 841 21162 1026 21196
rect 603 21140 1026 21162
rect 603 21106 632 21140
rect 666 21124 1026 21140
rect 666 21106 807 21124
rect 603 21090 807 21106
rect 841 21090 1026 21124
rect 603 21072 1026 21090
rect 603 21038 632 21072
rect 666 21052 1026 21072
rect 666 21038 807 21052
rect 603 21018 807 21038
rect 841 21018 1026 21052
rect 603 21004 1026 21018
rect 603 20970 632 21004
rect 666 20980 1026 21004
rect 666 20970 807 20980
rect 603 20946 807 20970
rect 841 20946 1026 20980
rect 603 20936 1026 20946
rect 603 20902 632 20936
rect 666 20908 1026 20936
rect 666 20902 807 20908
rect 603 20874 807 20902
rect 841 20874 1026 20908
rect 603 20868 1026 20874
rect 603 20834 632 20868
rect 666 20836 1026 20868
rect 666 20834 807 20836
rect 603 20802 807 20834
rect 841 20802 1026 20836
rect 603 20800 1026 20802
rect 603 20766 632 20800
rect 666 20766 1026 20800
rect 603 20764 1026 20766
rect 603 20732 807 20764
rect 603 20698 632 20732
rect 666 20730 807 20732
rect 841 20730 1026 20764
rect 666 20698 1026 20730
rect 603 20692 1026 20698
rect 603 20664 807 20692
rect 603 20630 632 20664
rect 666 20658 807 20664
rect 841 20658 1026 20692
rect 666 20630 1026 20658
rect 603 20620 1026 20630
rect 603 20596 807 20620
rect 603 20562 632 20596
rect 666 20586 807 20596
rect 841 20586 1026 20620
rect 666 20562 1026 20586
rect 603 20548 1026 20562
rect 603 20528 807 20548
rect 603 20494 632 20528
rect 666 20514 807 20528
rect 841 20514 1026 20548
rect 666 20494 1026 20514
rect 603 20476 1026 20494
rect 603 20460 807 20476
rect 603 20426 632 20460
rect 666 20442 807 20460
rect 841 20442 1026 20476
rect 666 20426 1026 20442
rect 603 20404 1026 20426
rect 603 20392 807 20404
rect 603 20358 632 20392
rect 666 20370 807 20392
rect 841 20370 1026 20404
rect 666 20358 1026 20370
rect 603 20332 1026 20358
rect 603 20324 807 20332
rect 603 20290 632 20324
rect 666 20298 807 20324
rect 841 20298 1026 20332
rect 666 20290 1026 20298
rect 603 20260 1026 20290
rect 603 20256 807 20260
rect 603 20222 632 20256
rect 666 20226 807 20256
rect 841 20226 1026 20260
rect 666 20222 1026 20226
rect 603 20188 1026 20222
rect 603 20154 632 20188
rect 666 20154 807 20188
rect 841 20154 1026 20188
rect 603 20120 1026 20154
rect 603 20086 632 20120
rect 666 20116 1026 20120
rect 666 20086 807 20116
rect 603 20082 807 20086
rect 841 20082 1026 20116
rect 603 20052 1026 20082
rect 603 20018 632 20052
rect 666 20044 1026 20052
rect 666 20018 807 20044
rect 603 20010 807 20018
rect 841 20010 1026 20044
rect 603 19984 1026 20010
rect 603 19950 632 19984
rect 666 19972 1026 19984
rect 666 19950 807 19972
rect 603 19938 807 19950
rect 841 19938 1026 19972
rect 603 19916 1026 19938
rect 603 19882 632 19916
rect 666 19900 1026 19916
rect 666 19882 807 19900
rect 603 19866 807 19882
rect 841 19866 1026 19900
rect 603 19848 1026 19866
rect 603 19814 632 19848
rect 666 19828 1026 19848
rect 666 19814 807 19828
rect 603 19794 807 19814
rect 841 19794 1026 19828
rect 603 19780 1026 19794
rect 603 19746 632 19780
rect 666 19756 1026 19780
rect 666 19746 807 19756
rect 603 19722 807 19746
rect 841 19722 1026 19756
rect 603 19712 1026 19722
rect 603 19678 632 19712
rect 666 19684 1026 19712
rect 666 19678 807 19684
rect 603 19650 807 19678
rect 841 19650 1026 19684
rect 603 19644 1026 19650
rect 603 19610 632 19644
rect 666 19612 1026 19644
rect 666 19610 807 19612
rect 603 19578 807 19610
rect 841 19578 1026 19612
rect 603 19576 1026 19578
rect 603 19542 632 19576
rect 666 19542 1026 19576
rect 603 19540 1026 19542
rect 603 19508 807 19540
rect 603 19474 632 19508
rect 666 19506 807 19508
rect 841 19506 1026 19540
rect 666 19474 1026 19506
rect 603 19468 1026 19474
rect 603 19440 807 19468
rect 603 19406 632 19440
rect 666 19434 807 19440
rect 841 19434 1026 19468
rect 666 19406 1026 19434
rect 603 19396 1026 19406
rect 603 19372 807 19396
rect 603 19338 632 19372
rect 666 19362 807 19372
rect 841 19362 1026 19396
rect 666 19338 1026 19362
rect 603 19324 1026 19338
rect 603 19304 807 19324
rect 603 19270 632 19304
rect 666 19290 807 19304
rect 841 19290 1026 19324
rect 666 19270 1026 19290
rect 603 19252 1026 19270
rect 603 19236 807 19252
rect 603 19202 632 19236
rect 666 19218 807 19236
rect 841 19218 1026 19252
rect 666 19202 1026 19218
rect 603 19180 1026 19202
rect 603 19168 807 19180
rect 603 19134 632 19168
rect 666 19146 807 19168
rect 841 19146 1026 19180
rect 666 19134 1026 19146
rect 603 19108 1026 19134
rect 603 19100 807 19108
rect 603 19066 632 19100
rect 666 19074 807 19100
rect 841 19074 1026 19108
rect 666 19066 1026 19074
rect 603 19036 1026 19066
rect 603 19032 807 19036
rect 603 18998 632 19032
rect 666 19002 807 19032
rect 841 19002 1026 19036
rect 666 18998 1026 19002
rect 603 18964 1026 18998
rect 603 18930 632 18964
rect 666 18930 807 18964
rect 841 18930 1026 18964
rect 603 18896 1026 18930
rect 603 18862 632 18896
rect 666 18892 1026 18896
rect 666 18862 807 18892
rect 603 18858 807 18862
rect 841 18858 1026 18892
rect 603 18828 1026 18858
rect 603 18794 632 18828
rect 666 18820 1026 18828
rect 666 18794 807 18820
rect 603 18786 807 18794
rect 841 18786 1026 18820
rect 603 18760 1026 18786
rect 603 18726 632 18760
rect 666 18748 1026 18760
rect 666 18726 807 18748
rect 603 18714 807 18726
rect 841 18714 1026 18748
rect 603 18692 1026 18714
rect 603 18658 632 18692
rect 666 18676 1026 18692
rect 666 18658 807 18676
rect 603 18642 807 18658
rect 841 18642 1026 18676
rect 603 18624 1026 18642
rect 603 18590 632 18624
rect 666 18604 1026 18624
rect 666 18590 807 18604
rect 603 18570 807 18590
rect 841 18570 1026 18604
rect 603 18556 1026 18570
rect 603 18522 632 18556
rect 666 18532 1026 18556
rect 666 18522 807 18532
rect 603 18498 807 18522
rect 841 18498 1026 18532
rect 603 18488 1026 18498
rect 603 18454 632 18488
rect 666 18460 1026 18488
rect 666 18454 807 18460
rect 603 18426 807 18454
rect 841 18426 1026 18460
rect 603 18420 1026 18426
rect 603 18386 632 18420
rect 666 18388 1026 18420
rect 666 18386 807 18388
rect 603 18354 807 18386
rect 841 18354 1026 18388
rect 603 18352 1026 18354
rect 603 18318 632 18352
rect 666 18318 1026 18352
rect 603 18316 1026 18318
rect 603 18284 807 18316
rect 603 18250 632 18284
rect 666 18282 807 18284
rect 841 18282 1026 18316
rect 666 18250 1026 18282
rect 603 18244 1026 18250
rect 603 18216 807 18244
rect 603 18182 632 18216
rect 666 18210 807 18216
rect 841 18210 1026 18244
rect 666 18182 1026 18210
rect 603 18172 1026 18182
rect 603 18148 807 18172
rect 603 18114 632 18148
rect 666 18138 807 18148
rect 841 18138 1026 18172
rect 666 18114 1026 18138
rect 603 18100 1026 18114
rect 603 18080 807 18100
rect 603 18046 632 18080
rect 666 18066 807 18080
rect 841 18066 1026 18100
rect 666 18046 1026 18066
rect 603 18028 1026 18046
rect 603 18012 807 18028
rect 603 17978 632 18012
rect 666 17994 807 18012
rect 841 17994 1026 18028
rect 666 17978 1026 17994
rect 603 17956 1026 17978
rect 603 17944 807 17956
rect 603 17910 632 17944
rect 666 17922 807 17944
rect 841 17922 1026 17956
rect 666 17910 1026 17922
rect 603 17884 1026 17910
rect 603 17876 807 17884
rect 603 17842 632 17876
rect 666 17850 807 17876
rect 841 17850 1026 17884
rect 666 17842 1026 17850
rect 603 17812 1026 17842
rect 603 17808 807 17812
rect 603 17774 632 17808
rect 666 17778 807 17808
rect 841 17778 1026 17812
rect 666 17774 1026 17778
rect 603 17740 1026 17774
rect 603 17706 632 17740
rect 666 17706 807 17740
rect 841 17706 1026 17740
rect 603 17672 1026 17706
rect 603 17638 632 17672
rect 666 17668 1026 17672
rect 666 17638 807 17668
rect 603 17634 807 17638
rect 841 17634 1026 17668
rect 603 17604 1026 17634
rect 603 17570 632 17604
rect 666 17596 1026 17604
rect 666 17570 807 17596
rect 603 17562 807 17570
rect 841 17562 1026 17596
rect 603 17536 1026 17562
rect 603 17502 632 17536
rect 666 17524 1026 17536
rect 666 17502 807 17524
rect 603 17490 807 17502
rect 841 17490 1026 17524
rect 603 17468 1026 17490
rect 603 17434 632 17468
rect 666 17452 1026 17468
rect 666 17434 807 17452
rect 603 17418 807 17434
rect 841 17418 1026 17452
rect 603 17400 1026 17418
rect 603 17366 632 17400
rect 666 17380 1026 17400
rect 666 17366 807 17380
rect 603 17346 807 17366
rect 841 17346 1026 17380
rect 603 17332 1026 17346
rect 603 17298 632 17332
rect 666 17308 1026 17332
rect 666 17298 807 17308
rect 603 17274 807 17298
rect 841 17274 1026 17308
rect 603 17264 1026 17274
rect 603 17230 632 17264
rect 666 17236 1026 17264
rect 666 17230 807 17236
rect 603 17202 807 17230
rect 841 17202 1026 17236
rect 603 17196 1026 17202
rect 603 17162 632 17196
rect 666 17164 1026 17196
rect 666 17162 807 17164
rect 603 17130 807 17162
rect 841 17130 1026 17164
rect 603 17128 1026 17130
rect 603 17094 632 17128
rect 666 17094 1026 17128
rect 603 17092 1026 17094
rect 603 17060 807 17092
rect 603 17026 632 17060
rect 666 17058 807 17060
rect 841 17058 1026 17092
rect 666 17026 1026 17058
rect 603 17020 1026 17026
rect 603 16992 807 17020
rect 603 16958 632 16992
rect 666 16986 807 16992
rect 841 16986 1026 17020
rect 666 16958 1026 16986
rect 603 16948 1026 16958
rect 603 16924 807 16948
rect 603 16890 632 16924
rect 666 16914 807 16924
rect 841 16914 1026 16948
rect 666 16890 1026 16914
rect 603 16876 1026 16890
rect 603 16856 807 16876
rect 603 16822 632 16856
rect 666 16842 807 16856
rect 841 16842 1026 16876
rect 666 16822 1026 16842
rect 603 16804 1026 16822
rect 603 16788 807 16804
rect 603 16754 632 16788
rect 666 16770 807 16788
rect 841 16770 1026 16804
rect 666 16754 1026 16770
rect 603 16732 1026 16754
rect 603 16720 807 16732
rect 603 16686 632 16720
rect 666 16698 807 16720
rect 841 16698 1026 16732
rect 666 16686 1026 16698
rect 603 16660 1026 16686
rect 603 16652 807 16660
rect 603 16618 632 16652
rect 666 16626 807 16652
rect 841 16626 1026 16660
rect 666 16618 1026 16626
rect 603 16588 1026 16618
rect 603 16584 807 16588
rect 603 16550 632 16584
rect 666 16554 807 16584
rect 841 16554 1026 16588
rect 666 16550 1026 16554
rect 603 16516 1026 16550
rect 603 16482 632 16516
rect 666 16482 807 16516
rect 841 16482 1026 16516
rect 603 16448 1026 16482
rect 603 16414 632 16448
rect 666 16444 1026 16448
rect 666 16414 807 16444
rect 603 16410 807 16414
rect 841 16410 1026 16444
rect 603 16380 1026 16410
rect 603 16346 632 16380
rect 666 16372 1026 16380
rect 666 16346 807 16372
rect 603 16338 807 16346
rect 841 16338 1026 16372
rect 603 16312 1026 16338
rect 603 16278 632 16312
rect 666 16300 1026 16312
rect 666 16278 807 16300
rect 603 16266 807 16278
rect 841 16266 1026 16300
rect 603 16244 1026 16266
rect 603 16210 632 16244
rect 666 16228 1026 16244
rect 666 16210 807 16228
rect 603 16194 807 16210
rect 841 16194 1026 16228
rect 603 16176 1026 16194
rect 603 16142 632 16176
rect 666 16156 1026 16176
rect 666 16142 807 16156
rect 603 16122 807 16142
rect 841 16122 1026 16156
rect 603 16108 1026 16122
rect 603 16074 632 16108
rect 666 16084 1026 16108
rect 666 16074 807 16084
rect 603 16050 807 16074
rect 841 16050 1026 16084
rect 603 16040 1026 16050
rect 603 16006 632 16040
rect 666 16012 1026 16040
rect 666 16006 807 16012
rect 603 15978 807 16006
rect 841 15978 1026 16012
rect 603 15972 1026 15978
rect 603 15938 632 15972
rect 666 15940 1026 15972
rect 666 15938 807 15940
rect 603 15906 807 15938
rect 841 15906 1026 15940
rect 603 15904 1026 15906
rect 603 15870 632 15904
rect 666 15870 1026 15904
rect 603 15868 1026 15870
rect 603 15836 807 15868
rect 603 15802 632 15836
rect 666 15834 807 15836
rect 841 15834 1026 15868
rect 666 15802 1026 15834
rect 603 15796 1026 15802
rect 603 15768 807 15796
rect 603 15734 632 15768
rect 666 15762 807 15768
rect 841 15762 1026 15796
rect 666 15734 1026 15762
rect 603 15724 1026 15734
rect 603 15700 807 15724
rect 603 15666 632 15700
rect 666 15690 807 15700
rect 841 15690 1026 15724
rect 666 15666 1026 15690
rect 603 15652 1026 15666
rect 603 15632 807 15652
rect 603 15598 632 15632
rect 666 15618 807 15632
rect 841 15618 1026 15652
rect 666 15598 1026 15618
rect 603 15580 1026 15598
rect 603 15564 807 15580
rect 603 15530 632 15564
rect 666 15546 807 15564
rect 841 15546 1026 15580
rect 666 15530 1026 15546
rect 603 15508 1026 15530
rect 603 15496 807 15508
rect 603 15462 632 15496
rect 666 15474 807 15496
rect 841 15474 1026 15508
rect 666 15462 1026 15474
rect 603 15436 1026 15462
rect 603 15428 807 15436
rect 603 15394 632 15428
rect 666 15402 807 15428
rect 841 15402 1026 15436
rect 666 15394 1026 15402
rect 603 15364 1026 15394
rect 603 15360 807 15364
rect 603 15326 632 15360
rect 666 15330 807 15360
rect 841 15330 1026 15364
rect 666 15326 1026 15330
rect 603 15292 1026 15326
rect 603 15258 632 15292
rect 666 15258 807 15292
rect 841 15258 1026 15292
rect 603 15224 1026 15258
rect 603 15190 632 15224
rect 666 15220 1026 15224
rect 666 15190 807 15220
rect 603 15186 807 15190
rect 841 15186 1026 15220
rect 603 15156 1026 15186
rect 603 15122 632 15156
rect 666 15148 1026 15156
rect 666 15122 807 15148
rect 603 15114 807 15122
rect 841 15114 1026 15148
rect 603 15088 1026 15114
rect 603 15054 632 15088
rect 666 15076 1026 15088
rect 666 15054 807 15076
rect 603 15042 807 15054
rect 841 15042 1026 15076
rect 603 15020 1026 15042
rect 603 14986 632 15020
rect 666 15004 1026 15020
rect 666 14986 807 15004
rect 603 14970 807 14986
rect 841 14970 1026 15004
rect 603 14952 1026 14970
rect 603 14918 632 14952
rect 666 14932 1026 14952
rect 666 14918 807 14932
rect 603 14898 807 14918
rect 841 14898 1026 14932
rect 603 14884 1026 14898
rect 603 14850 632 14884
rect 666 14860 1026 14884
rect 666 14850 807 14860
rect 603 14826 807 14850
rect 841 14826 1026 14860
rect 603 14816 1026 14826
rect 603 14782 632 14816
rect 666 14788 1026 14816
rect 666 14782 807 14788
rect 603 14754 807 14782
rect 841 14754 1026 14788
rect 603 14748 1026 14754
rect 603 14714 632 14748
rect 666 14716 1026 14748
rect 666 14714 807 14716
rect 603 14682 807 14714
rect 841 14682 1026 14716
rect 603 14680 1026 14682
rect 603 14646 632 14680
rect 666 14646 1026 14680
rect 603 14644 1026 14646
rect 603 14612 807 14644
rect 603 14578 632 14612
rect 666 14610 807 14612
rect 841 14610 1026 14644
rect 666 14578 1026 14610
rect 603 14572 1026 14578
rect 603 14544 807 14572
rect 603 14510 632 14544
rect 666 14538 807 14544
rect 841 14538 1026 14572
rect 666 14510 1026 14538
rect 603 14500 1026 14510
rect 603 14476 807 14500
rect 603 14442 632 14476
rect 666 14466 807 14476
rect 841 14466 1026 14500
rect 666 14442 1026 14466
rect 603 14428 1026 14442
rect 603 14408 807 14428
rect 603 14374 632 14408
rect 666 14394 807 14408
rect 841 14394 1026 14428
rect 666 14374 1026 14394
rect 603 14356 1026 14374
rect 603 14340 807 14356
rect 603 14306 632 14340
rect 666 14322 807 14340
rect 841 14322 1026 14356
rect 666 14306 1026 14322
rect 603 14284 1026 14306
rect 603 14272 807 14284
rect 603 14238 632 14272
rect 666 14250 807 14272
rect 841 14250 1026 14284
rect 666 14238 1026 14250
rect 603 14212 1026 14238
rect 603 14204 807 14212
rect 603 14170 632 14204
rect 666 14178 807 14204
rect 841 14178 1026 14212
rect 666 14170 1026 14178
rect 603 14140 1026 14170
rect 603 14136 807 14140
rect 603 14102 632 14136
rect 666 14106 807 14136
rect 841 14106 1026 14140
rect 666 14102 1026 14106
rect 603 14068 1026 14102
rect 603 14034 632 14068
rect 666 14034 807 14068
rect 841 14034 1026 14068
rect 603 14000 1026 14034
rect 603 13966 632 14000
rect 666 13996 1026 14000
rect 666 13966 807 13996
rect 603 13962 807 13966
rect 841 13962 1026 13996
rect 603 13932 1026 13962
rect 603 13898 632 13932
rect 666 13924 1026 13932
rect 666 13898 807 13924
rect 603 13890 807 13898
rect 841 13890 1026 13924
rect 603 13864 1026 13890
rect 603 13830 632 13864
rect 666 13852 1026 13864
rect 666 13830 807 13852
rect 603 13818 807 13830
rect 841 13818 1026 13852
rect 603 13796 1026 13818
rect 603 13762 632 13796
rect 666 13780 1026 13796
rect 666 13762 807 13780
rect 603 13746 807 13762
rect 841 13746 1026 13780
rect 603 13728 1026 13746
rect 603 13694 632 13728
rect 666 13708 1026 13728
rect 666 13694 807 13708
rect 603 13674 807 13694
rect 841 13674 1026 13708
rect 603 13660 1026 13674
rect 603 13626 632 13660
rect 666 13636 1026 13660
rect 666 13626 807 13636
rect 603 13602 807 13626
rect 841 13602 1026 13636
rect 603 13592 1026 13602
rect 603 13558 632 13592
rect 666 13564 1026 13592
rect 666 13558 807 13564
rect 603 13530 807 13558
rect 841 13530 1026 13564
rect 603 13524 1026 13530
rect 603 13490 632 13524
rect 666 13492 1026 13524
rect 666 13490 807 13492
rect 603 13458 807 13490
rect 841 13458 1026 13492
rect 603 13456 1026 13458
rect 603 13422 632 13456
rect 666 13422 1026 13456
rect 603 13420 1026 13422
rect 603 13388 807 13420
rect 603 13354 632 13388
rect 666 13386 807 13388
rect 841 13386 1026 13420
rect 666 13354 1026 13386
rect 603 13348 1026 13354
rect 603 13320 807 13348
rect 603 13286 632 13320
rect 666 13314 807 13320
rect 841 13314 1026 13348
rect 666 13286 1026 13314
rect 603 13276 1026 13286
rect 603 13252 807 13276
rect 603 13218 632 13252
rect 666 13242 807 13252
rect 841 13242 1026 13276
rect 666 13218 1026 13242
rect 603 13204 1026 13218
rect 603 13184 807 13204
rect 603 13150 632 13184
rect 666 13170 807 13184
rect 841 13170 1026 13204
rect 666 13150 1026 13170
rect 603 13132 1026 13150
rect 603 13116 807 13132
rect 603 13082 632 13116
rect 666 13098 807 13116
rect 841 13098 1026 13132
rect 666 13082 1026 13098
rect 603 13060 1026 13082
rect 603 13048 807 13060
rect 603 13014 632 13048
rect 666 13026 807 13048
rect 841 13026 1026 13060
rect 666 13014 1026 13026
rect 603 12988 1026 13014
rect 603 12980 807 12988
rect 603 12946 632 12980
rect 666 12954 807 12980
rect 841 12954 1026 12988
rect 666 12946 1026 12954
rect 603 12916 1026 12946
rect 603 12912 807 12916
rect 603 12878 632 12912
rect 666 12882 807 12912
rect 841 12882 1026 12916
rect 666 12878 1026 12882
rect 603 12844 1026 12878
rect 603 12810 632 12844
rect 666 12810 807 12844
rect 841 12810 1026 12844
rect 603 12776 1026 12810
rect 603 12742 632 12776
rect 666 12772 1026 12776
rect 666 12742 807 12772
rect 603 12738 807 12742
rect 841 12738 1026 12772
rect 603 12708 1026 12738
rect 603 12674 632 12708
rect 666 12700 1026 12708
rect 666 12674 807 12700
rect 603 12666 807 12674
rect 841 12666 1026 12700
rect 603 12640 1026 12666
rect 603 12606 632 12640
rect 666 12628 1026 12640
rect 666 12606 807 12628
rect 603 12594 807 12606
rect 841 12594 1026 12628
rect 603 12572 1026 12594
rect 603 12538 632 12572
rect 666 12556 1026 12572
rect 666 12538 807 12556
rect 603 12522 807 12538
rect 841 12522 1026 12556
rect 603 12504 1026 12522
rect 603 12470 632 12504
rect 666 12484 1026 12504
rect 666 12470 807 12484
rect 603 12450 807 12470
rect 841 12450 1026 12484
rect 603 12436 1026 12450
rect 603 12402 632 12436
rect 666 12412 1026 12436
rect 666 12402 807 12412
rect 603 12378 807 12402
rect 841 12378 1026 12412
rect 603 12368 1026 12378
rect 603 12334 632 12368
rect 666 12340 1026 12368
rect 666 12334 807 12340
rect 603 12306 807 12334
rect 841 12306 1026 12340
rect 603 12300 1026 12306
rect 603 12266 632 12300
rect 666 12268 1026 12300
rect 666 12266 807 12268
rect 603 12234 807 12266
rect 841 12234 1026 12268
rect 603 12232 1026 12234
rect 603 12198 632 12232
rect 666 12198 1026 12232
rect 603 12196 1026 12198
rect 603 12164 807 12196
rect 603 12130 632 12164
rect 666 12162 807 12164
rect 841 12162 1026 12196
rect 666 12130 1026 12162
rect 603 12124 1026 12130
rect 603 12096 807 12124
rect 603 12062 632 12096
rect 666 12090 807 12096
rect 841 12090 1026 12124
rect 666 12062 1026 12090
rect 603 12052 1026 12062
rect 603 12028 807 12052
rect 603 11994 632 12028
rect 666 12018 807 12028
rect 841 12018 1026 12052
rect 666 11994 1026 12018
rect 603 11980 1026 11994
rect 603 11960 807 11980
rect 603 11926 632 11960
rect 666 11946 807 11960
rect 841 11946 1026 11980
rect 666 11926 1026 11946
rect 603 11908 1026 11926
rect 603 11892 807 11908
rect 603 11858 632 11892
rect 666 11874 807 11892
rect 841 11874 1026 11908
rect 666 11858 1026 11874
rect 603 11836 1026 11858
rect 603 11824 807 11836
rect 603 11790 632 11824
rect 666 11802 807 11824
rect 841 11802 1026 11836
rect 666 11790 1026 11802
rect 603 11764 1026 11790
rect 603 11756 807 11764
rect 603 11722 632 11756
rect 666 11730 807 11756
rect 841 11730 1026 11764
rect 666 11722 1026 11730
rect 603 11692 1026 11722
rect 603 11688 807 11692
rect 603 11654 632 11688
rect 666 11658 807 11688
rect 841 11658 1026 11692
rect 666 11654 1026 11658
rect 603 11620 1026 11654
rect 603 11586 632 11620
rect 666 11586 807 11620
rect 841 11586 1026 11620
rect 603 11552 1026 11586
rect 603 11518 632 11552
rect 666 11548 1026 11552
rect 666 11518 807 11548
rect 603 11514 807 11518
rect 841 11514 1026 11548
rect 603 11484 1026 11514
rect 603 11450 632 11484
rect 666 11476 1026 11484
rect 666 11450 807 11476
rect 603 11442 807 11450
rect 841 11442 1026 11476
rect 603 11416 1026 11442
rect 603 11382 632 11416
rect 666 11404 1026 11416
rect 666 11382 807 11404
rect 603 11370 807 11382
rect 841 11370 1026 11404
rect 603 11348 1026 11370
rect 603 11314 632 11348
rect 666 11332 1026 11348
rect 666 11314 807 11332
rect 603 11298 807 11314
rect 841 11298 1026 11332
rect 603 11280 1026 11298
rect 603 11246 632 11280
rect 666 11260 1026 11280
rect 666 11246 807 11260
rect 603 11226 807 11246
rect 841 11226 1026 11260
rect 603 11212 1026 11226
rect 603 11178 632 11212
rect 666 11188 1026 11212
rect 666 11178 807 11188
rect 603 11154 807 11178
rect 841 11154 1026 11188
rect 603 11144 1026 11154
rect 603 11110 632 11144
rect 666 11116 1026 11144
rect 666 11110 807 11116
rect 603 11082 807 11110
rect 841 11082 1026 11116
rect 603 11076 1026 11082
rect 603 11042 632 11076
rect 666 11044 1026 11076
rect 666 11042 807 11044
rect 603 11010 807 11042
rect 841 11010 1026 11044
rect 603 11008 1026 11010
rect 603 10974 632 11008
rect 666 10974 1026 11008
rect 603 10972 1026 10974
rect 603 10940 807 10972
rect 603 10906 632 10940
rect 666 10938 807 10940
rect 841 10938 1026 10972
rect 666 10906 1026 10938
rect 603 10900 1026 10906
rect 603 10872 807 10900
rect 603 10838 632 10872
rect 666 10866 807 10872
rect 841 10866 1026 10900
rect 666 10838 1026 10866
rect 603 10828 1026 10838
rect 603 10804 807 10828
rect 603 10770 632 10804
rect 666 10794 807 10804
rect 841 10794 1026 10828
rect 666 10770 1026 10794
rect 603 10756 1026 10770
rect 603 10736 807 10756
rect 603 10702 632 10736
rect 666 10722 807 10736
rect 841 10722 1026 10756
rect 666 10702 1026 10722
rect 603 10684 1026 10702
rect 603 10668 807 10684
rect 603 10634 632 10668
rect 666 10650 807 10668
rect 841 10650 1026 10684
rect 666 10634 1026 10650
rect 603 10612 1026 10634
rect 603 10600 807 10612
rect 603 10566 632 10600
rect 666 10578 807 10600
rect 841 10578 1026 10612
rect 666 10566 1026 10578
rect 603 10540 1026 10566
rect 603 10532 807 10540
rect 603 10498 632 10532
rect 666 10506 807 10532
rect 841 10506 1026 10540
rect 666 10498 1026 10506
rect 603 10468 1026 10498
rect 603 10464 807 10468
rect 603 10430 632 10464
rect 666 10434 807 10464
rect 841 10434 1026 10468
rect 666 10430 1026 10434
rect 603 10396 1026 10430
rect 603 10362 632 10396
rect 666 10362 807 10396
rect 841 10362 1026 10396
rect 603 10328 1026 10362
rect 603 10294 632 10328
rect 666 10324 1026 10328
rect 666 10294 807 10324
rect 603 10290 807 10294
rect 841 10290 1026 10324
rect 603 10260 1026 10290
rect 603 10226 632 10260
rect 666 10252 1026 10260
rect 666 10226 807 10252
rect 603 10218 807 10226
rect 841 10218 1026 10252
rect 1148 34650 13844 34694
rect 1148 34616 1325 34650
rect 1361 34616 1395 34650
rect 1431 34616 1463 34650
rect 1503 34616 1531 34650
rect 1575 34616 1599 34650
rect 1647 34616 1667 34650
rect 1719 34616 1735 34650
rect 1791 34616 1803 34650
rect 1863 34616 1871 34650
rect 1935 34616 1939 34650
rect 2041 34616 2045 34650
rect 2109 34616 2117 34650
rect 2177 34616 2189 34650
rect 2245 34616 2261 34650
rect 2313 34616 2333 34650
rect 2381 34616 2405 34650
rect 2449 34616 2477 34650
rect 2517 34616 2549 34650
rect 2585 34616 2619 34650
rect 2655 34616 2687 34650
rect 2727 34616 2755 34650
rect 2799 34616 2823 34650
rect 2871 34616 2891 34650
rect 2943 34616 2959 34650
rect 3015 34616 3027 34650
rect 3087 34616 3095 34650
rect 3159 34616 3163 34650
rect 3265 34616 3269 34650
rect 3333 34616 3341 34650
rect 3401 34616 3413 34650
rect 3469 34616 3485 34650
rect 3537 34616 3557 34650
rect 3605 34616 3629 34650
rect 3673 34616 3701 34650
rect 3741 34616 3773 34650
rect 3809 34616 3843 34650
rect 3879 34616 3911 34650
rect 3951 34616 3979 34650
rect 4023 34616 4047 34650
rect 4095 34616 4115 34650
rect 4167 34616 4183 34650
rect 4239 34616 4251 34650
rect 4311 34616 4319 34650
rect 4383 34616 4387 34650
rect 4489 34616 4493 34650
rect 4557 34616 4565 34650
rect 4625 34616 4637 34650
rect 4693 34616 4709 34650
rect 4761 34616 4781 34650
rect 4829 34616 4853 34650
rect 4897 34616 4925 34650
rect 4965 34616 4997 34650
rect 5033 34616 5067 34650
rect 5103 34616 5135 34650
rect 5175 34616 5203 34650
rect 5247 34616 5271 34650
rect 5319 34616 5339 34650
rect 5391 34616 5407 34650
rect 5463 34616 5475 34650
rect 5535 34616 5543 34650
rect 5607 34616 5611 34650
rect 5713 34616 5717 34650
rect 5781 34616 5789 34650
rect 5849 34616 5861 34650
rect 5917 34616 5933 34650
rect 5985 34616 6005 34650
rect 6053 34616 6077 34650
rect 6121 34616 6149 34650
rect 6189 34616 6221 34650
rect 6257 34616 6291 34650
rect 6327 34616 6359 34650
rect 6399 34616 6427 34650
rect 6471 34616 6495 34650
rect 6543 34616 6563 34650
rect 6615 34616 6631 34650
rect 6687 34616 6699 34650
rect 6759 34616 6767 34650
rect 6831 34616 6835 34650
rect 6937 34616 6941 34650
rect 7005 34616 7013 34650
rect 7073 34616 7085 34650
rect 7141 34616 7157 34650
rect 7209 34616 7229 34650
rect 7277 34616 7301 34650
rect 7345 34616 7373 34650
rect 7413 34616 7445 34650
rect 7481 34616 7515 34650
rect 7551 34616 7583 34650
rect 7623 34616 7651 34650
rect 7695 34616 7719 34650
rect 7767 34616 7787 34650
rect 7839 34616 7855 34650
rect 7911 34616 7923 34650
rect 7983 34616 7991 34650
rect 8055 34616 8059 34650
rect 8161 34616 8165 34650
rect 8229 34616 8237 34650
rect 8297 34616 8309 34650
rect 8365 34616 8381 34650
rect 8433 34616 8453 34650
rect 8501 34616 8525 34650
rect 8569 34616 8597 34650
rect 8637 34616 8669 34650
rect 8705 34616 8739 34650
rect 8775 34616 8807 34650
rect 8847 34616 8875 34650
rect 8919 34616 8943 34650
rect 8991 34616 9011 34650
rect 9063 34616 9079 34650
rect 9135 34616 9147 34650
rect 9207 34616 9215 34650
rect 9279 34616 9283 34650
rect 9385 34616 9389 34650
rect 9453 34616 9461 34650
rect 9521 34616 9533 34650
rect 9589 34616 9605 34650
rect 9657 34616 9677 34650
rect 9725 34616 9749 34650
rect 9793 34616 9821 34650
rect 9861 34616 9893 34650
rect 9929 34616 9963 34650
rect 9999 34616 10031 34650
rect 10071 34616 10099 34650
rect 10143 34616 10167 34650
rect 10215 34616 10235 34650
rect 10287 34616 10303 34650
rect 10359 34616 10371 34650
rect 10431 34616 10439 34650
rect 10503 34616 10507 34650
rect 10609 34616 10613 34650
rect 10677 34616 10685 34650
rect 10745 34616 10757 34650
rect 10813 34616 10829 34650
rect 10881 34616 10901 34650
rect 10949 34616 10973 34650
rect 11017 34616 11045 34650
rect 11085 34616 11117 34650
rect 11153 34616 11187 34650
rect 11223 34616 11255 34650
rect 11295 34616 11323 34650
rect 11367 34616 11391 34650
rect 11439 34616 11459 34650
rect 11511 34616 11527 34650
rect 11583 34616 11595 34650
rect 11655 34616 11663 34650
rect 11727 34616 11731 34650
rect 11833 34616 11837 34650
rect 11901 34616 11909 34650
rect 11969 34616 11981 34650
rect 12037 34616 12053 34650
rect 12105 34616 12125 34650
rect 12173 34616 12197 34650
rect 12241 34616 12269 34650
rect 12309 34616 12341 34650
rect 12377 34616 12411 34650
rect 12447 34616 12479 34650
rect 12519 34616 12547 34650
rect 12591 34616 12615 34650
rect 12663 34616 12683 34650
rect 12735 34616 12751 34650
rect 12807 34616 12819 34650
rect 12879 34616 12887 34650
rect 12951 34616 12955 34650
rect 13057 34616 13061 34650
rect 13125 34616 13133 34650
rect 13193 34616 13205 34650
rect 13261 34616 13277 34650
rect 13329 34616 13349 34650
rect 13397 34616 13421 34650
rect 13465 34616 13493 34650
rect 13533 34616 13565 34650
rect 13601 34616 13635 34650
rect 13671 34616 13844 34650
rect 1148 34574 13844 34616
rect 1148 34521 1268 34574
rect 1148 34475 1192 34521
rect 1226 34475 1268 34521
rect 1148 34453 1268 34475
rect 1148 34403 1192 34453
rect 1226 34403 1268 34453
rect 1148 34385 1268 34403
rect 1148 34331 1192 34385
rect 1226 34331 1268 34385
rect 1148 34317 1268 34331
rect 1148 34259 1192 34317
rect 1226 34259 1268 34317
rect 1148 34249 1268 34259
rect 1148 34187 1192 34249
rect 1226 34187 1268 34249
rect 1148 34181 1268 34187
rect 1148 34115 1192 34181
rect 1226 34115 1268 34181
rect 1148 34113 1268 34115
rect 1148 34079 1192 34113
rect 1226 34079 1268 34113
rect 1148 34077 1268 34079
rect 1148 34011 1192 34077
rect 1226 34011 1268 34077
rect 1148 34005 1268 34011
rect 1148 33943 1192 34005
rect 1226 33943 1268 34005
rect 1148 33933 1268 33943
rect 1148 33875 1192 33933
rect 1226 33875 1268 33933
rect 1148 33861 1268 33875
rect 1148 33807 1192 33861
rect 1226 33807 1268 33861
rect 1148 33789 1268 33807
rect 1148 33739 1192 33789
rect 1226 33739 1268 33789
rect 1148 33717 1268 33739
rect 1148 33671 1192 33717
rect 1226 33671 1268 33717
rect 1148 33645 1268 33671
rect 1148 33603 1192 33645
rect 1226 33603 1268 33645
rect 1148 33573 1268 33603
rect 1148 33535 1192 33573
rect 1226 33535 1268 33573
rect 1148 33501 1268 33535
rect 1148 33467 1192 33501
rect 1226 33467 1268 33501
rect 1148 33433 1268 33467
rect 1148 33395 1192 33433
rect 1226 33395 1268 33433
rect 1148 33365 1268 33395
rect 1148 33323 1192 33365
rect 1226 33323 1268 33365
rect 1148 33297 1268 33323
rect 1148 33251 1192 33297
rect 1226 33251 1268 33297
rect 1148 33229 1268 33251
rect 1148 33179 1192 33229
rect 1226 33179 1268 33229
rect 1148 33161 1268 33179
rect 1148 33107 1192 33161
rect 1226 33107 1268 33161
rect 1148 33093 1268 33107
rect 1148 33035 1192 33093
rect 1226 33035 1268 33093
rect 1148 33025 1268 33035
rect 1148 32963 1192 33025
rect 1226 32963 1268 33025
rect 1148 32957 1268 32963
rect 1148 32891 1192 32957
rect 1226 32891 1268 32957
rect 1148 32889 1268 32891
rect 1148 32855 1192 32889
rect 1226 32855 1268 32889
rect 1148 32853 1268 32855
rect 1148 32787 1192 32853
rect 1226 32787 1268 32853
rect 1148 32781 1268 32787
rect 1148 32719 1192 32781
rect 1226 32719 1268 32781
rect 1148 32709 1268 32719
rect 1148 32651 1192 32709
rect 1226 32651 1268 32709
rect 1148 32637 1268 32651
rect 1148 32583 1192 32637
rect 1226 32583 1268 32637
rect 1148 32565 1268 32583
rect 1148 32515 1192 32565
rect 1226 32515 1268 32565
rect 1148 32493 1268 32515
rect 1148 32447 1192 32493
rect 1226 32447 1268 32493
rect 1148 32421 1268 32447
rect 1148 32379 1192 32421
rect 1226 32379 1268 32421
rect 1148 32349 1268 32379
rect 1148 32311 1192 32349
rect 1226 32311 1268 32349
rect 1148 32277 1268 32311
rect 1148 32243 1192 32277
rect 1226 32243 1268 32277
rect 1148 32209 1268 32243
rect 1148 32171 1192 32209
rect 1226 32171 1268 32209
rect 1148 32141 1268 32171
rect 1148 32099 1192 32141
rect 1226 32099 1268 32141
rect 1148 32073 1268 32099
rect 1148 32027 1192 32073
rect 1226 32027 1268 32073
rect 1148 32005 1268 32027
rect 1148 31955 1192 32005
rect 1226 31955 1268 32005
rect 1148 31937 1268 31955
rect 1148 31883 1192 31937
rect 1226 31883 1268 31937
rect 1148 31869 1268 31883
rect 1148 31811 1192 31869
rect 1226 31811 1268 31869
rect 1148 31801 1268 31811
rect 1148 31739 1192 31801
rect 1226 31739 1268 31801
rect 1148 31733 1268 31739
rect 1148 31667 1192 31733
rect 1226 31667 1268 31733
rect 1148 31665 1268 31667
rect 1148 31631 1192 31665
rect 1226 31631 1268 31665
rect 1148 31629 1268 31631
rect 1148 31563 1192 31629
rect 1226 31563 1268 31629
rect 1148 31557 1268 31563
rect 1148 31495 1192 31557
rect 1226 31495 1268 31557
rect 1148 31485 1268 31495
rect 1148 31427 1192 31485
rect 1226 31427 1268 31485
rect 1148 31413 1268 31427
rect 1148 31359 1192 31413
rect 1226 31359 1268 31413
rect 13724 34534 13844 34574
rect 13724 34474 13768 34534
rect 13802 34474 13844 34534
rect 13724 34466 13844 34474
rect 13724 34402 13768 34466
rect 13802 34402 13844 34466
rect 13724 34398 13844 34402
rect 13724 34296 13768 34398
rect 13802 34296 13844 34398
rect 13724 34292 13844 34296
rect 13724 34228 13768 34292
rect 13802 34228 13844 34292
rect 13724 34220 13844 34228
rect 13724 34160 13768 34220
rect 13802 34160 13844 34220
rect 13724 34148 13844 34160
rect 13724 34092 13768 34148
rect 13802 34092 13844 34148
rect 13724 34076 13844 34092
rect 13724 34024 13768 34076
rect 13802 34024 13844 34076
rect 13724 34004 13844 34024
rect 13724 33956 13768 34004
rect 13802 33956 13844 34004
rect 13724 33932 13844 33956
rect 13724 33888 13768 33932
rect 13802 33888 13844 33932
rect 13724 33860 13844 33888
rect 13724 33820 13768 33860
rect 13802 33820 13844 33860
rect 13724 33788 13844 33820
rect 13724 33752 13768 33788
rect 13802 33752 13844 33788
rect 13724 33718 13844 33752
rect 13724 33682 13768 33718
rect 13802 33682 13844 33718
rect 13724 33650 13844 33682
rect 13724 33610 13768 33650
rect 13802 33610 13844 33650
rect 13724 33582 13844 33610
rect 13724 33538 13768 33582
rect 13802 33538 13844 33582
rect 13724 33514 13844 33538
rect 13724 33466 13768 33514
rect 13802 33466 13844 33514
rect 13724 33446 13844 33466
rect 13724 33394 13768 33446
rect 13802 33394 13844 33446
rect 13724 33378 13844 33394
rect 13724 33322 13768 33378
rect 13802 33322 13844 33378
rect 13724 33310 13844 33322
rect 13724 33250 13768 33310
rect 13802 33250 13844 33310
rect 13724 33242 13844 33250
rect 13724 33178 13768 33242
rect 13802 33178 13844 33242
rect 13724 33174 13844 33178
rect 13724 33072 13768 33174
rect 13802 33072 13844 33174
rect 13724 33068 13844 33072
rect 13724 33004 13768 33068
rect 13802 33004 13844 33068
rect 13724 32996 13844 33004
rect 13724 32936 13768 32996
rect 13802 32936 13844 32996
rect 13724 32924 13844 32936
rect 13724 32868 13768 32924
rect 13802 32868 13844 32924
rect 13724 32852 13844 32868
rect 13724 32800 13768 32852
rect 13802 32800 13844 32852
rect 13724 32780 13844 32800
rect 13724 32732 13768 32780
rect 13802 32732 13844 32780
rect 13724 32708 13844 32732
rect 13724 32664 13768 32708
rect 13802 32664 13844 32708
rect 13724 32636 13844 32664
rect 13724 32596 13768 32636
rect 13802 32596 13844 32636
rect 13724 32564 13844 32596
rect 13724 32528 13768 32564
rect 13802 32528 13844 32564
rect 13724 32494 13844 32528
rect 13724 32458 13768 32494
rect 13802 32458 13844 32494
rect 13724 32426 13844 32458
rect 13724 32386 13768 32426
rect 13802 32386 13844 32426
rect 13724 32358 13844 32386
rect 13724 32314 13768 32358
rect 13802 32314 13844 32358
rect 13724 32290 13844 32314
rect 13724 32242 13768 32290
rect 13802 32242 13844 32290
rect 13724 32222 13844 32242
rect 13724 32170 13768 32222
rect 13802 32170 13844 32222
rect 13724 32154 13844 32170
rect 13724 32098 13768 32154
rect 13802 32098 13844 32154
rect 13724 32086 13844 32098
rect 13724 32026 13768 32086
rect 13802 32026 13844 32086
rect 13724 32018 13844 32026
rect 13724 31954 13768 32018
rect 13802 31954 13844 32018
rect 13724 31950 13844 31954
rect 13724 31848 13768 31950
rect 13802 31848 13844 31950
rect 13724 31844 13844 31848
rect 13724 31780 13768 31844
rect 13802 31780 13844 31844
rect 13724 31772 13844 31780
rect 13724 31712 13768 31772
rect 13802 31712 13844 31772
rect 13724 31700 13844 31712
rect 13724 31644 13768 31700
rect 13802 31644 13844 31700
rect 13724 31628 13844 31644
rect 13724 31576 13768 31628
rect 13802 31576 13844 31628
rect 13724 31556 13844 31576
rect 13724 31508 13768 31556
rect 13802 31508 13844 31556
rect 13724 31484 13844 31508
rect 13724 31440 13768 31484
rect 13802 31440 13844 31484
rect 13724 31412 13844 31440
rect 1148 31341 1268 31359
rect 1148 31291 1192 31341
rect 1226 31291 1268 31341
rect 1148 31269 1268 31291
rect 1148 31223 1192 31269
rect 1226 31223 1268 31269
rect 1148 31197 1268 31223
rect 1148 31155 1192 31197
rect 1226 31155 1268 31197
rect 1148 31125 1268 31155
rect 1148 31087 1192 31125
rect 1226 31087 1268 31125
rect 1148 31053 1268 31087
rect 1148 31019 1192 31053
rect 1226 31019 1268 31053
rect 1148 30985 1268 31019
rect 1148 30947 1192 30985
rect 1226 30947 1268 30985
rect 1148 30917 1268 30947
rect 1148 30875 1192 30917
rect 1226 30875 1268 30917
rect 1148 30849 1268 30875
rect 1148 30803 1192 30849
rect 1226 30803 1268 30849
rect 1148 30781 1268 30803
rect 1148 30731 1192 30781
rect 1226 30731 1268 30781
rect 1148 30713 1268 30731
rect 1148 30659 1192 30713
rect 1226 30659 1268 30713
rect 1148 30645 1268 30659
rect 1148 30587 1192 30645
rect 1226 30587 1268 30645
rect 1148 30577 1268 30587
rect 1148 30515 1192 30577
rect 1226 30515 1268 30577
rect 1148 30509 1268 30515
rect 1148 30443 1192 30509
rect 1226 30443 1268 30509
rect 1148 30441 1268 30443
rect 1148 30407 1192 30441
rect 1226 30407 1268 30441
rect 1148 30405 1268 30407
rect 1148 30339 1192 30405
rect 1226 30339 1268 30405
rect 1148 30333 1268 30339
rect 1148 30271 1192 30333
rect 1226 30271 1268 30333
rect 1148 30261 1268 30271
rect 1148 30203 1192 30261
rect 1226 30203 1268 30261
rect 1148 30189 1268 30203
rect 1148 30135 1192 30189
rect 1226 30135 1268 30189
rect 1148 30117 1268 30135
rect 1148 30067 1192 30117
rect 1226 30067 1268 30117
rect 1148 30045 1268 30067
rect 1148 29999 1192 30045
rect 1226 29999 1268 30045
rect 1148 29973 1268 29999
rect 1148 29931 1192 29973
rect 1226 29931 1268 29973
rect 1148 29901 1268 29931
rect 1148 29863 1192 29901
rect 1226 29863 1268 29901
rect 1148 29829 1268 29863
rect 1148 29795 1192 29829
rect 1226 29795 1268 29829
rect 1148 29761 1268 29795
rect 1148 29723 1192 29761
rect 1226 29723 1268 29761
rect 1148 29693 1268 29723
rect 1148 29651 1192 29693
rect 1226 29651 1268 29693
rect 1148 29625 1268 29651
rect 1148 29579 1192 29625
rect 1226 29579 1268 29625
rect 1148 29557 1268 29579
rect 1148 29507 1192 29557
rect 1226 29507 1268 29557
rect 1148 29489 1268 29507
rect 1148 29435 1192 29489
rect 1226 29435 1268 29489
rect 1148 29421 1268 29435
rect 1148 29363 1192 29421
rect 1226 29363 1268 29421
rect 1148 29353 1268 29363
rect 1148 29291 1192 29353
rect 1226 29291 1268 29353
rect 1148 29285 1268 29291
rect 1148 29219 1192 29285
rect 1226 29219 1268 29285
rect 1148 29217 1268 29219
rect 1148 29183 1192 29217
rect 1226 29183 1268 29217
rect 1148 29181 1268 29183
rect 1148 29115 1192 29181
rect 1226 29115 1268 29181
rect 1148 29109 1268 29115
rect 1148 29047 1192 29109
rect 1226 29047 1268 29109
rect 1148 29037 1268 29047
rect 1148 28979 1192 29037
rect 1226 28979 1268 29037
rect 1148 28965 1268 28979
rect 1148 28911 1192 28965
rect 1226 28911 1268 28965
rect 1148 28893 1268 28911
rect 1148 28843 1192 28893
rect 1226 28843 1268 28893
rect 1148 28821 1268 28843
rect 1148 28775 1192 28821
rect 1226 28775 1268 28821
rect 1148 28749 1268 28775
rect 1148 28707 1192 28749
rect 1226 28707 1268 28749
rect 1148 28677 1268 28707
rect 1148 28639 1192 28677
rect 1226 28639 1268 28677
rect 1148 28605 1268 28639
rect 1148 28571 1192 28605
rect 1226 28571 1268 28605
rect 1148 28537 1268 28571
rect 1148 28499 1192 28537
rect 1226 28499 1268 28537
rect 1148 28469 1268 28499
rect 1148 28427 1192 28469
rect 1226 28427 1268 28469
rect 1148 28401 1268 28427
rect 1148 28355 1192 28401
rect 1226 28355 1268 28401
rect 1148 28333 1268 28355
rect 1148 28283 1192 28333
rect 1226 28283 1268 28333
rect 1148 28265 1268 28283
rect 1148 28211 1192 28265
rect 1226 28211 1268 28265
rect 1148 28197 1268 28211
rect 1148 28139 1192 28197
rect 1226 28139 1268 28197
rect 1148 28129 1268 28139
rect 1148 28067 1192 28129
rect 1226 28067 1268 28129
rect 1148 28061 1268 28067
rect 1148 27995 1192 28061
rect 1226 27995 1268 28061
rect 1148 27993 1268 27995
rect 1148 27959 1192 27993
rect 1226 27959 1268 27993
rect 1148 27957 1268 27959
rect 1148 27891 1192 27957
rect 1226 27891 1268 27957
rect 1148 27885 1268 27891
rect 1148 27823 1192 27885
rect 1226 27823 1268 27885
rect 1148 27813 1268 27823
rect 1148 27755 1192 27813
rect 1226 27755 1268 27813
rect 1148 27741 1268 27755
rect 1148 27687 1192 27741
rect 1226 27687 1268 27741
rect 1148 27669 1268 27687
rect 1148 27619 1192 27669
rect 1226 27619 1268 27669
rect 1148 27597 1268 27619
rect 1148 27551 1192 27597
rect 1226 27551 1268 27597
rect 1148 27525 1268 27551
rect 1148 27483 1192 27525
rect 1226 27483 1268 27525
rect 1148 27453 1268 27483
rect 1148 27415 1192 27453
rect 1226 27415 1268 27453
rect 1148 27381 1268 27415
rect 1148 27347 1192 27381
rect 1226 27347 1268 27381
rect 1148 27313 1268 27347
rect 1148 27275 1192 27313
rect 1226 27275 1268 27313
rect 1148 27245 1268 27275
rect 1148 27203 1192 27245
rect 1226 27203 1268 27245
rect 1148 27177 1268 27203
rect 1148 27131 1192 27177
rect 1226 27131 1268 27177
rect 1148 27109 1268 27131
rect 1148 27059 1192 27109
rect 1226 27059 1268 27109
rect 1148 27041 1268 27059
rect 1148 26987 1192 27041
rect 1226 26987 1268 27041
rect 1659 31349 13357 31379
rect 1659 31345 2119 31349
rect 12897 31345 13357 31349
rect 1659 31023 1982 31345
rect 13032 31023 13357 31345
rect 1659 30975 2119 31023
rect 12897 30975 13357 31023
rect 1659 30948 13357 30975
rect 1659 30915 1726 30948
rect 1976 30945 13357 30948
rect 1976 30915 2093 30945
rect 1659 27481 1689 30915
rect 2063 27481 2093 30915
rect 12923 30941 13357 30945
rect 12923 30915 13031 30941
rect 13281 30915 13357 30941
rect 2156 30636 12840 30838
rect 2156 30222 2382 30636
rect 12614 30222 12840 30636
rect 2156 30020 12840 30222
rect 2156 29606 2382 30020
rect 12614 29606 12840 30020
rect 2156 29404 12840 29606
rect 2156 28990 2382 29404
rect 12614 28990 12840 29404
rect 2156 28788 12840 28990
rect 2156 28374 2382 28788
rect 12614 28374 12840 28788
rect 2156 28172 12840 28374
rect 2156 27758 2382 28172
rect 12614 27758 12840 28172
rect 2156 27556 12840 27758
rect 1659 27458 1726 27481
rect 1976 27458 2093 27481
rect 1659 27451 2093 27458
rect 12923 27481 12953 30915
rect 13327 27481 13357 30915
rect 12923 27451 13031 27481
rect 13281 27451 13357 27481
rect 1659 27421 13357 27451
rect 1659 27334 2119 27421
rect 12897 27334 13357 27421
rect 1659 27084 1985 27334
rect 13035 27084 13357 27334
rect 1659 27047 2119 27084
rect 12897 27047 13357 27084
rect 1659 27017 13357 27047
rect 13724 31372 13768 31412
rect 13802 31372 13844 31412
rect 13724 31338 13844 31372
rect 13724 31304 13768 31338
rect 13802 31304 13844 31338
rect 13724 31270 13844 31304
rect 13724 31236 13768 31270
rect 13802 31236 13844 31270
rect 13724 31202 13844 31236
rect 13724 31168 13768 31202
rect 13802 31168 13844 31202
rect 13724 31134 13844 31168
rect 13724 31100 13768 31134
rect 13802 31100 13844 31134
rect 13724 31066 13844 31100
rect 13724 31032 13768 31066
rect 13802 31032 13844 31066
rect 13724 30998 13844 31032
rect 13724 30964 13768 30998
rect 13802 30964 13844 30998
rect 13724 30930 13844 30964
rect 13724 30896 13768 30930
rect 13802 30896 13844 30930
rect 13724 30862 13844 30896
rect 13724 30828 13768 30862
rect 13802 30828 13844 30862
rect 13724 30794 13844 30828
rect 13724 30760 13768 30794
rect 13802 30760 13844 30794
rect 13724 30726 13844 30760
rect 13724 30692 13768 30726
rect 13802 30692 13844 30726
rect 13724 30658 13844 30692
rect 13724 30624 13768 30658
rect 13802 30624 13844 30658
rect 13724 30590 13844 30624
rect 13724 30556 13768 30590
rect 13802 30556 13844 30590
rect 13724 30522 13844 30556
rect 13724 30488 13768 30522
rect 13802 30488 13844 30522
rect 13724 30454 13844 30488
rect 13724 30420 13768 30454
rect 13802 30420 13844 30454
rect 13724 30386 13844 30420
rect 13724 30352 13768 30386
rect 13802 30352 13844 30386
rect 13724 30318 13844 30352
rect 13724 30284 13768 30318
rect 13802 30284 13844 30318
rect 13724 30250 13844 30284
rect 13724 30216 13768 30250
rect 13802 30216 13844 30250
rect 13724 30182 13844 30216
rect 13724 30148 13768 30182
rect 13802 30148 13844 30182
rect 13724 30114 13844 30148
rect 13724 30080 13768 30114
rect 13802 30080 13844 30114
rect 13724 30046 13844 30080
rect 13724 30012 13768 30046
rect 13802 30012 13844 30046
rect 13724 29978 13844 30012
rect 13724 29944 13768 29978
rect 13802 29944 13844 29978
rect 13724 29910 13844 29944
rect 13724 29876 13768 29910
rect 13802 29876 13844 29910
rect 13724 29842 13844 29876
rect 13724 29808 13768 29842
rect 13802 29808 13844 29842
rect 13724 29774 13844 29808
rect 13724 29740 13768 29774
rect 13802 29740 13844 29774
rect 13724 29706 13844 29740
rect 13724 29672 13768 29706
rect 13802 29672 13844 29706
rect 13724 29638 13844 29672
rect 13724 29604 13768 29638
rect 13802 29604 13844 29638
rect 13724 29570 13844 29604
rect 13724 29536 13768 29570
rect 13802 29536 13844 29570
rect 13724 29502 13844 29536
rect 13724 29468 13768 29502
rect 13802 29468 13844 29502
rect 13724 29434 13844 29468
rect 13724 29400 13768 29434
rect 13802 29400 13844 29434
rect 13724 29366 13844 29400
rect 13724 29332 13768 29366
rect 13802 29332 13844 29366
rect 13724 29298 13844 29332
rect 13724 29264 13768 29298
rect 13802 29264 13844 29298
rect 13724 29230 13844 29264
rect 13724 29196 13768 29230
rect 13802 29196 13844 29230
rect 13724 29162 13844 29196
rect 13724 29128 13768 29162
rect 13802 29128 13844 29162
rect 13724 29094 13844 29128
rect 13724 29060 13768 29094
rect 13802 29060 13844 29094
rect 13724 29026 13844 29060
rect 13724 28992 13768 29026
rect 13802 28992 13844 29026
rect 13724 28958 13844 28992
rect 13724 28924 13768 28958
rect 13802 28924 13844 28958
rect 13724 28890 13844 28924
rect 13724 28856 13768 28890
rect 13802 28856 13844 28890
rect 13724 28822 13844 28856
rect 13724 28788 13768 28822
rect 13802 28788 13844 28822
rect 13724 28754 13844 28788
rect 13724 28720 13768 28754
rect 13802 28720 13844 28754
rect 13724 28686 13844 28720
rect 13724 28652 13768 28686
rect 13802 28652 13844 28686
rect 13724 28618 13844 28652
rect 13724 28584 13768 28618
rect 13802 28584 13844 28618
rect 13724 28550 13844 28584
rect 13724 28516 13768 28550
rect 13802 28516 13844 28550
rect 13724 28482 13844 28516
rect 13724 28448 13768 28482
rect 13802 28448 13844 28482
rect 13724 28414 13844 28448
rect 13724 28380 13768 28414
rect 13802 28380 13844 28414
rect 13724 28346 13844 28380
rect 13724 28312 13768 28346
rect 13802 28312 13844 28346
rect 13724 28278 13844 28312
rect 13724 28244 13768 28278
rect 13802 28244 13844 28278
rect 13724 28210 13844 28244
rect 13724 28176 13768 28210
rect 13802 28176 13844 28210
rect 13724 28142 13844 28176
rect 13724 28108 13768 28142
rect 13802 28108 13844 28142
rect 13724 28074 13844 28108
rect 13724 28040 13768 28074
rect 13802 28040 13844 28074
rect 13724 28006 13844 28040
rect 13724 27972 13768 28006
rect 13802 27972 13844 28006
rect 13724 27938 13844 27972
rect 13724 27904 13768 27938
rect 13802 27904 13844 27938
rect 13724 27870 13844 27904
rect 13724 27836 13768 27870
rect 13802 27836 13844 27870
rect 13724 27802 13844 27836
rect 13724 27768 13768 27802
rect 13802 27768 13844 27802
rect 13724 27734 13844 27768
rect 13724 27700 13768 27734
rect 13802 27700 13844 27734
rect 13724 27666 13844 27700
rect 13724 27632 13768 27666
rect 13802 27632 13844 27666
rect 13724 27598 13844 27632
rect 13724 27564 13768 27598
rect 13802 27564 13844 27598
rect 13724 27530 13844 27564
rect 13724 27496 13768 27530
rect 13802 27496 13844 27530
rect 13724 27462 13844 27496
rect 13724 27428 13768 27462
rect 13802 27428 13844 27462
rect 13724 27394 13844 27428
rect 13724 27360 13768 27394
rect 13802 27360 13844 27394
rect 13724 27326 13844 27360
rect 13724 27292 13768 27326
rect 13802 27292 13844 27326
rect 13724 27258 13844 27292
rect 13724 27224 13768 27258
rect 13802 27224 13844 27258
rect 13724 27190 13844 27224
rect 13724 27156 13768 27190
rect 13802 27156 13844 27190
rect 13724 27122 13844 27156
rect 13724 27088 13768 27122
rect 13802 27088 13844 27122
rect 13724 27054 13844 27088
rect 13724 27020 13768 27054
rect 13802 27020 13844 27054
rect 1148 26973 1268 26987
rect 1148 26915 1192 26973
rect 1226 26915 1268 26973
rect 1148 26905 1268 26915
rect 1148 26843 1192 26905
rect 1226 26843 1268 26905
rect 1148 26837 1268 26843
rect 1148 26771 1192 26837
rect 1226 26771 1268 26837
rect 1148 26769 1268 26771
rect 1148 26735 1192 26769
rect 1226 26735 1268 26769
rect 1148 26733 1268 26735
rect 1148 26667 1192 26733
rect 1226 26667 1268 26733
rect 13724 26986 13844 27020
rect 13724 26952 13768 26986
rect 13802 26952 13844 26986
rect 13724 26918 13844 26952
rect 13724 26884 13768 26918
rect 13802 26884 13844 26918
rect 13724 26850 13844 26884
rect 13724 26816 13768 26850
rect 13802 26816 13844 26850
rect 13724 26782 13844 26816
rect 13724 26748 13768 26782
rect 13802 26748 13844 26782
rect 13724 26714 13844 26748
rect 13724 26680 13768 26714
rect 13802 26680 13844 26714
rect 13724 26673 13844 26680
rect 1148 26661 1268 26667
rect 1148 26599 1192 26661
rect 1226 26599 1268 26661
rect 1148 26589 1268 26599
rect 1148 26531 1192 26589
rect 1226 26531 1268 26589
rect 1148 26517 1268 26531
rect 1148 26463 1192 26517
rect 1226 26463 1268 26517
rect 1148 26445 1268 26463
rect 1148 26395 1192 26445
rect 1226 26395 1268 26445
rect 1148 26373 1268 26395
rect 1148 26327 1192 26373
rect 1226 26327 1268 26373
rect 1148 26301 1268 26327
rect 1148 26259 1192 26301
rect 1226 26259 1268 26301
rect 1148 26229 1268 26259
rect 1148 26191 1192 26229
rect 1226 26191 1268 26229
rect 1148 26157 1268 26191
rect 1148 26123 1192 26157
rect 1226 26123 1268 26157
rect 1148 26089 1268 26123
rect 1148 26051 1192 26089
rect 1226 26051 1268 26089
rect 1148 26021 1268 26051
rect 1148 25979 1192 26021
rect 1226 25979 1268 26021
rect 1148 25953 1268 25979
rect 1148 25907 1192 25953
rect 1226 25907 1268 25953
rect 1148 25885 1268 25907
rect 1148 25835 1192 25885
rect 1226 25835 1268 25885
rect 1148 25817 1268 25835
rect 1148 25763 1192 25817
rect 1226 25763 1268 25817
rect 1148 25749 1268 25763
rect 1148 25691 1192 25749
rect 1226 25691 1268 25749
rect 1148 25681 1268 25691
rect 1148 25619 1192 25681
rect 1226 25619 1268 25681
rect 1148 25613 1268 25619
rect 1148 25547 1192 25613
rect 1226 25547 1268 25613
rect 1148 25545 1268 25547
rect 1148 25511 1192 25545
rect 1226 25511 1268 25545
rect 1148 25509 1268 25511
rect 1148 25443 1192 25509
rect 1226 25443 1268 25509
rect 1148 25437 1268 25443
rect 1148 25375 1192 25437
rect 1226 25375 1268 25437
rect 1148 25365 1268 25375
rect 1148 25307 1192 25365
rect 1226 25307 1268 25365
rect 1148 25293 1268 25307
rect 1148 25239 1192 25293
rect 1226 25239 1268 25293
rect 1148 25221 1268 25239
rect 1148 25171 1192 25221
rect 1226 25171 1268 25221
rect 1148 25149 1268 25171
rect 1148 25103 1192 25149
rect 1226 25103 1268 25149
rect 1148 25077 1268 25103
rect 1148 25035 1192 25077
rect 1226 25035 1268 25077
rect 1148 25005 1268 25035
rect 1148 24967 1192 25005
rect 1226 24967 1268 25005
rect 1148 24933 1268 24967
rect 1148 24899 1192 24933
rect 1226 24899 1268 24933
rect 1148 24865 1268 24899
rect 1148 24827 1192 24865
rect 1226 24827 1268 24865
rect 1148 24797 1268 24827
rect 1148 24755 1192 24797
rect 1226 24755 1268 24797
rect 1148 24729 1268 24755
rect 1148 24683 1192 24729
rect 1226 24683 1268 24729
rect 1148 24661 1268 24683
rect 1148 24611 1192 24661
rect 1226 24611 1268 24661
rect 1148 24593 1268 24611
rect 1148 24539 1192 24593
rect 1226 24539 1268 24593
rect 1148 24525 1268 24539
rect 1148 24467 1192 24525
rect 1226 24467 1268 24525
rect 1148 24457 1268 24467
rect 1148 24395 1192 24457
rect 1226 24395 1268 24457
rect 1148 24389 1268 24395
rect 1148 24323 1192 24389
rect 1226 24323 1268 24389
rect 1148 24321 1268 24323
rect 1148 24287 1192 24321
rect 1226 24287 1268 24321
rect 1148 24285 1268 24287
rect 1148 24219 1192 24285
rect 1226 24219 1268 24285
rect 1148 24213 1268 24219
rect 1148 24151 1192 24213
rect 1226 24151 1268 24213
rect 1148 24141 1268 24151
rect 1148 24083 1192 24141
rect 1226 24083 1268 24141
rect 1148 24069 1268 24083
rect 1148 24015 1192 24069
rect 1226 24015 1268 24069
rect 1148 23997 1268 24015
rect 1148 23947 1192 23997
rect 1226 23947 1268 23997
rect 1148 23925 1268 23947
rect 1148 23879 1192 23925
rect 1226 23879 1268 23925
rect 1148 23853 1268 23879
rect 1148 23811 1192 23853
rect 1226 23811 1268 23853
rect 1148 23781 1268 23811
rect 1148 23743 1192 23781
rect 1226 23743 1268 23781
rect 1148 23709 1268 23743
rect 1148 23675 1192 23709
rect 1226 23675 1268 23709
rect 1148 23641 1268 23675
rect 1148 23603 1192 23641
rect 1226 23603 1268 23641
rect 1148 23573 1268 23603
rect 1148 23531 1192 23573
rect 1226 23531 1268 23573
rect 1148 23505 1268 23531
rect 1148 23459 1192 23505
rect 1226 23459 1268 23505
rect 1148 23437 1268 23459
rect 1148 23387 1192 23437
rect 1226 23387 1268 23437
rect 1148 23369 1268 23387
rect 1148 23315 1192 23369
rect 1226 23315 1268 23369
rect 1148 23301 1268 23315
rect 1148 23243 1192 23301
rect 1226 23243 1268 23301
rect 1148 23233 1268 23243
rect 1148 23171 1192 23233
rect 1226 23171 1268 23233
rect 1148 23165 1268 23171
rect 1148 23099 1192 23165
rect 1226 23099 1268 23165
rect 1148 23097 1268 23099
rect 1148 23063 1192 23097
rect 1226 23063 1268 23097
rect 1148 23061 1268 23063
rect 1148 22995 1192 23061
rect 1226 22995 1268 23061
rect 1148 22989 1268 22995
rect 1148 22927 1192 22989
rect 1226 22927 1268 22989
rect 1148 22917 1268 22927
rect 1148 22859 1192 22917
rect 1226 22859 1268 22917
rect 1148 22845 1268 22859
rect 1148 22791 1192 22845
rect 1226 22791 1268 22845
rect 1698 26646 13844 26673
rect 1698 26612 13768 26646
rect 13802 26612 13844 26646
rect 1698 26578 13844 26612
rect 1698 26544 13768 26578
rect 13802 26544 13844 26578
rect 1698 26510 13844 26544
rect 1698 26476 13768 26510
rect 13802 26476 13844 26510
rect 1698 26442 13844 26476
rect 1698 26408 13768 26442
rect 13802 26408 13844 26442
rect 1698 26374 13844 26408
rect 1698 26340 13768 26374
rect 13802 26340 13844 26374
rect 1698 26306 13844 26340
rect 1698 26272 13768 26306
rect 13802 26272 13844 26306
rect 1698 26238 13844 26272
rect 1698 26204 13768 26238
rect 13802 26204 13844 26238
rect 1698 26170 13844 26204
rect 1698 26140 13768 26170
rect 1698 23373 2270 26140
rect 12712 26136 13768 26140
rect 13802 26136 13844 26170
rect 12712 26102 13844 26136
rect 12712 26068 13768 26102
rect 13802 26068 13844 26102
rect 12712 26034 13844 26068
rect 12712 26000 13768 26034
rect 13802 26000 13844 26034
rect 12712 25966 13844 26000
rect 12712 25932 13768 25966
rect 13802 25932 13844 25966
rect 12712 25898 13844 25932
rect 12712 25864 13768 25898
rect 13802 25864 13844 25898
rect 12712 25830 13844 25864
rect 12712 25796 13768 25830
rect 13802 25796 13844 25830
rect 12712 25762 13844 25796
rect 12712 25728 13768 25762
rect 13802 25728 13844 25762
rect 12712 25694 13844 25728
rect 12712 25660 13768 25694
rect 13802 25660 13844 25694
rect 2398 25480 12594 25660
rect 12712 25626 13844 25660
rect 12712 25592 13768 25626
rect 13802 25592 13844 25626
rect 12712 25558 13844 25592
rect 12712 25524 13768 25558
rect 13802 25524 13844 25558
rect 12712 25490 13844 25524
rect 12712 25456 13768 25490
rect 13802 25456 13844 25490
rect 12712 25422 13844 25456
rect 12712 25388 13768 25422
rect 13802 25388 13844 25422
rect 12712 25354 13844 25388
rect 12712 25320 13768 25354
rect 13802 25320 13844 25354
rect 12712 25286 13844 25320
rect 12712 25252 13768 25286
rect 13802 25252 13844 25286
rect 12712 25218 13844 25252
rect 12712 25184 13768 25218
rect 13802 25184 13844 25218
rect 12712 25150 13844 25184
rect 2398 24948 12594 25128
rect 12712 25116 13768 25150
rect 13802 25116 13844 25150
rect 12712 25082 13844 25116
rect 12712 25048 13768 25082
rect 13802 25048 13844 25082
rect 12712 25014 13844 25048
rect 12712 24980 13768 25014
rect 13802 24980 13844 25014
rect 12712 24946 13844 24980
rect 12712 24912 13768 24946
rect 13802 24912 13844 24946
rect 12712 24878 13844 24912
rect 12712 24844 13768 24878
rect 13802 24844 13844 24878
rect 12712 24810 13844 24844
rect 12712 24776 13768 24810
rect 13802 24776 13844 24810
rect 12712 24742 13844 24776
rect 12712 24708 13768 24742
rect 13802 24708 13844 24742
rect 12712 24674 13844 24708
rect 12712 24640 13768 24674
rect 13802 24640 13844 24674
rect 12712 24606 13844 24640
rect 2398 24416 12594 24596
rect 12712 24572 13768 24606
rect 13802 24572 13844 24606
rect 12712 24538 13844 24572
rect 12712 24504 13768 24538
rect 13802 24504 13844 24538
rect 12712 24470 13844 24504
rect 12712 24436 13768 24470
rect 13802 24436 13844 24470
rect 12712 24402 13844 24436
rect 12712 24368 13768 24402
rect 13802 24368 13844 24402
rect 12712 24334 13844 24368
rect 12712 24300 13768 24334
rect 13802 24300 13844 24334
rect 12712 24266 13844 24300
rect 12712 24232 13768 24266
rect 13802 24232 13844 24266
rect 12712 24198 13844 24232
rect 12712 24164 13768 24198
rect 13802 24164 13844 24198
rect 12712 24130 13844 24164
rect 12712 24096 13768 24130
rect 13802 24096 13844 24130
rect 2398 23884 12594 24064
rect 12712 24062 13844 24096
rect 12712 24028 13768 24062
rect 13802 24028 13844 24062
rect 12712 23994 13844 24028
rect 12712 23960 13768 23994
rect 13802 23960 13844 23994
rect 12712 23926 13844 23960
rect 12712 23892 13768 23926
rect 13802 23892 13844 23926
rect 12712 23858 13844 23892
rect 12712 23824 13768 23858
rect 13802 23824 13844 23858
rect 12712 23790 13844 23824
rect 12712 23756 13768 23790
rect 13802 23756 13844 23790
rect 12712 23722 13844 23756
rect 12712 23688 13768 23722
rect 13802 23688 13844 23722
rect 12712 23654 13844 23688
rect 12712 23620 13768 23654
rect 13802 23620 13844 23654
rect 12712 23586 13844 23620
rect 12712 23552 13768 23586
rect 13802 23552 13844 23586
rect 12712 23518 13844 23552
rect 12712 23484 13768 23518
rect 13802 23484 13844 23518
rect 12712 23450 13844 23484
rect 12712 23416 13768 23450
rect 13802 23416 13844 23450
rect 12712 23382 13844 23416
rect 12712 23373 13768 23382
rect 1698 23348 13768 23373
rect 13802 23348 13844 23382
rect 1698 23314 13844 23348
rect 1698 23280 13768 23314
rect 13802 23280 13844 23314
rect 1698 23246 13844 23280
rect 1698 23212 13768 23246
rect 13802 23212 13844 23246
rect 1698 23178 13844 23212
rect 1698 23144 13768 23178
rect 13802 23144 13844 23178
rect 1698 23110 13844 23144
rect 1698 23076 13768 23110
rect 13802 23076 13844 23110
rect 1698 23042 13844 23076
rect 1698 23008 13768 23042
rect 13802 23008 13844 23042
rect 1698 22974 13844 23008
rect 1698 22940 13768 22974
rect 13802 22940 13844 22974
rect 1698 22906 13844 22940
rect 1698 22872 13768 22906
rect 13802 22872 13844 22906
rect 1698 22840 13844 22872
rect 1148 22773 1268 22791
rect 1148 22723 1192 22773
rect 1226 22723 1268 22773
rect 1148 22701 1268 22723
rect 1148 22655 1192 22701
rect 1226 22655 1268 22701
rect 1148 22629 1268 22655
rect 1148 22587 1192 22629
rect 1226 22587 1268 22629
rect 1148 22557 1268 22587
rect 1148 22519 1192 22557
rect 1226 22519 1268 22557
rect 1148 22485 1268 22519
rect 1148 22451 1192 22485
rect 1226 22451 1268 22485
rect 1148 22417 1268 22451
rect 1148 22379 1192 22417
rect 1226 22379 1268 22417
rect 1148 22349 1268 22379
rect 1148 22307 1192 22349
rect 1226 22307 1268 22349
rect 1148 22281 1268 22307
rect 1148 22235 1192 22281
rect 1226 22235 1268 22281
rect 1148 22213 1268 22235
rect 1148 22163 1192 22213
rect 1226 22163 1268 22213
rect 1148 22145 1268 22163
rect 1148 22091 1192 22145
rect 1226 22091 1268 22145
rect 1148 22077 1268 22091
rect 1148 22019 1192 22077
rect 1226 22019 1268 22077
rect 1148 22009 1268 22019
rect 1148 21947 1192 22009
rect 1226 21947 1268 22009
rect 1148 21941 1268 21947
rect 1148 21875 1192 21941
rect 1226 21875 1268 21941
rect 1148 21873 1268 21875
rect 1148 21839 1192 21873
rect 1226 21839 1268 21873
rect 1148 21837 1268 21839
rect 1148 21771 1192 21837
rect 1226 21771 1268 21837
rect 1148 21765 1268 21771
rect 1148 21703 1192 21765
rect 1226 21703 1268 21765
rect 1148 21693 1268 21703
rect 1148 21635 1192 21693
rect 1226 21635 1268 21693
rect 1148 21621 1268 21635
rect 1148 21567 1192 21621
rect 1226 21567 1268 21621
rect 1148 21549 1268 21567
rect 1148 21499 1192 21549
rect 1226 21499 1268 21549
rect 1148 21477 1268 21499
rect 1148 21431 1192 21477
rect 1226 21431 1268 21477
rect 1148 21405 1268 21431
rect 1148 21363 1192 21405
rect 1226 21363 1268 21405
rect 1148 21333 1268 21363
rect 1148 21295 1192 21333
rect 1226 21295 1268 21333
rect 1148 21261 1268 21295
rect 1148 21227 1192 21261
rect 1226 21227 1268 21261
rect 1148 21193 1268 21227
rect 1148 21155 1192 21193
rect 1226 21155 1268 21193
rect 1148 21125 1268 21155
rect 1148 21083 1192 21125
rect 1226 21083 1268 21125
rect 1148 21057 1268 21083
rect 1148 21011 1192 21057
rect 1226 21011 1268 21057
rect 1148 20989 1268 21011
rect 1148 20939 1192 20989
rect 1226 20939 1268 20989
rect 1148 20921 1268 20939
rect 1148 20867 1192 20921
rect 1226 20867 1268 20921
rect 1148 20853 1268 20867
rect 1148 20795 1192 20853
rect 1226 20795 1268 20853
rect 1148 20785 1268 20795
rect 1148 20723 1192 20785
rect 1226 20723 1268 20785
rect 1148 20717 1268 20723
rect 1148 20651 1192 20717
rect 1226 20651 1268 20717
rect 1148 20649 1268 20651
rect 1148 20615 1192 20649
rect 1226 20615 1268 20649
rect 1148 20613 1268 20615
rect 1148 20547 1192 20613
rect 1226 20547 1268 20613
rect 1148 20541 1268 20547
rect 1148 20479 1192 20541
rect 1226 20479 1268 20541
rect 1148 20469 1268 20479
rect 1148 20411 1192 20469
rect 1226 20411 1268 20469
rect 1148 20397 1268 20411
rect 1148 20343 1192 20397
rect 1226 20343 1268 20397
rect 1148 20325 1268 20343
rect 1148 20275 1192 20325
rect 1226 20275 1268 20325
rect 1148 20253 1268 20275
rect 1148 20207 1192 20253
rect 1226 20207 1268 20253
rect 1148 20181 1268 20207
rect 1148 20139 1192 20181
rect 1226 20139 1268 20181
rect 1148 20109 1268 20139
rect 1148 20071 1192 20109
rect 1226 20071 1268 20109
rect 1148 20037 1268 20071
rect 1148 20003 1192 20037
rect 1226 20003 1268 20037
rect 1148 19969 1268 20003
rect 1148 19931 1192 19969
rect 1226 19931 1268 19969
rect 1148 19901 1268 19931
rect 1148 19859 1192 19901
rect 1226 19859 1268 19901
rect 1148 19833 1268 19859
rect 1148 19787 1192 19833
rect 1226 19787 1268 19833
rect 1148 19765 1268 19787
rect 1148 19715 1192 19765
rect 1226 19715 1268 19765
rect 1148 19697 1268 19715
rect 1148 19643 1192 19697
rect 1226 19643 1268 19697
rect 1148 19629 1268 19643
rect 1148 19571 1192 19629
rect 1226 19571 1268 19629
rect 1148 19561 1268 19571
rect 1148 19499 1192 19561
rect 1226 19499 1268 19561
rect 1148 19493 1268 19499
rect 1148 19427 1192 19493
rect 1226 19427 1268 19493
rect 1148 19425 1268 19427
rect 1148 19391 1192 19425
rect 1226 19391 1268 19425
rect 1148 19389 1268 19391
rect 1148 19323 1192 19389
rect 1226 19323 1268 19389
rect 1148 19317 1268 19323
rect 1148 19255 1192 19317
rect 1226 19255 1268 19317
rect 1148 19245 1268 19255
rect 1148 19187 1192 19245
rect 1226 19187 1268 19245
rect 1148 19173 1268 19187
rect 1148 19119 1192 19173
rect 1226 19119 1268 19173
rect 1148 19101 1268 19119
rect 1148 19051 1192 19101
rect 1226 19051 1268 19101
rect 1148 19029 1268 19051
rect 1148 18983 1192 19029
rect 1226 18983 1268 19029
rect 1148 18957 1268 18983
rect 1148 18915 1192 18957
rect 1226 18915 1268 18957
rect 1148 18885 1268 18915
rect 1148 18847 1192 18885
rect 1226 18847 1268 18885
rect 1148 18813 1268 18847
rect 1148 18779 1192 18813
rect 1226 18779 1268 18813
rect 1148 18745 1268 18779
rect 1148 18707 1192 18745
rect 1226 18707 1268 18745
rect 1148 18677 1268 18707
rect 1148 18635 1192 18677
rect 1226 18635 1268 18677
rect 1148 18609 1268 18635
rect 1148 18563 1192 18609
rect 1226 18563 1268 18609
rect 1148 18541 1268 18563
rect 1148 18491 1192 18541
rect 1226 18491 1268 18541
rect 1148 18473 1268 18491
rect 1148 18419 1192 18473
rect 1226 18419 1268 18473
rect 1148 18405 1268 18419
rect 1148 18347 1192 18405
rect 1226 18347 1268 18405
rect 1148 18337 1268 18347
rect 1148 18275 1192 18337
rect 1226 18275 1268 18337
rect 1148 18269 1268 18275
rect 1148 18203 1192 18269
rect 1226 18203 1268 18269
rect 1148 18201 1268 18203
rect 1148 18167 1192 18201
rect 1226 18167 1268 18201
rect 1148 18165 1268 18167
rect 1148 18099 1192 18165
rect 1226 18099 1268 18165
rect 1148 18093 1268 18099
rect 1148 18031 1192 18093
rect 1226 18031 1268 18093
rect 1148 18021 1268 18031
rect 1148 17963 1192 18021
rect 1226 17963 1268 18021
rect 1148 17949 1268 17963
rect 1148 17895 1192 17949
rect 1226 17895 1268 17949
rect 1148 17877 1268 17895
rect 1148 17827 1192 17877
rect 1226 17827 1268 17877
rect 1148 17805 1268 17827
rect 1148 17759 1192 17805
rect 1226 17759 1268 17805
rect 1148 17733 1268 17759
rect 1148 17691 1192 17733
rect 1226 17691 1268 17733
rect 1148 17661 1268 17691
rect 1148 17623 1192 17661
rect 1226 17623 1268 17661
rect 1148 17589 1268 17623
rect 1148 17555 1192 17589
rect 1226 17555 1268 17589
rect 1148 17521 1268 17555
rect 1148 17483 1192 17521
rect 1226 17483 1268 17521
rect 1148 17453 1268 17483
rect 1148 17411 1192 17453
rect 1226 17411 1268 17453
rect 1148 17385 1268 17411
rect 1148 17339 1192 17385
rect 1226 17339 1268 17385
rect 1148 17317 1268 17339
rect 1148 17267 1192 17317
rect 1226 17267 1268 17317
rect 1148 17249 1268 17267
rect 1148 17195 1192 17249
rect 1226 17195 1268 17249
rect 1148 17181 1268 17195
rect 1148 17123 1192 17181
rect 1226 17123 1268 17181
rect 1148 17113 1268 17123
rect 1148 17051 1192 17113
rect 1226 17051 1268 17113
rect 1148 17045 1268 17051
rect 1148 16979 1192 17045
rect 1226 16979 1268 17045
rect 1148 16977 1268 16979
rect 1148 16943 1192 16977
rect 1226 16943 1268 16977
rect 1148 16941 1268 16943
rect 1148 16875 1192 16941
rect 1226 16875 1268 16941
rect 1148 16869 1268 16875
rect 1148 16807 1192 16869
rect 1226 16807 1268 16869
rect 1148 16797 1268 16807
rect 1148 16739 1192 16797
rect 1226 16739 1268 16797
rect 1148 16725 1268 16739
rect 1148 16671 1192 16725
rect 1226 16671 1268 16725
rect 1148 16653 1268 16671
rect 1148 16603 1192 16653
rect 1226 16603 1268 16653
rect 1148 16581 1268 16603
rect 1148 16535 1192 16581
rect 1226 16535 1268 16581
rect 1148 16509 1268 16535
rect 1148 16467 1192 16509
rect 1226 16467 1268 16509
rect 1148 16437 1268 16467
rect 1148 16399 1192 16437
rect 1226 16399 1268 16437
rect 1148 16365 1268 16399
rect 1148 16331 1192 16365
rect 1226 16331 1268 16365
rect 1148 16297 1268 16331
rect 1148 16259 1192 16297
rect 1226 16259 1268 16297
rect 1148 16229 1268 16259
rect 1148 16187 1192 16229
rect 1226 16187 1268 16229
rect 1148 16161 1268 16187
rect 1148 16115 1192 16161
rect 1226 16115 1268 16161
rect 1148 16093 1268 16115
rect 1148 16043 1192 16093
rect 1226 16043 1268 16093
rect 1148 16025 1268 16043
rect 1148 15971 1192 16025
rect 1226 15971 1268 16025
rect 1148 15957 1268 15971
rect 1148 15899 1192 15957
rect 1226 15899 1268 15957
rect 1148 15889 1268 15899
rect 1148 15827 1192 15889
rect 1226 15827 1268 15889
rect 1148 15821 1268 15827
rect 1148 15755 1192 15821
rect 1226 15755 1268 15821
rect 1148 15753 1268 15755
rect 1148 15719 1192 15753
rect 1226 15719 1268 15753
rect 1148 15717 1268 15719
rect 1148 15651 1192 15717
rect 1226 15651 1268 15717
rect 1148 15645 1268 15651
rect 1148 15583 1192 15645
rect 1226 15583 1268 15645
rect 1148 15573 1268 15583
rect 1148 15515 1192 15573
rect 1226 15515 1268 15573
rect 1148 15501 1268 15515
rect 1148 15447 1192 15501
rect 1226 15447 1268 15501
rect 1148 15429 1268 15447
rect 1148 15379 1192 15429
rect 1226 15379 1268 15429
rect 1148 15357 1268 15379
rect 1148 15311 1192 15357
rect 1226 15311 1268 15357
rect 1148 15285 1268 15311
rect 1148 15243 1192 15285
rect 1226 15243 1268 15285
rect 1148 15213 1268 15243
rect 1148 15175 1192 15213
rect 1226 15175 1268 15213
rect 1148 15141 1268 15175
rect 1148 15107 1192 15141
rect 1226 15107 1268 15141
rect 1148 15073 1268 15107
rect 1148 15035 1192 15073
rect 1226 15035 1268 15073
rect 1148 15005 1268 15035
rect 1148 14963 1192 15005
rect 1226 14963 1268 15005
rect 1148 14937 1268 14963
rect 1148 14891 1192 14937
rect 1226 14891 1268 14937
rect 1148 14869 1268 14891
rect 1148 14819 1192 14869
rect 1226 14819 1268 14869
rect 1148 14801 1268 14819
rect 1148 14747 1192 14801
rect 1226 14747 1268 14801
rect 1148 14733 1268 14747
rect 1148 14675 1192 14733
rect 1226 14675 1268 14733
rect 1148 14665 1268 14675
rect 1148 14603 1192 14665
rect 1226 14603 1268 14665
rect 1148 14597 1268 14603
rect 1148 14531 1192 14597
rect 1226 14531 1268 14597
rect 1148 14529 1268 14531
rect 1148 14495 1192 14529
rect 1226 14495 1268 14529
rect 1148 14493 1268 14495
rect 1148 14427 1192 14493
rect 1226 14427 1268 14493
rect 1148 14421 1268 14427
rect 1148 14359 1192 14421
rect 1226 14359 1268 14421
rect 1148 14349 1268 14359
rect 1148 14291 1192 14349
rect 1226 14291 1268 14349
rect 1148 14277 1268 14291
rect 1148 14223 1192 14277
rect 1226 14223 1268 14277
rect 1148 14205 1268 14223
rect 1148 14155 1192 14205
rect 1226 14155 1268 14205
rect 1148 14133 1268 14155
rect 1148 14087 1192 14133
rect 1226 14087 1268 14133
rect 1148 14061 1268 14087
rect 1148 14019 1192 14061
rect 1226 14019 1268 14061
rect 1148 13989 1268 14019
rect 1148 13951 1192 13989
rect 1226 13951 1268 13989
rect 1148 13917 1268 13951
rect 1148 13883 1192 13917
rect 1226 13883 1268 13917
rect 1148 13849 1268 13883
rect 1148 13811 1192 13849
rect 1226 13811 1268 13849
rect 1148 13781 1268 13811
rect 1148 13739 1192 13781
rect 1226 13739 1268 13781
rect 1148 13713 1268 13739
rect 1148 13667 1192 13713
rect 1226 13667 1268 13713
rect 1148 13645 1268 13667
rect 1148 13595 1192 13645
rect 1226 13595 1268 13645
rect 1148 13577 1268 13595
rect 1148 13523 1192 13577
rect 1226 13523 1268 13577
rect 1148 13509 1268 13523
rect 1148 13451 1192 13509
rect 1226 13451 1268 13509
rect 1148 13441 1268 13451
rect 1148 13379 1192 13441
rect 1226 13379 1268 13441
rect 1148 13373 1268 13379
rect 1148 13307 1192 13373
rect 1226 13307 1268 13373
rect 1148 13305 1268 13307
rect 1148 13271 1192 13305
rect 1226 13271 1268 13305
rect 1148 13269 1268 13271
rect 1148 13203 1192 13269
rect 1226 13203 1268 13269
rect 1148 13197 1268 13203
rect 1148 13135 1192 13197
rect 1226 13135 1268 13197
rect 1148 13125 1268 13135
rect 1148 13067 1192 13125
rect 1226 13067 1268 13125
rect 1148 13053 1268 13067
rect 1148 12999 1192 13053
rect 1226 12999 1268 13053
rect 1148 12981 1268 12999
rect 1148 12931 1192 12981
rect 1226 12931 1268 12981
rect 1148 12909 1268 12931
rect 1148 12863 1192 12909
rect 1226 12863 1268 12909
rect 1148 12837 1268 12863
rect 1148 12795 1192 12837
rect 1226 12795 1268 12837
rect 1148 12765 1268 12795
rect 1148 12727 1192 12765
rect 1226 12727 1268 12765
rect 1148 12693 1268 12727
rect 1148 12659 1192 12693
rect 1226 12659 1268 12693
rect 1148 12625 1268 12659
rect 1148 12587 1192 12625
rect 1226 12587 1268 12625
rect 1148 12557 1268 12587
rect 1148 12515 1192 12557
rect 1226 12515 1268 12557
rect 1148 12489 1268 12515
rect 1148 12443 1192 12489
rect 1226 12443 1268 12489
rect 1148 12421 1268 12443
rect 1148 12371 1192 12421
rect 1226 12371 1268 12421
rect 1148 12353 1268 12371
rect 1148 12299 1192 12353
rect 1226 12299 1268 12353
rect 1148 12285 1268 12299
rect 1148 12227 1192 12285
rect 1226 12227 1268 12285
rect 1148 12217 1268 12227
rect 1148 12155 1192 12217
rect 1226 12155 1268 12217
rect 1148 12149 1268 12155
rect 1148 12083 1192 12149
rect 1226 12083 1268 12149
rect 1148 12081 1268 12083
rect 1148 12047 1192 12081
rect 1226 12047 1268 12081
rect 1148 12045 1268 12047
rect 1148 11979 1192 12045
rect 1226 11979 1268 12045
rect 1148 11973 1268 11979
rect 1148 11911 1192 11973
rect 1226 11911 1268 11973
rect 1148 11901 1268 11911
rect 1148 11843 1192 11901
rect 1226 11843 1268 11901
rect 1148 11829 1268 11843
rect 1148 11775 1192 11829
rect 1226 11775 1268 11829
rect 1148 11757 1268 11775
rect 1148 11707 1192 11757
rect 1226 11707 1268 11757
rect 1148 11685 1268 11707
rect 1148 11639 1192 11685
rect 1226 11639 1268 11685
rect 1148 11613 1268 11639
rect 1148 11571 1192 11613
rect 1226 11571 1268 11613
rect 1148 11541 1268 11571
rect 1148 11503 1192 11541
rect 1226 11503 1268 11541
rect 1148 11469 1268 11503
rect 1148 11435 1192 11469
rect 1226 11435 1268 11469
rect 1148 11401 1268 11435
rect 1148 11363 1192 11401
rect 1226 11363 1268 11401
rect 1148 11333 1268 11363
rect 1148 11291 1192 11333
rect 1226 11291 1268 11333
rect 1148 11265 1268 11291
rect 1148 11219 1192 11265
rect 1226 11219 1268 11265
rect 1148 11197 1268 11219
rect 1148 11147 1192 11197
rect 1226 11147 1268 11197
rect 1148 11129 1268 11147
rect 1148 11075 1192 11129
rect 1226 11075 1268 11129
rect 1148 11061 1268 11075
rect 1148 11003 1192 11061
rect 1226 11003 1268 11061
rect 1148 10993 1268 11003
rect 1148 10931 1192 10993
rect 1226 10931 1268 10993
rect 1148 10925 1268 10931
rect 1148 10859 1192 10925
rect 1226 10859 1268 10925
rect 1148 10857 1268 10859
rect 1148 10823 1192 10857
rect 1226 10823 1268 10857
rect 1148 10821 1268 10823
rect 1148 10755 1192 10821
rect 1226 10755 1268 10821
rect 1148 10749 1268 10755
rect 1148 10687 1192 10749
rect 1226 10687 1268 10749
rect 1148 10677 1268 10687
rect 1148 10619 1192 10677
rect 1226 10619 1268 10677
rect 1148 10605 1268 10619
rect 1148 10551 1192 10605
rect 1226 10551 1268 10605
rect 1148 10533 1268 10551
rect 1148 10483 1192 10533
rect 1226 10483 1268 10533
rect 1148 10461 1268 10483
rect 1148 10415 1192 10461
rect 1226 10415 1268 10461
rect 1148 10362 1268 10415
rect 13724 22838 13844 22840
rect 13724 22804 13768 22838
rect 13802 22804 13844 22838
rect 13724 22770 13844 22804
rect 13724 22736 13768 22770
rect 13802 22736 13844 22770
rect 13724 22702 13844 22736
rect 13724 22668 13768 22702
rect 13802 22668 13844 22702
rect 13724 22634 13844 22668
rect 13724 22600 13768 22634
rect 13802 22600 13844 22634
rect 13724 22566 13844 22600
rect 13724 22532 13768 22566
rect 13802 22532 13844 22566
rect 13724 22498 13844 22532
rect 13724 22464 13768 22498
rect 13802 22464 13844 22498
rect 13724 22430 13844 22464
rect 13724 22396 13768 22430
rect 13802 22396 13844 22430
rect 13724 22362 13844 22396
rect 13724 22328 13768 22362
rect 13802 22328 13844 22362
rect 13724 22294 13844 22328
rect 13724 22260 13768 22294
rect 13802 22260 13844 22294
rect 13724 22226 13844 22260
rect 13724 22192 13768 22226
rect 13802 22192 13844 22226
rect 13724 22158 13844 22192
rect 13724 22124 13768 22158
rect 13802 22124 13844 22158
rect 13724 22090 13844 22124
rect 13724 22056 13768 22090
rect 13802 22056 13844 22090
rect 13724 22022 13844 22056
rect 13724 21988 13768 22022
rect 13802 21988 13844 22022
rect 13724 21954 13844 21988
rect 13724 21920 13768 21954
rect 13802 21920 13844 21954
rect 13724 21886 13844 21920
rect 13724 21852 13768 21886
rect 13802 21852 13844 21886
rect 13724 21818 13844 21852
rect 13724 21784 13768 21818
rect 13802 21784 13844 21818
rect 13724 21750 13844 21784
rect 13724 21716 13768 21750
rect 13802 21716 13844 21750
rect 13724 21682 13844 21716
rect 13724 21648 13768 21682
rect 13802 21648 13844 21682
rect 13724 21614 13844 21648
rect 13724 21580 13768 21614
rect 13802 21580 13844 21614
rect 13724 21546 13844 21580
rect 13724 21512 13768 21546
rect 13802 21512 13844 21546
rect 13724 21478 13844 21512
rect 13724 21444 13768 21478
rect 13802 21444 13844 21478
rect 13724 21410 13844 21444
rect 13724 21376 13768 21410
rect 13802 21376 13844 21410
rect 13724 21342 13844 21376
rect 13724 21308 13768 21342
rect 13802 21308 13844 21342
rect 13724 21274 13844 21308
rect 13724 21240 13768 21274
rect 13802 21240 13844 21274
rect 13724 21219 13844 21240
rect 13724 21172 13768 21219
rect 13802 21172 13844 21219
rect 13724 21147 13844 21172
rect 13724 21104 13768 21147
rect 13802 21104 13844 21147
rect 13724 21075 13844 21104
rect 13724 21036 13768 21075
rect 13802 21036 13844 21075
rect 13724 21003 13844 21036
rect 13724 20968 13768 21003
rect 13802 20968 13844 21003
rect 13724 20934 13844 20968
rect 13724 20897 13768 20934
rect 13802 20897 13844 20934
rect 13724 20866 13844 20897
rect 13724 20825 13768 20866
rect 13802 20825 13844 20866
rect 13724 20798 13844 20825
rect 13724 20753 13768 20798
rect 13802 20753 13844 20798
rect 13724 20730 13844 20753
rect 13724 20681 13768 20730
rect 13802 20681 13844 20730
rect 13724 20662 13844 20681
rect 13724 20609 13768 20662
rect 13802 20609 13844 20662
rect 13724 20594 13844 20609
rect 13724 20537 13768 20594
rect 13802 20537 13844 20594
rect 13724 20526 13844 20537
rect 13724 20465 13768 20526
rect 13802 20465 13844 20526
rect 13724 20458 13844 20465
rect 13724 20393 13768 20458
rect 13802 20393 13844 20458
rect 13724 20390 13844 20393
rect 13724 20356 13768 20390
rect 13802 20356 13844 20390
rect 13724 20355 13844 20356
rect 13724 20288 13768 20355
rect 13802 20288 13844 20355
rect 13724 20283 13844 20288
rect 13724 20220 13768 20283
rect 13802 20220 13844 20283
rect 13724 20211 13844 20220
rect 13724 20152 13768 20211
rect 13802 20152 13844 20211
rect 13724 20139 13844 20152
rect 13724 20084 13768 20139
rect 13802 20084 13844 20139
rect 13724 20067 13844 20084
rect 13724 20016 13768 20067
rect 13802 20016 13844 20067
rect 13724 19995 13844 20016
rect 13724 19948 13768 19995
rect 13802 19948 13844 19995
rect 13724 19923 13844 19948
rect 13724 19880 13768 19923
rect 13802 19880 13844 19923
rect 13724 19851 13844 19880
rect 13724 19812 13768 19851
rect 13802 19812 13844 19851
rect 13724 19779 13844 19812
rect 13724 19744 13768 19779
rect 13802 19744 13844 19779
rect 13724 19710 13844 19744
rect 13724 19673 13768 19710
rect 13802 19673 13844 19710
rect 13724 19642 13844 19673
rect 13724 19601 13768 19642
rect 13802 19601 13844 19642
rect 13724 19574 13844 19601
rect 13724 19529 13768 19574
rect 13802 19529 13844 19574
rect 13724 19506 13844 19529
rect 13724 19457 13768 19506
rect 13802 19457 13844 19506
rect 13724 19438 13844 19457
rect 13724 19385 13768 19438
rect 13802 19385 13844 19438
rect 13724 19370 13844 19385
rect 13724 19313 13768 19370
rect 13802 19313 13844 19370
rect 13724 19302 13844 19313
rect 13724 19241 13768 19302
rect 13802 19241 13844 19302
rect 13724 19234 13844 19241
rect 13724 19169 13768 19234
rect 13802 19169 13844 19234
rect 13724 19166 13844 19169
rect 13724 19132 13768 19166
rect 13802 19132 13844 19166
rect 13724 19131 13844 19132
rect 13724 19064 13768 19131
rect 13802 19064 13844 19131
rect 13724 19059 13844 19064
rect 13724 18996 13768 19059
rect 13802 18996 13844 19059
rect 13724 18987 13844 18996
rect 13724 18928 13768 18987
rect 13802 18928 13844 18987
rect 13724 18915 13844 18928
rect 13724 18860 13768 18915
rect 13802 18860 13844 18915
rect 13724 18843 13844 18860
rect 13724 18792 13768 18843
rect 13802 18792 13844 18843
rect 13724 18771 13844 18792
rect 13724 18724 13768 18771
rect 13802 18724 13844 18771
rect 13724 18699 13844 18724
rect 13724 18656 13768 18699
rect 13802 18656 13844 18699
rect 13724 18627 13844 18656
rect 13724 18588 13768 18627
rect 13802 18588 13844 18627
rect 13724 18555 13844 18588
rect 13724 18520 13768 18555
rect 13802 18520 13844 18555
rect 13724 18486 13844 18520
rect 13724 18449 13768 18486
rect 13802 18449 13844 18486
rect 13724 18418 13844 18449
rect 13724 18377 13768 18418
rect 13802 18377 13844 18418
rect 13724 18350 13844 18377
rect 13724 18305 13768 18350
rect 13802 18305 13844 18350
rect 13724 18282 13844 18305
rect 13724 18233 13768 18282
rect 13802 18233 13844 18282
rect 13724 18214 13844 18233
rect 13724 18161 13768 18214
rect 13802 18161 13844 18214
rect 13724 18146 13844 18161
rect 13724 18089 13768 18146
rect 13802 18089 13844 18146
rect 13724 18078 13844 18089
rect 13724 18017 13768 18078
rect 13802 18017 13844 18078
rect 13724 18010 13844 18017
rect 13724 17945 13768 18010
rect 13802 17945 13844 18010
rect 13724 17942 13844 17945
rect 13724 17908 13768 17942
rect 13802 17908 13844 17942
rect 13724 17907 13844 17908
rect 13724 17840 13768 17907
rect 13802 17840 13844 17907
rect 13724 17835 13844 17840
rect 13724 17772 13768 17835
rect 13802 17772 13844 17835
rect 13724 17763 13844 17772
rect 13724 17704 13768 17763
rect 13802 17704 13844 17763
rect 13724 17691 13844 17704
rect 13724 17636 13768 17691
rect 13802 17636 13844 17691
rect 13724 17619 13844 17636
rect 13724 17568 13768 17619
rect 13802 17568 13844 17619
rect 13724 17547 13844 17568
rect 13724 17500 13768 17547
rect 13802 17500 13844 17547
rect 13724 17475 13844 17500
rect 13724 17432 13768 17475
rect 13802 17432 13844 17475
rect 13724 17403 13844 17432
rect 13724 17364 13768 17403
rect 13802 17364 13844 17403
rect 13724 17331 13844 17364
rect 13724 17296 13768 17331
rect 13802 17296 13844 17331
rect 13724 17262 13844 17296
rect 13724 17225 13768 17262
rect 13802 17225 13844 17262
rect 13724 17194 13844 17225
rect 13724 17153 13768 17194
rect 13802 17153 13844 17194
rect 13724 17126 13844 17153
rect 13724 17081 13768 17126
rect 13802 17081 13844 17126
rect 13724 17058 13844 17081
rect 13724 17009 13768 17058
rect 13802 17009 13844 17058
rect 13724 16990 13844 17009
rect 13724 16937 13768 16990
rect 13802 16937 13844 16990
rect 13724 16922 13844 16937
rect 13724 16865 13768 16922
rect 13802 16865 13844 16922
rect 13724 16854 13844 16865
rect 13724 16793 13768 16854
rect 13802 16793 13844 16854
rect 13724 16786 13844 16793
rect 13724 16721 13768 16786
rect 13802 16721 13844 16786
rect 13724 16718 13844 16721
rect 13724 16684 13768 16718
rect 13802 16684 13844 16718
rect 13724 16683 13844 16684
rect 13724 16616 13768 16683
rect 13802 16616 13844 16683
rect 13724 16611 13844 16616
rect 13724 16548 13768 16611
rect 13802 16548 13844 16611
rect 13724 16539 13844 16548
rect 13724 16480 13768 16539
rect 13802 16480 13844 16539
rect 13724 16467 13844 16480
rect 13724 16412 13768 16467
rect 13802 16412 13844 16467
rect 13724 16395 13844 16412
rect 13724 16344 13768 16395
rect 13802 16344 13844 16395
rect 13724 16323 13844 16344
rect 13724 16276 13768 16323
rect 13802 16276 13844 16323
rect 13724 16251 13844 16276
rect 13724 16208 13768 16251
rect 13802 16208 13844 16251
rect 13724 16179 13844 16208
rect 13724 16140 13768 16179
rect 13802 16140 13844 16179
rect 13724 16107 13844 16140
rect 13724 16072 13768 16107
rect 13802 16072 13844 16107
rect 13724 16038 13844 16072
rect 13724 16001 13768 16038
rect 13802 16001 13844 16038
rect 13724 15970 13844 16001
rect 13724 15929 13768 15970
rect 13802 15929 13844 15970
rect 13724 15902 13844 15929
rect 13724 15857 13768 15902
rect 13802 15857 13844 15902
rect 13724 15834 13844 15857
rect 13724 15785 13768 15834
rect 13802 15785 13844 15834
rect 13724 15766 13844 15785
rect 13724 15713 13768 15766
rect 13802 15713 13844 15766
rect 13724 15698 13844 15713
rect 13724 15641 13768 15698
rect 13802 15641 13844 15698
rect 13724 15630 13844 15641
rect 13724 15569 13768 15630
rect 13802 15569 13844 15630
rect 13724 15562 13844 15569
rect 13724 15497 13768 15562
rect 13802 15497 13844 15562
rect 13724 15494 13844 15497
rect 13724 15460 13768 15494
rect 13802 15460 13844 15494
rect 13724 15459 13844 15460
rect 13724 15392 13768 15459
rect 13802 15392 13844 15459
rect 13724 15387 13844 15392
rect 13724 15324 13768 15387
rect 13802 15324 13844 15387
rect 13724 15315 13844 15324
rect 13724 15256 13768 15315
rect 13802 15256 13844 15315
rect 13724 15243 13844 15256
rect 13724 15188 13768 15243
rect 13802 15188 13844 15243
rect 13724 15171 13844 15188
rect 13724 15120 13768 15171
rect 13802 15120 13844 15171
rect 13724 15099 13844 15120
rect 13724 15052 13768 15099
rect 13802 15052 13844 15099
rect 13724 15027 13844 15052
rect 13724 14984 13768 15027
rect 13802 14984 13844 15027
rect 13724 14955 13844 14984
rect 13724 14916 13768 14955
rect 13802 14916 13844 14955
rect 13724 14883 13844 14916
rect 13724 14848 13768 14883
rect 13802 14848 13844 14883
rect 13724 14814 13844 14848
rect 13724 14777 13768 14814
rect 13802 14777 13844 14814
rect 13724 14746 13844 14777
rect 13724 14705 13768 14746
rect 13802 14705 13844 14746
rect 13724 14678 13844 14705
rect 13724 14633 13768 14678
rect 13802 14633 13844 14678
rect 13724 14610 13844 14633
rect 13724 14561 13768 14610
rect 13802 14561 13844 14610
rect 13724 14542 13844 14561
rect 13724 14489 13768 14542
rect 13802 14489 13844 14542
rect 13724 14474 13844 14489
rect 13724 14417 13768 14474
rect 13802 14417 13844 14474
rect 13724 14406 13844 14417
rect 13724 14345 13768 14406
rect 13802 14345 13844 14406
rect 13724 14338 13844 14345
rect 13724 14273 13768 14338
rect 13802 14273 13844 14338
rect 13724 14270 13844 14273
rect 13724 14236 13768 14270
rect 13802 14236 13844 14270
rect 13724 14235 13844 14236
rect 13724 14168 13768 14235
rect 13802 14168 13844 14235
rect 13724 14163 13844 14168
rect 13724 14100 13768 14163
rect 13802 14100 13844 14163
rect 13724 14091 13844 14100
rect 13724 14032 13768 14091
rect 13802 14032 13844 14091
rect 13724 14019 13844 14032
rect 13724 13964 13768 14019
rect 13802 13964 13844 14019
rect 13724 13947 13844 13964
rect 13724 13896 13768 13947
rect 13802 13896 13844 13947
rect 13724 13875 13844 13896
rect 13724 13828 13768 13875
rect 13802 13828 13844 13875
rect 13724 13803 13844 13828
rect 13724 13760 13768 13803
rect 13802 13760 13844 13803
rect 13724 13731 13844 13760
rect 13724 13692 13768 13731
rect 13802 13692 13844 13731
rect 13724 13659 13844 13692
rect 13724 13624 13768 13659
rect 13802 13624 13844 13659
rect 13724 13590 13844 13624
rect 13724 13553 13768 13590
rect 13802 13553 13844 13590
rect 13724 13522 13844 13553
rect 13724 13481 13768 13522
rect 13802 13481 13844 13522
rect 13724 13454 13844 13481
rect 13724 13409 13768 13454
rect 13802 13409 13844 13454
rect 13724 13386 13844 13409
rect 13724 13337 13768 13386
rect 13802 13337 13844 13386
rect 13724 13318 13844 13337
rect 13724 13265 13768 13318
rect 13802 13265 13844 13318
rect 13724 13250 13844 13265
rect 13724 13193 13768 13250
rect 13802 13193 13844 13250
rect 13724 13182 13844 13193
rect 13724 13121 13768 13182
rect 13802 13121 13844 13182
rect 13724 13114 13844 13121
rect 13724 13049 13768 13114
rect 13802 13049 13844 13114
rect 13724 13046 13844 13049
rect 13724 13012 13768 13046
rect 13802 13012 13844 13046
rect 13724 13011 13844 13012
rect 13724 12944 13768 13011
rect 13802 12944 13844 13011
rect 13724 12939 13844 12944
rect 13724 12876 13768 12939
rect 13802 12876 13844 12939
rect 13724 12867 13844 12876
rect 13724 12808 13768 12867
rect 13802 12808 13844 12867
rect 13724 12795 13844 12808
rect 13724 12740 13768 12795
rect 13802 12740 13844 12795
rect 13724 12723 13844 12740
rect 13724 12672 13768 12723
rect 13802 12672 13844 12723
rect 13724 12651 13844 12672
rect 13724 12604 13768 12651
rect 13802 12604 13844 12651
rect 13724 12579 13844 12604
rect 13724 12536 13768 12579
rect 13802 12536 13844 12579
rect 13724 12507 13844 12536
rect 13724 12468 13768 12507
rect 13802 12468 13844 12507
rect 13724 12435 13844 12468
rect 13724 12400 13768 12435
rect 13802 12400 13844 12435
rect 13724 12366 13844 12400
rect 13724 12329 13768 12366
rect 13802 12329 13844 12366
rect 13724 12298 13844 12329
rect 13724 12257 13768 12298
rect 13802 12257 13844 12298
rect 13724 12230 13844 12257
rect 13724 12185 13768 12230
rect 13802 12185 13844 12230
rect 13724 12162 13844 12185
rect 13724 12113 13768 12162
rect 13802 12113 13844 12162
rect 13724 12094 13844 12113
rect 13724 12041 13768 12094
rect 13802 12041 13844 12094
rect 13724 12026 13844 12041
rect 13724 11969 13768 12026
rect 13802 11969 13844 12026
rect 13724 11958 13844 11969
rect 13724 11897 13768 11958
rect 13802 11897 13844 11958
rect 13724 11890 13844 11897
rect 13724 11825 13768 11890
rect 13802 11825 13844 11890
rect 13724 11822 13844 11825
rect 13724 11788 13768 11822
rect 13802 11788 13844 11822
rect 13724 11787 13844 11788
rect 13724 11720 13768 11787
rect 13802 11720 13844 11787
rect 13724 11715 13844 11720
rect 13724 11652 13768 11715
rect 13802 11652 13844 11715
rect 13724 11643 13844 11652
rect 13724 11584 13768 11643
rect 13802 11584 13844 11643
rect 13724 11571 13844 11584
rect 13724 11516 13768 11571
rect 13802 11516 13844 11571
rect 13724 11499 13844 11516
rect 13724 11448 13768 11499
rect 13802 11448 13844 11499
rect 13724 11427 13844 11448
rect 13724 11380 13768 11427
rect 13802 11380 13844 11427
rect 13724 11355 13844 11380
rect 13724 11312 13768 11355
rect 13802 11312 13844 11355
rect 13724 11283 13844 11312
rect 13724 11244 13768 11283
rect 13802 11244 13844 11283
rect 13724 11211 13844 11244
rect 13724 11176 13768 11211
rect 13802 11176 13844 11211
rect 13724 11142 13844 11176
rect 13724 11105 13768 11142
rect 13802 11105 13844 11142
rect 13724 11074 13844 11105
rect 13724 11033 13768 11074
rect 13802 11033 13844 11074
rect 13724 11006 13844 11033
rect 13724 10961 13768 11006
rect 13802 10961 13844 11006
rect 13724 10938 13844 10961
rect 13724 10889 13768 10938
rect 13802 10889 13844 10938
rect 13724 10870 13844 10889
rect 13724 10817 13768 10870
rect 13802 10817 13844 10870
rect 13724 10802 13844 10817
rect 13724 10745 13768 10802
rect 13802 10745 13844 10802
rect 13724 10734 13844 10745
rect 13724 10673 13768 10734
rect 13802 10673 13844 10734
rect 13724 10666 13844 10673
rect 13724 10601 13768 10666
rect 13802 10601 13844 10666
rect 13724 10598 13844 10601
rect 13724 10564 13768 10598
rect 13802 10564 13844 10598
rect 13724 10563 13844 10564
rect 13724 10496 13768 10563
rect 13802 10496 13844 10563
rect 13724 10491 13844 10496
rect 13724 10428 13768 10491
rect 13802 10428 13844 10491
rect 13724 10419 13844 10428
rect 13724 10362 13768 10419
rect 1148 10360 13768 10362
rect 13802 10360 13844 10419
rect 1148 10318 13844 10360
rect 1148 10284 1327 10318
rect 1363 10284 1397 10318
rect 1433 10284 1465 10318
rect 1505 10284 1533 10318
rect 1577 10284 1601 10318
rect 1649 10284 1669 10318
rect 1721 10284 1737 10318
rect 1793 10284 1805 10318
rect 1865 10284 1873 10318
rect 1937 10284 1941 10318
rect 2043 10284 2047 10318
rect 2111 10284 2119 10318
rect 2179 10284 2191 10318
rect 2247 10284 2263 10318
rect 2315 10284 2335 10318
rect 2383 10284 2407 10318
rect 2451 10284 2479 10318
rect 2519 10284 2551 10318
rect 2587 10284 2621 10318
rect 2657 10284 2689 10318
rect 2729 10284 2757 10318
rect 2801 10284 2825 10318
rect 2873 10284 2893 10318
rect 2945 10284 2961 10318
rect 3017 10284 3029 10318
rect 3089 10284 3097 10318
rect 3161 10284 3165 10318
rect 3267 10284 3271 10318
rect 3335 10284 3343 10318
rect 3403 10284 3415 10318
rect 3471 10284 3487 10318
rect 3539 10284 3559 10318
rect 3607 10284 3631 10318
rect 3675 10284 3703 10318
rect 3743 10284 3775 10318
rect 3811 10284 3845 10318
rect 3881 10284 3913 10318
rect 3953 10284 3981 10318
rect 4025 10284 4049 10318
rect 4097 10284 4117 10318
rect 4169 10284 4185 10318
rect 4241 10284 4253 10318
rect 4313 10284 4321 10318
rect 4385 10284 4389 10318
rect 4491 10284 4495 10318
rect 4559 10284 4567 10318
rect 4627 10284 4639 10318
rect 4695 10284 4711 10318
rect 4763 10284 4783 10318
rect 4831 10284 4855 10318
rect 4899 10284 4927 10318
rect 4967 10284 4999 10318
rect 5035 10284 5069 10318
rect 5105 10284 5137 10318
rect 5177 10284 5205 10318
rect 5249 10284 5273 10318
rect 5321 10284 5341 10318
rect 5393 10284 5409 10318
rect 5465 10284 5477 10318
rect 5537 10284 5545 10318
rect 5609 10284 5613 10318
rect 5715 10284 5719 10318
rect 5783 10284 5791 10318
rect 5851 10284 5863 10318
rect 5919 10284 5935 10318
rect 5987 10284 6007 10318
rect 6055 10284 6079 10318
rect 6123 10284 6151 10318
rect 6191 10284 6223 10318
rect 6259 10284 6293 10318
rect 6329 10284 6361 10318
rect 6401 10284 6429 10318
rect 6473 10284 6497 10318
rect 6545 10284 6565 10318
rect 6617 10284 6633 10318
rect 6689 10284 6701 10318
rect 6761 10284 6769 10318
rect 6833 10284 6837 10318
rect 6939 10284 6943 10318
rect 7007 10284 7015 10318
rect 7075 10284 7087 10318
rect 7143 10284 7159 10318
rect 7211 10284 7231 10318
rect 7279 10284 7303 10318
rect 7347 10284 7375 10318
rect 7415 10284 7447 10318
rect 7483 10284 7517 10318
rect 7553 10284 7585 10318
rect 7625 10284 7653 10318
rect 7697 10284 7721 10318
rect 7769 10284 7789 10318
rect 7841 10284 7857 10318
rect 7913 10284 7925 10318
rect 7985 10284 7993 10318
rect 8057 10284 8061 10318
rect 8163 10284 8167 10318
rect 8231 10284 8239 10318
rect 8299 10284 8311 10318
rect 8367 10284 8383 10318
rect 8435 10284 8455 10318
rect 8503 10284 8527 10318
rect 8571 10284 8599 10318
rect 8639 10284 8671 10318
rect 8707 10284 8741 10318
rect 8777 10284 8809 10318
rect 8849 10284 8877 10318
rect 8921 10284 8945 10318
rect 8993 10284 9013 10318
rect 9065 10284 9081 10318
rect 9137 10284 9149 10318
rect 9209 10284 9217 10318
rect 9281 10284 9285 10318
rect 9387 10284 9391 10318
rect 9455 10284 9463 10318
rect 9523 10284 9535 10318
rect 9591 10284 9607 10318
rect 9659 10284 9679 10318
rect 9727 10284 9751 10318
rect 9795 10284 9823 10318
rect 9863 10284 9895 10318
rect 9931 10284 9965 10318
rect 10001 10284 10033 10318
rect 10073 10284 10101 10318
rect 10145 10284 10169 10318
rect 10217 10284 10237 10318
rect 10289 10284 10305 10318
rect 10361 10284 10373 10318
rect 10433 10284 10441 10318
rect 10505 10284 10509 10318
rect 10611 10284 10615 10318
rect 10679 10284 10687 10318
rect 10747 10284 10759 10318
rect 10815 10284 10831 10318
rect 10883 10284 10903 10318
rect 10951 10284 10975 10318
rect 11019 10284 11047 10318
rect 11087 10284 11119 10318
rect 11155 10284 11189 10318
rect 11225 10284 11257 10318
rect 11297 10284 11325 10318
rect 11369 10284 11393 10318
rect 11441 10284 11461 10318
rect 11513 10284 11529 10318
rect 11585 10284 11597 10318
rect 11657 10284 11665 10318
rect 11729 10284 11733 10318
rect 11835 10284 11839 10318
rect 11903 10284 11911 10318
rect 11971 10284 11983 10318
rect 12039 10284 12055 10318
rect 12107 10284 12127 10318
rect 12175 10284 12199 10318
rect 12243 10284 12271 10318
rect 12311 10284 12343 10318
rect 12379 10284 12413 10318
rect 12449 10284 12481 10318
rect 12521 10284 12549 10318
rect 12593 10284 12617 10318
rect 12665 10284 12685 10318
rect 12737 10284 12753 10318
rect 12809 10284 12821 10318
rect 12881 10284 12889 10318
rect 12953 10284 12957 10318
rect 13059 10284 13063 10318
rect 13127 10284 13135 10318
rect 13195 10284 13207 10318
rect 13263 10284 13279 10318
rect 13331 10284 13351 10318
rect 13399 10284 13423 10318
rect 13467 10284 13495 10318
rect 13535 10284 13567 10318
rect 13603 10284 13637 10318
rect 13673 10284 13844 10318
rect 1148 10242 13844 10284
rect 13968 34691 14142 34725
rect 14176 34706 14297 34725
rect 14331 34706 14361 34740
rect 14176 34691 14361 34706
rect 13968 34672 14361 34691
rect 13968 34653 14297 34672
rect 13968 34619 14142 34653
rect 14176 34638 14297 34653
rect 14331 34638 14361 34672
rect 14176 34619 14361 34638
rect 13968 34604 14361 34619
rect 13968 34581 14297 34604
rect 13968 34547 14142 34581
rect 14176 34570 14297 34581
rect 14331 34570 14361 34604
rect 14176 34547 14361 34570
rect 13968 34536 14361 34547
rect 13968 34509 14297 34536
rect 13968 34475 14142 34509
rect 14176 34502 14297 34509
rect 14331 34502 14361 34536
rect 14176 34475 14361 34502
rect 13968 34468 14361 34475
rect 13968 34437 14297 34468
rect 13968 34403 14142 34437
rect 14176 34434 14297 34437
rect 14331 34434 14361 34468
rect 14176 34403 14361 34434
rect 13968 34400 14361 34403
rect 13968 34366 14297 34400
rect 14331 34366 14361 34400
rect 13968 34365 14361 34366
rect 13968 34331 14142 34365
rect 14176 34332 14361 34365
rect 14176 34331 14297 34332
rect 13968 34298 14297 34331
rect 14331 34298 14361 34332
rect 13968 34293 14361 34298
rect 13968 34259 14142 34293
rect 14176 34264 14361 34293
rect 14176 34259 14297 34264
rect 13968 34230 14297 34259
rect 14331 34230 14361 34264
rect 13968 34221 14361 34230
rect 13968 34187 14142 34221
rect 14176 34196 14361 34221
rect 14176 34187 14297 34196
rect 13968 34162 14297 34187
rect 14331 34162 14361 34196
rect 13968 34149 14361 34162
rect 13968 34115 14142 34149
rect 14176 34128 14361 34149
rect 14176 34115 14297 34128
rect 13968 34094 14297 34115
rect 14331 34094 14361 34128
rect 13968 34077 14361 34094
rect 13968 34043 14142 34077
rect 14176 34060 14361 34077
rect 14176 34043 14297 34060
rect 13968 34026 14297 34043
rect 14331 34026 14361 34060
rect 13968 34005 14361 34026
rect 13968 33971 14142 34005
rect 14176 33992 14361 34005
rect 14176 33971 14297 33992
rect 13968 33958 14297 33971
rect 14331 33958 14361 33992
rect 13968 33933 14361 33958
rect 13968 33899 14142 33933
rect 14176 33924 14361 33933
rect 14176 33899 14297 33924
rect 13968 33890 14297 33899
rect 14331 33890 14361 33924
rect 13968 33861 14361 33890
rect 13968 33827 14142 33861
rect 14176 33856 14361 33861
rect 14176 33827 14297 33856
rect 13968 33822 14297 33827
rect 14331 33822 14361 33856
rect 13968 33789 14361 33822
rect 13968 33755 14142 33789
rect 14176 33788 14361 33789
rect 14176 33755 14297 33788
rect 13968 33754 14297 33755
rect 14331 33754 14361 33788
rect 13968 33720 14361 33754
rect 13968 33717 14297 33720
rect 13968 33683 14142 33717
rect 14176 33686 14297 33717
rect 14331 33686 14361 33720
rect 14176 33683 14361 33686
rect 13968 33652 14361 33683
rect 13968 33645 14297 33652
rect 13968 33611 14142 33645
rect 14176 33618 14297 33645
rect 14331 33618 14361 33652
rect 14176 33611 14361 33618
rect 13968 33584 14361 33611
rect 13968 33573 14297 33584
rect 13968 33539 14142 33573
rect 14176 33550 14297 33573
rect 14331 33550 14361 33584
rect 14176 33539 14361 33550
rect 13968 33516 14361 33539
rect 13968 33501 14297 33516
rect 13968 33467 14142 33501
rect 14176 33482 14297 33501
rect 14331 33482 14361 33516
rect 14176 33467 14361 33482
rect 13968 33448 14361 33467
rect 13968 33429 14297 33448
rect 13968 33395 14142 33429
rect 14176 33414 14297 33429
rect 14331 33414 14361 33448
rect 14176 33395 14361 33414
rect 13968 33380 14361 33395
rect 13968 33357 14297 33380
rect 13968 33323 14142 33357
rect 14176 33346 14297 33357
rect 14331 33346 14361 33380
rect 14176 33323 14361 33346
rect 13968 33312 14361 33323
rect 13968 33285 14297 33312
rect 13968 33251 14142 33285
rect 14176 33278 14297 33285
rect 14331 33278 14361 33312
rect 14176 33251 14361 33278
rect 13968 33244 14361 33251
rect 13968 33213 14297 33244
rect 13968 33179 14142 33213
rect 14176 33210 14297 33213
rect 14331 33210 14361 33244
rect 14176 33179 14361 33210
rect 13968 33176 14361 33179
rect 13968 33142 14297 33176
rect 14331 33142 14361 33176
rect 13968 33141 14361 33142
rect 13968 33107 14142 33141
rect 14176 33108 14361 33141
rect 14176 33107 14297 33108
rect 13968 33074 14297 33107
rect 14331 33074 14361 33108
rect 13968 33069 14361 33074
rect 13968 33035 14142 33069
rect 14176 33040 14361 33069
rect 14176 33035 14297 33040
rect 13968 33006 14297 33035
rect 14331 33006 14361 33040
rect 13968 32997 14361 33006
rect 13968 32963 14142 32997
rect 14176 32972 14361 32997
rect 14176 32963 14297 32972
rect 13968 32938 14297 32963
rect 14331 32938 14361 32972
rect 13968 32925 14361 32938
rect 13968 32891 14142 32925
rect 14176 32904 14361 32925
rect 14176 32891 14297 32904
rect 13968 32870 14297 32891
rect 14331 32870 14361 32904
rect 13968 32853 14361 32870
rect 13968 32819 14142 32853
rect 14176 32836 14361 32853
rect 14176 32819 14297 32836
rect 13968 32802 14297 32819
rect 14331 32802 14361 32836
rect 13968 32781 14361 32802
rect 13968 32747 14142 32781
rect 14176 32768 14361 32781
rect 14176 32747 14297 32768
rect 13968 32734 14297 32747
rect 14331 32734 14361 32768
rect 13968 32709 14361 32734
rect 13968 32675 14142 32709
rect 14176 32700 14361 32709
rect 14176 32675 14297 32700
rect 13968 32666 14297 32675
rect 14331 32666 14361 32700
rect 13968 32637 14361 32666
rect 13968 32603 14142 32637
rect 14176 32632 14361 32637
rect 14176 32603 14297 32632
rect 13968 32598 14297 32603
rect 14331 32598 14361 32632
rect 13968 32565 14361 32598
rect 13968 32531 14142 32565
rect 14176 32564 14361 32565
rect 14176 32531 14297 32564
rect 13968 32530 14297 32531
rect 14331 32530 14361 32564
rect 13968 32496 14361 32530
rect 13968 32493 14297 32496
rect 13968 32459 14142 32493
rect 14176 32462 14297 32493
rect 14331 32462 14361 32496
rect 14176 32459 14361 32462
rect 13968 32428 14361 32459
rect 13968 32421 14297 32428
rect 13968 32387 14142 32421
rect 14176 32394 14297 32421
rect 14331 32394 14361 32428
rect 14176 32387 14361 32394
rect 13968 32360 14361 32387
rect 13968 32349 14297 32360
rect 13968 32315 14142 32349
rect 14176 32326 14297 32349
rect 14331 32326 14361 32360
rect 14176 32315 14361 32326
rect 13968 32292 14361 32315
rect 13968 32277 14297 32292
rect 13968 32243 14142 32277
rect 14176 32258 14297 32277
rect 14331 32258 14361 32292
rect 14176 32243 14361 32258
rect 13968 32224 14361 32243
rect 13968 32205 14297 32224
rect 13968 32171 14142 32205
rect 14176 32190 14297 32205
rect 14331 32190 14361 32224
rect 14176 32171 14361 32190
rect 13968 32156 14361 32171
rect 13968 32133 14297 32156
rect 13968 32099 14142 32133
rect 14176 32122 14297 32133
rect 14331 32122 14361 32156
rect 14176 32099 14361 32122
rect 13968 32088 14361 32099
rect 13968 32061 14297 32088
rect 13968 32027 14142 32061
rect 14176 32054 14297 32061
rect 14331 32054 14361 32088
rect 14176 32027 14361 32054
rect 13968 32020 14361 32027
rect 13968 31989 14297 32020
rect 13968 31955 14142 31989
rect 14176 31986 14297 31989
rect 14331 31986 14361 32020
rect 14176 31955 14361 31986
rect 13968 31952 14361 31955
rect 13968 31918 14297 31952
rect 14331 31918 14361 31952
rect 13968 31917 14361 31918
rect 13968 31883 14142 31917
rect 14176 31884 14361 31917
rect 14176 31883 14297 31884
rect 13968 31850 14297 31883
rect 14331 31850 14361 31884
rect 13968 31845 14361 31850
rect 13968 31811 14142 31845
rect 14176 31816 14361 31845
rect 14176 31811 14297 31816
rect 13968 31782 14297 31811
rect 14331 31782 14361 31816
rect 13968 31773 14361 31782
rect 13968 31739 14142 31773
rect 14176 31748 14361 31773
rect 14176 31739 14297 31748
rect 13968 31714 14297 31739
rect 14331 31714 14361 31748
rect 13968 31701 14361 31714
rect 13968 31667 14142 31701
rect 14176 31680 14361 31701
rect 14176 31667 14297 31680
rect 13968 31646 14297 31667
rect 14331 31646 14361 31680
rect 13968 31629 14361 31646
rect 13968 31595 14142 31629
rect 14176 31612 14361 31629
rect 14176 31595 14297 31612
rect 13968 31578 14297 31595
rect 14331 31578 14361 31612
rect 13968 31557 14361 31578
rect 13968 31523 14142 31557
rect 14176 31544 14361 31557
rect 14176 31523 14297 31544
rect 13968 31510 14297 31523
rect 14331 31510 14361 31544
rect 13968 31485 14361 31510
rect 13968 31451 14142 31485
rect 14176 31476 14361 31485
rect 14176 31451 14297 31476
rect 13968 31442 14297 31451
rect 14331 31442 14361 31476
rect 13968 31413 14361 31442
rect 13968 31379 14142 31413
rect 14176 31408 14361 31413
rect 14176 31379 14297 31408
rect 13968 31374 14297 31379
rect 14331 31374 14361 31408
rect 13968 31341 14361 31374
rect 13968 31307 14142 31341
rect 14176 31340 14361 31341
rect 14176 31307 14297 31340
rect 13968 31306 14297 31307
rect 14331 31306 14361 31340
rect 13968 31272 14361 31306
rect 13968 31269 14297 31272
rect 13968 31235 14142 31269
rect 14176 31238 14297 31269
rect 14331 31238 14361 31272
rect 14176 31235 14361 31238
rect 13968 31204 14361 31235
rect 13968 31197 14297 31204
rect 13968 31163 14142 31197
rect 14176 31170 14297 31197
rect 14331 31170 14361 31204
rect 14176 31163 14361 31170
rect 13968 31136 14361 31163
rect 13968 31125 14297 31136
rect 13968 31091 14142 31125
rect 14176 31102 14297 31125
rect 14331 31102 14361 31136
rect 14176 31091 14361 31102
rect 13968 31068 14361 31091
rect 13968 31053 14297 31068
rect 13968 31019 14142 31053
rect 14176 31034 14297 31053
rect 14331 31034 14361 31068
rect 14176 31019 14361 31034
rect 13968 31000 14361 31019
rect 13968 30981 14297 31000
rect 13968 30947 14142 30981
rect 14176 30966 14297 30981
rect 14331 30966 14361 31000
rect 14176 30947 14361 30966
rect 13968 30932 14361 30947
rect 13968 30909 14297 30932
rect 13968 30875 14142 30909
rect 14176 30898 14297 30909
rect 14331 30898 14361 30932
rect 14176 30875 14361 30898
rect 13968 30864 14361 30875
rect 13968 30837 14297 30864
rect 13968 30803 14142 30837
rect 14176 30830 14297 30837
rect 14331 30830 14361 30864
rect 14176 30803 14361 30830
rect 13968 30796 14361 30803
rect 13968 30765 14297 30796
rect 13968 30731 14142 30765
rect 14176 30762 14297 30765
rect 14331 30762 14361 30796
rect 14176 30731 14361 30762
rect 13968 30728 14361 30731
rect 13968 30694 14297 30728
rect 14331 30694 14361 30728
rect 13968 30693 14361 30694
rect 13968 30659 14142 30693
rect 14176 30660 14361 30693
rect 14176 30659 14297 30660
rect 13968 30626 14297 30659
rect 14331 30626 14361 30660
rect 13968 30621 14361 30626
rect 13968 30587 14142 30621
rect 14176 30592 14361 30621
rect 14176 30587 14297 30592
rect 13968 30558 14297 30587
rect 14331 30558 14361 30592
rect 13968 30549 14361 30558
rect 13968 30515 14142 30549
rect 14176 30524 14361 30549
rect 14176 30515 14297 30524
rect 13968 30490 14297 30515
rect 14331 30490 14361 30524
rect 13968 30477 14361 30490
rect 13968 30443 14142 30477
rect 14176 30456 14361 30477
rect 14176 30443 14297 30456
rect 13968 30422 14297 30443
rect 14331 30422 14361 30456
rect 13968 30405 14361 30422
rect 13968 30371 14142 30405
rect 14176 30388 14361 30405
rect 14176 30371 14297 30388
rect 13968 30354 14297 30371
rect 14331 30354 14361 30388
rect 13968 30333 14361 30354
rect 13968 30299 14142 30333
rect 14176 30320 14361 30333
rect 14176 30299 14297 30320
rect 13968 30286 14297 30299
rect 14331 30286 14361 30320
rect 13968 30261 14361 30286
rect 13968 30227 14142 30261
rect 14176 30252 14361 30261
rect 14176 30227 14297 30252
rect 13968 30218 14297 30227
rect 14331 30218 14361 30252
rect 13968 30189 14361 30218
rect 13968 30155 14142 30189
rect 14176 30184 14361 30189
rect 14176 30155 14297 30184
rect 13968 30150 14297 30155
rect 14331 30150 14361 30184
rect 13968 30117 14361 30150
rect 13968 30083 14142 30117
rect 14176 30116 14361 30117
rect 14176 30083 14297 30116
rect 13968 30082 14297 30083
rect 14331 30082 14361 30116
rect 13968 30048 14361 30082
rect 13968 30045 14297 30048
rect 13968 30011 14142 30045
rect 14176 30014 14297 30045
rect 14331 30014 14361 30048
rect 14176 30011 14361 30014
rect 13968 29980 14361 30011
rect 13968 29973 14297 29980
rect 13968 29939 14142 29973
rect 14176 29946 14297 29973
rect 14331 29946 14361 29980
rect 14176 29939 14361 29946
rect 13968 29912 14361 29939
rect 13968 29901 14297 29912
rect 13968 29867 14142 29901
rect 14176 29878 14297 29901
rect 14331 29878 14361 29912
rect 14176 29867 14361 29878
rect 13968 29844 14361 29867
rect 13968 29829 14297 29844
rect 13968 29795 14142 29829
rect 14176 29810 14297 29829
rect 14331 29810 14361 29844
rect 14176 29795 14361 29810
rect 13968 29776 14361 29795
rect 13968 29757 14297 29776
rect 13968 29723 14142 29757
rect 14176 29742 14297 29757
rect 14331 29742 14361 29776
rect 14176 29723 14361 29742
rect 13968 29708 14361 29723
rect 13968 29685 14297 29708
rect 13968 29651 14142 29685
rect 14176 29674 14297 29685
rect 14331 29674 14361 29708
rect 14176 29651 14361 29674
rect 13968 29640 14361 29651
rect 13968 29613 14297 29640
rect 13968 29579 14142 29613
rect 14176 29606 14297 29613
rect 14331 29606 14361 29640
rect 14176 29579 14361 29606
rect 13968 29572 14361 29579
rect 13968 29541 14297 29572
rect 13968 29507 14142 29541
rect 14176 29538 14297 29541
rect 14331 29538 14361 29572
rect 14176 29507 14361 29538
rect 13968 29504 14361 29507
rect 13968 29470 14297 29504
rect 14331 29470 14361 29504
rect 13968 29469 14361 29470
rect 13968 29435 14142 29469
rect 14176 29436 14361 29469
rect 14176 29435 14297 29436
rect 13968 29402 14297 29435
rect 14331 29402 14361 29436
rect 13968 29397 14361 29402
rect 13968 29363 14142 29397
rect 14176 29368 14361 29397
rect 14176 29363 14297 29368
rect 13968 29334 14297 29363
rect 14331 29334 14361 29368
rect 13968 29325 14361 29334
rect 13968 29291 14142 29325
rect 14176 29300 14361 29325
rect 14176 29291 14297 29300
rect 13968 29266 14297 29291
rect 14331 29266 14361 29300
rect 13968 29253 14361 29266
rect 13968 29219 14142 29253
rect 14176 29232 14361 29253
rect 14176 29219 14297 29232
rect 13968 29198 14297 29219
rect 14331 29198 14361 29232
rect 13968 29181 14361 29198
rect 13968 29147 14142 29181
rect 14176 29164 14361 29181
rect 14176 29147 14297 29164
rect 13968 29130 14297 29147
rect 14331 29130 14361 29164
rect 13968 29109 14361 29130
rect 13968 29075 14142 29109
rect 14176 29096 14361 29109
rect 14176 29075 14297 29096
rect 13968 29062 14297 29075
rect 14331 29062 14361 29096
rect 13968 29037 14361 29062
rect 13968 29003 14142 29037
rect 14176 29028 14361 29037
rect 14176 29003 14297 29028
rect 13968 28994 14297 29003
rect 14331 28994 14361 29028
rect 13968 28965 14361 28994
rect 13968 28931 14142 28965
rect 14176 28960 14361 28965
rect 14176 28931 14297 28960
rect 13968 28926 14297 28931
rect 14331 28926 14361 28960
rect 13968 28893 14361 28926
rect 13968 28859 14142 28893
rect 14176 28892 14361 28893
rect 14176 28859 14297 28892
rect 13968 28858 14297 28859
rect 14331 28858 14361 28892
rect 13968 28824 14361 28858
rect 13968 28821 14297 28824
rect 13968 28787 14142 28821
rect 14176 28790 14297 28821
rect 14331 28790 14361 28824
rect 14176 28787 14361 28790
rect 13968 28756 14361 28787
rect 13968 28749 14297 28756
rect 13968 28715 14142 28749
rect 14176 28722 14297 28749
rect 14331 28722 14361 28756
rect 14176 28715 14361 28722
rect 13968 28688 14361 28715
rect 13968 28677 14297 28688
rect 13968 28643 14142 28677
rect 14176 28654 14297 28677
rect 14331 28654 14361 28688
rect 14176 28643 14361 28654
rect 13968 28620 14361 28643
rect 13968 28605 14297 28620
rect 13968 28571 14142 28605
rect 14176 28586 14297 28605
rect 14331 28586 14361 28620
rect 14176 28571 14361 28586
rect 13968 28552 14361 28571
rect 13968 28533 14297 28552
rect 13968 28499 14142 28533
rect 14176 28518 14297 28533
rect 14331 28518 14361 28552
rect 14176 28499 14361 28518
rect 13968 28484 14361 28499
rect 13968 28461 14297 28484
rect 13968 28427 14142 28461
rect 14176 28450 14297 28461
rect 14331 28450 14361 28484
rect 14176 28427 14361 28450
rect 13968 28416 14361 28427
rect 13968 28389 14297 28416
rect 13968 28355 14142 28389
rect 14176 28382 14297 28389
rect 14331 28382 14361 28416
rect 14176 28355 14361 28382
rect 13968 28348 14361 28355
rect 13968 28317 14297 28348
rect 13968 28283 14142 28317
rect 14176 28314 14297 28317
rect 14331 28314 14361 28348
rect 14176 28283 14361 28314
rect 13968 28280 14361 28283
rect 13968 28246 14297 28280
rect 14331 28246 14361 28280
rect 13968 28245 14361 28246
rect 13968 28211 14142 28245
rect 14176 28212 14361 28245
rect 14176 28211 14297 28212
rect 13968 28178 14297 28211
rect 14331 28178 14361 28212
rect 13968 28173 14361 28178
rect 13968 28139 14142 28173
rect 14176 28144 14361 28173
rect 14176 28139 14297 28144
rect 13968 28110 14297 28139
rect 14331 28110 14361 28144
rect 13968 28101 14361 28110
rect 13968 28067 14142 28101
rect 14176 28076 14361 28101
rect 14176 28067 14297 28076
rect 13968 28042 14297 28067
rect 14331 28042 14361 28076
rect 13968 28029 14361 28042
rect 13968 27995 14142 28029
rect 14176 28008 14361 28029
rect 14176 27995 14297 28008
rect 13968 27974 14297 27995
rect 14331 27974 14361 28008
rect 13968 27957 14361 27974
rect 13968 27923 14142 27957
rect 14176 27940 14361 27957
rect 14176 27923 14297 27940
rect 13968 27906 14297 27923
rect 14331 27906 14361 27940
rect 13968 27885 14361 27906
rect 13968 27851 14142 27885
rect 14176 27872 14361 27885
rect 14176 27851 14297 27872
rect 13968 27838 14297 27851
rect 14331 27838 14361 27872
rect 13968 27813 14361 27838
rect 13968 27779 14142 27813
rect 14176 27804 14361 27813
rect 14176 27779 14297 27804
rect 13968 27770 14297 27779
rect 14331 27770 14361 27804
rect 13968 27741 14361 27770
rect 13968 27707 14142 27741
rect 14176 27736 14361 27741
rect 14176 27707 14297 27736
rect 13968 27702 14297 27707
rect 14331 27702 14361 27736
rect 13968 27669 14361 27702
rect 13968 27635 14142 27669
rect 14176 27668 14361 27669
rect 14176 27635 14297 27668
rect 13968 27634 14297 27635
rect 14331 27634 14361 27668
rect 13968 27600 14361 27634
rect 13968 27597 14297 27600
rect 13968 27563 14142 27597
rect 14176 27566 14297 27597
rect 14331 27566 14361 27600
rect 14176 27563 14361 27566
rect 13968 27532 14361 27563
rect 13968 27525 14297 27532
rect 13968 27491 14142 27525
rect 14176 27498 14297 27525
rect 14331 27498 14361 27532
rect 14176 27491 14361 27498
rect 13968 27464 14361 27491
rect 13968 27453 14297 27464
rect 13968 27419 14142 27453
rect 14176 27430 14297 27453
rect 14331 27430 14361 27464
rect 14176 27419 14361 27430
rect 13968 27396 14361 27419
rect 13968 27381 14297 27396
rect 13968 27347 14142 27381
rect 14176 27362 14297 27381
rect 14331 27362 14361 27396
rect 14176 27347 14361 27362
rect 13968 27328 14361 27347
rect 13968 27309 14297 27328
rect 13968 27275 14142 27309
rect 14176 27294 14297 27309
rect 14331 27294 14361 27328
rect 14176 27275 14361 27294
rect 13968 27260 14361 27275
rect 13968 27237 14297 27260
rect 13968 27203 14142 27237
rect 14176 27226 14297 27237
rect 14331 27226 14361 27260
rect 14176 27203 14361 27226
rect 13968 27192 14361 27203
rect 13968 27165 14297 27192
rect 13968 27131 14142 27165
rect 14176 27158 14297 27165
rect 14331 27158 14361 27192
rect 14176 27131 14361 27158
rect 13968 27124 14361 27131
rect 13968 27093 14297 27124
rect 13968 27059 14142 27093
rect 14176 27090 14297 27093
rect 14331 27090 14361 27124
rect 14176 27059 14361 27090
rect 13968 27056 14361 27059
rect 13968 27022 14297 27056
rect 14331 27022 14361 27056
rect 13968 27021 14361 27022
rect 13968 26987 14142 27021
rect 14176 26988 14361 27021
rect 14176 26987 14297 26988
rect 13968 26954 14297 26987
rect 14331 26954 14361 26988
rect 13968 26949 14361 26954
rect 13968 26915 14142 26949
rect 14176 26920 14361 26949
rect 14176 26915 14297 26920
rect 13968 26886 14297 26915
rect 14331 26886 14361 26920
rect 13968 26877 14361 26886
rect 13968 26843 14142 26877
rect 14176 26852 14361 26877
rect 14176 26843 14297 26852
rect 13968 26818 14297 26843
rect 14331 26818 14361 26852
rect 13968 26805 14361 26818
rect 13968 26771 14142 26805
rect 14176 26784 14361 26805
rect 14176 26771 14297 26784
rect 13968 26750 14297 26771
rect 14331 26750 14361 26784
rect 13968 26733 14361 26750
rect 13968 26699 14142 26733
rect 14176 26716 14361 26733
rect 14176 26699 14297 26716
rect 13968 26682 14297 26699
rect 14331 26682 14361 26716
rect 13968 26661 14361 26682
rect 13968 26627 14142 26661
rect 14176 26648 14361 26661
rect 14176 26627 14297 26648
rect 13968 26614 14297 26627
rect 14331 26614 14361 26648
rect 13968 26589 14361 26614
rect 13968 26555 14142 26589
rect 14176 26580 14361 26589
rect 14176 26555 14297 26580
rect 13968 26546 14297 26555
rect 14331 26546 14361 26580
rect 13968 26517 14361 26546
rect 13968 26483 14142 26517
rect 14176 26512 14361 26517
rect 14176 26483 14297 26512
rect 13968 26478 14297 26483
rect 14331 26478 14361 26512
rect 13968 26445 14361 26478
rect 13968 26411 14142 26445
rect 14176 26444 14361 26445
rect 14176 26411 14297 26444
rect 13968 26410 14297 26411
rect 14331 26410 14361 26444
rect 13968 26376 14361 26410
rect 13968 26373 14297 26376
rect 13968 26339 14142 26373
rect 14176 26342 14297 26373
rect 14331 26342 14361 26376
rect 14176 26339 14361 26342
rect 13968 26308 14361 26339
rect 13968 26301 14297 26308
rect 13968 26267 14142 26301
rect 14176 26274 14297 26301
rect 14331 26274 14361 26308
rect 14176 26267 14361 26274
rect 13968 26240 14361 26267
rect 13968 26229 14297 26240
rect 13968 26195 14142 26229
rect 14176 26206 14297 26229
rect 14331 26206 14361 26240
rect 14176 26195 14361 26206
rect 13968 26172 14361 26195
rect 13968 26157 14297 26172
rect 13968 26123 14142 26157
rect 14176 26138 14297 26157
rect 14331 26138 14361 26172
rect 14176 26123 14361 26138
rect 13968 26104 14361 26123
rect 13968 26085 14297 26104
rect 13968 26051 14142 26085
rect 14176 26070 14297 26085
rect 14331 26070 14361 26104
rect 14176 26051 14361 26070
rect 13968 26036 14361 26051
rect 13968 26013 14297 26036
rect 13968 25979 14142 26013
rect 14176 26002 14297 26013
rect 14331 26002 14361 26036
rect 14176 25979 14361 26002
rect 13968 25968 14361 25979
rect 13968 25941 14297 25968
rect 13968 25907 14142 25941
rect 14176 25934 14297 25941
rect 14331 25934 14361 25968
rect 14176 25907 14361 25934
rect 13968 25900 14361 25907
rect 13968 25869 14297 25900
rect 13968 25835 14142 25869
rect 14176 25866 14297 25869
rect 14331 25866 14361 25900
rect 14176 25835 14361 25866
rect 13968 25832 14361 25835
rect 13968 25798 14297 25832
rect 14331 25798 14361 25832
rect 13968 25797 14361 25798
rect 13968 25763 14142 25797
rect 14176 25764 14361 25797
rect 14176 25763 14297 25764
rect 13968 25730 14297 25763
rect 14331 25730 14361 25764
rect 13968 25725 14361 25730
rect 13968 25691 14142 25725
rect 14176 25696 14361 25725
rect 14176 25691 14297 25696
rect 13968 25662 14297 25691
rect 14331 25662 14361 25696
rect 13968 25653 14361 25662
rect 13968 25619 14142 25653
rect 14176 25628 14361 25653
rect 14176 25619 14297 25628
rect 13968 25594 14297 25619
rect 14331 25594 14361 25628
rect 13968 25581 14361 25594
rect 13968 25547 14142 25581
rect 14176 25560 14361 25581
rect 14176 25547 14297 25560
rect 13968 25526 14297 25547
rect 14331 25526 14361 25560
rect 13968 25509 14361 25526
rect 13968 25475 14142 25509
rect 14176 25492 14361 25509
rect 14176 25475 14297 25492
rect 13968 25458 14297 25475
rect 14331 25458 14361 25492
rect 13968 25437 14361 25458
rect 13968 25403 14142 25437
rect 14176 25424 14361 25437
rect 14176 25403 14297 25424
rect 13968 25390 14297 25403
rect 14331 25390 14361 25424
rect 13968 25365 14361 25390
rect 13968 25331 14142 25365
rect 14176 25356 14361 25365
rect 14176 25331 14297 25356
rect 13968 25322 14297 25331
rect 14331 25322 14361 25356
rect 13968 25293 14361 25322
rect 13968 25259 14142 25293
rect 14176 25288 14361 25293
rect 14176 25259 14297 25288
rect 13968 25254 14297 25259
rect 14331 25254 14361 25288
rect 13968 25221 14361 25254
rect 13968 25187 14142 25221
rect 14176 25220 14361 25221
rect 14176 25187 14297 25220
rect 13968 25186 14297 25187
rect 14331 25186 14361 25220
rect 13968 25152 14361 25186
rect 13968 25149 14297 25152
rect 13968 25115 14142 25149
rect 14176 25118 14297 25149
rect 14331 25118 14361 25152
rect 14176 25115 14361 25118
rect 13968 25084 14361 25115
rect 13968 25077 14297 25084
rect 13968 25043 14142 25077
rect 14176 25050 14297 25077
rect 14331 25050 14361 25084
rect 14176 25043 14361 25050
rect 13968 25016 14361 25043
rect 13968 25005 14297 25016
rect 13968 24971 14142 25005
rect 14176 24982 14297 25005
rect 14331 24982 14361 25016
rect 14176 24971 14361 24982
rect 13968 24948 14361 24971
rect 13968 24933 14297 24948
rect 13968 24899 14142 24933
rect 14176 24914 14297 24933
rect 14331 24914 14361 24948
rect 14176 24899 14361 24914
rect 13968 24880 14361 24899
rect 13968 24861 14297 24880
rect 13968 24827 14142 24861
rect 14176 24846 14297 24861
rect 14331 24846 14361 24880
rect 14176 24827 14361 24846
rect 13968 24812 14361 24827
rect 13968 24789 14297 24812
rect 13968 24755 14142 24789
rect 14176 24778 14297 24789
rect 14331 24778 14361 24812
rect 14176 24755 14361 24778
rect 13968 24744 14361 24755
rect 13968 24717 14297 24744
rect 13968 24683 14142 24717
rect 14176 24710 14297 24717
rect 14331 24710 14361 24744
rect 14176 24683 14361 24710
rect 13968 24676 14361 24683
rect 13968 24645 14297 24676
rect 13968 24611 14142 24645
rect 14176 24642 14297 24645
rect 14331 24642 14361 24676
rect 14176 24611 14361 24642
rect 13968 24608 14361 24611
rect 13968 24574 14297 24608
rect 14331 24574 14361 24608
rect 13968 24573 14361 24574
rect 13968 24539 14142 24573
rect 14176 24540 14361 24573
rect 14176 24539 14297 24540
rect 13968 24506 14297 24539
rect 14331 24506 14361 24540
rect 13968 24501 14361 24506
rect 13968 24467 14142 24501
rect 14176 24472 14361 24501
rect 14176 24467 14297 24472
rect 13968 24438 14297 24467
rect 14331 24438 14361 24472
rect 13968 24429 14361 24438
rect 13968 24395 14142 24429
rect 14176 24404 14361 24429
rect 14176 24395 14297 24404
rect 13968 24370 14297 24395
rect 14331 24370 14361 24404
rect 13968 24357 14361 24370
rect 13968 24323 14142 24357
rect 14176 24336 14361 24357
rect 14176 24323 14297 24336
rect 13968 24302 14297 24323
rect 14331 24302 14361 24336
rect 13968 24285 14361 24302
rect 13968 24251 14142 24285
rect 14176 24268 14361 24285
rect 14176 24251 14297 24268
rect 13968 24234 14297 24251
rect 14331 24234 14361 24268
rect 13968 24213 14361 24234
rect 13968 24179 14142 24213
rect 14176 24200 14361 24213
rect 14176 24179 14297 24200
rect 13968 24166 14297 24179
rect 14331 24166 14361 24200
rect 13968 24141 14361 24166
rect 13968 24107 14142 24141
rect 14176 24132 14361 24141
rect 14176 24107 14297 24132
rect 13968 24098 14297 24107
rect 14331 24098 14361 24132
rect 13968 24069 14361 24098
rect 13968 24035 14142 24069
rect 14176 24064 14361 24069
rect 14176 24035 14297 24064
rect 13968 24030 14297 24035
rect 14331 24030 14361 24064
rect 13968 23997 14361 24030
rect 13968 23963 14142 23997
rect 14176 23996 14361 23997
rect 14176 23963 14297 23996
rect 13968 23962 14297 23963
rect 14331 23962 14361 23996
rect 13968 23928 14361 23962
rect 13968 23925 14297 23928
rect 13968 23891 14142 23925
rect 14176 23894 14297 23925
rect 14331 23894 14361 23928
rect 14176 23891 14361 23894
rect 13968 23860 14361 23891
rect 13968 23853 14297 23860
rect 13968 23819 14142 23853
rect 14176 23826 14297 23853
rect 14331 23826 14361 23860
rect 14176 23819 14361 23826
rect 13968 23792 14361 23819
rect 13968 23781 14297 23792
rect 13968 23747 14142 23781
rect 14176 23758 14297 23781
rect 14331 23758 14361 23792
rect 14176 23747 14361 23758
rect 13968 23724 14361 23747
rect 13968 23709 14297 23724
rect 13968 23675 14142 23709
rect 14176 23690 14297 23709
rect 14331 23690 14361 23724
rect 14176 23675 14361 23690
rect 13968 23656 14361 23675
rect 13968 23637 14297 23656
rect 13968 23603 14142 23637
rect 14176 23622 14297 23637
rect 14331 23622 14361 23656
rect 14176 23603 14361 23622
rect 13968 23588 14361 23603
rect 13968 23565 14297 23588
rect 13968 23531 14142 23565
rect 14176 23554 14297 23565
rect 14331 23554 14361 23588
rect 14176 23531 14361 23554
rect 13968 23520 14361 23531
rect 13968 23493 14297 23520
rect 13968 23459 14142 23493
rect 14176 23486 14297 23493
rect 14331 23486 14361 23520
rect 14176 23459 14361 23486
rect 13968 23452 14361 23459
rect 13968 23421 14297 23452
rect 13968 23387 14142 23421
rect 14176 23418 14297 23421
rect 14331 23418 14361 23452
rect 14176 23387 14361 23418
rect 13968 23384 14361 23387
rect 13968 23350 14297 23384
rect 14331 23350 14361 23384
rect 13968 23349 14361 23350
rect 13968 23315 14142 23349
rect 14176 23316 14361 23349
rect 14176 23315 14297 23316
rect 13968 23282 14297 23315
rect 14331 23282 14361 23316
rect 13968 23277 14361 23282
rect 13968 23243 14142 23277
rect 14176 23248 14361 23277
rect 14176 23243 14297 23248
rect 13968 23214 14297 23243
rect 14331 23214 14361 23248
rect 13968 23205 14361 23214
rect 13968 23171 14142 23205
rect 14176 23180 14361 23205
rect 14176 23171 14297 23180
rect 13968 23146 14297 23171
rect 14331 23146 14361 23180
rect 13968 23133 14361 23146
rect 13968 23099 14142 23133
rect 14176 23112 14361 23133
rect 14176 23099 14297 23112
rect 13968 23078 14297 23099
rect 14331 23078 14361 23112
rect 13968 23061 14361 23078
rect 13968 23027 14142 23061
rect 14176 23044 14361 23061
rect 14176 23027 14297 23044
rect 13968 23010 14297 23027
rect 14331 23010 14361 23044
rect 13968 22989 14361 23010
rect 13968 22955 14142 22989
rect 14176 22976 14361 22989
rect 14176 22955 14297 22976
rect 13968 22942 14297 22955
rect 14331 22942 14361 22976
rect 13968 22917 14361 22942
rect 13968 22883 14142 22917
rect 14176 22908 14361 22917
rect 14176 22883 14297 22908
rect 13968 22874 14297 22883
rect 14331 22874 14361 22908
rect 13968 22845 14361 22874
rect 13968 22811 14142 22845
rect 14176 22840 14361 22845
rect 14176 22811 14297 22840
rect 13968 22806 14297 22811
rect 14331 22806 14361 22840
rect 13968 22773 14361 22806
rect 13968 22739 14142 22773
rect 14176 22772 14361 22773
rect 14176 22739 14297 22772
rect 13968 22738 14297 22739
rect 14331 22738 14361 22772
rect 13968 22704 14361 22738
rect 13968 22701 14297 22704
rect 13968 22667 14142 22701
rect 14176 22670 14297 22701
rect 14331 22670 14361 22704
rect 14176 22667 14361 22670
rect 13968 22636 14361 22667
rect 13968 22629 14297 22636
rect 13968 22595 14142 22629
rect 14176 22602 14297 22629
rect 14331 22602 14361 22636
rect 14176 22595 14361 22602
rect 13968 22568 14361 22595
rect 13968 22557 14297 22568
rect 13968 22523 14142 22557
rect 14176 22534 14297 22557
rect 14331 22534 14361 22568
rect 14176 22523 14361 22534
rect 13968 22500 14361 22523
rect 13968 22485 14297 22500
rect 13968 22451 14142 22485
rect 14176 22466 14297 22485
rect 14331 22466 14361 22500
rect 14176 22451 14361 22466
rect 13968 22432 14361 22451
rect 13968 22413 14297 22432
rect 13968 22379 14142 22413
rect 14176 22398 14297 22413
rect 14331 22398 14361 22432
rect 14176 22379 14361 22398
rect 13968 22364 14361 22379
rect 13968 22341 14297 22364
rect 13968 22307 14142 22341
rect 14176 22330 14297 22341
rect 14331 22330 14361 22364
rect 14176 22307 14361 22330
rect 13968 22296 14361 22307
rect 13968 22269 14297 22296
rect 13968 22235 14142 22269
rect 14176 22262 14297 22269
rect 14331 22262 14361 22296
rect 14176 22235 14361 22262
rect 13968 22228 14361 22235
rect 13968 22197 14297 22228
rect 13968 22163 14142 22197
rect 14176 22194 14297 22197
rect 14331 22194 14361 22228
rect 14176 22163 14361 22194
rect 13968 22160 14361 22163
rect 13968 22126 14297 22160
rect 14331 22126 14361 22160
rect 13968 22125 14361 22126
rect 13968 22091 14142 22125
rect 14176 22092 14361 22125
rect 14176 22091 14297 22092
rect 13968 22058 14297 22091
rect 14331 22058 14361 22092
rect 13968 22053 14361 22058
rect 13968 22019 14142 22053
rect 14176 22024 14361 22053
rect 14176 22019 14297 22024
rect 13968 21990 14297 22019
rect 14331 21990 14361 22024
rect 13968 21981 14361 21990
rect 13968 21947 14142 21981
rect 14176 21956 14361 21981
rect 14176 21947 14297 21956
rect 13968 21922 14297 21947
rect 14331 21922 14361 21956
rect 13968 21909 14361 21922
rect 13968 21875 14142 21909
rect 14176 21888 14361 21909
rect 14176 21875 14297 21888
rect 13968 21854 14297 21875
rect 14331 21854 14361 21888
rect 13968 21837 14361 21854
rect 13968 21803 14142 21837
rect 14176 21820 14361 21837
rect 14176 21803 14297 21820
rect 13968 21786 14297 21803
rect 14331 21786 14361 21820
rect 13968 21765 14361 21786
rect 13968 21731 14142 21765
rect 14176 21752 14361 21765
rect 14176 21731 14297 21752
rect 13968 21718 14297 21731
rect 14331 21718 14361 21752
rect 13968 21693 14361 21718
rect 13968 21659 14142 21693
rect 14176 21684 14361 21693
rect 14176 21659 14297 21684
rect 13968 21650 14297 21659
rect 14331 21650 14361 21684
rect 13968 21621 14361 21650
rect 13968 21587 14142 21621
rect 14176 21616 14361 21621
rect 14176 21587 14297 21616
rect 13968 21582 14297 21587
rect 14331 21582 14361 21616
rect 13968 21549 14361 21582
rect 13968 21515 14142 21549
rect 14176 21548 14361 21549
rect 14176 21515 14297 21548
rect 13968 21514 14297 21515
rect 14331 21514 14361 21548
rect 13968 21480 14361 21514
rect 13968 21477 14297 21480
rect 13968 21443 14142 21477
rect 14176 21446 14297 21477
rect 14331 21446 14361 21480
rect 14176 21443 14361 21446
rect 13968 21412 14361 21443
rect 13968 21405 14297 21412
rect 13968 21371 14142 21405
rect 14176 21378 14297 21405
rect 14331 21378 14361 21412
rect 14176 21371 14361 21378
rect 13968 21344 14361 21371
rect 13968 21333 14297 21344
rect 13968 21299 14142 21333
rect 14176 21310 14297 21333
rect 14331 21310 14361 21344
rect 14176 21299 14361 21310
rect 13968 21276 14361 21299
rect 13968 21261 14297 21276
rect 13968 21227 14142 21261
rect 14176 21242 14297 21261
rect 14331 21242 14361 21276
rect 14176 21227 14361 21242
rect 13968 21208 14361 21227
rect 13968 21189 14297 21208
rect 13968 21155 14142 21189
rect 14176 21174 14297 21189
rect 14331 21174 14361 21208
rect 14176 21155 14361 21174
rect 13968 21140 14361 21155
rect 13968 21117 14297 21140
rect 13968 21083 14142 21117
rect 14176 21106 14297 21117
rect 14331 21106 14361 21140
rect 14176 21083 14361 21106
rect 13968 21072 14361 21083
rect 13968 21045 14297 21072
rect 13968 21011 14142 21045
rect 14176 21038 14297 21045
rect 14331 21038 14361 21072
rect 14176 21011 14361 21038
rect 13968 21004 14361 21011
rect 13968 20973 14297 21004
rect 13968 20939 14142 20973
rect 14176 20970 14297 20973
rect 14331 20970 14361 21004
rect 14176 20939 14361 20970
rect 13968 20936 14361 20939
rect 13968 20902 14297 20936
rect 14331 20902 14361 20936
rect 13968 20901 14361 20902
rect 13968 20867 14142 20901
rect 14176 20868 14361 20901
rect 14176 20867 14297 20868
rect 13968 20834 14297 20867
rect 14331 20834 14361 20868
rect 13968 20829 14361 20834
rect 13968 20795 14142 20829
rect 14176 20800 14361 20829
rect 14176 20795 14297 20800
rect 13968 20766 14297 20795
rect 14331 20766 14361 20800
rect 13968 20757 14361 20766
rect 13968 20723 14142 20757
rect 14176 20732 14361 20757
rect 14176 20723 14297 20732
rect 13968 20698 14297 20723
rect 14331 20698 14361 20732
rect 13968 20685 14361 20698
rect 13968 20651 14142 20685
rect 14176 20664 14361 20685
rect 14176 20651 14297 20664
rect 13968 20630 14297 20651
rect 14331 20630 14361 20664
rect 13968 20613 14361 20630
rect 13968 20579 14142 20613
rect 14176 20596 14361 20613
rect 14176 20579 14297 20596
rect 13968 20562 14297 20579
rect 14331 20562 14361 20596
rect 13968 20541 14361 20562
rect 13968 20507 14142 20541
rect 14176 20528 14361 20541
rect 14176 20507 14297 20528
rect 13968 20494 14297 20507
rect 14331 20494 14361 20528
rect 13968 20469 14361 20494
rect 13968 20435 14142 20469
rect 14176 20460 14361 20469
rect 14176 20435 14297 20460
rect 13968 20426 14297 20435
rect 14331 20426 14361 20460
rect 13968 20397 14361 20426
rect 13968 20363 14142 20397
rect 14176 20392 14361 20397
rect 14176 20363 14297 20392
rect 13968 20358 14297 20363
rect 14331 20358 14361 20392
rect 13968 20325 14361 20358
rect 13968 20291 14142 20325
rect 14176 20324 14361 20325
rect 14176 20291 14297 20324
rect 13968 20290 14297 20291
rect 14331 20290 14361 20324
rect 13968 20256 14361 20290
rect 13968 20253 14297 20256
rect 13968 20219 14142 20253
rect 14176 20222 14297 20253
rect 14331 20222 14361 20256
rect 14176 20219 14361 20222
rect 13968 20188 14361 20219
rect 13968 20181 14297 20188
rect 13968 20147 14142 20181
rect 14176 20154 14297 20181
rect 14331 20154 14361 20188
rect 14176 20147 14361 20154
rect 13968 20120 14361 20147
rect 13968 20109 14297 20120
rect 13968 20075 14142 20109
rect 14176 20086 14297 20109
rect 14331 20086 14361 20120
rect 14176 20075 14361 20086
rect 13968 20052 14361 20075
rect 13968 20037 14297 20052
rect 13968 20003 14142 20037
rect 14176 20018 14297 20037
rect 14331 20018 14361 20052
rect 14176 20003 14361 20018
rect 13968 19984 14361 20003
rect 13968 19965 14297 19984
rect 13968 19931 14142 19965
rect 14176 19950 14297 19965
rect 14331 19950 14361 19984
rect 14176 19931 14361 19950
rect 13968 19916 14361 19931
rect 13968 19893 14297 19916
rect 13968 19859 14142 19893
rect 14176 19882 14297 19893
rect 14331 19882 14361 19916
rect 14176 19859 14361 19882
rect 13968 19848 14361 19859
rect 13968 19821 14297 19848
rect 13968 19787 14142 19821
rect 14176 19814 14297 19821
rect 14331 19814 14361 19848
rect 14176 19787 14361 19814
rect 13968 19780 14361 19787
rect 13968 19749 14297 19780
rect 13968 19715 14142 19749
rect 14176 19746 14297 19749
rect 14331 19746 14361 19780
rect 14176 19715 14361 19746
rect 13968 19712 14361 19715
rect 13968 19678 14297 19712
rect 14331 19678 14361 19712
rect 13968 19677 14361 19678
rect 13968 19643 14142 19677
rect 14176 19644 14361 19677
rect 14176 19643 14297 19644
rect 13968 19610 14297 19643
rect 14331 19610 14361 19644
rect 13968 19605 14361 19610
rect 13968 19571 14142 19605
rect 14176 19576 14361 19605
rect 14176 19571 14297 19576
rect 13968 19542 14297 19571
rect 14331 19542 14361 19576
rect 13968 19533 14361 19542
rect 13968 19499 14142 19533
rect 14176 19508 14361 19533
rect 14176 19499 14297 19508
rect 13968 19474 14297 19499
rect 14331 19474 14361 19508
rect 13968 19461 14361 19474
rect 13968 19427 14142 19461
rect 14176 19440 14361 19461
rect 14176 19427 14297 19440
rect 13968 19406 14297 19427
rect 14331 19406 14361 19440
rect 13968 19389 14361 19406
rect 13968 19355 14142 19389
rect 14176 19372 14361 19389
rect 14176 19355 14297 19372
rect 13968 19338 14297 19355
rect 14331 19338 14361 19372
rect 13968 19317 14361 19338
rect 13968 19283 14142 19317
rect 14176 19304 14361 19317
rect 14176 19283 14297 19304
rect 13968 19270 14297 19283
rect 14331 19270 14361 19304
rect 13968 19245 14361 19270
rect 13968 19211 14142 19245
rect 14176 19236 14361 19245
rect 14176 19211 14297 19236
rect 13968 19202 14297 19211
rect 14331 19202 14361 19236
rect 13968 19173 14361 19202
rect 13968 19139 14142 19173
rect 14176 19168 14361 19173
rect 14176 19139 14297 19168
rect 13968 19134 14297 19139
rect 14331 19134 14361 19168
rect 13968 19101 14361 19134
rect 13968 19067 14142 19101
rect 14176 19100 14361 19101
rect 14176 19067 14297 19100
rect 13968 19066 14297 19067
rect 14331 19066 14361 19100
rect 13968 19032 14361 19066
rect 13968 19029 14297 19032
rect 13968 18995 14142 19029
rect 14176 18998 14297 19029
rect 14331 18998 14361 19032
rect 14176 18995 14361 18998
rect 13968 18964 14361 18995
rect 13968 18957 14297 18964
rect 13968 18923 14142 18957
rect 14176 18930 14297 18957
rect 14331 18930 14361 18964
rect 14176 18923 14361 18930
rect 13968 18896 14361 18923
rect 13968 18885 14297 18896
rect 13968 18851 14142 18885
rect 14176 18862 14297 18885
rect 14331 18862 14361 18896
rect 14176 18851 14361 18862
rect 13968 18828 14361 18851
rect 13968 18813 14297 18828
rect 13968 18779 14142 18813
rect 14176 18794 14297 18813
rect 14331 18794 14361 18828
rect 14176 18779 14361 18794
rect 13968 18760 14361 18779
rect 13968 18741 14297 18760
rect 13968 18707 14142 18741
rect 14176 18726 14297 18741
rect 14331 18726 14361 18760
rect 14176 18707 14361 18726
rect 13968 18692 14361 18707
rect 13968 18669 14297 18692
rect 13968 18635 14142 18669
rect 14176 18658 14297 18669
rect 14331 18658 14361 18692
rect 14176 18635 14361 18658
rect 13968 18624 14361 18635
rect 13968 18597 14297 18624
rect 13968 18563 14142 18597
rect 14176 18590 14297 18597
rect 14331 18590 14361 18624
rect 14176 18563 14361 18590
rect 13968 18556 14361 18563
rect 13968 18525 14297 18556
rect 13968 18491 14142 18525
rect 14176 18522 14297 18525
rect 14331 18522 14361 18556
rect 14176 18491 14361 18522
rect 13968 18488 14361 18491
rect 13968 18454 14297 18488
rect 14331 18454 14361 18488
rect 13968 18453 14361 18454
rect 13968 18419 14142 18453
rect 14176 18420 14361 18453
rect 14176 18419 14297 18420
rect 13968 18386 14297 18419
rect 14331 18386 14361 18420
rect 13968 18381 14361 18386
rect 13968 18347 14142 18381
rect 14176 18352 14361 18381
rect 14176 18347 14297 18352
rect 13968 18318 14297 18347
rect 14331 18318 14361 18352
rect 13968 18309 14361 18318
rect 13968 18275 14142 18309
rect 14176 18284 14361 18309
rect 14176 18275 14297 18284
rect 13968 18250 14297 18275
rect 14331 18250 14361 18284
rect 13968 18237 14361 18250
rect 13968 18203 14142 18237
rect 14176 18216 14361 18237
rect 14176 18203 14297 18216
rect 13968 18182 14297 18203
rect 14331 18182 14361 18216
rect 13968 18165 14361 18182
rect 13968 18131 14142 18165
rect 14176 18148 14361 18165
rect 14176 18131 14297 18148
rect 13968 18114 14297 18131
rect 14331 18114 14361 18148
rect 13968 18093 14361 18114
rect 13968 18059 14142 18093
rect 14176 18080 14361 18093
rect 14176 18059 14297 18080
rect 13968 18046 14297 18059
rect 14331 18046 14361 18080
rect 13968 18021 14361 18046
rect 13968 17987 14142 18021
rect 14176 18012 14361 18021
rect 14176 17987 14297 18012
rect 13968 17978 14297 17987
rect 14331 17978 14361 18012
rect 13968 17949 14361 17978
rect 13968 17915 14142 17949
rect 14176 17944 14361 17949
rect 14176 17915 14297 17944
rect 13968 17910 14297 17915
rect 14331 17910 14361 17944
rect 13968 17877 14361 17910
rect 13968 17843 14142 17877
rect 14176 17876 14361 17877
rect 14176 17843 14297 17876
rect 13968 17842 14297 17843
rect 14331 17842 14361 17876
rect 13968 17808 14361 17842
rect 13968 17805 14297 17808
rect 13968 17771 14142 17805
rect 14176 17774 14297 17805
rect 14331 17774 14361 17808
rect 14176 17771 14361 17774
rect 13968 17740 14361 17771
rect 13968 17733 14297 17740
rect 13968 17699 14142 17733
rect 14176 17706 14297 17733
rect 14331 17706 14361 17740
rect 14176 17699 14361 17706
rect 13968 17672 14361 17699
rect 13968 17661 14297 17672
rect 13968 17627 14142 17661
rect 14176 17638 14297 17661
rect 14331 17638 14361 17672
rect 14176 17627 14361 17638
rect 13968 17604 14361 17627
rect 13968 17589 14297 17604
rect 13968 17555 14142 17589
rect 14176 17570 14297 17589
rect 14331 17570 14361 17604
rect 14176 17555 14361 17570
rect 13968 17536 14361 17555
rect 13968 17517 14297 17536
rect 13968 17483 14142 17517
rect 14176 17502 14297 17517
rect 14331 17502 14361 17536
rect 14176 17483 14361 17502
rect 13968 17468 14361 17483
rect 13968 17445 14297 17468
rect 13968 17411 14142 17445
rect 14176 17434 14297 17445
rect 14331 17434 14361 17468
rect 14176 17411 14361 17434
rect 13968 17400 14361 17411
rect 13968 17373 14297 17400
rect 13968 17339 14142 17373
rect 14176 17366 14297 17373
rect 14331 17366 14361 17400
rect 14176 17339 14361 17366
rect 13968 17332 14361 17339
rect 13968 17301 14297 17332
rect 13968 17267 14142 17301
rect 14176 17298 14297 17301
rect 14331 17298 14361 17332
rect 14176 17267 14361 17298
rect 13968 17264 14361 17267
rect 13968 17230 14297 17264
rect 14331 17230 14361 17264
rect 13968 17229 14361 17230
rect 13968 17195 14142 17229
rect 14176 17196 14361 17229
rect 14176 17195 14297 17196
rect 13968 17162 14297 17195
rect 14331 17162 14361 17196
rect 13968 17157 14361 17162
rect 13968 17123 14142 17157
rect 14176 17128 14361 17157
rect 14176 17123 14297 17128
rect 13968 17094 14297 17123
rect 14331 17094 14361 17128
rect 13968 17085 14361 17094
rect 13968 17051 14142 17085
rect 14176 17060 14361 17085
rect 14176 17051 14297 17060
rect 13968 17026 14297 17051
rect 14331 17026 14361 17060
rect 13968 17013 14361 17026
rect 13968 16979 14142 17013
rect 14176 16992 14361 17013
rect 14176 16979 14297 16992
rect 13968 16958 14297 16979
rect 14331 16958 14361 16992
rect 13968 16941 14361 16958
rect 13968 16907 14142 16941
rect 14176 16924 14361 16941
rect 14176 16907 14297 16924
rect 13968 16890 14297 16907
rect 14331 16890 14361 16924
rect 13968 16869 14361 16890
rect 13968 16835 14142 16869
rect 14176 16856 14361 16869
rect 14176 16835 14297 16856
rect 13968 16822 14297 16835
rect 14331 16822 14361 16856
rect 13968 16797 14361 16822
rect 13968 16763 14142 16797
rect 14176 16788 14361 16797
rect 14176 16763 14297 16788
rect 13968 16754 14297 16763
rect 14331 16754 14361 16788
rect 13968 16725 14361 16754
rect 13968 16691 14142 16725
rect 14176 16720 14361 16725
rect 14176 16691 14297 16720
rect 13968 16686 14297 16691
rect 14331 16686 14361 16720
rect 13968 16653 14361 16686
rect 13968 16619 14142 16653
rect 14176 16652 14361 16653
rect 14176 16619 14297 16652
rect 13968 16618 14297 16619
rect 14331 16618 14361 16652
rect 13968 16584 14361 16618
rect 13968 16581 14297 16584
rect 13968 16547 14142 16581
rect 14176 16550 14297 16581
rect 14331 16550 14361 16584
rect 14176 16547 14361 16550
rect 13968 16516 14361 16547
rect 13968 16509 14297 16516
rect 13968 16475 14142 16509
rect 14176 16482 14297 16509
rect 14331 16482 14361 16516
rect 14176 16475 14361 16482
rect 13968 16448 14361 16475
rect 13968 16437 14297 16448
rect 13968 16403 14142 16437
rect 14176 16414 14297 16437
rect 14331 16414 14361 16448
rect 14176 16403 14361 16414
rect 13968 16380 14361 16403
rect 13968 16365 14297 16380
rect 13968 16331 14142 16365
rect 14176 16346 14297 16365
rect 14331 16346 14361 16380
rect 14176 16331 14361 16346
rect 13968 16312 14361 16331
rect 13968 16293 14297 16312
rect 13968 16259 14142 16293
rect 14176 16278 14297 16293
rect 14331 16278 14361 16312
rect 14176 16259 14361 16278
rect 13968 16244 14361 16259
rect 13968 16221 14297 16244
rect 13968 16187 14142 16221
rect 14176 16210 14297 16221
rect 14331 16210 14361 16244
rect 14176 16187 14361 16210
rect 13968 16176 14361 16187
rect 13968 16149 14297 16176
rect 13968 16115 14142 16149
rect 14176 16142 14297 16149
rect 14331 16142 14361 16176
rect 14176 16115 14361 16142
rect 13968 16108 14361 16115
rect 13968 16077 14297 16108
rect 13968 16043 14142 16077
rect 14176 16074 14297 16077
rect 14331 16074 14361 16108
rect 14176 16043 14361 16074
rect 13968 16040 14361 16043
rect 13968 16006 14297 16040
rect 14331 16006 14361 16040
rect 13968 16005 14361 16006
rect 13968 15971 14142 16005
rect 14176 15972 14361 16005
rect 14176 15971 14297 15972
rect 13968 15938 14297 15971
rect 14331 15938 14361 15972
rect 13968 15933 14361 15938
rect 13968 15899 14142 15933
rect 14176 15904 14361 15933
rect 14176 15899 14297 15904
rect 13968 15870 14297 15899
rect 14331 15870 14361 15904
rect 13968 15861 14361 15870
rect 13968 15827 14142 15861
rect 14176 15836 14361 15861
rect 14176 15827 14297 15836
rect 13968 15802 14297 15827
rect 14331 15802 14361 15836
rect 13968 15789 14361 15802
rect 13968 15755 14142 15789
rect 14176 15768 14361 15789
rect 14176 15755 14297 15768
rect 13968 15734 14297 15755
rect 14331 15734 14361 15768
rect 13968 15717 14361 15734
rect 13968 15683 14142 15717
rect 14176 15700 14361 15717
rect 14176 15683 14297 15700
rect 13968 15666 14297 15683
rect 14331 15666 14361 15700
rect 13968 15645 14361 15666
rect 13968 15611 14142 15645
rect 14176 15632 14361 15645
rect 14176 15611 14297 15632
rect 13968 15598 14297 15611
rect 14331 15598 14361 15632
rect 13968 15573 14361 15598
rect 13968 15539 14142 15573
rect 14176 15564 14361 15573
rect 14176 15539 14297 15564
rect 13968 15530 14297 15539
rect 14331 15530 14361 15564
rect 13968 15501 14361 15530
rect 13968 15467 14142 15501
rect 14176 15496 14361 15501
rect 14176 15467 14297 15496
rect 13968 15462 14297 15467
rect 14331 15462 14361 15496
rect 13968 15429 14361 15462
rect 13968 15395 14142 15429
rect 14176 15428 14361 15429
rect 14176 15395 14297 15428
rect 13968 15394 14297 15395
rect 14331 15394 14361 15428
rect 13968 15360 14361 15394
rect 13968 15357 14297 15360
rect 13968 15323 14142 15357
rect 14176 15326 14297 15357
rect 14331 15326 14361 15360
rect 14176 15323 14361 15326
rect 13968 15292 14361 15323
rect 13968 15285 14297 15292
rect 13968 15251 14142 15285
rect 14176 15258 14297 15285
rect 14331 15258 14361 15292
rect 14176 15251 14361 15258
rect 13968 15224 14361 15251
rect 13968 15213 14297 15224
rect 13968 15179 14142 15213
rect 14176 15190 14297 15213
rect 14331 15190 14361 15224
rect 14176 15179 14361 15190
rect 13968 15156 14361 15179
rect 13968 15141 14297 15156
rect 13968 15107 14142 15141
rect 14176 15122 14297 15141
rect 14331 15122 14361 15156
rect 14176 15107 14361 15122
rect 13968 15088 14361 15107
rect 13968 15069 14297 15088
rect 13968 15035 14142 15069
rect 14176 15054 14297 15069
rect 14331 15054 14361 15088
rect 14176 15035 14361 15054
rect 13968 15020 14361 15035
rect 13968 14997 14297 15020
rect 13968 14963 14142 14997
rect 14176 14986 14297 14997
rect 14331 14986 14361 15020
rect 14176 14963 14361 14986
rect 13968 14952 14361 14963
rect 13968 14925 14297 14952
rect 13968 14891 14142 14925
rect 14176 14918 14297 14925
rect 14331 14918 14361 14952
rect 14176 14891 14361 14918
rect 13968 14884 14361 14891
rect 13968 14853 14297 14884
rect 13968 14819 14142 14853
rect 14176 14850 14297 14853
rect 14331 14850 14361 14884
rect 14176 14819 14361 14850
rect 13968 14816 14361 14819
rect 13968 14782 14297 14816
rect 14331 14782 14361 14816
rect 13968 14781 14361 14782
rect 13968 14747 14142 14781
rect 14176 14748 14361 14781
rect 14176 14747 14297 14748
rect 13968 14714 14297 14747
rect 14331 14714 14361 14748
rect 13968 14709 14361 14714
rect 13968 14675 14142 14709
rect 14176 14680 14361 14709
rect 14176 14675 14297 14680
rect 13968 14646 14297 14675
rect 14331 14646 14361 14680
rect 13968 14637 14361 14646
rect 13968 14603 14142 14637
rect 14176 14612 14361 14637
rect 14176 14603 14297 14612
rect 13968 14578 14297 14603
rect 14331 14578 14361 14612
rect 13968 14565 14361 14578
rect 13968 14531 14142 14565
rect 14176 14544 14361 14565
rect 14176 14531 14297 14544
rect 13968 14510 14297 14531
rect 14331 14510 14361 14544
rect 13968 14493 14361 14510
rect 13968 14459 14142 14493
rect 14176 14476 14361 14493
rect 14176 14459 14297 14476
rect 13968 14442 14297 14459
rect 14331 14442 14361 14476
rect 13968 14421 14361 14442
rect 13968 14387 14142 14421
rect 14176 14408 14361 14421
rect 14176 14387 14297 14408
rect 13968 14374 14297 14387
rect 14331 14374 14361 14408
rect 13968 14349 14361 14374
rect 13968 14315 14142 14349
rect 14176 14340 14361 14349
rect 14176 14315 14297 14340
rect 13968 14306 14297 14315
rect 14331 14306 14361 14340
rect 13968 14277 14361 14306
rect 13968 14243 14142 14277
rect 14176 14272 14361 14277
rect 14176 14243 14297 14272
rect 13968 14238 14297 14243
rect 14331 14238 14361 14272
rect 13968 14205 14361 14238
rect 13968 14171 14142 14205
rect 14176 14204 14361 14205
rect 14176 14171 14297 14204
rect 13968 14170 14297 14171
rect 14331 14170 14361 14204
rect 13968 14136 14361 14170
rect 13968 14133 14297 14136
rect 13968 14099 14142 14133
rect 14176 14102 14297 14133
rect 14331 14102 14361 14136
rect 14176 14099 14361 14102
rect 13968 14068 14361 14099
rect 13968 14061 14297 14068
rect 13968 14027 14142 14061
rect 14176 14034 14297 14061
rect 14331 14034 14361 14068
rect 14176 14027 14361 14034
rect 13968 14000 14361 14027
rect 13968 13989 14297 14000
rect 13968 13955 14142 13989
rect 14176 13966 14297 13989
rect 14331 13966 14361 14000
rect 14176 13955 14361 13966
rect 13968 13932 14361 13955
rect 13968 13917 14297 13932
rect 13968 13883 14142 13917
rect 14176 13898 14297 13917
rect 14331 13898 14361 13932
rect 14176 13883 14361 13898
rect 13968 13864 14361 13883
rect 13968 13845 14297 13864
rect 13968 13811 14142 13845
rect 14176 13830 14297 13845
rect 14331 13830 14361 13864
rect 14176 13811 14361 13830
rect 13968 13796 14361 13811
rect 13968 13773 14297 13796
rect 13968 13739 14142 13773
rect 14176 13762 14297 13773
rect 14331 13762 14361 13796
rect 14176 13739 14361 13762
rect 13968 13728 14361 13739
rect 13968 13701 14297 13728
rect 13968 13667 14142 13701
rect 14176 13694 14297 13701
rect 14331 13694 14361 13728
rect 14176 13667 14361 13694
rect 13968 13660 14361 13667
rect 13968 13629 14297 13660
rect 13968 13595 14142 13629
rect 14176 13626 14297 13629
rect 14331 13626 14361 13660
rect 14176 13595 14361 13626
rect 13968 13592 14361 13595
rect 13968 13558 14297 13592
rect 14331 13558 14361 13592
rect 13968 13557 14361 13558
rect 13968 13523 14142 13557
rect 14176 13524 14361 13557
rect 14176 13523 14297 13524
rect 13968 13490 14297 13523
rect 14331 13490 14361 13524
rect 13968 13485 14361 13490
rect 13968 13451 14142 13485
rect 14176 13456 14361 13485
rect 14176 13451 14297 13456
rect 13968 13422 14297 13451
rect 14331 13422 14361 13456
rect 13968 13413 14361 13422
rect 13968 13379 14142 13413
rect 14176 13388 14361 13413
rect 14176 13379 14297 13388
rect 13968 13354 14297 13379
rect 14331 13354 14361 13388
rect 13968 13341 14361 13354
rect 13968 13307 14142 13341
rect 14176 13320 14361 13341
rect 14176 13307 14297 13320
rect 13968 13286 14297 13307
rect 14331 13286 14361 13320
rect 13968 13269 14361 13286
rect 13968 13235 14142 13269
rect 14176 13252 14361 13269
rect 14176 13235 14297 13252
rect 13968 13218 14297 13235
rect 14331 13218 14361 13252
rect 13968 13197 14361 13218
rect 13968 13163 14142 13197
rect 14176 13184 14361 13197
rect 14176 13163 14297 13184
rect 13968 13150 14297 13163
rect 14331 13150 14361 13184
rect 13968 13125 14361 13150
rect 13968 13091 14142 13125
rect 14176 13116 14361 13125
rect 14176 13091 14297 13116
rect 13968 13082 14297 13091
rect 14331 13082 14361 13116
rect 13968 13053 14361 13082
rect 13968 13019 14142 13053
rect 14176 13048 14361 13053
rect 14176 13019 14297 13048
rect 13968 13014 14297 13019
rect 14331 13014 14361 13048
rect 13968 12981 14361 13014
rect 13968 12947 14142 12981
rect 14176 12980 14361 12981
rect 14176 12947 14297 12980
rect 13968 12946 14297 12947
rect 14331 12946 14361 12980
rect 13968 12912 14361 12946
rect 13968 12909 14297 12912
rect 13968 12875 14142 12909
rect 14176 12878 14297 12909
rect 14331 12878 14361 12912
rect 14176 12875 14361 12878
rect 13968 12844 14361 12875
rect 13968 12837 14297 12844
rect 13968 12803 14142 12837
rect 14176 12810 14297 12837
rect 14331 12810 14361 12844
rect 14176 12803 14361 12810
rect 13968 12776 14361 12803
rect 13968 12765 14297 12776
rect 13968 12731 14142 12765
rect 14176 12742 14297 12765
rect 14331 12742 14361 12776
rect 14176 12731 14361 12742
rect 13968 12708 14361 12731
rect 13968 12693 14297 12708
rect 13968 12659 14142 12693
rect 14176 12674 14297 12693
rect 14331 12674 14361 12708
rect 14176 12659 14361 12674
rect 13968 12640 14361 12659
rect 13968 12621 14297 12640
rect 13968 12587 14142 12621
rect 14176 12606 14297 12621
rect 14331 12606 14361 12640
rect 14176 12587 14361 12606
rect 13968 12572 14361 12587
rect 13968 12549 14297 12572
rect 13968 12515 14142 12549
rect 14176 12538 14297 12549
rect 14331 12538 14361 12572
rect 14176 12515 14361 12538
rect 13968 12504 14361 12515
rect 13968 12477 14297 12504
rect 13968 12443 14142 12477
rect 14176 12470 14297 12477
rect 14331 12470 14361 12504
rect 14176 12443 14361 12470
rect 13968 12436 14361 12443
rect 13968 12405 14297 12436
rect 13968 12371 14142 12405
rect 14176 12402 14297 12405
rect 14331 12402 14361 12436
rect 14176 12371 14361 12402
rect 13968 12368 14361 12371
rect 13968 12334 14297 12368
rect 14331 12334 14361 12368
rect 13968 12333 14361 12334
rect 13968 12299 14142 12333
rect 14176 12300 14361 12333
rect 14176 12299 14297 12300
rect 13968 12266 14297 12299
rect 14331 12266 14361 12300
rect 13968 12261 14361 12266
rect 13968 12227 14142 12261
rect 14176 12232 14361 12261
rect 14176 12227 14297 12232
rect 13968 12198 14297 12227
rect 14331 12198 14361 12232
rect 13968 12189 14361 12198
rect 13968 12155 14142 12189
rect 14176 12164 14361 12189
rect 14176 12155 14297 12164
rect 13968 12130 14297 12155
rect 14331 12130 14361 12164
rect 13968 12117 14361 12130
rect 13968 12083 14142 12117
rect 14176 12096 14361 12117
rect 14176 12083 14297 12096
rect 13968 12062 14297 12083
rect 14331 12062 14361 12096
rect 13968 12045 14361 12062
rect 13968 12011 14142 12045
rect 14176 12028 14361 12045
rect 14176 12011 14297 12028
rect 13968 11994 14297 12011
rect 14331 11994 14361 12028
rect 13968 11973 14361 11994
rect 13968 11939 14142 11973
rect 14176 11960 14361 11973
rect 14176 11939 14297 11960
rect 13968 11926 14297 11939
rect 14331 11926 14361 11960
rect 13968 11901 14361 11926
rect 13968 11867 14142 11901
rect 14176 11892 14361 11901
rect 14176 11867 14297 11892
rect 13968 11858 14297 11867
rect 14331 11858 14361 11892
rect 13968 11829 14361 11858
rect 13968 11795 14142 11829
rect 14176 11824 14361 11829
rect 14176 11795 14297 11824
rect 13968 11790 14297 11795
rect 14331 11790 14361 11824
rect 13968 11757 14361 11790
rect 13968 11723 14142 11757
rect 14176 11756 14361 11757
rect 14176 11723 14297 11756
rect 13968 11722 14297 11723
rect 14331 11722 14361 11756
rect 13968 11688 14361 11722
rect 13968 11685 14297 11688
rect 13968 11651 14142 11685
rect 14176 11654 14297 11685
rect 14331 11654 14361 11688
rect 14176 11651 14361 11654
rect 13968 11620 14361 11651
rect 13968 11613 14297 11620
rect 13968 11579 14142 11613
rect 14176 11586 14297 11613
rect 14331 11586 14361 11620
rect 14176 11579 14361 11586
rect 13968 11552 14361 11579
rect 13968 11541 14297 11552
rect 13968 11507 14142 11541
rect 14176 11518 14297 11541
rect 14331 11518 14361 11552
rect 14176 11507 14361 11518
rect 13968 11484 14361 11507
rect 13968 11469 14297 11484
rect 13968 11435 14142 11469
rect 14176 11450 14297 11469
rect 14331 11450 14361 11484
rect 14176 11435 14361 11450
rect 13968 11416 14361 11435
rect 13968 11397 14297 11416
rect 13968 11363 14142 11397
rect 14176 11382 14297 11397
rect 14331 11382 14361 11416
rect 14176 11363 14361 11382
rect 13968 11348 14361 11363
rect 13968 11325 14297 11348
rect 13968 11291 14142 11325
rect 14176 11314 14297 11325
rect 14331 11314 14361 11348
rect 14176 11291 14361 11314
rect 13968 11280 14361 11291
rect 13968 11253 14297 11280
rect 13968 11219 14142 11253
rect 14176 11246 14297 11253
rect 14331 11246 14361 11280
rect 14176 11219 14361 11246
rect 13968 11212 14361 11219
rect 13968 11181 14297 11212
rect 13968 11147 14142 11181
rect 14176 11178 14297 11181
rect 14331 11178 14361 11212
rect 14176 11147 14361 11178
rect 13968 11144 14361 11147
rect 13968 11110 14297 11144
rect 14331 11110 14361 11144
rect 13968 11109 14361 11110
rect 13968 11075 14142 11109
rect 14176 11076 14361 11109
rect 14176 11075 14297 11076
rect 13968 11042 14297 11075
rect 14331 11042 14361 11076
rect 13968 11037 14361 11042
rect 13968 11003 14142 11037
rect 14176 11008 14361 11037
rect 14176 11003 14297 11008
rect 13968 10974 14297 11003
rect 14331 10974 14361 11008
rect 13968 10965 14361 10974
rect 13968 10931 14142 10965
rect 14176 10940 14361 10965
rect 14176 10931 14297 10940
rect 13968 10906 14297 10931
rect 14331 10906 14361 10940
rect 13968 10893 14361 10906
rect 13968 10859 14142 10893
rect 14176 10872 14361 10893
rect 14176 10859 14297 10872
rect 13968 10838 14297 10859
rect 14331 10838 14361 10872
rect 13968 10821 14361 10838
rect 13968 10787 14142 10821
rect 14176 10804 14361 10821
rect 14176 10787 14297 10804
rect 13968 10770 14297 10787
rect 14331 10770 14361 10804
rect 13968 10749 14361 10770
rect 13968 10715 14142 10749
rect 14176 10736 14361 10749
rect 14176 10715 14297 10736
rect 13968 10702 14297 10715
rect 14331 10702 14361 10736
rect 13968 10677 14361 10702
rect 13968 10643 14142 10677
rect 14176 10668 14361 10677
rect 14176 10643 14297 10668
rect 13968 10634 14297 10643
rect 14331 10634 14361 10668
rect 13968 10605 14361 10634
rect 13968 10571 14142 10605
rect 14176 10600 14361 10605
rect 14176 10571 14297 10600
rect 13968 10566 14297 10571
rect 14331 10566 14361 10600
rect 13968 10533 14361 10566
rect 13968 10499 14142 10533
rect 14176 10532 14361 10533
rect 14176 10499 14297 10532
rect 13968 10498 14297 10499
rect 14331 10498 14361 10532
rect 13968 10464 14361 10498
rect 13968 10461 14297 10464
rect 13968 10427 14142 10461
rect 14176 10430 14297 10461
rect 14331 10430 14361 10464
rect 14176 10427 14361 10430
rect 13968 10396 14361 10427
rect 13968 10389 14297 10396
rect 13968 10355 14142 10389
rect 14176 10362 14297 10389
rect 14331 10362 14361 10396
rect 14176 10355 14361 10362
rect 13968 10328 14361 10355
rect 13968 10317 14297 10328
rect 13968 10283 14142 10317
rect 14176 10294 14297 10317
rect 14331 10294 14361 10328
rect 14176 10283 14361 10294
rect 13968 10260 14361 10283
rect 13968 10245 14297 10260
rect 603 10192 1026 10218
rect 603 10158 632 10192
rect 666 10180 1026 10192
rect 666 10158 807 10180
rect 603 10146 807 10158
rect 841 10146 1026 10180
rect 603 10124 1026 10146
rect 603 10090 632 10124
rect 666 10108 1026 10124
rect 666 10090 807 10108
rect 603 10074 807 10090
rect 841 10088 1026 10108
rect 13968 10211 14142 10245
rect 14176 10226 14297 10245
rect 14331 10226 14361 10260
rect 14176 10211 14361 10226
rect 13968 10192 14361 10211
rect 13968 10173 14297 10192
rect 13968 10139 14142 10173
rect 14176 10158 14297 10173
rect 14331 10158 14361 10192
rect 14176 10139 14361 10158
rect 13968 10124 14361 10139
rect 13968 10101 14297 10124
rect 13968 10088 14142 10101
rect 841 10074 14142 10088
rect 603 10067 14142 10074
rect 14176 10090 14297 10101
rect 14331 10090 14361 10124
rect 14176 10067 14361 10090
rect 603 10056 14361 10067
rect 603 10022 632 10056
rect 666 10022 14297 10056
rect 14331 10022 14361 10056
rect 603 9988 14361 10022
rect 603 9954 632 9988
rect 666 9954 14297 9988
rect 14331 9954 14361 9988
rect 603 9942 14361 9954
rect 603 9920 891 9942
rect 603 9886 632 9920
rect 666 9908 891 9920
rect 925 9908 963 9942
rect 997 9908 1035 9942
rect 1069 9908 1107 9942
rect 1141 9908 1179 9942
rect 1213 9908 1251 9942
rect 1285 9908 1323 9942
rect 1357 9908 1395 9942
rect 1429 9908 1467 9942
rect 1501 9908 1539 9942
rect 1573 9908 1611 9942
rect 1645 9908 1683 9942
rect 1717 9908 1755 9942
rect 1789 9908 1827 9942
rect 1861 9908 1899 9942
rect 1933 9908 1971 9942
rect 2005 9908 2043 9942
rect 2077 9908 2115 9942
rect 2149 9908 2187 9942
rect 2221 9908 2259 9942
rect 2293 9908 2331 9942
rect 2365 9908 2403 9942
rect 2437 9908 2475 9942
rect 2509 9908 2547 9942
rect 2581 9908 2619 9942
rect 2653 9908 2691 9942
rect 2725 9908 2763 9942
rect 2797 9908 2835 9942
rect 2869 9908 2907 9942
rect 2941 9908 2979 9942
rect 3013 9908 3051 9942
rect 3085 9908 3123 9942
rect 3157 9908 3195 9942
rect 3229 9908 3267 9942
rect 3301 9908 3339 9942
rect 3373 9908 3411 9942
rect 3445 9908 3483 9942
rect 3517 9908 3555 9942
rect 3589 9908 3627 9942
rect 3661 9908 3699 9942
rect 3733 9908 3771 9942
rect 3805 9908 3843 9942
rect 3877 9908 3915 9942
rect 3949 9908 3987 9942
rect 4021 9908 4059 9942
rect 4093 9908 4131 9942
rect 4165 9908 4203 9942
rect 4237 9908 4275 9942
rect 4309 9908 4347 9942
rect 4381 9908 4419 9942
rect 4453 9908 4491 9942
rect 4525 9908 4563 9942
rect 4597 9908 4635 9942
rect 4669 9908 4707 9942
rect 4741 9908 4779 9942
rect 4813 9908 4851 9942
rect 4885 9908 4923 9942
rect 4957 9908 4995 9942
rect 5029 9908 5067 9942
rect 5101 9908 5139 9942
rect 5173 9908 5211 9942
rect 5245 9908 5283 9942
rect 5317 9908 5355 9942
rect 5389 9908 5427 9942
rect 5461 9908 5499 9942
rect 5533 9908 5571 9942
rect 5605 9908 5643 9942
rect 5677 9908 5715 9942
rect 5749 9908 5787 9942
rect 5821 9908 5859 9942
rect 5893 9908 5931 9942
rect 5965 9908 6003 9942
rect 6037 9908 6075 9942
rect 6109 9908 6147 9942
rect 6181 9908 6219 9942
rect 6253 9908 6291 9942
rect 6325 9908 6363 9942
rect 6397 9908 6435 9942
rect 6469 9908 6507 9942
rect 6541 9908 6579 9942
rect 6613 9908 6651 9942
rect 6685 9908 6723 9942
rect 6757 9908 6795 9942
rect 6829 9908 6867 9942
rect 6901 9908 6939 9942
rect 6973 9908 7011 9942
rect 7045 9908 7083 9942
rect 7117 9908 7155 9942
rect 7189 9908 7227 9942
rect 7261 9908 7299 9942
rect 7333 9908 7371 9942
rect 7405 9908 7443 9942
rect 7477 9908 7515 9942
rect 7549 9908 7587 9942
rect 7621 9908 7659 9942
rect 7693 9908 7731 9942
rect 7765 9908 7803 9942
rect 7837 9908 7875 9942
rect 7909 9908 7947 9942
rect 7981 9908 8019 9942
rect 8053 9908 8091 9942
rect 8125 9908 8163 9942
rect 8197 9908 8235 9942
rect 8269 9908 8307 9942
rect 8341 9908 8379 9942
rect 8413 9908 8451 9942
rect 8485 9908 8523 9942
rect 8557 9908 8595 9942
rect 8629 9908 8667 9942
rect 8701 9908 8739 9942
rect 8773 9908 8811 9942
rect 8845 9908 8883 9942
rect 8917 9908 8955 9942
rect 8989 9908 9027 9942
rect 9061 9908 9099 9942
rect 9133 9908 9171 9942
rect 9205 9908 9243 9942
rect 9277 9908 9315 9942
rect 9349 9908 9387 9942
rect 9421 9908 9459 9942
rect 9493 9908 9531 9942
rect 9565 9908 9603 9942
rect 9637 9908 9675 9942
rect 9709 9908 9747 9942
rect 9781 9908 9819 9942
rect 9853 9908 9891 9942
rect 9925 9908 9963 9942
rect 9997 9908 10035 9942
rect 10069 9908 10107 9942
rect 10141 9908 10179 9942
rect 10213 9908 10251 9942
rect 10285 9908 10323 9942
rect 10357 9908 10395 9942
rect 10429 9908 10467 9942
rect 10501 9908 10539 9942
rect 10573 9908 10611 9942
rect 10645 9908 10683 9942
rect 10717 9908 10755 9942
rect 10789 9908 10827 9942
rect 10861 9908 10899 9942
rect 10933 9908 10971 9942
rect 11005 9908 11043 9942
rect 11077 9908 11115 9942
rect 11149 9908 11187 9942
rect 11221 9908 11259 9942
rect 11293 9908 11331 9942
rect 11365 9908 11403 9942
rect 11437 9908 11475 9942
rect 11509 9908 11547 9942
rect 11581 9908 11619 9942
rect 11653 9908 11691 9942
rect 11725 9908 11763 9942
rect 11797 9908 11835 9942
rect 11869 9908 11907 9942
rect 11941 9908 11979 9942
rect 12013 9908 12051 9942
rect 12085 9908 12123 9942
rect 12157 9908 12195 9942
rect 12229 9908 12267 9942
rect 12301 9908 12339 9942
rect 12373 9908 12411 9942
rect 12445 9908 12483 9942
rect 12517 9908 12555 9942
rect 12589 9908 12627 9942
rect 12661 9908 12699 9942
rect 12733 9908 12771 9942
rect 12805 9908 12843 9942
rect 12877 9908 12915 9942
rect 12949 9908 12987 9942
rect 13021 9908 13059 9942
rect 13093 9908 13131 9942
rect 13165 9908 13203 9942
rect 13237 9908 13275 9942
rect 13309 9908 13347 9942
rect 13381 9908 13419 9942
rect 13453 9908 13491 9942
rect 13525 9908 13563 9942
rect 13597 9908 13635 9942
rect 13669 9908 13707 9942
rect 13741 9908 13779 9942
rect 13813 9908 13851 9942
rect 13885 9908 13923 9942
rect 13957 9908 13995 9942
rect 14029 9920 14361 9942
rect 14029 9908 14297 9920
rect 666 9886 14297 9908
rect 14331 9886 14361 9920
rect 603 9775 14361 9886
rect 603 9741 740 9775
rect 774 9741 808 9775
rect 842 9741 883 9775
rect 949 9741 955 9775
rect 1017 9741 1027 9775
rect 1085 9741 1099 9775
rect 1153 9741 1171 9775
rect 1221 9741 1243 9775
rect 1289 9741 1315 9775
rect 1357 9741 1387 9775
rect 1425 9741 1459 9775
rect 1493 9741 1527 9775
rect 1565 9741 1595 9775
rect 1637 9741 1663 9775
rect 1709 9741 1731 9775
rect 1781 9741 1799 9775
rect 1853 9741 1867 9775
rect 1925 9741 1935 9775
rect 1997 9741 2003 9775
rect 2069 9741 2121 9775
rect 2155 9741 2189 9775
rect 2223 9741 2257 9775
rect 2291 9741 2325 9775
rect 2359 9741 2393 9775
rect 2427 9741 2461 9775
rect 2495 9741 2529 9775
rect 2563 9741 2597 9775
rect 2631 9741 2665 9775
rect 2699 9741 2733 9775
rect 2767 9741 2801 9775
rect 2835 9741 2869 9775
rect 2903 9741 2937 9775
rect 2971 9741 3005 9775
rect 3039 9741 3073 9775
rect 3107 9741 3141 9775
rect 3175 9741 3209 9775
rect 3243 9741 3277 9775
rect 3311 9741 3345 9775
rect 3379 9741 3413 9775
rect 3447 9741 3481 9775
rect 3515 9741 3549 9775
rect 3583 9741 3617 9775
rect 3651 9741 3685 9775
rect 3719 9741 3753 9775
rect 3787 9741 3821 9775
rect 3855 9741 3889 9775
rect 3923 9741 3957 9775
rect 3991 9741 4025 9775
rect 4059 9741 4093 9775
rect 4127 9741 4161 9775
rect 4195 9741 4229 9775
rect 4263 9741 4297 9775
rect 4331 9741 4365 9775
rect 4399 9741 4433 9775
rect 4467 9741 4501 9775
rect 4535 9741 4569 9775
rect 4603 9741 4637 9775
rect 4671 9741 4705 9775
rect 4739 9741 4773 9775
rect 4807 9741 4841 9775
rect 4875 9741 4909 9775
rect 4943 9741 4977 9775
rect 5011 9741 5045 9775
rect 5079 9741 5113 9775
rect 5147 9741 5181 9775
rect 5215 9741 5249 9775
rect 5283 9741 5317 9775
rect 5351 9741 5385 9775
rect 5419 9741 5453 9775
rect 5487 9741 5521 9775
rect 5555 9741 5589 9775
rect 5623 9741 5657 9775
rect 5691 9741 5725 9775
rect 5759 9741 5793 9775
rect 5827 9741 5861 9775
rect 5895 9741 5929 9775
rect 5963 9741 5997 9775
rect 6031 9741 6065 9775
rect 6099 9741 6133 9775
rect 6167 9741 6201 9775
rect 6235 9741 6269 9775
rect 6303 9741 6337 9775
rect 6371 9741 6405 9775
rect 6439 9741 6473 9775
rect 6507 9741 6541 9775
rect 6575 9741 6609 9775
rect 6643 9741 6677 9775
rect 6711 9741 6745 9775
rect 6779 9741 6813 9775
rect 6847 9741 6881 9775
rect 6915 9741 6949 9775
rect 6983 9741 7017 9775
rect 7051 9741 7085 9775
rect 7119 9741 7153 9775
rect 7187 9741 7221 9775
rect 7255 9741 7289 9775
rect 7323 9741 7357 9775
rect 7391 9741 7425 9775
rect 7459 9741 7493 9775
rect 7527 9741 7561 9775
rect 7595 9741 7629 9775
rect 7663 9741 7697 9775
rect 7731 9741 7765 9775
rect 7799 9741 7833 9775
rect 7867 9741 7901 9775
rect 7935 9741 7969 9775
rect 8003 9741 8037 9775
rect 8071 9741 8105 9775
rect 8139 9741 8173 9775
rect 8207 9741 8241 9775
rect 8275 9741 8309 9775
rect 8343 9741 8377 9775
rect 8411 9741 8445 9775
rect 8479 9741 8513 9775
rect 8547 9741 8581 9775
rect 8615 9741 8649 9775
rect 8683 9741 8717 9775
rect 8751 9741 8785 9775
rect 8819 9741 8853 9775
rect 8887 9741 8921 9775
rect 8955 9741 8989 9775
rect 9023 9741 9057 9775
rect 9091 9741 9125 9775
rect 9159 9741 9193 9775
rect 9227 9741 9261 9775
rect 9295 9741 9329 9775
rect 9363 9741 9397 9775
rect 9431 9741 9465 9775
rect 9499 9741 9533 9775
rect 9567 9741 9601 9775
rect 9635 9741 9669 9775
rect 9703 9741 9737 9775
rect 9771 9741 9805 9775
rect 9839 9741 9873 9775
rect 9907 9741 9941 9775
rect 9975 9741 10009 9775
rect 10043 9741 10077 9775
rect 10111 9741 10145 9775
rect 10179 9741 10213 9775
rect 10247 9741 10281 9775
rect 10315 9741 10349 9775
rect 10383 9741 10417 9775
rect 10451 9741 10485 9775
rect 10519 9741 10553 9775
rect 10587 9741 10621 9775
rect 10655 9741 10689 9775
rect 10723 9741 10757 9775
rect 10791 9741 10825 9775
rect 10859 9741 10893 9775
rect 10927 9741 10961 9775
rect 10995 9741 11029 9775
rect 11063 9741 11097 9775
rect 11131 9741 11165 9775
rect 11199 9741 11233 9775
rect 11267 9741 11301 9775
rect 11335 9741 11369 9775
rect 11403 9741 11437 9775
rect 11471 9741 11505 9775
rect 11539 9741 11573 9775
rect 11607 9741 11641 9775
rect 11675 9741 11709 9775
rect 11743 9741 11777 9775
rect 11811 9741 11845 9775
rect 11879 9741 11913 9775
rect 11947 9741 11981 9775
rect 12015 9741 12049 9775
rect 12083 9741 12117 9775
rect 12151 9741 12185 9775
rect 12219 9741 12253 9775
rect 12287 9741 12321 9775
rect 12355 9741 12389 9775
rect 12423 9741 12457 9775
rect 12491 9741 12525 9775
rect 12559 9741 12593 9775
rect 12627 9741 12661 9775
rect 12695 9741 12729 9775
rect 12763 9741 12797 9775
rect 12831 9774 14115 9775
rect 12831 9741 12883 9774
rect 603 9740 12883 9741
rect 12949 9740 12955 9774
rect 13017 9740 13027 9774
rect 13085 9740 13099 9774
rect 13153 9740 13171 9774
rect 13221 9740 13243 9774
rect 13289 9740 13315 9774
rect 13357 9740 13387 9774
rect 13425 9740 13459 9774
rect 13493 9740 13527 9774
rect 13565 9740 13595 9774
rect 13637 9740 13663 9774
rect 13709 9740 13731 9774
rect 13781 9740 13799 9774
rect 13853 9740 13867 9774
rect 13925 9740 13935 9774
rect 13997 9740 14003 9774
rect 14069 9741 14115 9774
rect 14149 9741 14183 9775
rect 14217 9741 14361 9775
rect 14069 9740 14361 9741
rect 603 9711 14361 9740
rect 882 9710 2070 9711
rect 12882 9710 14361 9711
rect 14539 36190 14724 36207
rect 14539 36173 14614 36190
rect 14539 36139 14611 36173
rect 14648 36156 14724 36190
rect 14645 36139 14724 36156
rect 14539 36118 14724 36139
rect 14539 36105 14614 36118
rect 14539 36071 14611 36105
rect 14648 36084 14724 36118
rect 14645 36071 14724 36084
rect 14539 36046 14724 36071
rect 14539 36037 14614 36046
rect 14539 36003 14611 36037
rect 14648 36012 14724 36046
rect 14645 36003 14724 36012
rect 14539 35974 14724 36003
rect 14539 35969 14614 35974
rect 14539 35935 14611 35969
rect 14648 35940 14724 35974
rect 14645 35935 14724 35940
rect 14539 35902 14724 35935
rect 14539 35901 14614 35902
rect 14539 35867 14611 35901
rect 14648 35868 14724 35902
rect 14645 35867 14724 35868
rect 14539 35833 14724 35867
rect 14539 35799 14611 35833
rect 14645 35830 14724 35833
rect 14539 35796 14614 35799
rect 14648 35796 14724 35830
rect 14539 35765 14724 35796
rect 14539 35731 14611 35765
rect 14645 35758 14724 35765
rect 14539 35724 14614 35731
rect 14648 35724 14724 35758
rect 14539 35697 14724 35724
rect 14539 35663 14611 35697
rect 14645 35686 14724 35697
rect 14539 35652 14614 35663
rect 14648 35652 14724 35686
rect 14539 35629 14724 35652
rect 14539 35595 14611 35629
rect 14645 35614 14724 35629
rect 14539 35580 14614 35595
rect 14648 35580 14724 35614
rect 14539 35561 14724 35580
rect 14539 35527 14611 35561
rect 14645 35542 14724 35561
rect 14539 35508 14614 35527
rect 14648 35508 14724 35542
rect 14539 35493 14724 35508
rect 14539 35459 14611 35493
rect 14645 35470 14724 35493
rect 14539 35436 14614 35459
rect 14648 35436 14724 35470
rect 14539 35425 14724 35436
rect 14539 35391 14611 35425
rect 14645 35398 14724 35425
rect 14539 35364 14614 35391
rect 14648 35364 14724 35398
rect 14539 35357 14724 35364
rect 14539 35323 14611 35357
rect 14645 35326 14724 35357
rect 14539 35292 14614 35323
rect 14648 35292 14724 35326
rect 14539 35289 14724 35292
rect 14539 35255 14611 35289
rect 14645 35255 14724 35289
rect 14539 35254 14724 35255
rect 14539 35221 14614 35254
rect 14539 35187 14611 35221
rect 14648 35220 14724 35254
rect 14645 35187 14724 35220
rect 14539 35182 14724 35187
rect 14539 35153 14614 35182
rect 14539 35119 14611 35153
rect 14648 35148 14724 35182
rect 14645 35119 14724 35148
rect 14539 35110 14724 35119
rect 14539 35085 14614 35110
rect 14539 35051 14611 35085
rect 14648 35076 14724 35110
rect 14645 35051 14724 35076
rect 14539 35038 14724 35051
rect 14539 35017 14614 35038
rect 14539 34983 14611 35017
rect 14648 35004 14724 35038
rect 14645 34983 14724 35004
rect 14539 34966 14724 34983
rect 14539 34949 14614 34966
rect 14539 34915 14611 34949
rect 14648 34932 14724 34966
rect 14645 34915 14724 34932
rect 14539 34894 14724 34915
rect 14539 34881 14614 34894
rect 14539 34847 14611 34881
rect 14648 34860 14724 34894
rect 14645 34847 14724 34860
rect 14539 34822 14724 34847
rect 14539 34813 14614 34822
rect 14539 34779 14611 34813
rect 14648 34788 14724 34822
rect 14645 34779 14724 34788
rect 14539 34750 14724 34779
rect 14539 34745 14614 34750
rect 14539 34711 14611 34745
rect 14648 34716 14724 34750
rect 14645 34711 14724 34716
rect 14539 34678 14724 34711
rect 14539 34677 14614 34678
rect 14539 34643 14611 34677
rect 14648 34644 14724 34678
rect 14645 34643 14724 34644
rect 14539 34609 14724 34643
rect 14539 34575 14611 34609
rect 14645 34606 14724 34609
rect 14539 34572 14614 34575
rect 14648 34572 14724 34606
rect 14539 34541 14724 34572
rect 14539 34507 14611 34541
rect 14645 34534 14724 34541
rect 14539 34500 14614 34507
rect 14648 34500 14724 34534
rect 14539 34473 14724 34500
rect 14539 34439 14611 34473
rect 14645 34462 14724 34473
rect 14539 34428 14614 34439
rect 14648 34428 14724 34462
rect 14539 34405 14724 34428
rect 14539 34371 14611 34405
rect 14645 34390 14724 34405
rect 14539 34356 14614 34371
rect 14648 34356 14724 34390
rect 14539 34337 14724 34356
rect 14539 34303 14611 34337
rect 14645 34318 14724 34337
rect 14539 34284 14614 34303
rect 14648 34284 14724 34318
rect 14539 34269 14724 34284
rect 14539 34235 14611 34269
rect 14645 34246 14724 34269
rect 14539 34212 14614 34235
rect 14648 34212 14724 34246
rect 14539 34201 14724 34212
rect 14539 34167 14611 34201
rect 14645 34174 14724 34201
rect 14539 34140 14614 34167
rect 14648 34140 14724 34174
rect 14539 34133 14724 34140
rect 14539 34099 14611 34133
rect 14645 34102 14724 34133
rect 14539 34068 14614 34099
rect 14648 34068 14724 34102
rect 14539 34065 14724 34068
rect 14539 34031 14611 34065
rect 14645 34031 14724 34065
rect 14539 34030 14724 34031
rect 14539 33997 14614 34030
rect 14539 33963 14611 33997
rect 14648 33996 14724 34030
rect 14645 33963 14724 33996
rect 14539 33958 14724 33963
rect 14539 33929 14614 33958
rect 14539 33895 14611 33929
rect 14648 33924 14724 33958
rect 14645 33895 14724 33924
rect 14539 33886 14724 33895
rect 14539 33861 14614 33886
rect 14539 33827 14611 33861
rect 14648 33852 14724 33886
rect 14645 33827 14724 33852
rect 14539 33814 14724 33827
rect 14539 33793 14614 33814
rect 14539 33759 14611 33793
rect 14648 33780 14724 33814
rect 14645 33759 14724 33780
rect 14539 33742 14724 33759
rect 14539 33725 14614 33742
rect 14539 33691 14611 33725
rect 14648 33708 14724 33742
rect 14645 33691 14724 33708
rect 14539 33670 14724 33691
rect 14539 33657 14614 33670
rect 14539 33623 14611 33657
rect 14648 33636 14724 33670
rect 14645 33623 14724 33636
rect 14539 33598 14724 33623
rect 14539 33589 14614 33598
rect 14539 33555 14611 33589
rect 14648 33564 14724 33598
rect 14645 33555 14724 33564
rect 14539 33526 14724 33555
rect 14539 33521 14614 33526
rect 14539 33487 14611 33521
rect 14648 33492 14724 33526
rect 14645 33487 14724 33492
rect 14539 33454 14724 33487
rect 14539 33453 14614 33454
rect 14539 33419 14611 33453
rect 14648 33420 14724 33454
rect 14645 33419 14724 33420
rect 14539 33385 14724 33419
rect 14539 33351 14611 33385
rect 14645 33382 14724 33385
rect 14539 33348 14614 33351
rect 14648 33348 14724 33382
rect 14539 33317 14724 33348
rect 14539 33283 14611 33317
rect 14645 33310 14724 33317
rect 14539 33276 14614 33283
rect 14648 33276 14724 33310
rect 14539 33249 14724 33276
rect 14539 33215 14611 33249
rect 14645 33238 14724 33249
rect 14539 33204 14614 33215
rect 14648 33204 14724 33238
rect 14539 33181 14724 33204
rect 14539 33147 14611 33181
rect 14645 33166 14724 33181
rect 14539 33132 14614 33147
rect 14648 33132 14724 33166
rect 14539 33113 14724 33132
rect 14539 33079 14611 33113
rect 14645 33094 14724 33113
rect 14539 33060 14614 33079
rect 14648 33060 14724 33094
rect 14539 33045 14724 33060
rect 14539 33011 14611 33045
rect 14645 33022 14724 33045
rect 14539 32988 14614 33011
rect 14648 32988 14724 33022
rect 14539 32977 14724 32988
rect 14539 32943 14611 32977
rect 14645 32950 14724 32977
rect 14539 32916 14614 32943
rect 14648 32916 14724 32950
rect 14539 32909 14724 32916
rect 14539 32875 14611 32909
rect 14645 32878 14724 32909
rect 14539 32844 14614 32875
rect 14648 32844 14724 32878
rect 14539 32841 14724 32844
rect 14539 32807 14611 32841
rect 14645 32807 14724 32841
rect 14539 32806 14724 32807
rect 14539 32773 14614 32806
rect 14539 32739 14611 32773
rect 14648 32772 14724 32806
rect 14645 32739 14724 32772
rect 14539 32734 14724 32739
rect 14539 32705 14614 32734
rect 14539 32671 14611 32705
rect 14648 32700 14724 32734
rect 14645 32671 14724 32700
rect 14539 32662 14724 32671
rect 14539 32637 14614 32662
rect 14539 32603 14611 32637
rect 14648 32628 14724 32662
rect 14645 32603 14724 32628
rect 14539 32590 14724 32603
rect 14539 32569 14614 32590
rect 14539 32535 14611 32569
rect 14648 32556 14724 32590
rect 14645 32535 14724 32556
rect 14539 32518 14724 32535
rect 14539 32501 14614 32518
rect 14539 32467 14611 32501
rect 14648 32484 14724 32518
rect 14645 32467 14724 32484
rect 14539 32446 14724 32467
rect 14539 32433 14614 32446
rect 14539 32399 14611 32433
rect 14648 32412 14724 32446
rect 14645 32399 14724 32412
rect 14539 32374 14724 32399
rect 14539 32365 14614 32374
rect 14539 32331 14611 32365
rect 14648 32340 14724 32374
rect 14645 32331 14724 32340
rect 14539 32302 14724 32331
rect 14539 32297 14614 32302
rect 14539 32263 14611 32297
rect 14648 32268 14724 32302
rect 14645 32263 14724 32268
rect 14539 32230 14724 32263
rect 14539 32229 14614 32230
rect 14539 32195 14611 32229
rect 14648 32196 14724 32230
rect 14645 32195 14724 32196
rect 14539 32161 14724 32195
rect 14539 32127 14611 32161
rect 14645 32158 14724 32161
rect 14539 32124 14614 32127
rect 14648 32124 14724 32158
rect 14539 32093 14724 32124
rect 14539 32059 14611 32093
rect 14645 32086 14724 32093
rect 14539 32052 14614 32059
rect 14648 32052 14724 32086
rect 14539 32025 14724 32052
rect 14539 31991 14611 32025
rect 14645 32014 14724 32025
rect 14539 31980 14614 31991
rect 14648 31980 14724 32014
rect 14539 31957 14724 31980
rect 14539 31923 14611 31957
rect 14645 31942 14724 31957
rect 14539 31908 14614 31923
rect 14648 31908 14724 31942
rect 14539 31889 14724 31908
rect 14539 31855 14611 31889
rect 14645 31870 14724 31889
rect 14539 31836 14614 31855
rect 14648 31836 14724 31870
rect 14539 31821 14724 31836
rect 14539 31787 14611 31821
rect 14645 31798 14724 31821
rect 14539 31764 14614 31787
rect 14648 31764 14724 31798
rect 14539 31753 14724 31764
rect 14539 31719 14611 31753
rect 14645 31726 14724 31753
rect 14539 31692 14614 31719
rect 14648 31692 14724 31726
rect 14539 31685 14724 31692
rect 14539 31651 14611 31685
rect 14645 31654 14724 31685
rect 14539 31620 14614 31651
rect 14648 31620 14724 31654
rect 14539 31617 14724 31620
rect 14539 31583 14611 31617
rect 14645 31583 14724 31617
rect 14539 31582 14724 31583
rect 14539 31549 14614 31582
rect 14539 31515 14611 31549
rect 14648 31548 14724 31582
rect 14645 31515 14724 31548
rect 14539 31510 14724 31515
rect 14539 31481 14614 31510
rect 14539 31447 14611 31481
rect 14648 31476 14724 31510
rect 14645 31447 14724 31476
rect 14539 31438 14724 31447
rect 14539 31413 14614 31438
rect 14539 31379 14611 31413
rect 14648 31404 14724 31438
rect 14645 31379 14724 31404
rect 14539 31366 14724 31379
rect 14539 31345 14614 31366
rect 14539 31311 14611 31345
rect 14648 31332 14724 31366
rect 14645 31311 14724 31332
rect 14539 31294 14724 31311
rect 14539 31277 14614 31294
rect 14539 31243 14611 31277
rect 14648 31260 14724 31294
rect 14645 31243 14724 31260
rect 14539 31222 14724 31243
rect 14539 31209 14614 31222
rect 14539 31175 14611 31209
rect 14648 31188 14724 31222
rect 14645 31175 14724 31188
rect 14539 31150 14724 31175
rect 14539 31141 14614 31150
rect 14539 31107 14611 31141
rect 14648 31116 14724 31150
rect 14645 31107 14724 31116
rect 14539 31078 14724 31107
rect 14539 31073 14614 31078
rect 14539 31039 14611 31073
rect 14648 31044 14724 31078
rect 14645 31039 14724 31044
rect 14539 31006 14724 31039
rect 14539 31005 14614 31006
rect 14539 30971 14611 31005
rect 14648 30972 14724 31006
rect 14645 30971 14724 30972
rect 14539 30937 14724 30971
rect 14539 30903 14611 30937
rect 14645 30934 14724 30937
rect 14539 30900 14614 30903
rect 14648 30900 14724 30934
rect 14539 30869 14724 30900
rect 14539 30835 14611 30869
rect 14645 30862 14724 30869
rect 14539 30828 14614 30835
rect 14648 30828 14724 30862
rect 14539 30801 14724 30828
rect 14539 30767 14611 30801
rect 14645 30790 14724 30801
rect 14539 30756 14614 30767
rect 14648 30756 14724 30790
rect 14539 30733 14724 30756
rect 14539 30699 14611 30733
rect 14645 30718 14724 30733
rect 14539 30684 14614 30699
rect 14648 30684 14724 30718
rect 14539 30665 14724 30684
rect 14539 30631 14611 30665
rect 14645 30646 14724 30665
rect 14539 30612 14614 30631
rect 14648 30612 14724 30646
rect 14539 30597 14724 30612
rect 14539 30563 14611 30597
rect 14645 30574 14724 30597
rect 14539 30540 14614 30563
rect 14648 30540 14724 30574
rect 14539 30529 14724 30540
rect 14539 30495 14611 30529
rect 14645 30502 14724 30529
rect 14539 30468 14614 30495
rect 14648 30468 14724 30502
rect 14539 30461 14724 30468
rect 14539 30427 14611 30461
rect 14645 30430 14724 30461
rect 14539 30396 14614 30427
rect 14648 30396 14724 30430
rect 14539 30393 14724 30396
rect 14539 30359 14611 30393
rect 14645 30359 14724 30393
rect 14539 30358 14724 30359
rect 14539 30325 14614 30358
rect 14539 30291 14611 30325
rect 14648 30324 14724 30358
rect 14645 30291 14724 30324
rect 14539 30286 14724 30291
rect 14539 30257 14614 30286
rect 14539 30223 14611 30257
rect 14648 30252 14724 30286
rect 14645 30223 14724 30252
rect 14539 30214 14724 30223
rect 14539 30189 14614 30214
rect 14539 30155 14611 30189
rect 14648 30180 14724 30214
rect 14645 30155 14724 30180
rect 14539 30142 14724 30155
rect 14539 30121 14614 30142
rect 14539 30087 14611 30121
rect 14648 30108 14724 30142
rect 14645 30087 14724 30108
rect 14539 30070 14724 30087
rect 14539 30053 14614 30070
rect 14539 30019 14611 30053
rect 14648 30036 14724 30070
rect 14645 30019 14724 30036
rect 14539 29998 14724 30019
rect 14539 29985 14614 29998
rect 14539 29951 14611 29985
rect 14648 29964 14724 29998
rect 14645 29951 14724 29964
rect 14539 29926 14724 29951
rect 14539 29917 14614 29926
rect 14539 29883 14611 29917
rect 14648 29892 14724 29926
rect 14645 29883 14724 29892
rect 14539 29854 14724 29883
rect 14539 29849 14614 29854
rect 14539 29815 14611 29849
rect 14648 29820 14724 29854
rect 14645 29815 14724 29820
rect 14539 29782 14724 29815
rect 14539 29781 14614 29782
rect 14539 29747 14611 29781
rect 14648 29748 14724 29782
rect 14645 29747 14724 29748
rect 14539 29713 14724 29747
rect 14539 29679 14611 29713
rect 14645 29710 14724 29713
rect 14539 29676 14614 29679
rect 14648 29676 14724 29710
rect 14539 29645 14724 29676
rect 14539 29611 14611 29645
rect 14645 29638 14724 29645
rect 14539 29604 14614 29611
rect 14648 29604 14724 29638
rect 14539 29577 14724 29604
rect 14539 29543 14611 29577
rect 14645 29566 14724 29577
rect 14539 29532 14614 29543
rect 14648 29532 14724 29566
rect 14539 29509 14724 29532
rect 14539 29475 14611 29509
rect 14645 29494 14724 29509
rect 14539 29460 14614 29475
rect 14648 29460 14724 29494
rect 14539 29441 14724 29460
rect 14539 29407 14611 29441
rect 14645 29422 14724 29441
rect 14539 29388 14614 29407
rect 14648 29388 14724 29422
rect 14539 29373 14724 29388
rect 14539 29339 14611 29373
rect 14645 29350 14724 29373
rect 14539 29316 14614 29339
rect 14648 29316 14724 29350
rect 14539 29305 14724 29316
rect 14539 29271 14611 29305
rect 14645 29278 14724 29305
rect 14539 29244 14614 29271
rect 14648 29244 14724 29278
rect 14539 29237 14724 29244
rect 14539 29203 14611 29237
rect 14645 29206 14724 29237
rect 14539 29172 14614 29203
rect 14648 29172 14724 29206
rect 14539 29169 14724 29172
rect 14539 29135 14611 29169
rect 14645 29135 14724 29169
rect 14539 29134 14724 29135
rect 14539 29101 14614 29134
rect 14539 29067 14611 29101
rect 14648 29100 14724 29134
rect 14645 29067 14724 29100
rect 14539 29062 14724 29067
rect 14539 29033 14614 29062
rect 14539 28999 14611 29033
rect 14648 29028 14724 29062
rect 14645 28999 14724 29028
rect 14539 28990 14724 28999
rect 14539 28965 14614 28990
rect 14539 28931 14611 28965
rect 14648 28956 14724 28990
rect 14645 28931 14724 28956
rect 14539 28918 14724 28931
rect 14539 28897 14614 28918
rect 14539 28863 14611 28897
rect 14648 28884 14724 28918
rect 14645 28863 14724 28884
rect 14539 28846 14724 28863
rect 14539 28829 14614 28846
rect 14539 28795 14611 28829
rect 14648 28812 14724 28846
rect 14645 28795 14724 28812
rect 14539 28774 14724 28795
rect 14539 28761 14614 28774
rect 14539 28727 14611 28761
rect 14648 28740 14724 28774
rect 14645 28727 14724 28740
rect 14539 28702 14724 28727
rect 14539 28693 14614 28702
rect 14539 28659 14611 28693
rect 14648 28668 14724 28702
rect 14645 28659 14724 28668
rect 14539 28630 14724 28659
rect 14539 28625 14614 28630
rect 14539 28591 14611 28625
rect 14648 28596 14724 28630
rect 14645 28591 14724 28596
rect 14539 28558 14724 28591
rect 14539 28557 14614 28558
rect 14539 28523 14611 28557
rect 14648 28524 14724 28558
rect 14645 28523 14724 28524
rect 14539 28489 14724 28523
rect 14539 28455 14611 28489
rect 14645 28486 14724 28489
rect 14539 28452 14614 28455
rect 14648 28452 14724 28486
rect 14539 28421 14724 28452
rect 14539 28387 14611 28421
rect 14645 28414 14724 28421
rect 14539 28380 14614 28387
rect 14648 28380 14724 28414
rect 14539 28353 14724 28380
rect 14539 28319 14611 28353
rect 14645 28342 14724 28353
rect 14539 28308 14614 28319
rect 14648 28308 14724 28342
rect 14539 28285 14724 28308
rect 14539 28251 14611 28285
rect 14645 28270 14724 28285
rect 14539 28236 14614 28251
rect 14648 28236 14724 28270
rect 14539 28217 14724 28236
rect 14539 28183 14611 28217
rect 14645 28198 14724 28217
rect 14539 28164 14614 28183
rect 14648 28164 14724 28198
rect 14539 28149 14724 28164
rect 14539 28115 14611 28149
rect 14645 28126 14724 28149
rect 14539 28092 14614 28115
rect 14648 28092 14724 28126
rect 14539 28081 14724 28092
rect 14539 28047 14611 28081
rect 14645 28054 14724 28081
rect 14539 28020 14614 28047
rect 14648 28020 14724 28054
rect 14539 28013 14724 28020
rect 14539 27979 14611 28013
rect 14645 27982 14724 28013
rect 14539 27948 14614 27979
rect 14648 27948 14724 27982
rect 14539 27945 14724 27948
rect 14539 27911 14611 27945
rect 14645 27911 14724 27945
rect 14539 27910 14724 27911
rect 14539 27877 14614 27910
rect 14539 27843 14611 27877
rect 14648 27876 14724 27910
rect 14645 27843 14724 27876
rect 14539 27838 14724 27843
rect 14539 27809 14614 27838
rect 14539 27775 14611 27809
rect 14648 27804 14724 27838
rect 14645 27775 14724 27804
rect 14539 27766 14724 27775
rect 14539 27741 14614 27766
rect 14539 27707 14611 27741
rect 14648 27732 14724 27766
rect 14645 27707 14724 27732
rect 14539 27694 14724 27707
rect 14539 27673 14614 27694
rect 14539 27639 14611 27673
rect 14648 27660 14724 27694
rect 14645 27639 14724 27660
rect 14539 27622 14724 27639
rect 14539 27605 14614 27622
rect 14539 27571 14611 27605
rect 14648 27588 14724 27622
rect 14645 27571 14724 27588
rect 14539 27550 14724 27571
rect 14539 27537 14614 27550
rect 14539 27503 14611 27537
rect 14648 27516 14724 27550
rect 14645 27503 14724 27516
rect 14539 27478 14724 27503
rect 14539 27469 14614 27478
rect 14539 27435 14611 27469
rect 14648 27444 14724 27478
rect 14645 27435 14724 27444
rect 14539 27406 14724 27435
rect 14539 27401 14614 27406
rect 14539 27367 14611 27401
rect 14648 27372 14724 27406
rect 14645 27367 14724 27372
rect 14539 27334 14724 27367
rect 14539 27333 14614 27334
rect 14539 27299 14611 27333
rect 14648 27300 14724 27334
rect 14645 27299 14724 27300
rect 14539 27265 14724 27299
rect 14539 27231 14611 27265
rect 14645 27262 14724 27265
rect 14539 27228 14614 27231
rect 14648 27228 14724 27262
rect 14539 27197 14724 27228
rect 14539 27163 14611 27197
rect 14645 27190 14724 27197
rect 14539 27156 14614 27163
rect 14648 27156 14724 27190
rect 14539 27129 14724 27156
rect 14539 27095 14611 27129
rect 14645 27118 14724 27129
rect 14539 27084 14614 27095
rect 14648 27084 14724 27118
rect 14539 27061 14724 27084
rect 14539 27027 14611 27061
rect 14645 27046 14724 27061
rect 14539 27012 14614 27027
rect 14648 27012 14724 27046
rect 14539 26993 14724 27012
rect 14539 26959 14611 26993
rect 14645 26974 14724 26993
rect 14539 26940 14614 26959
rect 14648 26940 14724 26974
rect 14539 26925 14724 26940
rect 14539 26891 14611 26925
rect 14645 26902 14724 26925
rect 14539 26868 14614 26891
rect 14648 26868 14724 26902
rect 14539 26857 14724 26868
rect 14539 26823 14611 26857
rect 14645 26830 14724 26857
rect 14539 26796 14614 26823
rect 14648 26796 14724 26830
rect 14539 26789 14724 26796
rect 14539 26755 14611 26789
rect 14645 26758 14724 26789
rect 14539 26724 14614 26755
rect 14648 26724 14724 26758
rect 14539 26721 14724 26724
rect 14539 26687 14611 26721
rect 14645 26687 14724 26721
rect 14539 26686 14724 26687
rect 14539 26653 14614 26686
rect 14539 26619 14611 26653
rect 14648 26652 14724 26686
rect 14645 26619 14724 26652
rect 14539 26614 14724 26619
rect 14539 26585 14614 26614
rect 14539 26551 14611 26585
rect 14648 26580 14724 26614
rect 14645 26551 14724 26580
rect 14539 26542 14724 26551
rect 14539 26517 14614 26542
rect 14539 26483 14611 26517
rect 14648 26508 14724 26542
rect 14645 26483 14724 26508
rect 14539 26470 14724 26483
rect 14539 26449 14614 26470
rect 14539 26415 14611 26449
rect 14648 26436 14724 26470
rect 14645 26415 14724 26436
rect 14539 26398 14724 26415
rect 14539 26381 14614 26398
rect 14539 26347 14611 26381
rect 14648 26364 14724 26398
rect 14645 26347 14724 26364
rect 14539 26326 14724 26347
rect 14539 26313 14614 26326
rect 14539 26279 14611 26313
rect 14648 26292 14724 26326
rect 14645 26279 14724 26292
rect 14539 26254 14724 26279
rect 14539 26245 14614 26254
rect 14539 26211 14611 26245
rect 14648 26220 14724 26254
rect 14645 26211 14724 26220
rect 14539 26182 14724 26211
rect 14539 26177 14614 26182
rect 14539 26143 14611 26177
rect 14648 26148 14724 26182
rect 14645 26143 14724 26148
rect 14539 26110 14724 26143
rect 14539 26109 14614 26110
rect 14539 26075 14611 26109
rect 14648 26076 14724 26110
rect 14645 26075 14724 26076
rect 14539 26041 14724 26075
rect 14539 26007 14611 26041
rect 14645 26038 14724 26041
rect 14539 26004 14614 26007
rect 14648 26004 14724 26038
rect 14539 25973 14724 26004
rect 14539 25939 14611 25973
rect 14645 25966 14724 25973
rect 14539 25932 14614 25939
rect 14648 25932 14724 25966
rect 14539 25905 14724 25932
rect 14539 25871 14611 25905
rect 14645 25894 14724 25905
rect 14539 25860 14614 25871
rect 14648 25860 14724 25894
rect 14539 25837 14724 25860
rect 14539 25803 14611 25837
rect 14645 25822 14724 25837
rect 14539 25788 14614 25803
rect 14648 25788 14724 25822
rect 14539 25769 14724 25788
rect 14539 25735 14611 25769
rect 14645 25750 14724 25769
rect 14539 25716 14614 25735
rect 14648 25716 14724 25750
rect 14539 25701 14724 25716
rect 14539 25667 14611 25701
rect 14645 25678 14724 25701
rect 14539 25644 14614 25667
rect 14648 25644 14724 25678
rect 14539 25633 14724 25644
rect 14539 25599 14611 25633
rect 14645 25606 14724 25633
rect 14539 25572 14614 25599
rect 14648 25572 14724 25606
rect 14539 25565 14724 25572
rect 14539 25531 14611 25565
rect 14645 25534 14724 25565
rect 14539 25500 14614 25531
rect 14648 25500 14724 25534
rect 14539 25497 14724 25500
rect 14539 25463 14611 25497
rect 14645 25463 14724 25497
rect 14539 25462 14724 25463
rect 14539 25429 14614 25462
rect 14539 25395 14611 25429
rect 14648 25428 14724 25462
rect 14645 25395 14724 25428
rect 14539 25390 14724 25395
rect 14539 25361 14614 25390
rect 14539 25327 14611 25361
rect 14648 25356 14724 25390
rect 14645 25327 14724 25356
rect 14539 25318 14724 25327
rect 14539 25293 14614 25318
rect 14539 25259 14611 25293
rect 14648 25284 14724 25318
rect 14645 25259 14724 25284
rect 14539 25246 14724 25259
rect 14539 25225 14614 25246
rect 14539 25191 14611 25225
rect 14648 25212 14724 25246
rect 14645 25191 14724 25212
rect 14539 25174 14724 25191
rect 14539 25157 14614 25174
rect 14539 25123 14611 25157
rect 14648 25140 14724 25174
rect 14645 25123 14724 25140
rect 14539 25102 14724 25123
rect 14539 25089 14614 25102
rect 14539 25055 14611 25089
rect 14648 25068 14724 25102
rect 14645 25055 14724 25068
rect 14539 25030 14724 25055
rect 14539 25021 14614 25030
rect 14539 24987 14611 25021
rect 14648 24996 14724 25030
rect 14645 24987 14724 24996
rect 14539 24958 14724 24987
rect 14539 24953 14614 24958
rect 14539 24919 14611 24953
rect 14648 24924 14724 24958
rect 14645 24919 14724 24924
rect 14539 24886 14724 24919
rect 14539 24885 14614 24886
rect 14539 24851 14611 24885
rect 14648 24852 14724 24886
rect 14645 24851 14724 24852
rect 14539 24817 14724 24851
rect 14539 24783 14611 24817
rect 14645 24814 14724 24817
rect 14539 24780 14614 24783
rect 14648 24780 14724 24814
rect 14539 24749 14724 24780
rect 14539 24715 14611 24749
rect 14645 24742 14724 24749
rect 14539 24708 14614 24715
rect 14648 24708 14724 24742
rect 14539 24681 14724 24708
rect 14539 24647 14611 24681
rect 14645 24670 14724 24681
rect 14539 24636 14614 24647
rect 14648 24636 14724 24670
rect 14539 24613 14724 24636
rect 14539 24579 14611 24613
rect 14645 24598 14724 24613
rect 14539 24564 14614 24579
rect 14648 24564 14724 24598
rect 14539 24545 14724 24564
rect 14539 24511 14611 24545
rect 14645 24526 14724 24545
rect 14539 24492 14614 24511
rect 14648 24492 14724 24526
rect 14539 24477 14724 24492
rect 14539 24443 14611 24477
rect 14645 24454 14724 24477
rect 14539 24420 14614 24443
rect 14648 24420 14724 24454
rect 14539 24409 14724 24420
rect 14539 24375 14611 24409
rect 14645 24382 14724 24409
rect 14539 24348 14614 24375
rect 14648 24348 14724 24382
rect 14539 24341 14724 24348
rect 14539 24307 14611 24341
rect 14645 24310 14724 24341
rect 14539 24276 14614 24307
rect 14648 24276 14724 24310
rect 14539 24273 14724 24276
rect 14539 24239 14611 24273
rect 14645 24239 14724 24273
rect 14539 24238 14724 24239
rect 14539 24205 14614 24238
rect 14539 24171 14611 24205
rect 14648 24204 14724 24238
rect 14645 24171 14724 24204
rect 14539 24166 14724 24171
rect 14539 24137 14614 24166
rect 14539 24103 14611 24137
rect 14648 24132 14724 24166
rect 14645 24103 14724 24132
rect 14539 24094 14724 24103
rect 14539 24069 14614 24094
rect 14539 24035 14611 24069
rect 14648 24060 14724 24094
rect 14645 24035 14724 24060
rect 14539 24022 14724 24035
rect 14539 24001 14614 24022
rect 14539 23967 14611 24001
rect 14648 23988 14724 24022
rect 14645 23967 14724 23988
rect 14539 23950 14724 23967
rect 14539 23933 14614 23950
rect 14539 23899 14611 23933
rect 14648 23916 14724 23950
rect 14645 23899 14724 23916
rect 14539 23878 14724 23899
rect 14539 23865 14614 23878
rect 14539 23831 14611 23865
rect 14648 23844 14724 23878
rect 14645 23831 14724 23844
rect 14539 23806 14724 23831
rect 14539 23797 14614 23806
rect 14539 23763 14611 23797
rect 14648 23772 14724 23806
rect 14645 23763 14724 23772
rect 14539 23734 14724 23763
rect 14539 23729 14614 23734
rect 14539 23695 14611 23729
rect 14648 23700 14724 23734
rect 14645 23695 14724 23700
rect 14539 23662 14724 23695
rect 14539 23661 14614 23662
rect 14539 23627 14611 23661
rect 14648 23628 14724 23662
rect 14645 23627 14724 23628
rect 14539 23593 14724 23627
rect 14539 23559 14611 23593
rect 14645 23590 14724 23593
rect 14539 23556 14614 23559
rect 14648 23556 14724 23590
rect 14539 23525 14724 23556
rect 14539 23491 14611 23525
rect 14645 23518 14724 23525
rect 14539 23484 14614 23491
rect 14648 23484 14724 23518
rect 14539 23457 14724 23484
rect 14539 23423 14611 23457
rect 14645 23446 14724 23457
rect 14539 23412 14614 23423
rect 14648 23412 14724 23446
rect 14539 23389 14724 23412
rect 14539 23355 14611 23389
rect 14645 23374 14724 23389
rect 14539 23340 14614 23355
rect 14648 23340 14724 23374
rect 14539 23321 14724 23340
rect 14539 23287 14611 23321
rect 14645 23302 14724 23321
rect 14539 23268 14614 23287
rect 14648 23268 14724 23302
rect 14539 23253 14724 23268
rect 14539 23219 14611 23253
rect 14645 23230 14724 23253
rect 14539 23196 14614 23219
rect 14648 23196 14724 23230
rect 14539 23185 14724 23196
rect 14539 23151 14611 23185
rect 14645 23158 14724 23185
rect 14539 23124 14614 23151
rect 14648 23124 14724 23158
rect 14539 23117 14724 23124
rect 14539 23083 14611 23117
rect 14645 23086 14724 23117
rect 14539 23052 14614 23083
rect 14648 23052 14724 23086
rect 14539 23049 14724 23052
rect 14539 23015 14611 23049
rect 14645 23015 14724 23049
rect 14539 23014 14724 23015
rect 14539 22981 14614 23014
rect 14539 22947 14611 22981
rect 14648 22980 14724 23014
rect 14645 22947 14724 22980
rect 14539 22942 14724 22947
rect 14539 22913 14614 22942
rect 14539 22879 14611 22913
rect 14648 22908 14724 22942
rect 14645 22879 14724 22908
rect 14539 22870 14724 22879
rect 14539 22845 14614 22870
rect 14539 22811 14611 22845
rect 14648 22836 14724 22870
rect 14645 22811 14724 22836
rect 14539 22798 14724 22811
rect 14539 22777 14614 22798
rect 14539 22743 14611 22777
rect 14648 22764 14724 22798
rect 14645 22743 14724 22764
rect 14539 22726 14724 22743
rect 14539 22709 14614 22726
rect 14539 22675 14611 22709
rect 14648 22692 14724 22726
rect 14645 22675 14724 22692
rect 14539 22654 14724 22675
rect 14539 22641 14614 22654
rect 14539 22607 14611 22641
rect 14648 22620 14724 22654
rect 14645 22607 14724 22620
rect 14539 22582 14724 22607
rect 14539 22573 14614 22582
rect 14539 22539 14611 22573
rect 14648 22548 14724 22582
rect 14645 22539 14724 22548
rect 14539 22510 14724 22539
rect 14539 22505 14614 22510
rect 14539 22471 14611 22505
rect 14648 22476 14724 22510
rect 14645 22471 14724 22476
rect 14539 22438 14724 22471
rect 14539 22437 14614 22438
rect 14539 22403 14611 22437
rect 14648 22404 14724 22438
rect 14645 22403 14724 22404
rect 14539 22369 14724 22403
rect 14539 22335 14611 22369
rect 14645 22366 14724 22369
rect 14539 22332 14614 22335
rect 14648 22332 14724 22366
rect 14539 22301 14724 22332
rect 14539 22267 14611 22301
rect 14645 22294 14724 22301
rect 14539 22260 14614 22267
rect 14648 22260 14724 22294
rect 14539 22233 14724 22260
rect 14539 22199 14611 22233
rect 14645 22222 14724 22233
rect 14539 22188 14614 22199
rect 14648 22188 14724 22222
rect 14539 22165 14724 22188
rect 14539 22131 14611 22165
rect 14645 22150 14724 22165
rect 14539 22116 14614 22131
rect 14648 22116 14724 22150
rect 14539 22097 14724 22116
rect 14539 22063 14611 22097
rect 14645 22078 14724 22097
rect 14539 22044 14614 22063
rect 14648 22044 14724 22078
rect 14539 22029 14724 22044
rect 14539 21995 14611 22029
rect 14645 22006 14724 22029
rect 14539 21972 14614 21995
rect 14648 21972 14724 22006
rect 14539 21961 14724 21972
rect 14539 21927 14611 21961
rect 14645 21934 14724 21961
rect 14539 21900 14614 21927
rect 14648 21900 14724 21934
rect 14539 21893 14724 21900
rect 14539 21859 14611 21893
rect 14645 21862 14724 21893
rect 14539 21828 14614 21859
rect 14648 21828 14724 21862
rect 14539 21825 14724 21828
rect 14539 21791 14611 21825
rect 14645 21791 14724 21825
rect 14539 21790 14724 21791
rect 14539 21757 14614 21790
rect 14539 21723 14611 21757
rect 14648 21756 14724 21790
rect 14645 21723 14724 21756
rect 14539 21718 14724 21723
rect 14539 21689 14614 21718
rect 14539 21655 14611 21689
rect 14648 21684 14724 21718
rect 14645 21655 14724 21684
rect 14539 21646 14724 21655
rect 14539 21621 14614 21646
rect 14539 21587 14611 21621
rect 14648 21612 14724 21646
rect 14645 21587 14724 21612
rect 14539 21574 14724 21587
rect 14539 21553 14614 21574
rect 14539 21519 14611 21553
rect 14648 21540 14724 21574
rect 14645 21519 14724 21540
rect 14539 21502 14724 21519
rect 14539 21485 14614 21502
rect 14539 21451 14611 21485
rect 14648 21468 14724 21502
rect 14645 21451 14724 21468
rect 14539 21430 14724 21451
rect 14539 21417 14614 21430
rect 14539 21383 14611 21417
rect 14648 21396 14724 21430
rect 14645 21383 14724 21396
rect 14539 21358 14724 21383
rect 14539 21349 14614 21358
rect 14539 21315 14611 21349
rect 14648 21324 14724 21358
rect 14645 21315 14724 21324
rect 14539 21286 14724 21315
rect 14539 21281 14614 21286
rect 14539 21247 14611 21281
rect 14648 21252 14724 21286
rect 14645 21247 14724 21252
rect 14539 21214 14724 21247
rect 14539 21213 14614 21214
rect 14539 21179 14611 21213
rect 14648 21180 14724 21214
rect 14645 21179 14724 21180
rect 14539 21145 14724 21179
rect 14539 21111 14611 21145
rect 14645 21142 14724 21145
rect 14539 21108 14614 21111
rect 14648 21108 14724 21142
rect 14539 21077 14724 21108
rect 14539 21043 14611 21077
rect 14645 21070 14724 21077
rect 14539 21036 14614 21043
rect 14648 21036 14724 21070
rect 14539 21009 14724 21036
rect 14539 20975 14611 21009
rect 14645 20998 14724 21009
rect 14539 20964 14614 20975
rect 14648 20964 14724 20998
rect 14539 20941 14724 20964
rect 14539 20907 14611 20941
rect 14645 20926 14724 20941
rect 14539 20892 14614 20907
rect 14648 20892 14724 20926
rect 14539 20873 14724 20892
rect 14539 20839 14611 20873
rect 14645 20854 14724 20873
rect 14539 20820 14614 20839
rect 14648 20820 14724 20854
rect 14539 20805 14724 20820
rect 14539 20771 14611 20805
rect 14645 20782 14724 20805
rect 14539 20748 14614 20771
rect 14648 20748 14724 20782
rect 14539 20737 14724 20748
rect 14539 20703 14611 20737
rect 14645 20710 14724 20737
rect 14539 20676 14614 20703
rect 14648 20676 14724 20710
rect 14539 20669 14724 20676
rect 14539 20635 14611 20669
rect 14645 20638 14724 20669
rect 14539 20604 14614 20635
rect 14648 20604 14724 20638
rect 14539 20601 14724 20604
rect 14539 20567 14611 20601
rect 14645 20567 14724 20601
rect 14539 20566 14724 20567
rect 14539 20533 14614 20566
rect 14539 20499 14611 20533
rect 14648 20532 14724 20566
rect 14645 20499 14724 20532
rect 14539 20494 14724 20499
rect 14539 20465 14614 20494
rect 14539 20431 14611 20465
rect 14648 20460 14724 20494
rect 14645 20431 14724 20460
rect 14539 20422 14724 20431
rect 14539 20397 14614 20422
rect 14539 20363 14611 20397
rect 14648 20388 14724 20422
rect 14645 20363 14724 20388
rect 14539 20350 14724 20363
rect 14539 20329 14614 20350
rect 14539 20295 14611 20329
rect 14648 20316 14724 20350
rect 14645 20295 14724 20316
rect 14539 20278 14724 20295
rect 14539 20261 14614 20278
rect 14539 20227 14611 20261
rect 14648 20244 14724 20278
rect 14645 20227 14724 20244
rect 14539 20206 14724 20227
rect 14539 20193 14614 20206
rect 14539 20159 14611 20193
rect 14648 20172 14724 20206
rect 14645 20159 14724 20172
rect 14539 20134 14724 20159
rect 14539 20125 14614 20134
rect 14539 20091 14611 20125
rect 14648 20100 14724 20134
rect 14645 20091 14724 20100
rect 14539 20062 14724 20091
rect 14539 20057 14614 20062
rect 14539 20023 14611 20057
rect 14648 20028 14724 20062
rect 14645 20023 14724 20028
rect 14539 19990 14724 20023
rect 14539 19989 14614 19990
rect 14539 19955 14611 19989
rect 14648 19956 14724 19990
rect 14645 19955 14724 19956
rect 14539 19921 14724 19955
rect 14539 19887 14611 19921
rect 14645 19918 14724 19921
rect 14539 19884 14614 19887
rect 14648 19884 14724 19918
rect 14539 19853 14724 19884
rect 14539 19819 14611 19853
rect 14645 19846 14724 19853
rect 14539 19812 14614 19819
rect 14648 19812 14724 19846
rect 14539 19785 14724 19812
rect 14539 19751 14611 19785
rect 14645 19774 14724 19785
rect 14539 19740 14614 19751
rect 14648 19740 14724 19774
rect 14539 19717 14724 19740
rect 14539 19683 14611 19717
rect 14645 19702 14724 19717
rect 14539 19668 14614 19683
rect 14648 19668 14724 19702
rect 14539 19649 14724 19668
rect 14539 19615 14611 19649
rect 14645 19630 14724 19649
rect 14539 19596 14614 19615
rect 14648 19596 14724 19630
rect 14539 19581 14724 19596
rect 14539 19547 14611 19581
rect 14645 19558 14724 19581
rect 14539 19524 14614 19547
rect 14648 19524 14724 19558
rect 14539 19513 14724 19524
rect 14539 19479 14611 19513
rect 14645 19486 14724 19513
rect 14539 19452 14614 19479
rect 14648 19452 14724 19486
rect 14539 19445 14724 19452
rect 14539 19411 14611 19445
rect 14645 19414 14724 19445
rect 14539 19380 14614 19411
rect 14648 19380 14724 19414
rect 14539 19377 14724 19380
rect 14539 19343 14611 19377
rect 14645 19343 14724 19377
rect 14539 19342 14724 19343
rect 14539 19309 14614 19342
rect 14539 19275 14611 19309
rect 14648 19308 14724 19342
rect 14645 19275 14724 19308
rect 14539 19270 14724 19275
rect 14539 19241 14614 19270
rect 14539 19207 14611 19241
rect 14648 19236 14724 19270
rect 14645 19207 14724 19236
rect 14539 19198 14724 19207
rect 14539 19173 14614 19198
rect 14539 19139 14611 19173
rect 14648 19164 14724 19198
rect 14645 19139 14724 19164
rect 14539 19126 14724 19139
rect 14539 19105 14614 19126
rect 14539 19071 14611 19105
rect 14648 19092 14724 19126
rect 14645 19071 14724 19092
rect 14539 19054 14724 19071
rect 14539 19037 14614 19054
rect 14539 19003 14611 19037
rect 14648 19020 14724 19054
rect 14645 19003 14724 19020
rect 14539 18982 14724 19003
rect 14539 18969 14614 18982
rect 14539 18935 14611 18969
rect 14648 18948 14724 18982
rect 14645 18935 14724 18948
rect 14539 18910 14724 18935
rect 14539 18901 14614 18910
rect 14539 18867 14611 18901
rect 14648 18876 14724 18910
rect 14645 18867 14724 18876
rect 14539 18838 14724 18867
rect 14539 18833 14614 18838
rect 14539 18799 14611 18833
rect 14648 18804 14724 18838
rect 14645 18799 14724 18804
rect 14539 18766 14724 18799
rect 14539 18765 14614 18766
rect 14539 18731 14611 18765
rect 14648 18732 14724 18766
rect 14645 18731 14724 18732
rect 14539 18697 14724 18731
rect 14539 18663 14611 18697
rect 14645 18694 14724 18697
rect 14539 18660 14614 18663
rect 14648 18660 14724 18694
rect 14539 18629 14724 18660
rect 14539 18595 14611 18629
rect 14645 18622 14724 18629
rect 14539 18588 14614 18595
rect 14648 18588 14724 18622
rect 14539 18561 14724 18588
rect 14539 18527 14611 18561
rect 14645 18550 14724 18561
rect 14539 18516 14614 18527
rect 14648 18516 14724 18550
rect 14539 18493 14724 18516
rect 14539 18459 14611 18493
rect 14645 18478 14724 18493
rect 14539 18444 14614 18459
rect 14648 18444 14724 18478
rect 14539 18425 14724 18444
rect 14539 18391 14611 18425
rect 14645 18406 14724 18425
rect 14539 18372 14614 18391
rect 14648 18372 14724 18406
rect 14539 18357 14724 18372
rect 14539 18323 14611 18357
rect 14645 18334 14724 18357
rect 14539 18300 14614 18323
rect 14648 18300 14724 18334
rect 14539 18289 14724 18300
rect 14539 18255 14611 18289
rect 14645 18262 14724 18289
rect 14539 18228 14614 18255
rect 14648 18228 14724 18262
rect 14539 18221 14724 18228
rect 14539 18187 14611 18221
rect 14645 18190 14724 18221
rect 14539 18156 14614 18187
rect 14648 18156 14724 18190
rect 14539 18153 14724 18156
rect 14539 18119 14611 18153
rect 14645 18119 14724 18153
rect 14539 18118 14724 18119
rect 14539 18085 14614 18118
rect 14539 18051 14611 18085
rect 14648 18084 14724 18118
rect 14645 18051 14724 18084
rect 14539 18046 14724 18051
rect 14539 18017 14614 18046
rect 14539 17983 14611 18017
rect 14648 18012 14724 18046
rect 14645 17983 14724 18012
rect 14539 17974 14724 17983
rect 14539 17949 14614 17974
rect 14539 17915 14611 17949
rect 14648 17940 14724 17974
rect 14645 17915 14724 17940
rect 14539 17902 14724 17915
rect 14539 17881 14614 17902
rect 14539 17847 14611 17881
rect 14648 17868 14724 17902
rect 14645 17847 14724 17868
rect 14539 17830 14724 17847
rect 14539 17813 14614 17830
rect 14539 17779 14611 17813
rect 14648 17796 14724 17830
rect 14645 17779 14724 17796
rect 14539 17758 14724 17779
rect 14539 17745 14614 17758
rect 14539 17711 14611 17745
rect 14648 17724 14724 17758
rect 14645 17711 14724 17724
rect 14539 17686 14724 17711
rect 14539 17677 14614 17686
rect 14539 17643 14611 17677
rect 14648 17652 14724 17686
rect 14645 17643 14724 17652
rect 14539 17614 14724 17643
rect 14539 17609 14614 17614
rect 14539 17575 14611 17609
rect 14648 17580 14724 17614
rect 14645 17575 14724 17580
rect 14539 17542 14724 17575
rect 14539 17541 14614 17542
rect 14539 17507 14611 17541
rect 14648 17508 14724 17542
rect 14645 17507 14724 17508
rect 14539 17473 14724 17507
rect 14539 17439 14611 17473
rect 14645 17470 14724 17473
rect 14539 17436 14614 17439
rect 14648 17436 14724 17470
rect 14539 17405 14724 17436
rect 14539 17371 14611 17405
rect 14645 17398 14724 17405
rect 14539 17364 14614 17371
rect 14648 17364 14724 17398
rect 14539 17337 14724 17364
rect 14539 17303 14611 17337
rect 14645 17326 14724 17337
rect 14539 17292 14614 17303
rect 14648 17292 14724 17326
rect 14539 17269 14724 17292
rect 14539 17235 14611 17269
rect 14645 17254 14724 17269
rect 14539 17220 14614 17235
rect 14648 17220 14724 17254
rect 14539 17201 14724 17220
rect 14539 17167 14611 17201
rect 14645 17182 14724 17201
rect 14539 17148 14614 17167
rect 14648 17148 14724 17182
rect 14539 17133 14724 17148
rect 14539 17099 14611 17133
rect 14645 17110 14724 17133
rect 14539 17076 14614 17099
rect 14648 17076 14724 17110
rect 14539 17065 14724 17076
rect 14539 17031 14611 17065
rect 14645 17038 14724 17065
rect 14539 17004 14614 17031
rect 14648 17004 14724 17038
rect 14539 16997 14724 17004
rect 14539 16963 14611 16997
rect 14645 16966 14724 16997
rect 14539 16932 14614 16963
rect 14648 16932 14724 16966
rect 14539 16929 14724 16932
rect 14539 16895 14611 16929
rect 14645 16895 14724 16929
rect 14539 16894 14724 16895
rect 14539 16861 14614 16894
rect 14539 16827 14611 16861
rect 14648 16860 14724 16894
rect 14645 16827 14724 16860
rect 14539 16822 14724 16827
rect 14539 16793 14614 16822
rect 14539 16759 14611 16793
rect 14648 16788 14724 16822
rect 14645 16759 14724 16788
rect 14539 16750 14724 16759
rect 14539 16725 14614 16750
rect 14539 16691 14611 16725
rect 14648 16716 14724 16750
rect 14645 16691 14724 16716
rect 14539 16678 14724 16691
rect 14539 16657 14614 16678
rect 14539 16623 14611 16657
rect 14648 16644 14724 16678
rect 14645 16623 14724 16644
rect 14539 16606 14724 16623
rect 14539 16589 14614 16606
rect 14539 16555 14611 16589
rect 14648 16572 14724 16606
rect 14645 16555 14724 16572
rect 14539 16534 14724 16555
rect 14539 16521 14614 16534
rect 14539 16487 14611 16521
rect 14648 16500 14724 16534
rect 14645 16487 14724 16500
rect 14539 16462 14724 16487
rect 14539 16453 14614 16462
rect 14539 16419 14611 16453
rect 14648 16428 14724 16462
rect 14645 16419 14724 16428
rect 14539 16390 14724 16419
rect 14539 16385 14614 16390
rect 14539 16351 14611 16385
rect 14648 16356 14724 16390
rect 14645 16351 14724 16356
rect 14539 16318 14724 16351
rect 14539 16317 14614 16318
rect 14539 16283 14611 16317
rect 14648 16284 14724 16318
rect 14645 16283 14724 16284
rect 14539 16249 14724 16283
rect 14539 16215 14611 16249
rect 14645 16246 14724 16249
rect 14539 16212 14614 16215
rect 14648 16212 14724 16246
rect 14539 16181 14724 16212
rect 14539 16147 14611 16181
rect 14645 16174 14724 16181
rect 14539 16140 14614 16147
rect 14648 16140 14724 16174
rect 14539 16113 14724 16140
rect 14539 16079 14611 16113
rect 14645 16102 14724 16113
rect 14539 16068 14614 16079
rect 14648 16068 14724 16102
rect 14539 16045 14724 16068
rect 14539 16011 14611 16045
rect 14645 16030 14724 16045
rect 14539 15996 14614 16011
rect 14648 15996 14724 16030
rect 14539 15977 14724 15996
rect 14539 15943 14611 15977
rect 14645 15958 14724 15977
rect 14539 15924 14614 15943
rect 14648 15924 14724 15958
rect 14539 15909 14724 15924
rect 14539 15875 14611 15909
rect 14645 15886 14724 15909
rect 14539 15852 14614 15875
rect 14648 15852 14724 15886
rect 14539 15841 14724 15852
rect 14539 15807 14611 15841
rect 14645 15814 14724 15841
rect 14539 15780 14614 15807
rect 14648 15780 14724 15814
rect 14539 15773 14724 15780
rect 14539 15739 14611 15773
rect 14645 15742 14724 15773
rect 14539 15708 14614 15739
rect 14648 15708 14724 15742
rect 14539 15705 14724 15708
rect 14539 15671 14611 15705
rect 14645 15671 14724 15705
rect 14539 15670 14724 15671
rect 14539 15637 14614 15670
rect 14539 15603 14611 15637
rect 14648 15636 14724 15670
rect 14645 15603 14724 15636
rect 14539 15598 14724 15603
rect 14539 15569 14614 15598
rect 14539 15535 14611 15569
rect 14648 15564 14724 15598
rect 14645 15535 14724 15564
rect 14539 15526 14724 15535
rect 14539 15501 14614 15526
rect 14539 15467 14611 15501
rect 14648 15492 14724 15526
rect 14645 15467 14724 15492
rect 14539 15454 14724 15467
rect 14539 15433 14614 15454
rect 14539 15399 14611 15433
rect 14648 15420 14724 15454
rect 14645 15399 14724 15420
rect 14539 15382 14724 15399
rect 14539 15365 14614 15382
rect 14539 15331 14611 15365
rect 14648 15348 14724 15382
rect 14645 15331 14724 15348
rect 14539 15310 14724 15331
rect 14539 15297 14614 15310
rect 14539 15263 14611 15297
rect 14648 15276 14724 15310
rect 14645 15263 14724 15276
rect 14539 15238 14724 15263
rect 14539 15229 14614 15238
rect 14539 15195 14611 15229
rect 14648 15204 14724 15238
rect 14645 15195 14724 15204
rect 14539 15166 14724 15195
rect 14539 15161 14614 15166
rect 14539 15127 14611 15161
rect 14648 15132 14724 15166
rect 14645 15127 14724 15132
rect 14539 15094 14724 15127
rect 14539 15093 14614 15094
rect 14539 15059 14611 15093
rect 14648 15060 14724 15094
rect 14645 15059 14724 15060
rect 14539 15025 14724 15059
rect 14539 14991 14611 15025
rect 14645 15022 14724 15025
rect 14539 14988 14614 14991
rect 14648 14988 14724 15022
rect 14539 14957 14724 14988
rect 14539 14923 14611 14957
rect 14645 14950 14724 14957
rect 14539 14916 14614 14923
rect 14648 14916 14724 14950
rect 14539 14889 14724 14916
rect 14539 14855 14611 14889
rect 14645 14878 14724 14889
rect 14539 14844 14614 14855
rect 14648 14844 14724 14878
rect 14539 14821 14724 14844
rect 14539 14787 14611 14821
rect 14645 14806 14724 14821
rect 14539 14772 14614 14787
rect 14648 14772 14724 14806
rect 14539 14753 14724 14772
rect 14539 14719 14611 14753
rect 14645 14734 14724 14753
rect 14539 14700 14614 14719
rect 14648 14700 14724 14734
rect 14539 14685 14724 14700
rect 14539 14651 14611 14685
rect 14645 14662 14724 14685
rect 14539 14628 14614 14651
rect 14648 14628 14724 14662
rect 14539 14617 14724 14628
rect 14539 14583 14611 14617
rect 14645 14590 14724 14617
rect 14539 14556 14614 14583
rect 14648 14556 14724 14590
rect 14539 14549 14724 14556
rect 14539 14515 14611 14549
rect 14645 14518 14724 14549
rect 14539 14484 14614 14515
rect 14648 14484 14724 14518
rect 14539 14481 14724 14484
rect 14539 14447 14611 14481
rect 14645 14447 14724 14481
rect 14539 14446 14724 14447
rect 14539 14413 14614 14446
rect 14539 14379 14611 14413
rect 14648 14412 14724 14446
rect 14645 14379 14724 14412
rect 14539 14374 14724 14379
rect 14539 14345 14614 14374
rect 14539 14311 14611 14345
rect 14648 14340 14724 14374
rect 14645 14311 14724 14340
rect 14539 14302 14724 14311
rect 14539 14277 14614 14302
rect 14539 14243 14611 14277
rect 14648 14268 14724 14302
rect 14645 14243 14724 14268
rect 14539 14230 14724 14243
rect 14539 14209 14614 14230
rect 14539 14175 14611 14209
rect 14648 14196 14724 14230
rect 14645 14175 14724 14196
rect 14539 14158 14724 14175
rect 14539 14141 14614 14158
rect 14539 14107 14611 14141
rect 14648 14124 14724 14158
rect 14645 14107 14724 14124
rect 14539 14086 14724 14107
rect 14539 14073 14614 14086
rect 14539 14039 14611 14073
rect 14648 14052 14724 14086
rect 14645 14039 14724 14052
rect 14539 14014 14724 14039
rect 14539 14005 14614 14014
rect 14539 13971 14611 14005
rect 14648 13980 14724 14014
rect 14645 13971 14724 13980
rect 14539 13942 14724 13971
rect 14539 13937 14614 13942
rect 14539 13903 14611 13937
rect 14648 13908 14724 13942
rect 14645 13903 14724 13908
rect 14539 13870 14724 13903
rect 14539 13869 14614 13870
rect 14539 13835 14611 13869
rect 14648 13836 14724 13870
rect 14645 13835 14724 13836
rect 14539 13801 14724 13835
rect 14539 13767 14611 13801
rect 14645 13798 14724 13801
rect 14539 13764 14614 13767
rect 14648 13764 14724 13798
rect 14539 13733 14724 13764
rect 14539 13699 14611 13733
rect 14645 13726 14724 13733
rect 14539 13692 14614 13699
rect 14648 13692 14724 13726
rect 14539 13665 14724 13692
rect 14539 13631 14611 13665
rect 14645 13654 14724 13665
rect 14539 13620 14614 13631
rect 14648 13620 14724 13654
rect 14539 13597 14724 13620
rect 14539 13563 14611 13597
rect 14645 13582 14724 13597
rect 14539 13548 14614 13563
rect 14648 13548 14724 13582
rect 14539 13529 14724 13548
rect 14539 13495 14611 13529
rect 14645 13510 14724 13529
rect 14539 13476 14614 13495
rect 14648 13476 14724 13510
rect 14539 13461 14724 13476
rect 14539 13427 14611 13461
rect 14645 13438 14724 13461
rect 14539 13404 14614 13427
rect 14648 13404 14724 13438
rect 14539 13393 14724 13404
rect 14539 13359 14611 13393
rect 14645 13366 14724 13393
rect 14539 13332 14614 13359
rect 14648 13332 14724 13366
rect 14539 13325 14724 13332
rect 14539 13291 14611 13325
rect 14645 13294 14724 13325
rect 14539 13260 14614 13291
rect 14648 13260 14724 13294
rect 14539 13257 14724 13260
rect 14539 13223 14611 13257
rect 14645 13223 14724 13257
rect 14539 13222 14724 13223
rect 14539 13189 14614 13222
rect 14539 13155 14611 13189
rect 14648 13188 14724 13222
rect 14645 13155 14724 13188
rect 14539 13150 14724 13155
rect 14539 13121 14614 13150
rect 14539 13087 14611 13121
rect 14648 13116 14724 13150
rect 14645 13087 14724 13116
rect 14539 13078 14724 13087
rect 14539 13053 14614 13078
rect 14539 13019 14611 13053
rect 14648 13044 14724 13078
rect 14645 13019 14724 13044
rect 14539 13006 14724 13019
rect 14539 12985 14614 13006
rect 14539 12951 14611 12985
rect 14648 12972 14724 13006
rect 14645 12951 14724 12972
rect 14539 12934 14724 12951
rect 14539 12917 14614 12934
rect 14539 12883 14611 12917
rect 14648 12900 14724 12934
rect 14645 12883 14724 12900
rect 14539 12862 14724 12883
rect 14539 12849 14614 12862
rect 14539 12815 14611 12849
rect 14648 12828 14724 12862
rect 14645 12815 14724 12828
rect 14539 12790 14724 12815
rect 14539 12781 14614 12790
rect 14539 12747 14611 12781
rect 14648 12756 14724 12790
rect 14645 12747 14724 12756
rect 14539 12718 14724 12747
rect 14539 12713 14614 12718
rect 14539 12679 14611 12713
rect 14648 12684 14724 12718
rect 14645 12679 14724 12684
rect 14539 12646 14724 12679
rect 14539 12645 14614 12646
rect 14539 12611 14611 12645
rect 14648 12612 14724 12646
rect 14645 12611 14724 12612
rect 14539 12577 14724 12611
rect 14539 12543 14611 12577
rect 14645 12574 14724 12577
rect 14539 12540 14614 12543
rect 14648 12540 14724 12574
rect 14539 12509 14724 12540
rect 14539 12475 14611 12509
rect 14645 12502 14724 12509
rect 14539 12468 14614 12475
rect 14648 12468 14724 12502
rect 14539 12441 14724 12468
rect 14539 12407 14611 12441
rect 14645 12430 14724 12441
rect 14539 12396 14614 12407
rect 14648 12396 14724 12430
rect 14539 12373 14724 12396
rect 14539 12339 14611 12373
rect 14645 12358 14724 12373
rect 14539 12324 14614 12339
rect 14648 12324 14724 12358
rect 14539 12305 14724 12324
rect 14539 12271 14611 12305
rect 14645 12286 14724 12305
rect 14539 12252 14614 12271
rect 14648 12252 14724 12286
rect 14539 12237 14724 12252
rect 14539 12203 14611 12237
rect 14645 12214 14724 12237
rect 14539 12180 14614 12203
rect 14648 12180 14724 12214
rect 14539 12169 14724 12180
rect 14539 12135 14611 12169
rect 14645 12142 14724 12169
rect 14539 12108 14614 12135
rect 14648 12108 14724 12142
rect 14539 12101 14724 12108
rect 14539 12067 14611 12101
rect 14645 12070 14724 12101
rect 14539 12036 14614 12067
rect 14648 12036 14724 12070
rect 14539 12033 14724 12036
rect 14539 11999 14611 12033
rect 14645 11999 14724 12033
rect 14539 11998 14724 11999
rect 14539 11965 14614 11998
rect 14539 11931 14611 11965
rect 14648 11964 14724 11998
rect 14645 11931 14724 11964
rect 14539 11926 14724 11931
rect 14539 11897 14614 11926
rect 14539 11863 14611 11897
rect 14648 11892 14724 11926
rect 14645 11863 14724 11892
rect 14539 11854 14724 11863
rect 14539 11829 14614 11854
rect 14539 11795 14611 11829
rect 14648 11820 14724 11854
rect 14645 11795 14724 11820
rect 14539 11782 14724 11795
rect 14539 11761 14614 11782
rect 14539 11727 14611 11761
rect 14648 11748 14724 11782
rect 14645 11727 14724 11748
rect 14539 11710 14724 11727
rect 14539 11693 14614 11710
rect 14539 11659 14611 11693
rect 14648 11676 14724 11710
rect 14645 11659 14724 11676
rect 14539 11638 14724 11659
rect 14539 11625 14614 11638
rect 14539 11591 14611 11625
rect 14648 11604 14724 11638
rect 14645 11591 14724 11604
rect 14539 11566 14724 11591
rect 14539 11557 14614 11566
rect 14539 11523 14611 11557
rect 14648 11532 14724 11566
rect 14645 11523 14724 11532
rect 14539 11494 14724 11523
rect 14539 11489 14614 11494
rect 14539 11455 14611 11489
rect 14648 11460 14724 11494
rect 14645 11455 14724 11460
rect 14539 11422 14724 11455
rect 14539 11421 14614 11422
rect 14539 11387 14611 11421
rect 14648 11388 14724 11422
rect 14645 11387 14724 11388
rect 14539 11353 14724 11387
rect 14539 11319 14611 11353
rect 14645 11350 14724 11353
rect 14539 11316 14614 11319
rect 14648 11316 14724 11350
rect 14539 11285 14724 11316
rect 14539 11251 14611 11285
rect 14645 11278 14724 11285
rect 14539 11244 14614 11251
rect 14648 11244 14724 11278
rect 14539 11217 14724 11244
rect 14539 11183 14611 11217
rect 14645 11206 14724 11217
rect 14539 11172 14614 11183
rect 14648 11172 14724 11206
rect 14539 11149 14724 11172
rect 14539 11115 14611 11149
rect 14645 11134 14724 11149
rect 14539 11100 14614 11115
rect 14648 11100 14724 11134
rect 14539 11081 14724 11100
rect 14539 11047 14611 11081
rect 14645 11062 14724 11081
rect 14539 11028 14614 11047
rect 14648 11028 14724 11062
rect 14539 11013 14724 11028
rect 14539 10979 14611 11013
rect 14645 10990 14724 11013
rect 14539 10956 14614 10979
rect 14648 10956 14724 10990
rect 14539 10945 14724 10956
rect 14539 10911 14611 10945
rect 14645 10918 14724 10945
rect 14539 10884 14614 10911
rect 14648 10884 14724 10918
rect 14539 10877 14724 10884
rect 14539 10843 14611 10877
rect 14645 10846 14724 10877
rect 14539 10812 14614 10843
rect 14648 10812 14724 10846
rect 14539 10809 14724 10812
rect 14539 10775 14611 10809
rect 14645 10775 14724 10809
rect 14539 10774 14724 10775
rect 14539 10741 14614 10774
rect 14539 10707 14611 10741
rect 14648 10740 14724 10774
rect 14645 10707 14724 10740
rect 14539 10702 14724 10707
rect 14539 10673 14614 10702
rect 14539 10639 14611 10673
rect 14648 10668 14724 10702
rect 14645 10639 14724 10668
rect 14539 10630 14724 10639
rect 14539 10605 14614 10630
rect 14539 10571 14611 10605
rect 14648 10596 14724 10630
rect 14645 10571 14724 10596
rect 14539 10558 14724 10571
rect 14539 10537 14614 10558
rect 14539 10503 14611 10537
rect 14648 10524 14724 10558
rect 14645 10503 14724 10524
rect 14539 10486 14724 10503
rect 14539 10469 14614 10486
rect 14539 10435 14611 10469
rect 14648 10452 14724 10486
rect 14645 10435 14724 10452
rect 14539 10414 14724 10435
rect 14539 10401 14614 10414
rect 14539 10367 14611 10401
rect 14648 10380 14724 10414
rect 14645 10367 14724 10380
rect 14539 10342 14724 10367
rect 14539 10333 14614 10342
rect 14539 10299 14611 10333
rect 14648 10308 14724 10342
rect 14645 10299 14724 10308
rect 14539 10270 14724 10299
rect 14539 10265 14614 10270
rect 14539 10231 14611 10265
rect 14648 10236 14724 10270
rect 14645 10231 14724 10236
rect 14539 10198 14724 10231
rect 14539 10197 14614 10198
rect 14539 10163 14611 10197
rect 14648 10164 14724 10198
rect 14645 10163 14724 10164
rect 14539 10129 14724 10163
rect 14539 10095 14611 10129
rect 14645 10126 14724 10129
rect 14539 10092 14614 10095
rect 14648 10092 14724 10126
rect 14539 10061 14724 10092
rect 14539 10027 14611 10061
rect 14645 10054 14724 10061
rect 14539 10020 14614 10027
rect 14648 10020 14724 10054
rect 14539 9993 14724 10020
rect 14539 9959 14611 9993
rect 14645 9982 14724 9993
rect 14539 9948 14614 9959
rect 14648 9948 14724 9982
rect 14539 9925 14724 9948
rect 14539 9891 14611 9925
rect 14645 9910 14724 9925
rect 14539 9876 14614 9891
rect 14648 9876 14724 9910
rect 14539 9857 14724 9876
rect 14539 9823 14611 9857
rect 14645 9838 14724 9857
rect 14539 9804 14614 9823
rect 14648 9804 14724 9838
rect 14539 9789 14724 9804
rect 14539 9755 14611 9789
rect 14645 9766 14724 9789
rect 14539 9732 14614 9755
rect 14648 9732 14724 9766
rect 14539 9721 14724 9732
rect 245 9663 320 9689
rect 354 9663 430 9697
rect 245 9655 430 9663
rect 245 9621 317 9655
rect 351 9621 430 9655
rect 245 9528 430 9621
rect 14539 9687 14611 9721
rect 14645 9694 14724 9721
rect 14539 9660 14614 9687
rect 14648 9660 14724 9694
rect 14539 9653 14724 9660
rect 14539 9619 14611 9653
rect 14645 9619 14724 9653
rect 14539 9528 14724 9619
rect 245 9452 14724 9528
rect 245 9418 320 9452
rect 354 9450 610 9452
rect 644 9450 2311 9452
rect 2345 9450 2383 9452
rect 2417 9450 2455 9452
rect 2489 9450 2527 9452
rect 2561 9450 2599 9452
rect 2633 9450 2671 9452
rect 2705 9450 2743 9452
rect 2777 9450 2815 9452
rect 2849 9450 2887 9452
rect 2921 9450 2959 9452
rect 2993 9450 3031 9452
rect 3065 9450 3103 9452
rect 3137 9450 3175 9452
rect 3209 9450 3247 9452
rect 3281 9450 3319 9452
rect 3353 9450 3391 9452
rect 3425 9450 3463 9452
rect 3497 9450 3535 9452
rect 3569 9450 3607 9452
rect 3641 9450 3679 9452
rect 3713 9450 3751 9452
rect 3785 9450 3823 9452
rect 3857 9450 3895 9452
rect 3929 9450 3967 9452
rect 4001 9450 4039 9452
rect 4073 9450 4111 9452
rect 4145 9450 4183 9452
rect 4217 9450 4255 9452
rect 4289 9450 4327 9452
rect 4361 9450 4399 9452
rect 4433 9450 4471 9452
rect 4505 9450 4543 9452
rect 4577 9450 4615 9452
rect 4649 9450 4687 9452
rect 4721 9450 4759 9452
rect 4793 9450 4831 9452
rect 4865 9450 4903 9452
rect 4937 9450 4975 9452
rect 5009 9450 5047 9452
rect 5081 9450 5119 9452
rect 5153 9450 5191 9452
rect 5225 9450 5263 9452
rect 5297 9450 5335 9452
rect 5369 9450 5407 9452
rect 5441 9450 5479 9452
rect 5513 9450 5551 9452
rect 5585 9450 5623 9452
rect 5657 9450 5695 9452
rect 5729 9450 5767 9452
rect 5801 9450 5839 9452
rect 5873 9450 5911 9452
rect 5945 9450 5983 9452
rect 6017 9450 6055 9452
rect 6089 9450 6127 9452
rect 6161 9450 6199 9452
rect 6233 9450 6271 9452
rect 6305 9450 6343 9452
rect 6377 9450 6415 9452
rect 6449 9450 6487 9452
rect 6521 9450 6559 9452
rect 6593 9450 6631 9452
rect 6665 9450 6703 9452
rect 6737 9450 6775 9452
rect 6809 9450 6847 9452
rect 6881 9450 6919 9452
rect 6953 9450 6991 9452
rect 7025 9450 7063 9452
rect 7097 9450 7135 9452
rect 7169 9450 7207 9452
rect 7241 9450 7279 9452
rect 7313 9450 7351 9452
rect 7385 9450 7423 9452
rect 7457 9450 7495 9452
rect 7529 9450 7567 9452
rect 7601 9450 7639 9452
rect 7673 9450 7711 9452
rect 7745 9450 7783 9452
rect 7817 9450 7855 9452
rect 7889 9450 7927 9452
rect 7961 9450 7999 9452
rect 8033 9450 8071 9452
rect 8105 9450 8143 9452
rect 8177 9450 8215 9452
rect 8249 9450 8287 9452
rect 8321 9450 8359 9452
rect 8393 9450 8431 9452
rect 8465 9450 8503 9452
rect 8537 9450 8575 9452
rect 8609 9450 8647 9452
rect 8681 9450 8719 9452
rect 8753 9450 8791 9452
rect 8825 9450 8863 9452
rect 8897 9450 8935 9452
rect 8969 9450 9007 9452
rect 9041 9450 9079 9452
rect 9113 9450 9151 9452
rect 9185 9450 9223 9452
rect 9257 9450 9295 9452
rect 9329 9450 9367 9452
rect 9401 9450 9439 9452
rect 9473 9450 9511 9452
rect 9545 9450 9583 9452
rect 9617 9450 9655 9452
rect 9689 9450 9727 9452
rect 9761 9450 9799 9452
rect 9833 9450 9871 9452
rect 9905 9450 9943 9452
rect 9977 9450 10015 9452
rect 10049 9450 10087 9452
rect 10121 9450 10159 9452
rect 10193 9450 10231 9452
rect 10265 9450 10303 9452
rect 10337 9450 10375 9452
rect 10409 9450 10447 9452
rect 10481 9450 10519 9452
rect 10553 9450 10591 9452
rect 10625 9450 10663 9452
rect 10697 9450 10735 9452
rect 10769 9450 10807 9452
rect 10841 9450 10879 9452
rect 10913 9450 10951 9452
rect 10985 9450 11023 9452
rect 11057 9450 11095 9452
rect 11129 9450 11167 9452
rect 11201 9450 11239 9452
rect 11273 9450 11311 9452
rect 11345 9450 11383 9452
rect 11417 9450 11455 9452
rect 11489 9450 11527 9452
rect 11561 9450 11599 9452
rect 11633 9450 11671 9452
rect 11705 9450 11743 9452
rect 11777 9450 11815 9452
rect 11849 9450 11887 9452
rect 11921 9450 11959 9452
rect 11993 9450 12031 9452
rect 12065 9450 12103 9452
rect 12137 9450 12175 9452
rect 12209 9450 12247 9452
rect 12281 9450 12319 9452
rect 12353 9450 12391 9452
rect 12425 9450 12463 9452
rect 12497 9450 12535 9452
rect 12569 9450 12607 9452
rect 12641 9450 14314 9452
rect 14348 9450 14614 9452
rect 354 9418 506 9450
rect 245 9416 506 9418
rect 540 9416 574 9450
rect 608 9418 610 9450
rect 608 9416 642 9418
rect 676 9416 710 9450
rect 744 9416 778 9450
rect 812 9416 846 9450
rect 880 9416 914 9450
rect 948 9416 982 9450
rect 1016 9416 1050 9450
rect 1084 9416 1118 9450
rect 1152 9416 1186 9450
rect 1220 9416 1254 9450
rect 1288 9416 1322 9450
rect 1356 9416 1390 9450
rect 1424 9416 1458 9450
rect 1492 9416 1526 9450
rect 1560 9416 1594 9450
rect 1628 9416 1662 9450
rect 1696 9416 1730 9450
rect 1764 9416 1798 9450
rect 1832 9416 1866 9450
rect 1900 9416 1934 9450
rect 1968 9416 2002 9450
rect 2036 9416 2070 9450
rect 2104 9416 2138 9450
rect 2172 9416 2206 9450
rect 2240 9416 2274 9450
rect 2308 9418 2311 9450
rect 2376 9418 2383 9450
rect 2444 9418 2455 9450
rect 2512 9418 2527 9450
rect 2580 9418 2599 9450
rect 2648 9418 2671 9450
rect 2716 9418 2743 9450
rect 2784 9418 2815 9450
rect 2308 9416 2342 9418
rect 2376 9416 2410 9418
rect 2444 9416 2478 9418
rect 2512 9416 2546 9418
rect 2580 9416 2614 9418
rect 2648 9416 2682 9418
rect 2716 9416 2750 9418
rect 2784 9416 2818 9418
rect 2852 9416 2886 9450
rect 2921 9418 2954 9450
rect 2993 9418 3022 9450
rect 3065 9418 3090 9450
rect 3137 9418 3158 9450
rect 3209 9418 3226 9450
rect 3281 9418 3294 9450
rect 3353 9418 3362 9450
rect 3425 9418 3430 9450
rect 3497 9418 3498 9450
rect 2920 9416 2954 9418
rect 2988 9416 3022 9418
rect 3056 9416 3090 9418
rect 3124 9416 3158 9418
rect 3192 9416 3226 9418
rect 3260 9416 3294 9418
rect 3328 9416 3362 9418
rect 3396 9416 3430 9418
rect 3464 9416 3498 9418
rect 3532 9418 3535 9450
rect 3600 9418 3607 9450
rect 3668 9418 3679 9450
rect 3736 9418 3751 9450
rect 3804 9418 3823 9450
rect 3872 9418 3895 9450
rect 3940 9418 3967 9450
rect 4008 9418 4039 9450
rect 3532 9416 3566 9418
rect 3600 9416 3634 9418
rect 3668 9416 3702 9418
rect 3736 9416 3770 9418
rect 3804 9416 3838 9418
rect 3872 9416 3906 9418
rect 3940 9416 3974 9418
rect 4008 9416 4042 9418
rect 4076 9416 4110 9450
rect 4145 9418 4178 9450
rect 4217 9418 4246 9450
rect 4289 9418 4314 9450
rect 4361 9418 4382 9450
rect 4433 9418 4450 9450
rect 4505 9418 4518 9450
rect 4577 9418 4586 9450
rect 4649 9418 4654 9450
rect 4721 9418 4722 9450
rect 4144 9416 4178 9418
rect 4212 9416 4246 9418
rect 4280 9416 4314 9418
rect 4348 9416 4382 9418
rect 4416 9416 4450 9418
rect 4484 9416 4518 9418
rect 4552 9416 4586 9418
rect 4620 9416 4654 9418
rect 4688 9416 4722 9418
rect 4756 9418 4759 9450
rect 4824 9418 4831 9450
rect 4892 9418 4903 9450
rect 4960 9418 4975 9450
rect 5028 9418 5047 9450
rect 5096 9418 5119 9450
rect 5164 9418 5191 9450
rect 5232 9418 5263 9450
rect 4756 9416 4790 9418
rect 4824 9416 4858 9418
rect 4892 9416 4926 9418
rect 4960 9416 4994 9418
rect 5028 9416 5062 9418
rect 5096 9416 5130 9418
rect 5164 9416 5198 9418
rect 5232 9416 5266 9418
rect 5300 9416 5334 9450
rect 5369 9418 5402 9450
rect 5441 9418 5470 9450
rect 5513 9418 5538 9450
rect 5585 9418 5606 9450
rect 5657 9418 5674 9450
rect 5729 9418 5742 9450
rect 5801 9418 5810 9450
rect 5873 9418 5878 9450
rect 5945 9418 5946 9450
rect 5368 9416 5402 9418
rect 5436 9416 5470 9418
rect 5504 9416 5538 9418
rect 5572 9416 5606 9418
rect 5640 9416 5674 9418
rect 5708 9416 5742 9418
rect 5776 9416 5810 9418
rect 5844 9416 5878 9418
rect 5912 9416 5946 9418
rect 5980 9418 5983 9450
rect 6048 9418 6055 9450
rect 6116 9418 6127 9450
rect 6184 9418 6199 9450
rect 6252 9418 6271 9450
rect 6320 9418 6343 9450
rect 6388 9418 6415 9450
rect 6456 9418 6487 9450
rect 5980 9416 6014 9418
rect 6048 9416 6082 9418
rect 6116 9416 6150 9418
rect 6184 9416 6218 9418
rect 6252 9416 6286 9418
rect 6320 9416 6354 9418
rect 6388 9416 6422 9418
rect 6456 9416 6490 9418
rect 6524 9416 6558 9450
rect 6593 9418 6626 9450
rect 6665 9418 6694 9450
rect 6737 9418 6762 9450
rect 6809 9418 6830 9450
rect 6881 9418 6898 9450
rect 6953 9418 6966 9450
rect 7025 9418 7034 9450
rect 7097 9418 7102 9450
rect 7169 9418 7170 9450
rect 6592 9416 6626 9418
rect 6660 9416 6694 9418
rect 6728 9416 6762 9418
rect 6796 9416 6830 9418
rect 6864 9416 6898 9418
rect 6932 9416 6966 9418
rect 7000 9416 7034 9418
rect 7068 9416 7102 9418
rect 7136 9416 7170 9418
rect 7204 9418 7207 9450
rect 7272 9418 7279 9450
rect 7340 9418 7351 9450
rect 7408 9418 7423 9450
rect 7476 9418 7495 9450
rect 7544 9418 7567 9450
rect 7612 9418 7639 9450
rect 7680 9418 7711 9450
rect 7204 9416 7238 9418
rect 7272 9416 7306 9418
rect 7340 9416 7374 9418
rect 7408 9416 7442 9418
rect 7476 9416 7510 9418
rect 7544 9416 7578 9418
rect 7612 9416 7646 9418
rect 7680 9416 7714 9418
rect 7748 9416 7782 9450
rect 7817 9418 7850 9450
rect 7889 9418 7918 9450
rect 7961 9418 7986 9450
rect 8033 9418 8054 9450
rect 8105 9418 8122 9450
rect 8177 9418 8190 9450
rect 8249 9418 8258 9450
rect 8321 9418 8326 9450
rect 8393 9418 8394 9450
rect 7816 9416 7850 9418
rect 7884 9416 7918 9418
rect 7952 9416 7986 9418
rect 8020 9416 8054 9418
rect 8088 9416 8122 9418
rect 8156 9416 8190 9418
rect 8224 9416 8258 9418
rect 8292 9416 8326 9418
rect 8360 9416 8394 9418
rect 8428 9418 8431 9450
rect 8496 9418 8503 9450
rect 8564 9418 8575 9450
rect 8632 9418 8647 9450
rect 8700 9418 8719 9450
rect 8768 9418 8791 9450
rect 8836 9418 8863 9450
rect 8904 9418 8935 9450
rect 8428 9416 8462 9418
rect 8496 9416 8530 9418
rect 8564 9416 8598 9418
rect 8632 9416 8666 9418
rect 8700 9416 8734 9418
rect 8768 9416 8802 9418
rect 8836 9416 8870 9418
rect 8904 9416 8938 9418
rect 8972 9416 9006 9450
rect 9041 9418 9074 9450
rect 9113 9418 9142 9450
rect 9185 9418 9210 9450
rect 9257 9418 9278 9450
rect 9329 9418 9346 9450
rect 9401 9418 9414 9450
rect 9473 9418 9482 9450
rect 9545 9418 9550 9450
rect 9617 9418 9618 9450
rect 9040 9416 9074 9418
rect 9108 9416 9142 9418
rect 9176 9416 9210 9418
rect 9244 9416 9278 9418
rect 9312 9416 9346 9418
rect 9380 9416 9414 9418
rect 9448 9416 9482 9418
rect 9516 9416 9550 9418
rect 9584 9416 9618 9418
rect 9652 9418 9655 9450
rect 9720 9418 9727 9450
rect 9788 9418 9799 9450
rect 9856 9418 9871 9450
rect 9924 9418 9943 9450
rect 9992 9418 10015 9450
rect 10060 9418 10087 9450
rect 10128 9418 10159 9450
rect 9652 9416 9686 9418
rect 9720 9416 9754 9418
rect 9788 9416 9822 9418
rect 9856 9416 9890 9418
rect 9924 9416 9958 9418
rect 9992 9416 10026 9418
rect 10060 9416 10094 9418
rect 10128 9416 10162 9418
rect 10196 9416 10230 9450
rect 10265 9418 10298 9450
rect 10337 9418 10366 9450
rect 10409 9418 10434 9450
rect 10481 9418 10502 9450
rect 10553 9418 10570 9450
rect 10625 9418 10638 9450
rect 10697 9418 10706 9450
rect 10769 9418 10774 9450
rect 10841 9418 10842 9450
rect 10264 9416 10298 9418
rect 10332 9416 10366 9418
rect 10400 9416 10434 9418
rect 10468 9416 10502 9418
rect 10536 9416 10570 9418
rect 10604 9416 10638 9418
rect 10672 9416 10706 9418
rect 10740 9416 10774 9418
rect 10808 9416 10842 9418
rect 10876 9418 10879 9450
rect 10944 9418 10951 9450
rect 11012 9418 11023 9450
rect 11080 9418 11095 9450
rect 11148 9418 11167 9450
rect 11216 9418 11239 9450
rect 11284 9418 11311 9450
rect 11352 9418 11383 9450
rect 10876 9416 10910 9418
rect 10944 9416 10978 9418
rect 11012 9416 11046 9418
rect 11080 9416 11114 9418
rect 11148 9416 11182 9418
rect 11216 9416 11250 9418
rect 11284 9416 11318 9418
rect 11352 9416 11386 9418
rect 11420 9416 11454 9450
rect 11489 9418 11522 9450
rect 11561 9418 11590 9450
rect 11633 9418 11658 9450
rect 11705 9418 11726 9450
rect 11777 9418 11794 9450
rect 11849 9418 11862 9450
rect 11921 9418 11930 9450
rect 11993 9418 11998 9450
rect 12065 9418 12066 9450
rect 11488 9416 11522 9418
rect 11556 9416 11590 9418
rect 11624 9416 11658 9418
rect 11692 9416 11726 9418
rect 11760 9416 11794 9418
rect 11828 9416 11862 9418
rect 11896 9416 11930 9418
rect 11964 9416 11998 9418
rect 12032 9416 12066 9418
rect 12100 9418 12103 9450
rect 12168 9418 12175 9450
rect 12236 9418 12247 9450
rect 12304 9418 12319 9450
rect 12372 9418 12391 9450
rect 12440 9418 12463 9450
rect 12508 9418 12535 9450
rect 12576 9418 12607 9450
rect 12100 9416 12134 9418
rect 12168 9416 12202 9418
rect 12236 9416 12270 9418
rect 12304 9416 12338 9418
rect 12372 9416 12406 9418
rect 12440 9416 12474 9418
rect 12508 9416 12542 9418
rect 12576 9416 12610 9418
rect 12644 9416 12678 9450
rect 12712 9416 12746 9450
rect 12780 9416 12814 9450
rect 12848 9416 12882 9450
rect 12916 9416 12950 9450
rect 12984 9416 13018 9450
rect 13052 9416 13086 9450
rect 13120 9416 13154 9450
rect 13188 9416 13222 9450
rect 13256 9416 13290 9450
rect 13324 9416 13358 9450
rect 13392 9416 13426 9450
rect 13460 9416 13494 9450
rect 13528 9416 13562 9450
rect 13596 9416 13630 9450
rect 13664 9416 13698 9450
rect 13732 9416 13766 9450
rect 13800 9416 13834 9450
rect 13868 9416 13902 9450
rect 13936 9416 13970 9450
rect 14004 9416 14038 9450
rect 14072 9416 14106 9450
rect 14140 9416 14174 9450
rect 14208 9416 14242 9450
rect 14276 9416 14310 9450
rect 14348 9418 14378 9450
rect 14344 9416 14378 9418
rect 14412 9416 14446 9450
rect 14480 9418 14614 9450
rect 14648 9418 14724 9452
rect 14480 9416 14724 9418
rect 245 9343 14724 9416
<< viali >>
rect 320 36500 354 36534
rect 14614 36499 14648 36533
rect 556 36464 566 36498
rect 566 36464 590 36498
rect 628 36464 634 36498
rect 634 36464 662 36498
rect 700 36464 702 36498
rect 702 36464 734 36498
rect 772 36464 804 36498
rect 804 36464 806 36498
rect 844 36464 872 36498
rect 872 36464 878 36498
rect 916 36464 940 36498
rect 940 36464 950 36498
rect 988 36464 1008 36498
rect 1008 36464 1022 36498
rect 1060 36464 1076 36498
rect 1076 36464 1094 36498
rect 1132 36464 1144 36498
rect 1144 36464 1166 36498
rect 1204 36464 1212 36498
rect 1212 36464 1238 36498
rect 1276 36464 1280 36498
rect 1280 36464 1310 36498
rect 1348 36464 1382 36498
rect 1420 36464 1450 36498
rect 1450 36464 1454 36498
rect 1492 36464 1518 36498
rect 1518 36464 1526 36498
rect 1564 36464 1586 36498
rect 1586 36464 1598 36498
rect 1636 36464 1654 36498
rect 1654 36464 1670 36498
rect 1708 36464 1722 36498
rect 1722 36464 1742 36498
rect 1780 36464 1790 36498
rect 1790 36464 1814 36498
rect 1852 36464 1858 36498
rect 1858 36464 1886 36498
rect 1924 36464 1926 36498
rect 1926 36464 1958 36498
rect 1996 36464 2028 36498
rect 2028 36464 2030 36498
rect 2068 36464 2096 36498
rect 2096 36464 2102 36498
rect 2140 36464 2164 36498
rect 2164 36464 2174 36498
rect 2212 36464 2232 36498
rect 2232 36464 2246 36498
rect 2284 36464 2300 36498
rect 2300 36464 2318 36498
rect 2356 36464 2368 36498
rect 2368 36464 2390 36498
rect 2428 36464 2436 36498
rect 2436 36464 2462 36498
rect 2500 36464 2504 36498
rect 2504 36464 2534 36498
rect 2572 36464 2606 36498
rect 2644 36464 2674 36498
rect 2674 36464 2678 36498
rect 2716 36464 2742 36498
rect 2742 36464 2750 36498
rect 2788 36464 2810 36498
rect 2810 36464 2822 36498
rect 2860 36464 2878 36498
rect 2878 36464 2894 36498
rect 2932 36464 2946 36498
rect 2946 36464 2966 36498
rect 3004 36464 3014 36498
rect 3014 36464 3038 36498
rect 3076 36464 3082 36498
rect 3082 36464 3110 36498
rect 3148 36464 3150 36498
rect 3150 36464 3182 36498
rect 3220 36464 3252 36498
rect 3252 36464 3254 36498
rect 3292 36464 3320 36498
rect 3320 36464 3326 36498
rect 3364 36464 3388 36498
rect 3388 36464 3398 36498
rect 3436 36464 3456 36498
rect 3456 36464 3470 36498
rect 3508 36464 3524 36498
rect 3524 36464 3542 36498
rect 3580 36464 3592 36498
rect 3592 36464 3614 36498
rect 3652 36464 3660 36498
rect 3660 36464 3686 36498
rect 3724 36464 3728 36498
rect 3728 36464 3758 36498
rect 3796 36464 3830 36498
rect 3868 36464 3898 36498
rect 3898 36464 3902 36498
rect 3940 36464 3966 36498
rect 3966 36464 3974 36498
rect 4012 36464 4034 36498
rect 4034 36464 4046 36498
rect 4084 36464 4102 36498
rect 4102 36464 4118 36498
rect 4156 36464 4170 36498
rect 4170 36464 4190 36498
rect 4228 36464 4238 36498
rect 4238 36464 4262 36498
rect 4300 36464 4306 36498
rect 4306 36464 4334 36498
rect 4372 36464 4374 36498
rect 4374 36464 4406 36498
rect 4444 36464 4476 36498
rect 4476 36464 4478 36498
rect 4516 36464 4544 36498
rect 4544 36464 4550 36498
rect 4588 36464 4612 36498
rect 4612 36464 4622 36498
rect 4660 36464 4680 36498
rect 4680 36464 4694 36498
rect 4732 36464 4748 36498
rect 4748 36464 4766 36498
rect 4804 36464 4816 36498
rect 4816 36464 4838 36498
rect 4876 36464 4884 36498
rect 4884 36464 4910 36498
rect 4948 36464 4952 36498
rect 4952 36464 4982 36498
rect 5020 36464 5054 36498
rect 5092 36464 5122 36498
rect 5122 36464 5126 36498
rect 5164 36464 5190 36498
rect 5190 36464 5198 36498
rect 5236 36464 5258 36498
rect 5258 36464 5270 36498
rect 5308 36464 5326 36498
rect 5326 36464 5342 36498
rect 5380 36464 5394 36498
rect 5394 36464 5414 36498
rect 5452 36464 5462 36498
rect 5462 36464 5486 36498
rect 5524 36464 5530 36498
rect 5530 36464 5558 36498
rect 5596 36464 5598 36498
rect 5598 36464 5630 36498
rect 5668 36464 5700 36498
rect 5700 36464 5702 36498
rect 5740 36464 5768 36498
rect 5768 36464 5774 36498
rect 5812 36464 5836 36498
rect 5836 36464 5846 36498
rect 5884 36464 5904 36498
rect 5904 36464 5918 36498
rect 5956 36464 5972 36498
rect 5972 36464 5990 36498
rect 6028 36464 6040 36498
rect 6040 36464 6062 36498
rect 6100 36464 6108 36498
rect 6108 36464 6134 36498
rect 6172 36464 6176 36498
rect 6176 36464 6206 36498
rect 6244 36464 6278 36498
rect 6316 36464 6346 36498
rect 6346 36464 6350 36498
rect 6388 36464 6414 36498
rect 6414 36464 6422 36498
rect 6460 36464 6482 36498
rect 6482 36464 6494 36498
rect 6532 36464 6550 36498
rect 6550 36464 6566 36498
rect 6604 36464 6618 36498
rect 6618 36464 6638 36498
rect 6676 36464 6686 36498
rect 6686 36464 6710 36498
rect 6748 36464 6754 36498
rect 6754 36464 6782 36498
rect 6820 36464 6822 36498
rect 6822 36464 6854 36498
rect 6892 36464 6924 36498
rect 6924 36464 6926 36498
rect 6964 36464 6992 36498
rect 6992 36464 6998 36498
rect 7036 36464 7060 36498
rect 7060 36464 7070 36498
rect 7108 36464 7128 36498
rect 7128 36464 7142 36498
rect 7180 36464 7196 36498
rect 7196 36464 7214 36498
rect 7252 36464 7264 36498
rect 7264 36464 7286 36498
rect 7324 36464 7332 36498
rect 7332 36464 7358 36498
rect 7396 36464 7400 36498
rect 7400 36464 7430 36498
rect 7468 36464 7502 36498
rect 7540 36464 7570 36498
rect 7570 36464 7574 36498
rect 7612 36464 7638 36498
rect 7638 36464 7646 36498
rect 7684 36464 7706 36498
rect 7706 36464 7718 36498
rect 7756 36464 7774 36498
rect 7774 36464 7790 36498
rect 7828 36464 7842 36498
rect 7842 36464 7862 36498
rect 7900 36464 7910 36498
rect 7910 36464 7934 36498
rect 7972 36464 7978 36498
rect 7978 36464 8006 36498
rect 8044 36464 8046 36498
rect 8046 36464 8078 36498
rect 8116 36464 8148 36498
rect 8148 36464 8150 36498
rect 8188 36464 8216 36498
rect 8216 36464 8222 36498
rect 8260 36464 8284 36498
rect 8284 36464 8294 36498
rect 8332 36464 8352 36498
rect 8352 36464 8366 36498
rect 8404 36464 8420 36498
rect 8420 36464 8438 36498
rect 8476 36464 8488 36498
rect 8488 36464 8510 36498
rect 8548 36464 8556 36498
rect 8556 36464 8582 36498
rect 8620 36464 8624 36498
rect 8624 36464 8654 36498
rect 8692 36464 8726 36498
rect 8764 36464 8794 36498
rect 8794 36464 8798 36498
rect 8836 36464 8862 36498
rect 8862 36464 8870 36498
rect 8908 36464 8930 36498
rect 8930 36464 8942 36498
rect 8980 36464 8998 36498
rect 8998 36464 9014 36498
rect 9052 36464 9066 36498
rect 9066 36464 9086 36498
rect 9124 36464 9134 36498
rect 9134 36464 9158 36498
rect 9196 36464 9202 36498
rect 9202 36464 9230 36498
rect 9268 36464 9270 36498
rect 9270 36464 9302 36498
rect 9340 36464 9372 36498
rect 9372 36464 9374 36498
rect 9412 36464 9440 36498
rect 9440 36464 9446 36498
rect 9484 36464 9508 36498
rect 9508 36464 9518 36498
rect 9556 36464 9576 36498
rect 9576 36464 9590 36498
rect 9628 36464 9644 36498
rect 9644 36464 9662 36498
rect 9700 36464 9712 36498
rect 9712 36464 9734 36498
rect 9772 36464 9780 36498
rect 9780 36464 9806 36498
rect 9844 36464 9848 36498
rect 9848 36464 9878 36498
rect 9916 36464 9950 36498
rect 9988 36464 10018 36498
rect 10018 36464 10022 36498
rect 10060 36464 10086 36498
rect 10086 36464 10094 36498
rect 10132 36464 10154 36498
rect 10154 36464 10166 36498
rect 10204 36464 10222 36498
rect 10222 36464 10238 36498
rect 10276 36464 10290 36498
rect 10290 36464 10310 36498
rect 10348 36464 10358 36498
rect 10358 36464 10382 36498
rect 10420 36464 10426 36498
rect 10426 36464 10454 36498
rect 10492 36464 10494 36498
rect 10494 36464 10526 36498
rect 10564 36464 10596 36498
rect 10596 36464 10598 36498
rect 10636 36464 10664 36498
rect 10664 36464 10670 36498
rect 10708 36464 10732 36498
rect 10732 36464 10742 36498
rect 10780 36464 10800 36498
rect 10800 36464 10814 36498
rect 10852 36464 10868 36498
rect 10868 36464 10886 36498
rect 10924 36464 10936 36498
rect 10936 36464 10958 36498
rect 10996 36464 11004 36498
rect 11004 36464 11030 36498
rect 11068 36464 11072 36498
rect 11072 36464 11102 36498
rect 11140 36464 11174 36498
rect 11212 36464 11242 36498
rect 11242 36464 11246 36498
rect 11284 36464 11310 36498
rect 11310 36464 11318 36498
rect 11356 36464 11378 36498
rect 11378 36464 11390 36498
rect 11428 36464 11446 36498
rect 11446 36464 11462 36498
rect 11500 36464 11514 36498
rect 11514 36464 11534 36498
rect 11572 36464 11582 36498
rect 11582 36464 11606 36498
rect 11644 36464 11650 36498
rect 11650 36464 11678 36498
rect 11716 36464 11718 36498
rect 11718 36464 11750 36498
rect 11788 36464 11820 36498
rect 11820 36464 11822 36498
rect 11860 36464 11888 36498
rect 11888 36464 11894 36498
rect 11932 36464 11956 36498
rect 11956 36464 11966 36498
rect 12004 36464 12024 36498
rect 12024 36464 12038 36498
rect 12076 36464 12092 36498
rect 12092 36464 12110 36498
rect 12148 36464 12160 36498
rect 12160 36464 12182 36498
rect 12220 36464 12228 36498
rect 12228 36464 12254 36498
rect 12292 36464 12296 36498
rect 12296 36464 12326 36498
rect 12364 36464 12398 36498
rect 12436 36464 12466 36498
rect 12466 36464 12470 36498
rect 12508 36464 12534 36498
rect 12534 36464 12542 36498
rect 12580 36464 12602 36498
rect 12602 36464 12614 36498
rect 12652 36464 12670 36498
rect 12670 36464 12686 36498
rect 12724 36464 12738 36498
rect 12738 36464 12758 36498
rect 12796 36464 12806 36498
rect 12806 36464 12830 36498
rect 12868 36464 12874 36498
rect 12874 36464 12902 36498
rect 12940 36464 12942 36498
rect 12942 36464 12974 36498
rect 13012 36464 13044 36498
rect 13044 36464 13046 36498
rect 13084 36464 13112 36498
rect 13112 36464 13118 36498
rect 13156 36464 13180 36498
rect 13180 36464 13190 36498
rect 13228 36464 13248 36498
rect 13248 36464 13262 36498
rect 13300 36464 13316 36498
rect 13316 36464 13334 36498
rect 13372 36464 13384 36498
rect 13384 36464 13406 36498
rect 13444 36464 13452 36498
rect 13452 36464 13478 36498
rect 13516 36464 13520 36498
rect 13520 36464 13550 36498
rect 13588 36464 13622 36498
rect 13660 36464 13690 36498
rect 13690 36464 13694 36498
rect 13732 36464 13758 36498
rect 13758 36464 13766 36498
rect 13804 36464 13826 36498
rect 13826 36464 13838 36498
rect 13876 36464 13894 36498
rect 13894 36464 13910 36498
rect 13948 36464 13962 36498
rect 13962 36464 13982 36498
rect 14020 36464 14030 36498
rect 14030 36464 14054 36498
rect 14092 36464 14098 36498
rect 14098 36464 14126 36498
rect 14164 36464 14166 36498
rect 14166 36464 14198 36498
rect 14236 36464 14268 36498
rect 14268 36464 14270 36498
rect 14308 36464 14336 36498
rect 14336 36464 14342 36498
rect 14380 36464 14404 36498
rect 14404 36464 14414 36498
rect 320 36428 354 36462
rect 14614 36427 14648 36461
rect 320 36243 354 36265
rect 320 36231 351 36243
rect 351 36231 354 36243
rect 14614 36241 14648 36262
rect 14614 36228 14645 36241
rect 14645 36228 14648 36241
rect 320 36175 354 36193
rect 320 36159 351 36175
rect 351 36159 354 36175
rect 320 36107 354 36121
rect 320 36087 351 36107
rect 351 36087 354 36107
rect 320 36039 354 36049
rect 320 36015 351 36039
rect 351 36015 354 36039
rect 320 35971 354 35977
rect 320 35943 351 35971
rect 351 35943 354 35971
rect 320 35903 354 35905
rect 320 35871 351 35903
rect 351 35871 354 35903
rect 320 35801 351 35833
rect 351 35801 354 35833
rect 320 35799 354 35801
rect 320 35733 351 35761
rect 351 35733 354 35761
rect 320 35727 354 35733
rect 320 35665 351 35689
rect 351 35665 354 35689
rect 320 35655 354 35665
rect 320 35597 351 35617
rect 351 35597 354 35617
rect 320 35583 354 35597
rect 320 35529 351 35545
rect 351 35529 354 35545
rect 320 35511 354 35529
rect 320 35461 351 35473
rect 351 35461 354 35473
rect 320 35439 354 35461
rect 320 35393 351 35401
rect 351 35393 354 35401
rect 320 35367 354 35393
rect 320 35325 351 35329
rect 351 35325 354 35329
rect 320 35295 354 35325
rect 320 35223 354 35257
rect 320 35155 354 35185
rect 320 35151 351 35155
rect 351 35151 354 35155
rect 320 35087 354 35113
rect 320 35079 351 35087
rect 351 35079 354 35087
rect 320 35019 354 35041
rect 320 35007 351 35019
rect 351 35007 354 35019
rect 320 34951 354 34969
rect 320 34935 351 34951
rect 351 34935 354 34951
rect 320 34883 354 34897
rect 320 34863 351 34883
rect 351 34863 354 34883
rect 320 34815 354 34825
rect 320 34791 351 34815
rect 351 34791 354 34815
rect 320 34747 354 34753
rect 320 34719 351 34747
rect 351 34719 354 34747
rect 320 34679 354 34681
rect 320 34647 351 34679
rect 351 34647 354 34679
rect 320 34577 351 34609
rect 351 34577 354 34609
rect 320 34575 354 34577
rect 320 34509 351 34537
rect 351 34509 354 34537
rect 320 34503 354 34509
rect 320 34441 351 34465
rect 351 34441 354 34465
rect 320 34431 354 34441
rect 320 34373 351 34393
rect 351 34373 354 34393
rect 320 34359 354 34373
rect 320 34305 351 34321
rect 351 34305 354 34321
rect 320 34287 354 34305
rect 320 34237 351 34249
rect 351 34237 354 34249
rect 320 34215 354 34237
rect 320 34169 351 34177
rect 351 34169 354 34177
rect 320 34143 354 34169
rect 320 34101 351 34105
rect 351 34101 354 34105
rect 320 34071 354 34101
rect 320 33999 354 34033
rect 320 33931 354 33961
rect 320 33927 351 33931
rect 351 33927 354 33931
rect 320 33863 354 33889
rect 320 33855 351 33863
rect 351 33855 354 33863
rect 320 33795 354 33817
rect 320 33783 351 33795
rect 351 33783 354 33795
rect 320 33727 354 33745
rect 320 33711 351 33727
rect 351 33711 354 33727
rect 320 33659 354 33673
rect 320 33639 351 33659
rect 351 33639 354 33659
rect 320 33591 354 33601
rect 320 33567 351 33591
rect 351 33567 354 33591
rect 320 33523 354 33529
rect 320 33495 351 33523
rect 351 33495 354 33523
rect 320 33455 354 33457
rect 320 33423 351 33455
rect 351 33423 354 33455
rect 320 33353 351 33385
rect 351 33353 354 33385
rect 320 33351 354 33353
rect 320 33285 351 33313
rect 351 33285 354 33313
rect 320 33279 354 33285
rect 320 33217 351 33241
rect 351 33217 354 33241
rect 320 33207 354 33217
rect 320 33149 351 33169
rect 351 33149 354 33169
rect 320 33135 354 33149
rect 320 33081 351 33097
rect 351 33081 354 33097
rect 320 33063 354 33081
rect 320 33013 351 33025
rect 351 33013 354 33025
rect 320 32991 354 33013
rect 320 32945 351 32953
rect 351 32945 354 32953
rect 320 32919 354 32945
rect 320 32877 351 32881
rect 351 32877 354 32881
rect 320 32847 354 32877
rect 320 32775 354 32809
rect 320 32707 354 32737
rect 320 32703 351 32707
rect 351 32703 354 32707
rect 320 32639 354 32665
rect 320 32631 351 32639
rect 351 32631 354 32639
rect 320 32571 354 32593
rect 320 32559 351 32571
rect 351 32559 354 32571
rect 320 32503 354 32521
rect 320 32487 351 32503
rect 351 32487 354 32503
rect 320 32435 354 32449
rect 320 32415 351 32435
rect 351 32415 354 32435
rect 320 32367 354 32377
rect 320 32343 351 32367
rect 351 32343 354 32367
rect 320 32299 354 32305
rect 320 32271 351 32299
rect 351 32271 354 32299
rect 320 32231 354 32233
rect 320 32199 351 32231
rect 351 32199 354 32231
rect 320 32129 351 32161
rect 351 32129 354 32161
rect 320 32127 354 32129
rect 320 32061 351 32089
rect 351 32061 354 32089
rect 320 32055 354 32061
rect 320 31993 351 32017
rect 351 31993 354 32017
rect 320 31983 354 31993
rect 320 31925 351 31945
rect 351 31925 354 31945
rect 320 31911 354 31925
rect 320 31857 351 31873
rect 351 31857 354 31873
rect 320 31839 354 31857
rect 320 31789 351 31801
rect 351 31789 354 31801
rect 320 31767 354 31789
rect 320 31721 351 31729
rect 351 31721 354 31729
rect 320 31695 354 31721
rect 320 31653 351 31657
rect 351 31653 354 31657
rect 320 31623 354 31653
rect 320 31551 354 31585
rect 320 31483 354 31513
rect 320 31479 351 31483
rect 351 31479 354 31483
rect 320 31415 354 31441
rect 320 31407 351 31415
rect 351 31407 354 31415
rect 320 31347 354 31369
rect 320 31335 351 31347
rect 351 31335 354 31347
rect 320 31279 354 31297
rect 320 31263 351 31279
rect 351 31263 354 31279
rect 320 31211 354 31225
rect 320 31191 351 31211
rect 351 31191 354 31211
rect 320 31143 354 31153
rect 320 31119 351 31143
rect 351 31119 354 31143
rect 320 31075 354 31081
rect 320 31047 351 31075
rect 351 31047 354 31075
rect 320 31007 354 31009
rect 320 30975 351 31007
rect 351 30975 354 31007
rect 320 30905 351 30937
rect 351 30905 354 30937
rect 320 30903 354 30905
rect 320 30837 351 30865
rect 351 30837 354 30865
rect 320 30831 354 30837
rect 320 30769 351 30793
rect 351 30769 354 30793
rect 320 30759 354 30769
rect 320 30701 351 30721
rect 351 30701 354 30721
rect 320 30687 354 30701
rect 320 30633 351 30649
rect 351 30633 354 30649
rect 320 30615 354 30633
rect 320 30565 351 30577
rect 351 30565 354 30577
rect 320 30543 354 30565
rect 320 30497 351 30505
rect 351 30497 354 30505
rect 320 30471 354 30497
rect 320 30429 351 30433
rect 351 30429 354 30433
rect 320 30399 354 30429
rect 320 30327 354 30361
rect 320 30259 354 30289
rect 320 30255 351 30259
rect 351 30255 354 30259
rect 320 30191 354 30217
rect 320 30183 351 30191
rect 351 30183 354 30191
rect 320 30123 354 30145
rect 320 30111 351 30123
rect 351 30111 354 30123
rect 320 30055 354 30073
rect 320 30039 351 30055
rect 351 30039 354 30055
rect 320 29987 354 30001
rect 320 29967 351 29987
rect 351 29967 354 29987
rect 320 29919 354 29929
rect 320 29895 351 29919
rect 351 29895 354 29919
rect 320 29851 354 29857
rect 320 29823 351 29851
rect 351 29823 354 29851
rect 320 29783 354 29785
rect 320 29751 351 29783
rect 351 29751 354 29783
rect 320 29681 351 29713
rect 351 29681 354 29713
rect 320 29679 354 29681
rect 320 29613 351 29641
rect 351 29613 354 29641
rect 320 29607 354 29613
rect 320 29545 351 29569
rect 351 29545 354 29569
rect 320 29535 354 29545
rect 320 29477 351 29497
rect 351 29477 354 29497
rect 320 29463 354 29477
rect 320 29409 351 29425
rect 351 29409 354 29425
rect 320 29391 354 29409
rect 320 29341 351 29353
rect 351 29341 354 29353
rect 320 29319 354 29341
rect 320 29273 351 29281
rect 351 29273 354 29281
rect 320 29247 354 29273
rect 320 29205 351 29209
rect 351 29205 354 29209
rect 320 29175 354 29205
rect 320 29103 354 29137
rect 320 29035 354 29065
rect 320 29031 351 29035
rect 351 29031 354 29035
rect 320 28967 354 28993
rect 320 28959 351 28967
rect 351 28959 354 28967
rect 320 28899 354 28921
rect 320 28887 351 28899
rect 351 28887 354 28899
rect 320 28831 354 28849
rect 320 28815 351 28831
rect 351 28815 354 28831
rect 320 28763 354 28777
rect 320 28743 351 28763
rect 351 28743 354 28763
rect 320 28695 354 28705
rect 320 28671 351 28695
rect 351 28671 354 28695
rect 320 28627 354 28633
rect 320 28599 351 28627
rect 351 28599 354 28627
rect 320 28559 354 28561
rect 320 28527 351 28559
rect 351 28527 354 28559
rect 320 28457 351 28489
rect 351 28457 354 28489
rect 320 28455 354 28457
rect 320 28389 351 28417
rect 351 28389 354 28417
rect 320 28383 354 28389
rect 320 28321 351 28345
rect 351 28321 354 28345
rect 320 28311 354 28321
rect 320 28253 351 28273
rect 351 28253 354 28273
rect 320 28239 354 28253
rect 320 28185 351 28201
rect 351 28185 354 28201
rect 320 28167 354 28185
rect 320 28117 351 28129
rect 351 28117 354 28129
rect 320 28095 354 28117
rect 320 28049 351 28057
rect 351 28049 354 28057
rect 320 28023 354 28049
rect 320 27981 351 27985
rect 351 27981 354 27985
rect 320 27951 354 27981
rect 320 27879 354 27913
rect 320 27811 354 27841
rect 320 27807 351 27811
rect 351 27807 354 27811
rect 320 27743 354 27769
rect 320 27735 351 27743
rect 351 27735 354 27743
rect 320 27675 354 27697
rect 320 27663 351 27675
rect 351 27663 354 27675
rect 320 27607 354 27625
rect 320 27591 351 27607
rect 351 27591 354 27607
rect 320 27539 354 27553
rect 320 27519 351 27539
rect 351 27519 354 27539
rect 320 27471 354 27481
rect 320 27447 351 27471
rect 351 27447 354 27471
rect 320 27403 354 27409
rect 320 27375 351 27403
rect 351 27375 354 27403
rect 320 27335 354 27337
rect 320 27303 351 27335
rect 351 27303 354 27335
rect 320 27233 351 27265
rect 351 27233 354 27265
rect 320 27231 354 27233
rect 320 27165 351 27193
rect 351 27165 354 27193
rect 320 27159 354 27165
rect 320 27097 351 27121
rect 351 27097 354 27121
rect 320 27087 354 27097
rect 320 27029 351 27049
rect 351 27029 354 27049
rect 320 27015 354 27029
rect 320 26961 351 26977
rect 351 26961 354 26977
rect 320 26943 354 26961
rect 320 26893 351 26905
rect 351 26893 354 26905
rect 320 26871 354 26893
rect 320 26825 351 26833
rect 351 26825 354 26833
rect 320 26799 354 26825
rect 320 26757 351 26761
rect 351 26757 354 26761
rect 320 26727 354 26757
rect 320 26655 354 26689
rect 320 26587 354 26617
rect 320 26583 351 26587
rect 351 26583 354 26587
rect 320 26519 354 26545
rect 320 26511 351 26519
rect 351 26511 354 26519
rect 320 26451 354 26473
rect 320 26439 351 26451
rect 351 26439 354 26451
rect 320 26383 354 26401
rect 320 26367 351 26383
rect 351 26367 354 26383
rect 320 26315 354 26329
rect 320 26295 351 26315
rect 351 26295 354 26315
rect 320 26247 354 26257
rect 320 26223 351 26247
rect 351 26223 354 26247
rect 320 26179 354 26185
rect 320 26151 351 26179
rect 351 26151 354 26179
rect 320 26111 354 26113
rect 320 26079 351 26111
rect 351 26079 354 26111
rect 320 26009 351 26041
rect 351 26009 354 26041
rect 320 26007 354 26009
rect 320 25941 351 25969
rect 351 25941 354 25969
rect 320 25935 354 25941
rect 320 25873 351 25897
rect 351 25873 354 25897
rect 320 25863 354 25873
rect 320 25805 351 25825
rect 351 25805 354 25825
rect 320 25791 354 25805
rect 320 25737 351 25753
rect 351 25737 354 25753
rect 320 25719 354 25737
rect 320 25669 351 25681
rect 351 25669 354 25681
rect 320 25647 354 25669
rect 320 25601 351 25609
rect 351 25601 354 25609
rect 320 25575 354 25601
rect 320 25533 351 25537
rect 351 25533 354 25537
rect 320 25503 354 25533
rect 320 25431 354 25465
rect 320 25363 354 25393
rect 320 25359 351 25363
rect 351 25359 354 25363
rect 320 25295 354 25321
rect 320 25287 351 25295
rect 351 25287 354 25295
rect 320 25227 354 25249
rect 320 25215 351 25227
rect 351 25215 354 25227
rect 320 25159 354 25177
rect 320 25143 351 25159
rect 351 25143 354 25159
rect 320 25091 354 25105
rect 320 25071 351 25091
rect 351 25071 354 25091
rect 320 25023 354 25033
rect 320 24999 351 25023
rect 351 24999 354 25023
rect 320 24955 354 24961
rect 320 24927 351 24955
rect 351 24927 354 24955
rect 320 24887 354 24889
rect 320 24855 351 24887
rect 351 24855 354 24887
rect 320 24785 351 24817
rect 351 24785 354 24817
rect 320 24783 354 24785
rect 320 24717 351 24745
rect 351 24717 354 24745
rect 320 24711 354 24717
rect 320 24649 351 24673
rect 351 24649 354 24673
rect 320 24639 354 24649
rect 320 24581 351 24601
rect 351 24581 354 24601
rect 320 24567 354 24581
rect 320 24513 351 24529
rect 351 24513 354 24529
rect 320 24495 354 24513
rect 320 24445 351 24457
rect 351 24445 354 24457
rect 320 24423 354 24445
rect 320 24377 351 24385
rect 351 24377 354 24385
rect 320 24351 354 24377
rect 320 24309 351 24313
rect 351 24309 354 24313
rect 320 24279 354 24309
rect 320 24207 354 24241
rect 320 24139 354 24169
rect 320 24135 351 24139
rect 351 24135 354 24139
rect 320 24071 354 24097
rect 320 24063 351 24071
rect 351 24063 354 24071
rect 320 24003 354 24025
rect 320 23991 351 24003
rect 351 23991 354 24003
rect 320 23935 354 23953
rect 320 23919 351 23935
rect 351 23919 354 23935
rect 320 23867 354 23881
rect 320 23847 351 23867
rect 351 23847 354 23867
rect 320 23799 354 23809
rect 320 23775 351 23799
rect 351 23775 354 23799
rect 320 23731 354 23737
rect 320 23703 351 23731
rect 351 23703 354 23731
rect 320 23663 354 23665
rect 320 23631 351 23663
rect 351 23631 354 23663
rect 320 23561 351 23593
rect 351 23561 354 23593
rect 320 23559 354 23561
rect 320 23493 351 23521
rect 351 23493 354 23521
rect 320 23487 354 23493
rect 320 23425 351 23449
rect 351 23425 354 23449
rect 320 23415 354 23425
rect 320 23357 351 23377
rect 351 23357 354 23377
rect 320 23343 354 23357
rect 320 23289 351 23305
rect 351 23289 354 23305
rect 320 23271 354 23289
rect 320 23221 351 23233
rect 351 23221 354 23233
rect 320 23199 354 23221
rect 320 23153 351 23161
rect 351 23153 354 23161
rect 320 23127 354 23153
rect 320 23085 351 23089
rect 351 23085 354 23089
rect 320 23055 354 23085
rect 320 22983 354 23017
rect 320 22915 354 22945
rect 320 22911 351 22915
rect 351 22911 354 22915
rect 320 22847 354 22873
rect 320 22839 351 22847
rect 351 22839 354 22847
rect 320 22779 354 22801
rect 320 22767 351 22779
rect 351 22767 354 22779
rect 320 22711 354 22729
rect 320 22695 351 22711
rect 351 22695 354 22711
rect 320 22643 354 22657
rect 320 22623 351 22643
rect 351 22623 354 22643
rect 320 22575 354 22585
rect 320 22551 351 22575
rect 351 22551 354 22575
rect 320 22507 354 22513
rect 320 22479 351 22507
rect 351 22479 354 22507
rect 320 22439 354 22441
rect 320 22407 351 22439
rect 351 22407 354 22439
rect 320 22337 351 22369
rect 351 22337 354 22369
rect 320 22335 354 22337
rect 320 22269 351 22297
rect 351 22269 354 22297
rect 320 22263 354 22269
rect 320 22201 351 22225
rect 351 22201 354 22225
rect 320 22191 354 22201
rect 320 22133 351 22153
rect 351 22133 354 22153
rect 320 22119 354 22133
rect 320 22065 351 22081
rect 351 22065 354 22081
rect 320 22047 354 22065
rect 320 21997 351 22009
rect 351 21997 354 22009
rect 320 21975 354 21997
rect 320 21929 351 21937
rect 351 21929 354 21937
rect 320 21903 354 21929
rect 320 21861 351 21865
rect 351 21861 354 21865
rect 320 21831 354 21861
rect 320 21759 354 21793
rect 320 21691 354 21721
rect 320 21687 351 21691
rect 351 21687 354 21691
rect 320 21623 354 21649
rect 320 21615 351 21623
rect 351 21615 354 21623
rect 320 21555 354 21577
rect 320 21543 351 21555
rect 351 21543 354 21555
rect 320 21487 354 21505
rect 320 21471 351 21487
rect 351 21471 354 21487
rect 320 21419 354 21433
rect 320 21399 351 21419
rect 351 21399 354 21419
rect 320 21351 354 21361
rect 320 21327 351 21351
rect 351 21327 354 21351
rect 320 21283 354 21289
rect 320 21255 351 21283
rect 351 21255 354 21283
rect 320 21215 354 21217
rect 320 21183 351 21215
rect 351 21183 354 21215
rect 320 21113 351 21145
rect 351 21113 354 21145
rect 320 21111 354 21113
rect 320 21045 351 21073
rect 351 21045 354 21073
rect 320 21039 354 21045
rect 320 20977 351 21001
rect 351 20977 354 21001
rect 320 20967 354 20977
rect 320 20909 351 20929
rect 351 20909 354 20929
rect 320 20895 354 20909
rect 320 20841 351 20857
rect 351 20841 354 20857
rect 320 20823 354 20841
rect 320 20773 351 20785
rect 351 20773 354 20785
rect 320 20751 354 20773
rect 320 20705 351 20713
rect 351 20705 354 20713
rect 320 20679 354 20705
rect 320 20637 351 20641
rect 351 20637 354 20641
rect 320 20607 354 20637
rect 320 20535 354 20569
rect 320 20467 354 20497
rect 320 20463 351 20467
rect 351 20463 354 20467
rect 320 20399 354 20425
rect 320 20391 351 20399
rect 351 20391 354 20399
rect 320 20331 354 20353
rect 320 20319 351 20331
rect 351 20319 354 20331
rect 320 20263 354 20281
rect 320 20247 351 20263
rect 351 20247 354 20263
rect 320 20195 354 20209
rect 320 20175 351 20195
rect 351 20175 354 20195
rect 320 20127 354 20137
rect 320 20103 351 20127
rect 351 20103 354 20127
rect 320 20059 354 20065
rect 320 20031 351 20059
rect 351 20031 354 20059
rect 320 19991 354 19993
rect 320 19959 351 19991
rect 351 19959 354 19991
rect 320 19889 351 19921
rect 351 19889 354 19921
rect 320 19887 354 19889
rect 320 19821 351 19849
rect 351 19821 354 19849
rect 320 19815 354 19821
rect 320 19753 351 19777
rect 351 19753 354 19777
rect 320 19743 354 19753
rect 320 19685 351 19705
rect 351 19685 354 19705
rect 320 19671 354 19685
rect 320 19617 351 19633
rect 351 19617 354 19633
rect 320 19599 354 19617
rect 320 19549 351 19561
rect 351 19549 354 19561
rect 320 19527 354 19549
rect 320 19481 351 19489
rect 351 19481 354 19489
rect 320 19455 354 19481
rect 320 19413 351 19417
rect 351 19413 354 19417
rect 320 19383 354 19413
rect 320 19311 354 19345
rect 320 19243 354 19273
rect 320 19239 351 19243
rect 351 19239 354 19243
rect 320 19175 354 19201
rect 320 19167 351 19175
rect 351 19167 354 19175
rect 320 19107 354 19129
rect 320 19095 351 19107
rect 351 19095 354 19107
rect 320 19039 354 19057
rect 320 19023 351 19039
rect 351 19023 354 19039
rect 320 18971 354 18985
rect 320 18951 351 18971
rect 351 18951 354 18971
rect 320 18903 354 18913
rect 320 18879 351 18903
rect 351 18879 354 18903
rect 320 18835 354 18841
rect 320 18807 351 18835
rect 351 18807 354 18835
rect 320 18767 354 18769
rect 320 18735 351 18767
rect 351 18735 354 18767
rect 320 18665 351 18697
rect 351 18665 354 18697
rect 320 18663 354 18665
rect 320 18597 351 18625
rect 351 18597 354 18625
rect 320 18591 354 18597
rect 320 18529 351 18553
rect 351 18529 354 18553
rect 320 18519 354 18529
rect 320 18461 351 18481
rect 351 18461 354 18481
rect 320 18447 354 18461
rect 320 18393 351 18409
rect 351 18393 354 18409
rect 320 18375 354 18393
rect 320 18325 351 18337
rect 351 18325 354 18337
rect 320 18303 354 18325
rect 320 18257 351 18265
rect 351 18257 354 18265
rect 320 18231 354 18257
rect 320 18189 351 18193
rect 351 18189 354 18193
rect 320 18159 354 18189
rect 320 18087 354 18121
rect 320 18019 354 18049
rect 320 18015 351 18019
rect 351 18015 354 18019
rect 320 17951 354 17977
rect 320 17943 351 17951
rect 351 17943 354 17951
rect 320 17883 354 17905
rect 320 17871 351 17883
rect 351 17871 354 17883
rect 320 17815 354 17833
rect 320 17799 351 17815
rect 351 17799 354 17815
rect 320 17747 354 17761
rect 320 17727 351 17747
rect 351 17727 354 17747
rect 320 17679 354 17689
rect 320 17655 351 17679
rect 351 17655 354 17679
rect 320 17611 354 17617
rect 320 17583 351 17611
rect 351 17583 354 17611
rect 320 17543 354 17545
rect 320 17511 351 17543
rect 351 17511 354 17543
rect 320 17441 351 17473
rect 351 17441 354 17473
rect 320 17439 354 17441
rect 320 17373 351 17401
rect 351 17373 354 17401
rect 320 17367 354 17373
rect 320 17305 351 17329
rect 351 17305 354 17329
rect 320 17295 354 17305
rect 320 17237 351 17257
rect 351 17237 354 17257
rect 320 17223 354 17237
rect 320 17169 351 17185
rect 351 17169 354 17185
rect 320 17151 354 17169
rect 320 17101 351 17113
rect 351 17101 354 17113
rect 320 17079 354 17101
rect 320 17033 351 17041
rect 351 17033 354 17041
rect 320 17007 354 17033
rect 320 16965 351 16969
rect 351 16965 354 16969
rect 320 16935 354 16965
rect 320 16863 354 16897
rect 320 16795 354 16825
rect 320 16791 351 16795
rect 351 16791 354 16795
rect 320 16727 354 16753
rect 320 16719 351 16727
rect 351 16719 354 16727
rect 320 16659 354 16681
rect 320 16647 351 16659
rect 351 16647 354 16659
rect 320 16591 354 16609
rect 320 16575 351 16591
rect 351 16575 354 16591
rect 320 16523 354 16537
rect 320 16503 351 16523
rect 351 16503 354 16523
rect 320 16455 354 16465
rect 320 16431 351 16455
rect 351 16431 354 16455
rect 320 16387 354 16393
rect 320 16359 351 16387
rect 351 16359 354 16387
rect 320 16319 354 16321
rect 320 16287 351 16319
rect 351 16287 354 16319
rect 320 16217 351 16249
rect 351 16217 354 16249
rect 320 16215 354 16217
rect 320 16149 351 16177
rect 351 16149 354 16177
rect 320 16143 354 16149
rect 320 16081 351 16105
rect 351 16081 354 16105
rect 320 16071 354 16081
rect 320 16013 351 16033
rect 351 16013 354 16033
rect 320 15999 354 16013
rect 320 15945 351 15961
rect 351 15945 354 15961
rect 320 15927 354 15945
rect 320 15877 351 15889
rect 351 15877 354 15889
rect 320 15855 354 15877
rect 320 15809 351 15817
rect 351 15809 354 15817
rect 320 15783 354 15809
rect 320 15741 351 15745
rect 351 15741 354 15745
rect 320 15711 354 15741
rect 320 15639 354 15673
rect 320 15571 354 15601
rect 320 15567 351 15571
rect 351 15567 354 15571
rect 320 15503 354 15529
rect 320 15495 351 15503
rect 351 15495 354 15503
rect 320 15435 354 15457
rect 320 15423 351 15435
rect 351 15423 354 15435
rect 320 15367 354 15385
rect 320 15351 351 15367
rect 351 15351 354 15367
rect 320 15299 354 15313
rect 320 15279 351 15299
rect 351 15279 354 15299
rect 320 15231 354 15241
rect 320 15207 351 15231
rect 351 15207 354 15231
rect 320 15163 354 15169
rect 320 15135 351 15163
rect 351 15135 354 15163
rect 320 15095 354 15097
rect 320 15063 351 15095
rect 351 15063 354 15095
rect 320 14993 351 15025
rect 351 14993 354 15025
rect 320 14991 354 14993
rect 320 14925 351 14953
rect 351 14925 354 14953
rect 320 14919 354 14925
rect 320 14857 351 14881
rect 351 14857 354 14881
rect 320 14847 354 14857
rect 320 14789 351 14809
rect 351 14789 354 14809
rect 320 14775 354 14789
rect 320 14721 351 14737
rect 351 14721 354 14737
rect 320 14703 354 14721
rect 320 14653 351 14665
rect 351 14653 354 14665
rect 320 14631 354 14653
rect 320 14585 351 14593
rect 351 14585 354 14593
rect 320 14559 354 14585
rect 320 14517 351 14521
rect 351 14517 354 14521
rect 320 14487 354 14517
rect 320 14415 354 14449
rect 320 14347 354 14377
rect 320 14343 351 14347
rect 351 14343 354 14347
rect 320 14279 354 14305
rect 320 14271 351 14279
rect 351 14271 354 14279
rect 320 14211 354 14233
rect 320 14199 351 14211
rect 351 14199 354 14211
rect 320 14143 354 14161
rect 320 14127 351 14143
rect 351 14127 354 14143
rect 320 14075 354 14089
rect 320 14055 351 14075
rect 351 14055 354 14075
rect 320 14007 354 14017
rect 320 13983 351 14007
rect 351 13983 354 14007
rect 320 13939 354 13945
rect 320 13911 351 13939
rect 351 13911 354 13939
rect 320 13871 354 13873
rect 320 13839 351 13871
rect 351 13839 354 13871
rect 320 13769 351 13801
rect 351 13769 354 13801
rect 320 13767 354 13769
rect 320 13701 351 13729
rect 351 13701 354 13729
rect 320 13695 354 13701
rect 320 13633 351 13657
rect 351 13633 354 13657
rect 320 13623 354 13633
rect 320 13565 351 13585
rect 351 13565 354 13585
rect 320 13551 354 13565
rect 320 13497 351 13513
rect 351 13497 354 13513
rect 320 13479 354 13497
rect 320 13429 351 13441
rect 351 13429 354 13441
rect 320 13407 354 13429
rect 320 13361 351 13369
rect 351 13361 354 13369
rect 320 13335 354 13361
rect 320 13293 351 13297
rect 351 13293 354 13297
rect 320 13263 354 13293
rect 320 13191 354 13225
rect 320 13123 354 13153
rect 320 13119 351 13123
rect 351 13119 354 13123
rect 320 13055 354 13081
rect 320 13047 351 13055
rect 351 13047 354 13055
rect 320 12987 354 13009
rect 320 12975 351 12987
rect 351 12975 354 12987
rect 320 12919 354 12937
rect 320 12903 351 12919
rect 351 12903 354 12919
rect 320 12851 354 12865
rect 320 12831 351 12851
rect 351 12831 354 12851
rect 320 12783 354 12793
rect 320 12759 351 12783
rect 351 12759 354 12783
rect 320 12715 354 12721
rect 320 12687 351 12715
rect 351 12687 354 12715
rect 320 12647 354 12649
rect 320 12615 351 12647
rect 351 12615 354 12647
rect 320 12545 351 12577
rect 351 12545 354 12577
rect 320 12543 354 12545
rect 320 12477 351 12505
rect 351 12477 354 12505
rect 320 12471 354 12477
rect 320 12409 351 12433
rect 351 12409 354 12433
rect 320 12399 354 12409
rect 320 12341 351 12361
rect 351 12341 354 12361
rect 320 12327 354 12341
rect 320 12273 351 12289
rect 351 12273 354 12289
rect 320 12255 354 12273
rect 320 12205 351 12217
rect 351 12205 354 12217
rect 320 12183 354 12205
rect 320 12137 351 12145
rect 351 12137 354 12145
rect 320 12111 354 12137
rect 320 12069 351 12073
rect 351 12069 354 12073
rect 320 12039 354 12069
rect 320 11967 354 12001
rect 320 11899 354 11929
rect 320 11895 351 11899
rect 351 11895 354 11899
rect 320 11831 354 11857
rect 320 11823 351 11831
rect 351 11823 354 11831
rect 320 11763 354 11785
rect 320 11751 351 11763
rect 351 11751 354 11763
rect 320 11695 354 11713
rect 320 11679 351 11695
rect 351 11679 354 11695
rect 320 11627 354 11641
rect 320 11607 351 11627
rect 351 11607 354 11627
rect 320 11559 354 11569
rect 320 11535 351 11559
rect 351 11535 354 11559
rect 320 11491 354 11497
rect 320 11463 351 11491
rect 351 11463 354 11491
rect 320 11423 354 11425
rect 320 11391 351 11423
rect 351 11391 354 11423
rect 320 11321 351 11353
rect 351 11321 354 11353
rect 320 11319 354 11321
rect 320 11253 351 11281
rect 351 11253 354 11281
rect 320 11247 354 11253
rect 320 11185 351 11209
rect 351 11185 354 11209
rect 320 11175 354 11185
rect 320 11117 351 11137
rect 351 11117 354 11137
rect 320 11103 354 11117
rect 320 11049 351 11065
rect 351 11049 354 11065
rect 320 11031 354 11049
rect 320 10981 351 10993
rect 351 10981 354 10993
rect 320 10959 354 10981
rect 320 10913 351 10921
rect 351 10913 354 10921
rect 320 10887 354 10913
rect 320 10845 351 10849
rect 351 10845 354 10849
rect 320 10815 354 10845
rect 320 10743 354 10777
rect 320 10675 354 10705
rect 320 10671 351 10675
rect 351 10671 354 10675
rect 320 10607 354 10633
rect 320 10599 351 10607
rect 351 10599 354 10607
rect 320 10539 354 10561
rect 320 10527 351 10539
rect 351 10527 354 10539
rect 320 10471 354 10489
rect 320 10455 351 10471
rect 351 10455 354 10471
rect 320 10403 354 10417
rect 320 10383 351 10403
rect 351 10383 354 10403
rect 320 10335 354 10345
rect 320 10311 351 10335
rect 351 10311 354 10335
rect 320 10267 354 10273
rect 320 10239 351 10267
rect 351 10239 354 10267
rect 320 10199 354 10201
rect 320 10167 351 10199
rect 351 10167 354 10199
rect 320 10097 351 10129
rect 351 10097 354 10129
rect 320 10095 354 10097
rect 320 10029 351 10057
rect 351 10029 354 10057
rect 320 10023 354 10029
rect 320 9961 351 9985
rect 351 9961 354 9985
rect 320 9951 354 9961
rect 320 9893 351 9913
rect 351 9893 354 9913
rect 320 9879 354 9893
rect 320 9825 351 9841
rect 351 9825 354 9841
rect 320 9807 354 9825
rect 320 9757 351 9769
rect 351 9757 354 9769
rect 320 9735 354 9757
rect 1007 35969 1041 36003
rect 1079 35969 1113 36003
rect 1151 35969 1185 36003
rect 1223 35969 1257 36003
rect 1295 35969 1329 36003
rect 1367 35969 1401 36003
rect 1439 35969 1473 36003
rect 1511 35969 1545 36003
rect 1583 35969 1617 36003
rect 1655 35969 1689 36003
rect 1727 35969 1761 36003
rect 1799 35969 1833 36003
rect 1871 35969 1905 36003
rect 1943 35969 1977 36003
rect 2015 35969 2049 36003
rect 2087 35969 2121 36003
rect 2159 35969 2193 36003
rect 2231 35969 2265 36003
rect 2303 35969 2337 36003
rect 2375 35969 2409 36003
rect 2447 35969 2481 36003
rect 2519 35969 2553 36003
rect 2591 35969 2625 36003
rect 2663 35969 2697 36003
rect 2735 35969 2769 36003
rect 2807 35969 2841 36003
rect 2879 35969 2913 36003
rect 2951 35969 2985 36003
rect 3023 35969 3057 36003
rect 3095 35969 3129 36003
rect 3167 35969 3201 36003
rect 3239 35969 3273 36003
rect 3311 35969 3345 36003
rect 3383 35969 3417 36003
rect 3455 35969 3489 36003
rect 3527 35969 3561 36003
rect 3599 35969 3633 36003
rect 3671 35969 3705 36003
rect 3743 35969 3777 36003
rect 3815 35969 3849 36003
rect 3887 35969 3921 36003
rect 3959 35969 3993 36003
rect 4031 35969 4065 36003
rect 4103 35969 4137 36003
rect 4175 35969 4209 36003
rect 4247 35969 4281 36003
rect 4319 35969 4353 36003
rect 4391 35969 4425 36003
rect 4463 35969 4497 36003
rect 4535 35969 4569 36003
rect 4607 35969 4641 36003
rect 4679 35969 4713 36003
rect 4751 35969 4785 36003
rect 4823 35969 4857 36003
rect 4895 35969 4929 36003
rect 4967 35969 5001 36003
rect 5039 35969 5073 36003
rect 5111 35969 5145 36003
rect 5183 35969 5217 36003
rect 5255 35969 5289 36003
rect 5327 35969 5361 36003
rect 5399 35969 5433 36003
rect 5471 35969 5505 36003
rect 5543 35969 5577 36003
rect 5615 35969 5649 36003
rect 5687 35969 5721 36003
rect 5759 35969 5793 36003
rect 5831 35969 5865 36003
rect 5903 35969 5937 36003
rect 5975 35969 6009 36003
rect 6047 35969 6081 36003
rect 6119 35969 6153 36003
rect 6191 35969 6225 36003
rect 6263 35969 6297 36003
rect 6335 35969 6369 36003
rect 6407 35969 6441 36003
rect 6479 35969 6513 36003
rect 6551 35969 6585 36003
rect 6623 35969 6657 36003
rect 6695 35969 6729 36003
rect 6767 35969 6801 36003
rect 6839 35969 6873 36003
rect 6911 35969 6945 36003
rect 6983 35969 7017 36003
rect 7055 35969 7089 36003
rect 7127 35969 7161 36003
rect 7199 35969 7233 36003
rect 7271 35969 7305 36003
rect 7343 35969 7377 36003
rect 7415 35969 7449 36003
rect 7487 35969 7521 36003
rect 7559 35969 7593 36003
rect 7631 35969 7665 36003
rect 7703 35969 7737 36003
rect 7775 35969 7809 36003
rect 7847 35969 7881 36003
rect 7919 35969 7953 36003
rect 7991 35969 8025 36003
rect 8063 35969 8097 36003
rect 8135 35969 8169 36003
rect 8207 35969 8241 36003
rect 8279 35969 8313 36003
rect 8351 35969 8385 36003
rect 8423 35969 8457 36003
rect 8495 35969 8529 36003
rect 8567 35969 8601 36003
rect 8639 35969 8673 36003
rect 8711 35969 8745 36003
rect 8783 35969 8817 36003
rect 8855 35969 8889 36003
rect 8927 35969 8961 36003
rect 8999 35969 9033 36003
rect 9071 35969 9105 36003
rect 9143 35969 9177 36003
rect 9215 35969 9249 36003
rect 9287 35969 9321 36003
rect 9359 35969 9393 36003
rect 9431 35969 9465 36003
rect 9503 35969 9537 36003
rect 9575 35969 9609 36003
rect 9647 35969 9681 36003
rect 9719 35969 9753 36003
rect 9791 35969 9825 36003
rect 9863 35969 9897 36003
rect 9935 35969 9969 36003
rect 10007 35969 10041 36003
rect 10079 35969 10113 36003
rect 10151 35969 10185 36003
rect 10223 35969 10257 36003
rect 10295 35969 10329 36003
rect 10367 35969 10401 36003
rect 10439 35969 10473 36003
rect 10511 35969 10545 36003
rect 10583 35969 10617 36003
rect 10655 35969 10689 36003
rect 10727 35969 10761 36003
rect 10799 35969 10833 36003
rect 10871 35969 10905 36003
rect 10943 35969 10977 36003
rect 11015 35969 11049 36003
rect 11087 35969 11121 36003
rect 11159 35969 11193 36003
rect 11231 35969 11265 36003
rect 11303 35969 11337 36003
rect 11375 35969 11409 36003
rect 11447 35969 11481 36003
rect 11519 35969 11553 36003
rect 11591 35969 11625 36003
rect 11663 35969 11697 36003
rect 11735 35969 11769 36003
rect 11807 35969 11841 36003
rect 11879 35969 11913 36003
rect 11951 35969 11985 36003
rect 12023 35969 12057 36003
rect 12095 35969 12129 36003
rect 12167 35969 12201 36003
rect 12239 35969 12273 36003
rect 12311 35969 12345 36003
rect 12383 35969 12417 36003
rect 12455 35969 12489 36003
rect 12527 35969 12561 36003
rect 12599 35969 12633 36003
rect 12671 35969 12705 36003
rect 12743 35969 12777 36003
rect 12815 35969 12849 36003
rect 12887 35969 12921 36003
rect 12959 35969 12993 36003
rect 13031 35969 13065 36003
rect 13103 35969 13137 36003
rect 13175 35969 13209 36003
rect 13247 35969 13281 36003
rect 13319 35969 13353 36003
rect 13391 35969 13425 36003
rect 13463 35969 13497 36003
rect 13535 35969 13569 36003
rect 13607 35969 13641 36003
rect 13679 35969 13713 36003
rect 13751 35969 13785 36003
rect 13823 35969 13857 36003
rect 13895 35969 13929 36003
rect 13967 35969 14001 36003
rect 807 35850 841 35884
rect 807 35778 841 35812
rect 14142 35771 14176 35805
rect 807 35706 841 35740
rect 14142 35699 14176 35733
rect 807 35634 841 35668
rect 14142 35627 14176 35661
rect 807 35562 841 35596
rect 14142 35555 14176 35589
rect 807 35490 841 35524
rect 14142 35483 14176 35517
rect 807 35418 841 35452
rect 14142 35411 14176 35445
rect 807 35346 841 35380
rect 14142 35339 14176 35373
rect 807 35274 841 35308
rect 14142 35267 14176 35301
rect 807 35202 841 35236
rect 14142 35195 14176 35229
rect 807 35130 841 35164
rect 14142 35123 14176 35157
rect 807 35058 841 35092
rect 14142 35051 14176 35085
rect 807 34986 841 35020
rect 14142 34979 14176 35013
rect 807 34914 841 34948
rect 14142 34907 14176 34941
rect 807 34842 841 34876
rect 14142 34835 14176 34869
rect 807 34770 841 34804
rect 807 34698 841 34732
rect 14142 34763 14176 34797
rect 807 34626 841 34660
rect 807 34554 841 34588
rect 807 34482 841 34516
rect 807 34410 841 34444
rect 807 34338 841 34372
rect 807 34266 841 34300
rect 807 34194 841 34228
rect 807 34122 841 34156
rect 807 34050 841 34084
rect 807 33978 841 34012
rect 807 33906 841 33940
rect 807 33834 841 33868
rect 807 33762 841 33796
rect 807 33690 841 33724
rect 807 33618 841 33652
rect 807 33546 841 33580
rect 807 33474 841 33508
rect 807 33402 841 33436
rect 807 33330 841 33364
rect 807 33258 841 33292
rect 807 33186 841 33220
rect 807 33114 841 33148
rect 807 33042 841 33076
rect 807 32970 841 33004
rect 807 32898 841 32932
rect 807 32826 841 32860
rect 807 32754 841 32788
rect 807 32682 841 32716
rect 807 32610 841 32644
rect 807 32538 841 32572
rect 807 32466 841 32500
rect 807 32394 841 32428
rect 807 32322 841 32356
rect 807 32250 841 32284
rect 807 32178 841 32212
rect 807 32106 841 32140
rect 807 32034 841 32068
rect 807 31962 841 31996
rect 807 31890 841 31924
rect 807 31818 841 31852
rect 807 31746 841 31780
rect 807 31674 841 31708
rect 807 31602 841 31636
rect 807 31530 841 31564
rect 807 31458 841 31492
rect 807 31386 841 31420
rect 807 31314 841 31348
rect 807 31242 841 31276
rect 807 31170 841 31204
rect 807 31098 841 31132
rect 807 31026 841 31060
rect 807 30954 841 30988
rect 807 30882 841 30916
rect 807 30810 841 30844
rect 807 30738 841 30772
rect 807 30666 841 30700
rect 807 30594 841 30628
rect 807 30522 841 30556
rect 807 30450 841 30484
rect 807 30378 841 30412
rect 807 30306 841 30340
rect 807 30234 841 30268
rect 807 30162 841 30196
rect 807 30090 841 30124
rect 807 30018 841 30052
rect 807 29946 841 29980
rect 807 29874 841 29908
rect 807 29802 841 29836
rect 807 29730 841 29764
rect 807 29658 841 29692
rect 807 29586 841 29620
rect 807 29514 841 29548
rect 807 29442 841 29476
rect 807 29370 841 29404
rect 807 29298 841 29332
rect 807 29226 841 29260
rect 807 29154 841 29188
rect 807 29082 841 29116
rect 807 29010 841 29044
rect 807 28938 841 28972
rect 807 28866 841 28900
rect 807 28794 841 28828
rect 807 28722 841 28756
rect 807 28650 841 28684
rect 807 28578 841 28612
rect 807 28506 841 28540
rect 807 28434 841 28468
rect 807 28362 841 28396
rect 807 28290 841 28324
rect 807 28218 841 28252
rect 807 28146 841 28180
rect 807 28074 841 28108
rect 807 28002 841 28036
rect 807 27930 841 27964
rect 807 27858 841 27892
rect 807 27786 841 27820
rect 807 27714 841 27748
rect 807 27642 841 27676
rect 807 27570 841 27604
rect 807 27498 841 27532
rect 807 27426 841 27460
rect 807 27354 841 27388
rect 807 27282 841 27316
rect 807 27210 841 27244
rect 807 27138 841 27172
rect 807 27066 841 27100
rect 807 26994 841 27028
rect 807 26922 841 26956
rect 807 26850 841 26884
rect 807 26778 841 26812
rect 807 26706 841 26740
rect 807 26634 841 26668
rect 807 26562 841 26596
rect 807 26490 841 26524
rect 807 26418 841 26452
rect 807 26346 841 26380
rect 807 26274 841 26308
rect 807 26202 841 26236
rect 807 26130 841 26164
rect 807 26058 841 26092
rect 807 25986 841 26020
rect 807 25914 841 25948
rect 807 25842 841 25876
rect 807 25770 841 25804
rect 807 25698 841 25732
rect 807 25626 841 25660
rect 807 25554 841 25588
rect 807 25482 841 25516
rect 807 25410 841 25444
rect 807 25338 841 25372
rect 807 25266 841 25300
rect 807 25194 841 25228
rect 807 25122 841 25156
rect 807 25050 841 25084
rect 807 24978 841 25012
rect 807 24906 841 24940
rect 807 24834 841 24868
rect 807 24762 841 24796
rect 807 24690 841 24724
rect 807 24618 841 24652
rect 807 24546 841 24580
rect 807 24474 841 24508
rect 807 24402 841 24436
rect 807 24330 841 24364
rect 807 24258 841 24292
rect 807 24186 841 24220
rect 807 24114 841 24148
rect 807 24042 841 24076
rect 807 23970 841 24004
rect 807 23898 841 23932
rect 807 23826 841 23860
rect 807 23754 841 23788
rect 807 23682 841 23716
rect 807 23610 841 23644
rect 807 23538 841 23572
rect 807 23466 841 23500
rect 807 23394 841 23428
rect 807 23322 841 23356
rect 807 23250 841 23284
rect 807 23178 841 23212
rect 807 23106 841 23140
rect 807 23034 841 23068
rect 807 22962 841 22996
rect 807 22890 841 22924
rect 807 22818 841 22852
rect 807 22746 841 22780
rect 807 22674 841 22708
rect 807 22602 841 22636
rect 807 22530 841 22564
rect 807 22458 841 22492
rect 807 22386 841 22420
rect 807 22314 841 22348
rect 807 22242 841 22276
rect 807 22170 841 22204
rect 807 22098 841 22132
rect 807 22026 841 22060
rect 807 21954 841 21988
rect 807 21882 841 21916
rect 807 21810 841 21844
rect 807 21738 841 21772
rect 807 21666 841 21700
rect 807 21594 841 21628
rect 807 21522 841 21556
rect 807 21450 841 21484
rect 807 21378 841 21412
rect 807 21306 841 21340
rect 807 21234 841 21268
rect 807 21162 841 21196
rect 807 21090 841 21124
rect 807 21018 841 21052
rect 807 20946 841 20980
rect 807 20874 841 20908
rect 807 20802 841 20836
rect 807 20730 841 20764
rect 807 20658 841 20692
rect 807 20586 841 20620
rect 807 20514 841 20548
rect 807 20442 841 20476
rect 807 20370 841 20404
rect 807 20298 841 20332
rect 807 20226 841 20260
rect 807 20154 841 20188
rect 807 20082 841 20116
rect 807 20010 841 20044
rect 807 19938 841 19972
rect 807 19866 841 19900
rect 807 19794 841 19828
rect 807 19722 841 19756
rect 807 19650 841 19684
rect 807 19578 841 19612
rect 807 19506 841 19540
rect 807 19434 841 19468
rect 807 19362 841 19396
rect 807 19290 841 19324
rect 807 19218 841 19252
rect 807 19146 841 19180
rect 807 19074 841 19108
rect 807 19002 841 19036
rect 807 18930 841 18964
rect 807 18858 841 18892
rect 807 18786 841 18820
rect 807 18714 841 18748
rect 807 18642 841 18676
rect 807 18570 841 18604
rect 807 18498 841 18532
rect 807 18426 841 18460
rect 807 18354 841 18388
rect 807 18282 841 18316
rect 807 18210 841 18244
rect 807 18138 841 18172
rect 807 18066 841 18100
rect 807 17994 841 18028
rect 807 17922 841 17956
rect 807 17850 841 17884
rect 807 17778 841 17812
rect 807 17706 841 17740
rect 807 17634 841 17668
rect 807 17562 841 17596
rect 807 17490 841 17524
rect 807 17418 841 17452
rect 807 17346 841 17380
rect 807 17274 841 17308
rect 807 17202 841 17236
rect 807 17130 841 17164
rect 807 17058 841 17092
rect 807 16986 841 17020
rect 807 16914 841 16948
rect 807 16842 841 16876
rect 807 16770 841 16804
rect 807 16698 841 16732
rect 807 16626 841 16660
rect 807 16554 841 16588
rect 807 16482 841 16516
rect 807 16410 841 16444
rect 807 16338 841 16372
rect 807 16266 841 16300
rect 807 16194 841 16228
rect 807 16122 841 16156
rect 807 16050 841 16084
rect 807 15978 841 16012
rect 807 15906 841 15940
rect 807 15834 841 15868
rect 807 15762 841 15796
rect 807 15690 841 15724
rect 807 15618 841 15652
rect 807 15546 841 15580
rect 807 15474 841 15508
rect 807 15402 841 15436
rect 807 15330 841 15364
rect 807 15258 841 15292
rect 807 15186 841 15220
rect 807 15114 841 15148
rect 807 15042 841 15076
rect 807 14970 841 15004
rect 807 14898 841 14932
rect 807 14826 841 14860
rect 807 14754 841 14788
rect 807 14682 841 14716
rect 807 14610 841 14644
rect 807 14538 841 14572
rect 807 14466 841 14500
rect 807 14394 841 14428
rect 807 14322 841 14356
rect 807 14250 841 14284
rect 807 14178 841 14212
rect 807 14106 841 14140
rect 807 14034 841 14068
rect 807 13962 841 13996
rect 807 13890 841 13924
rect 807 13818 841 13852
rect 807 13746 841 13780
rect 807 13674 841 13708
rect 807 13602 841 13636
rect 807 13530 841 13564
rect 807 13458 841 13492
rect 807 13386 841 13420
rect 807 13314 841 13348
rect 807 13242 841 13276
rect 807 13170 841 13204
rect 807 13098 841 13132
rect 807 13026 841 13060
rect 807 12954 841 12988
rect 807 12882 841 12916
rect 807 12810 841 12844
rect 807 12738 841 12772
rect 807 12666 841 12700
rect 807 12594 841 12628
rect 807 12522 841 12556
rect 807 12450 841 12484
rect 807 12378 841 12412
rect 807 12306 841 12340
rect 807 12234 841 12268
rect 807 12162 841 12196
rect 807 12090 841 12124
rect 807 12018 841 12052
rect 807 11946 841 11980
rect 807 11874 841 11908
rect 807 11802 841 11836
rect 807 11730 841 11764
rect 807 11658 841 11692
rect 807 11586 841 11620
rect 807 11514 841 11548
rect 807 11442 841 11476
rect 807 11370 841 11404
rect 807 11298 841 11332
rect 807 11226 841 11260
rect 807 11154 841 11188
rect 807 11082 841 11116
rect 807 11010 841 11044
rect 807 10938 841 10972
rect 807 10866 841 10900
rect 807 10794 841 10828
rect 807 10722 841 10756
rect 807 10650 841 10684
rect 807 10578 841 10612
rect 807 10506 841 10540
rect 807 10434 841 10468
rect 807 10362 841 10396
rect 807 10290 841 10324
rect 807 10218 841 10252
rect 1325 34616 1327 34650
rect 1327 34616 1359 34650
rect 1397 34616 1429 34650
rect 1429 34616 1431 34650
rect 1469 34616 1497 34650
rect 1497 34616 1503 34650
rect 1541 34616 1565 34650
rect 1565 34616 1575 34650
rect 1613 34616 1633 34650
rect 1633 34616 1647 34650
rect 1685 34616 1701 34650
rect 1701 34616 1719 34650
rect 1757 34616 1769 34650
rect 1769 34616 1791 34650
rect 1829 34616 1837 34650
rect 1837 34616 1863 34650
rect 1901 34616 1905 34650
rect 1905 34616 1935 34650
rect 1973 34616 2007 34650
rect 2045 34616 2075 34650
rect 2075 34616 2079 34650
rect 2117 34616 2143 34650
rect 2143 34616 2151 34650
rect 2189 34616 2211 34650
rect 2211 34616 2223 34650
rect 2261 34616 2279 34650
rect 2279 34616 2295 34650
rect 2333 34616 2347 34650
rect 2347 34616 2367 34650
rect 2405 34616 2415 34650
rect 2415 34616 2439 34650
rect 2477 34616 2483 34650
rect 2483 34616 2511 34650
rect 2549 34616 2551 34650
rect 2551 34616 2583 34650
rect 2621 34616 2653 34650
rect 2653 34616 2655 34650
rect 2693 34616 2721 34650
rect 2721 34616 2727 34650
rect 2765 34616 2789 34650
rect 2789 34616 2799 34650
rect 2837 34616 2857 34650
rect 2857 34616 2871 34650
rect 2909 34616 2925 34650
rect 2925 34616 2943 34650
rect 2981 34616 2993 34650
rect 2993 34616 3015 34650
rect 3053 34616 3061 34650
rect 3061 34616 3087 34650
rect 3125 34616 3129 34650
rect 3129 34616 3159 34650
rect 3197 34616 3231 34650
rect 3269 34616 3299 34650
rect 3299 34616 3303 34650
rect 3341 34616 3367 34650
rect 3367 34616 3375 34650
rect 3413 34616 3435 34650
rect 3435 34616 3447 34650
rect 3485 34616 3503 34650
rect 3503 34616 3519 34650
rect 3557 34616 3571 34650
rect 3571 34616 3591 34650
rect 3629 34616 3639 34650
rect 3639 34616 3663 34650
rect 3701 34616 3707 34650
rect 3707 34616 3735 34650
rect 3773 34616 3775 34650
rect 3775 34616 3807 34650
rect 3845 34616 3877 34650
rect 3877 34616 3879 34650
rect 3917 34616 3945 34650
rect 3945 34616 3951 34650
rect 3989 34616 4013 34650
rect 4013 34616 4023 34650
rect 4061 34616 4081 34650
rect 4081 34616 4095 34650
rect 4133 34616 4149 34650
rect 4149 34616 4167 34650
rect 4205 34616 4217 34650
rect 4217 34616 4239 34650
rect 4277 34616 4285 34650
rect 4285 34616 4311 34650
rect 4349 34616 4353 34650
rect 4353 34616 4383 34650
rect 4421 34616 4455 34650
rect 4493 34616 4523 34650
rect 4523 34616 4527 34650
rect 4565 34616 4591 34650
rect 4591 34616 4599 34650
rect 4637 34616 4659 34650
rect 4659 34616 4671 34650
rect 4709 34616 4727 34650
rect 4727 34616 4743 34650
rect 4781 34616 4795 34650
rect 4795 34616 4815 34650
rect 4853 34616 4863 34650
rect 4863 34616 4887 34650
rect 4925 34616 4931 34650
rect 4931 34616 4959 34650
rect 4997 34616 4999 34650
rect 4999 34616 5031 34650
rect 5069 34616 5101 34650
rect 5101 34616 5103 34650
rect 5141 34616 5169 34650
rect 5169 34616 5175 34650
rect 5213 34616 5237 34650
rect 5237 34616 5247 34650
rect 5285 34616 5305 34650
rect 5305 34616 5319 34650
rect 5357 34616 5373 34650
rect 5373 34616 5391 34650
rect 5429 34616 5441 34650
rect 5441 34616 5463 34650
rect 5501 34616 5509 34650
rect 5509 34616 5535 34650
rect 5573 34616 5577 34650
rect 5577 34616 5607 34650
rect 5645 34616 5679 34650
rect 5717 34616 5747 34650
rect 5747 34616 5751 34650
rect 5789 34616 5815 34650
rect 5815 34616 5823 34650
rect 5861 34616 5883 34650
rect 5883 34616 5895 34650
rect 5933 34616 5951 34650
rect 5951 34616 5967 34650
rect 6005 34616 6019 34650
rect 6019 34616 6039 34650
rect 6077 34616 6087 34650
rect 6087 34616 6111 34650
rect 6149 34616 6155 34650
rect 6155 34616 6183 34650
rect 6221 34616 6223 34650
rect 6223 34616 6255 34650
rect 6293 34616 6325 34650
rect 6325 34616 6327 34650
rect 6365 34616 6393 34650
rect 6393 34616 6399 34650
rect 6437 34616 6461 34650
rect 6461 34616 6471 34650
rect 6509 34616 6529 34650
rect 6529 34616 6543 34650
rect 6581 34616 6597 34650
rect 6597 34616 6615 34650
rect 6653 34616 6665 34650
rect 6665 34616 6687 34650
rect 6725 34616 6733 34650
rect 6733 34616 6759 34650
rect 6797 34616 6801 34650
rect 6801 34616 6831 34650
rect 6869 34616 6903 34650
rect 6941 34616 6971 34650
rect 6971 34616 6975 34650
rect 7013 34616 7039 34650
rect 7039 34616 7047 34650
rect 7085 34616 7107 34650
rect 7107 34616 7119 34650
rect 7157 34616 7175 34650
rect 7175 34616 7191 34650
rect 7229 34616 7243 34650
rect 7243 34616 7263 34650
rect 7301 34616 7311 34650
rect 7311 34616 7335 34650
rect 7373 34616 7379 34650
rect 7379 34616 7407 34650
rect 7445 34616 7447 34650
rect 7447 34616 7479 34650
rect 7517 34616 7549 34650
rect 7549 34616 7551 34650
rect 7589 34616 7617 34650
rect 7617 34616 7623 34650
rect 7661 34616 7685 34650
rect 7685 34616 7695 34650
rect 7733 34616 7753 34650
rect 7753 34616 7767 34650
rect 7805 34616 7821 34650
rect 7821 34616 7839 34650
rect 7877 34616 7889 34650
rect 7889 34616 7911 34650
rect 7949 34616 7957 34650
rect 7957 34616 7983 34650
rect 8021 34616 8025 34650
rect 8025 34616 8055 34650
rect 8093 34616 8127 34650
rect 8165 34616 8195 34650
rect 8195 34616 8199 34650
rect 8237 34616 8263 34650
rect 8263 34616 8271 34650
rect 8309 34616 8331 34650
rect 8331 34616 8343 34650
rect 8381 34616 8399 34650
rect 8399 34616 8415 34650
rect 8453 34616 8467 34650
rect 8467 34616 8487 34650
rect 8525 34616 8535 34650
rect 8535 34616 8559 34650
rect 8597 34616 8603 34650
rect 8603 34616 8631 34650
rect 8669 34616 8671 34650
rect 8671 34616 8703 34650
rect 8741 34616 8773 34650
rect 8773 34616 8775 34650
rect 8813 34616 8841 34650
rect 8841 34616 8847 34650
rect 8885 34616 8909 34650
rect 8909 34616 8919 34650
rect 8957 34616 8977 34650
rect 8977 34616 8991 34650
rect 9029 34616 9045 34650
rect 9045 34616 9063 34650
rect 9101 34616 9113 34650
rect 9113 34616 9135 34650
rect 9173 34616 9181 34650
rect 9181 34616 9207 34650
rect 9245 34616 9249 34650
rect 9249 34616 9279 34650
rect 9317 34616 9351 34650
rect 9389 34616 9419 34650
rect 9419 34616 9423 34650
rect 9461 34616 9487 34650
rect 9487 34616 9495 34650
rect 9533 34616 9555 34650
rect 9555 34616 9567 34650
rect 9605 34616 9623 34650
rect 9623 34616 9639 34650
rect 9677 34616 9691 34650
rect 9691 34616 9711 34650
rect 9749 34616 9759 34650
rect 9759 34616 9783 34650
rect 9821 34616 9827 34650
rect 9827 34616 9855 34650
rect 9893 34616 9895 34650
rect 9895 34616 9927 34650
rect 9965 34616 9997 34650
rect 9997 34616 9999 34650
rect 10037 34616 10065 34650
rect 10065 34616 10071 34650
rect 10109 34616 10133 34650
rect 10133 34616 10143 34650
rect 10181 34616 10201 34650
rect 10201 34616 10215 34650
rect 10253 34616 10269 34650
rect 10269 34616 10287 34650
rect 10325 34616 10337 34650
rect 10337 34616 10359 34650
rect 10397 34616 10405 34650
rect 10405 34616 10431 34650
rect 10469 34616 10473 34650
rect 10473 34616 10503 34650
rect 10541 34616 10575 34650
rect 10613 34616 10643 34650
rect 10643 34616 10647 34650
rect 10685 34616 10711 34650
rect 10711 34616 10719 34650
rect 10757 34616 10779 34650
rect 10779 34616 10791 34650
rect 10829 34616 10847 34650
rect 10847 34616 10863 34650
rect 10901 34616 10915 34650
rect 10915 34616 10935 34650
rect 10973 34616 10983 34650
rect 10983 34616 11007 34650
rect 11045 34616 11051 34650
rect 11051 34616 11079 34650
rect 11117 34616 11119 34650
rect 11119 34616 11151 34650
rect 11189 34616 11221 34650
rect 11221 34616 11223 34650
rect 11261 34616 11289 34650
rect 11289 34616 11295 34650
rect 11333 34616 11357 34650
rect 11357 34616 11367 34650
rect 11405 34616 11425 34650
rect 11425 34616 11439 34650
rect 11477 34616 11493 34650
rect 11493 34616 11511 34650
rect 11549 34616 11561 34650
rect 11561 34616 11583 34650
rect 11621 34616 11629 34650
rect 11629 34616 11655 34650
rect 11693 34616 11697 34650
rect 11697 34616 11727 34650
rect 11765 34616 11799 34650
rect 11837 34616 11867 34650
rect 11867 34616 11871 34650
rect 11909 34616 11935 34650
rect 11935 34616 11943 34650
rect 11981 34616 12003 34650
rect 12003 34616 12015 34650
rect 12053 34616 12071 34650
rect 12071 34616 12087 34650
rect 12125 34616 12139 34650
rect 12139 34616 12159 34650
rect 12197 34616 12207 34650
rect 12207 34616 12231 34650
rect 12269 34616 12275 34650
rect 12275 34616 12303 34650
rect 12341 34616 12343 34650
rect 12343 34616 12375 34650
rect 12413 34616 12445 34650
rect 12445 34616 12447 34650
rect 12485 34616 12513 34650
rect 12513 34616 12519 34650
rect 12557 34616 12581 34650
rect 12581 34616 12591 34650
rect 12629 34616 12649 34650
rect 12649 34616 12663 34650
rect 12701 34616 12717 34650
rect 12717 34616 12735 34650
rect 12773 34616 12785 34650
rect 12785 34616 12807 34650
rect 12845 34616 12853 34650
rect 12853 34616 12879 34650
rect 12917 34616 12921 34650
rect 12921 34616 12951 34650
rect 12989 34616 13023 34650
rect 13061 34616 13091 34650
rect 13091 34616 13095 34650
rect 13133 34616 13159 34650
rect 13159 34616 13167 34650
rect 13205 34616 13227 34650
rect 13227 34616 13239 34650
rect 13277 34616 13295 34650
rect 13295 34616 13311 34650
rect 13349 34616 13363 34650
rect 13363 34616 13383 34650
rect 13421 34616 13431 34650
rect 13431 34616 13455 34650
rect 13493 34616 13499 34650
rect 13499 34616 13527 34650
rect 13565 34616 13567 34650
rect 13567 34616 13599 34650
rect 13637 34616 13669 34650
rect 13669 34616 13671 34650
rect 1192 34487 1226 34509
rect 1192 34475 1226 34487
rect 1192 34419 1226 34437
rect 1192 34403 1226 34419
rect 1192 34351 1226 34365
rect 1192 34331 1226 34351
rect 1192 34283 1226 34293
rect 1192 34259 1226 34283
rect 1192 34215 1226 34221
rect 1192 34187 1226 34215
rect 1192 34147 1226 34149
rect 1192 34115 1226 34147
rect 1192 34045 1226 34077
rect 1192 34043 1226 34045
rect 1192 33977 1226 34005
rect 1192 33971 1226 33977
rect 1192 33909 1226 33933
rect 1192 33899 1226 33909
rect 1192 33841 1226 33861
rect 1192 33827 1226 33841
rect 1192 33773 1226 33789
rect 1192 33755 1226 33773
rect 1192 33705 1226 33717
rect 1192 33683 1226 33705
rect 1192 33637 1226 33645
rect 1192 33611 1226 33637
rect 1192 33569 1226 33573
rect 1192 33539 1226 33569
rect 1192 33467 1226 33501
rect 1192 33399 1226 33429
rect 1192 33395 1226 33399
rect 1192 33331 1226 33357
rect 1192 33323 1226 33331
rect 1192 33263 1226 33285
rect 1192 33251 1226 33263
rect 1192 33195 1226 33213
rect 1192 33179 1226 33195
rect 1192 33127 1226 33141
rect 1192 33107 1226 33127
rect 1192 33059 1226 33069
rect 1192 33035 1226 33059
rect 1192 32991 1226 32997
rect 1192 32963 1226 32991
rect 1192 32923 1226 32925
rect 1192 32891 1226 32923
rect 1192 32821 1226 32853
rect 1192 32819 1226 32821
rect 1192 32753 1226 32781
rect 1192 32747 1226 32753
rect 1192 32685 1226 32709
rect 1192 32675 1226 32685
rect 1192 32617 1226 32637
rect 1192 32603 1226 32617
rect 1192 32549 1226 32565
rect 1192 32531 1226 32549
rect 1192 32481 1226 32493
rect 1192 32459 1226 32481
rect 1192 32413 1226 32421
rect 1192 32387 1226 32413
rect 1192 32345 1226 32349
rect 1192 32315 1226 32345
rect 1192 32243 1226 32277
rect 1192 32175 1226 32205
rect 1192 32171 1226 32175
rect 1192 32107 1226 32133
rect 1192 32099 1226 32107
rect 1192 32039 1226 32061
rect 1192 32027 1226 32039
rect 1192 31971 1226 31989
rect 1192 31955 1226 31971
rect 1192 31903 1226 31917
rect 1192 31883 1226 31903
rect 1192 31835 1226 31845
rect 1192 31811 1226 31835
rect 1192 31767 1226 31773
rect 1192 31739 1226 31767
rect 1192 31699 1226 31701
rect 1192 31667 1226 31699
rect 1192 31597 1226 31629
rect 1192 31595 1226 31597
rect 1192 31529 1226 31557
rect 1192 31523 1226 31529
rect 1192 31461 1226 31485
rect 1192 31451 1226 31461
rect 1192 31393 1226 31413
rect 1192 31379 1226 31393
rect 13768 34500 13802 34508
rect 13768 34474 13802 34500
rect 13768 34432 13802 34436
rect 13768 34402 13802 34432
rect 13768 34330 13802 34364
rect 13768 34262 13802 34292
rect 13768 34258 13802 34262
rect 13768 34194 13802 34220
rect 13768 34186 13802 34194
rect 13768 34126 13802 34148
rect 13768 34114 13802 34126
rect 13768 34058 13802 34076
rect 13768 34042 13802 34058
rect 13768 33990 13802 34004
rect 13768 33970 13802 33990
rect 13768 33922 13802 33932
rect 13768 33898 13802 33922
rect 13768 33854 13802 33860
rect 13768 33826 13802 33854
rect 13768 33786 13802 33788
rect 13768 33754 13802 33786
rect 13768 33684 13802 33716
rect 13768 33682 13802 33684
rect 13768 33616 13802 33644
rect 13768 33610 13802 33616
rect 13768 33548 13802 33572
rect 13768 33538 13802 33548
rect 13768 33480 13802 33500
rect 13768 33466 13802 33480
rect 13768 33412 13802 33428
rect 13768 33394 13802 33412
rect 13768 33344 13802 33356
rect 13768 33322 13802 33344
rect 13768 33276 13802 33284
rect 13768 33250 13802 33276
rect 13768 33208 13802 33212
rect 13768 33178 13802 33208
rect 13768 33106 13802 33140
rect 13768 33038 13802 33068
rect 13768 33034 13802 33038
rect 13768 32970 13802 32996
rect 13768 32962 13802 32970
rect 13768 32902 13802 32924
rect 13768 32890 13802 32902
rect 13768 32834 13802 32852
rect 13768 32818 13802 32834
rect 13768 32766 13802 32780
rect 13768 32746 13802 32766
rect 13768 32698 13802 32708
rect 13768 32674 13802 32698
rect 13768 32630 13802 32636
rect 13768 32602 13802 32630
rect 13768 32562 13802 32564
rect 13768 32530 13802 32562
rect 13768 32460 13802 32492
rect 13768 32458 13802 32460
rect 13768 32392 13802 32420
rect 13768 32386 13802 32392
rect 13768 32324 13802 32348
rect 13768 32314 13802 32324
rect 13768 32256 13802 32276
rect 13768 32242 13802 32256
rect 13768 32188 13802 32204
rect 13768 32170 13802 32188
rect 13768 32120 13802 32132
rect 13768 32098 13802 32120
rect 13768 32052 13802 32060
rect 13768 32026 13802 32052
rect 13768 31984 13802 31988
rect 13768 31954 13802 31984
rect 13768 31882 13802 31916
rect 13768 31814 13802 31844
rect 13768 31810 13802 31814
rect 13768 31746 13802 31772
rect 13768 31738 13802 31746
rect 13768 31678 13802 31700
rect 13768 31666 13802 31678
rect 13768 31610 13802 31628
rect 13768 31594 13802 31610
rect 13768 31542 13802 31556
rect 13768 31522 13802 31542
rect 13768 31474 13802 31484
rect 13768 31450 13802 31474
rect 1192 31325 1226 31341
rect 1192 31307 1226 31325
rect 1192 31257 1226 31269
rect 1192 31235 1226 31257
rect 1192 31189 1226 31197
rect 1192 31163 1226 31189
rect 1192 31121 1226 31125
rect 1192 31091 1226 31121
rect 1192 31019 1226 31053
rect 1192 30951 1226 30981
rect 1192 30947 1226 30951
rect 1192 30883 1226 30909
rect 1192 30875 1226 30883
rect 1192 30815 1226 30837
rect 1192 30803 1226 30815
rect 1192 30747 1226 30765
rect 1192 30731 1226 30747
rect 1192 30679 1226 30693
rect 1192 30659 1226 30679
rect 1192 30611 1226 30621
rect 1192 30587 1226 30611
rect 1192 30543 1226 30549
rect 1192 30515 1226 30543
rect 1192 30475 1226 30477
rect 1192 30443 1226 30475
rect 1192 30373 1226 30405
rect 1192 30371 1226 30373
rect 1192 30305 1226 30333
rect 1192 30299 1226 30305
rect 1192 30237 1226 30261
rect 1192 30227 1226 30237
rect 1192 30169 1226 30189
rect 1192 30155 1226 30169
rect 1192 30101 1226 30117
rect 1192 30083 1226 30101
rect 1192 30033 1226 30045
rect 1192 30011 1226 30033
rect 1192 29965 1226 29973
rect 1192 29939 1226 29965
rect 1192 29897 1226 29901
rect 1192 29867 1226 29897
rect 1192 29795 1226 29829
rect 1192 29727 1226 29757
rect 1192 29723 1226 29727
rect 1192 29659 1226 29685
rect 1192 29651 1226 29659
rect 1192 29591 1226 29613
rect 1192 29579 1226 29591
rect 1192 29523 1226 29541
rect 1192 29507 1226 29523
rect 1192 29455 1226 29469
rect 1192 29435 1226 29455
rect 1192 29387 1226 29397
rect 1192 29363 1226 29387
rect 1192 29319 1226 29325
rect 1192 29291 1226 29319
rect 1192 29251 1226 29253
rect 1192 29219 1226 29251
rect 1192 29149 1226 29181
rect 1192 29147 1226 29149
rect 1192 29081 1226 29109
rect 1192 29075 1226 29081
rect 1192 29013 1226 29037
rect 1192 29003 1226 29013
rect 1192 28945 1226 28965
rect 1192 28931 1226 28945
rect 1192 28877 1226 28893
rect 1192 28859 1226 28877
rect 1192 28809 1226 28821
rect 1192 28787 1226 28809
rect 1192 28741 1226 28749
rect 1192 28715 1226 28741
rect 1192 28673 1226 28677
rect 1192 28643 1226 28673
rect 1192 28571 1226 28605
rect 1192 28503 1226 28533
rect 1192 28499 1226 28503
rect 1192 28435 1226 28461
rect 1192 28427 1226 28435
rect 1192 28367 1226 28389
rect 1192 28355 1226 28367
rect 1192 28299 1226 28317
rect 1192 28283 1226 28299
rect 1192 28231 1226 28245
rect 1192 28211 1226 28231
rect 1192 28163 1226 28173
rect 1192 28139 1226 28163
rect 1192 28095 1226 28101
rect 1192 28067 1226 28095
rect 1192 28027 1226 28029
rect 1192 27995 1226 28027
rect 1192 27925 1226 27957
rect 1192 27923 1226 27925
rect 1192 27857 1226 27885
rect 1192 27851 1226 27857
rect 1192 27789 1226 27813
rect 1192 27779 1226 27789
rect 1192 27721 1226 27741
rect 1192 27707 1226 27721
rect 1192 27653 1226 27669
rect 1192 27635 1226 27653
rect 1192 27585 1226 27597
rect 1192 27563 1226 27585
rect 1192 27517 1226 27525
rect 1192 27491 1226 27517
rect 1192 27449 1226 27453
rect 1192 27419 1226 27449
rect 1192 27347 1226 27381
rect 1192 27279 1226 27309
rect 1192 27275 1226 27279
rect 1192 27211 1226 27237
rect 1192 27203 1226 27211
rect 1192 27143 1226 27165
rect 1192 27131 1226 27143
rect 1192 27075 1226 27093
rect 1192 27059 1226 27075
rect 1192 27007 1226 27021
rect 1192 26987 1226 27007
rect 1982 31023 2119 31345
rect 2119 31023 12897 31345
rect 12897 31023 13032 31345
rect 1726 30915 1976 30948
rect 1726 27481 1976 30915
rect 13031 30915 13281 30941
rect 1726 27458 1976 27481
rect 13031 27481 13281 30915
rect 13031 27451 13281 27481
rect 1985 27084 2119 27334
rect 2119 27084 12897 27334
rect 12897 27084 13035 27334
rect 13768 31406 13802 31412
rect 13768 31378 13802 31406
rect 1192 26939 1226 26949
rect 1192 26915 1226 26939
rect 1192 26871 1226 26877
rect 1192 26843 1226 26871
rect 1192 26803 1226 26805
rect 1192 26771 1226 26803
rect 1192 26701 1226 26733
rect 1192 26699 1226 26701
rect 1192 26633 1226 26661
rect 1192 26627 1226 26633
rect 1192 26565 1226 26589
rect 1192 26555 1226 26565
rect 1192 26497 1226 26517
rect 1192 26483 1226 26497
rect 1192 26429 1226 26445
rect 1192 26411 1226 26429
rect 1192 26361 1226 26373
rect 1192 26339 1226 26361
rect 1192 26293 1226 26301
rect 1192 26267 1226 26293
rect 1192 26225 1226 26229
rect 1192 26195 1226 26225
rect 1192 26123 1226 26157
rect 1192 26055 1226 26085
rect 1192 26051 1226 26055
rect 1192 25987 1226 26013
rect 1192 25979 1226 25987
rect 1192 25919 1226 25941
rect 1192 25907 1226 25919
rect 1192 25851 1226 25869
rect 1192 25835 1226 25851
rect 1192 25783 1226 25797
rect 1192 25763 1226 25783
rect 1192 25715 1226 25725
rect 1192 25691 1226 25715
rect 1192 25647 1226 25653
rect 1192 25619 1226 25647
rect 1192 25579 1226 25581
rect 1192 25547 1226 25579
rect 1192 25477 1226 25509
rect 1192 25475 1226 25477
rect 1192 25409 1226 25437
rect 1192 25403 1226 25409
rect 1192 25341 1226 25365
rect 1192 25331 1226 25341
rect 1192 25273 1226 25293
rect 1192 25259 1226 25273
rect 1192 25205 1226 25221
rect 1192 25187 1226 25205
rect 1192 25137 1226 25149
rect 1192 25115 1226 25137
rect 1192 25069 1226 25077
rect 1192 25043 1226 25069
rect 1192 25001 1226 25005
rect 1192 24971 1226 25001
rect 1192 24899 1226 24933
rect 1192 24831 1226 24861
rect 1192 24827 1226 24831
rect 1192 24763 1226 24789
rect 1192 24755 1226 24763
rect 1192 24695 1226 24717
rect 1192 24683 1226 24695
rect 1192 24627 1226 24645
rect 1192 24611 1226 24627
rect 1192 24559 1226 24573
rect 1192 24539 1226 24559
rect 1192 24491 1226 24501
rect 1192 24467 1226 24491
rect 1192 24423 1226 24429
rect 1192 24395 1226 24423
rect 1192 24355 1226 24357
rect 1192 24323 1226 24355
rect 1192 24253 1226 24285
rect 1192 24251 1226 24253
rect 1192 24185 1226 24213
rect 1192 24179 1226 24185
rect 1192 24117 1226 24141
rect 1192 24107 1226 24117
rect 1192 24049 1226 24069
rect 1192 24035 1226 24049
rect 1192 23981 1226 23997
rect 1192 23963 1226 23981
rect 1192 23913 1226 23925
rect 1192 23891 1226 23913
rect 1192 23845 1226 23853
rect 1192 23819 1226 23845
rect 1192 23777 1226 23781
rect 1192 23747 1226 23777
rect 1192 23675 1226 23709
rect 1192 23607 1226 23637
rect 1192 23603 1226 23607
rect 1192 23539 1226 23565
rect 1192 23531 1226 23539
rect 1192 23471 1226 23493
rect 1192 23459 1226 23471
rect 1192 23403 1226 23421
rect 1192 23387 1226 23403
rect 1192 23335 1226 23349
rect 1192 23315 1226 23335
rect 1192 23267 1226 23277
rect 1192 23243 1226 23267
rect 1192 23199 1226 23205
rect 1192 23171 1226 23199
rect 1192 23131 1226 23133
rect 1192 23099 1226 23131
rect 1192 23029 1226 23061
rect 1192 23027 1226 23029
rect 1192 22961 1226 22989
rect 1192 22955 1226 22961
rect 1192 22893 1226 22917
rect 1192 22883 1226 22893
rect 1192 22825 1226 22845
rect 1192 22811 1226 22825
rect 1192 22757 1226 22773
rect 1192 22739 1226 22757
rect 1192 22689 1226 22701
rect 1192 22667 1226 22689
rect 1192 22621 1226 22629
rect 1192 22595 1226 22621
rect 1192 22553 1226 22557
rect 1192 22523 1226 22553
rect 1192 22451 1226 22485
rect 1192 22383 1226 22413
rect 1192 22379 1226 22383
rect 1192 22315 1226 22341
rect 1192 22307 1226 22315
rect 1192 22247 1226 22269
rect 1192 22235 1226 22247
rect 1192 22179 1226 22197
rect 1192 22163 1226 22179
rect 1192 22111 1226 22125
rect 1192 22091 1226 22111
rect 1192 22043 1226 22053
rect 1192 22019 1226 22043
rect 1192 21975 1226 21981
rect 1192 21947 1226 21975
rect 1192 21907 1226 21909
rect 1192 21875 1226 21907
rect 1192 21805 1226 21837
rect 1192 21803 1226 21805
rect 1192 21737 1226 21765
rect 1192 21731 1226 21737
rect 1192 21669 1226 21693
rect 1192 21659 1226 21669
rect 1192 21601 1226 21621
rect 1192 21587 1226 21601
rect 1192 21533 1226 21549
rect 1192 21515 1226 21533
rect 1192 21465 1226 21477
rect 1192 21443 1226 21465
rect 1192 21397 1226 21405
rect 1192 21371 1226 21397
rect 1192 21329 1226 21333
rect 1192 21299 1226 21329
rect 1192 21227 1226 21261
rect 1192 21159 1226 21189
rect 1192 21155 1226 21159
rect 1192 21091 1226 21117
rect 1192 21083 1226 21091
rect 1192 21023 1226 21045
rect 1192 21011 1226 21023
rect 1192 20955 1226 20973
rect 1192 20939 1226 20955
rect 1192 20887 1226 20901
rect 1192 20867 1226 20887
rect 1192 20819 1226 20829
rect 1192 20795 1226 20819
rect 1192 20751 1226 20757
rect 1192 20723 1226 20751
rect 1192 20683 1226 20685
rect 1192 20651 1226 20683
rect 1192 20581 1226 20613
rect 1192 20579 1226 20581
rect 1192 20513 1226 20541
rect 1192 20507 1226 20513
rect 1192 20445 1226 20469
rect 1192 20435 1226 20445
rect 1192 20377 1226 20397
rect 1192 20363 1226 20377
rect 1192 20309 1226 20325
rect 1192 20291 1226 20309
rect 1192 20241 1226 20253
rect 1192 20219 1226 20241
rect 1192 20173 1226 20181
rect 1192 20147 1226 20173
rect 1192 20105 1226 20109
rect 1192 20075 1226 20105
rect 1192 20003 1226 20037
rect 1192 19935 1226 19965
rect 1192 19931 1226 19935
rect 1192 19867 1226 19893
rect 1192 19859 1226 19867
rect 1192 19799 1226 19821
rect 1192 19787 1226 19799
rect 1192 19731 1226 19749
rect 1192 19715 1226 19731
rect 1192 19663 1226 19677
rect 1192 19643 1226 19663
rect 1192 19595 1226 19605
rect 1192 19571 1226 19595
rect 1192 19527 1226 19533
rect 1192 19499 1226 19527
rect 1192 19459 1226 19461
rect 1192 19427 1226 19459
rect 1192 19357 1226 19389
rect 1192 19355 1226 19357
rect 1192 19289 1226 19317
rect 1192 19283 1226 19289
rect 1192 19221 1226 19245
rect 1192 19211 1226 19221
rect 1192 19153 1226 19173
rect 1192 19139 1226 19153
rect 1192 19085 1226 19101
rect 1192 19067 1226 19085
rect 1192 19017 1226 19029
rect 1192 18995 1226 19017
rect 1192 18949 1226 18957
rect 1192 18923 1226 18949
rect 1192 18881 1226 18885
rect 1192 18851 1226 18881
rect 1192 18779 1226 18813
rect 1192 18711 1226 18741
rect 1192 18707 1226 18711
rect 1192 18643 1226 18669
rect 1192 18635 1226 18643
rect 1192 18575 1226 18597
rect 1192 18563 1226 18575
rect 1192 18507 1226 18525
rect 1192 18491 1226 18507
rect 1192 18439 1226 18453
rect 1192 18419 1226 18439
rect 1192 18371 1226 18381
rect 1192 18347 1226 18371
rect 1192 18303 1226 18309
rect 1192 18275 1226 18303
rect 1192 18235 1226 18237
rect 1192 18203 1226 18235
rect 1192 18133 1226 18165
rect 1192 18131 1226 18133
rect 1192 18065 1226 18093
rect 1192 18059 1226 18065
rect 1192 17997 1226 18021
rect 1192 17987 1226 17997
rect 1192 17929 1226 17949
rect 1192 17915 1226 17929
rect 1192 17861 1226 17877
rect 1192 17843 1226 17861
rect 1192 17793 1226 17805
rect 1192 17771 1226 17793
rect 1192 17725 1226 17733
rect 1192 17699 1226 17725
rect 1192 17657 1226 17661
rect 1192 17627 1226 17657
rect 1192 17555 1226 17589
rect 1192 17487 1226 17517
rect 1192 17483 1226 17487
rect 1192 17419 1226 17445
rect 1192 17411 1226 17419
rect 1192 17351 1226 17373
rect 1192 17339 1226 17351
rect 1192 17283 1226 17301
rect 1192 17267 1226 17283
rect 1192 17215 1226 17229
rect 1192 17195 1226 17215
rect 1192 17147 1226 17157
rect 1192 17123 1226 17147
rect 1192 17079 1226 17085
rect 1192 17051 1226 17079
rect 1192 17011 1226 17013
rect 1192 16979 1226 17011
rect 1192 16909 1226 16941
rect 1192 16907 1226 16909
rect 1192 16841 1226 16869
rect 1192 16835 1226 16841
rect 1192 16773 1226 16797
rect 1192 16763 1226 16773
rect 1192 16705 1226 16725
rect 1192 16691 1226 16705
rect 1192 16637 1226 16653
rect 1192 16619 1226 16637
rect 1192 16569 1226 16581
rect 1192 16547 1226 16569
rect 1192 16501 1226 16509
rect 1192 16475 1226 16501
rect 1192 16433 1226 16437
rect 1192 16403 1226 16433
rect 1192 16331 1226 16365
rect 1192 16263 1226 16293
rect 1192 16259 1226 16263
rect 1192 16195 1226 16221
rect 1192 16187 1226 16195
rect 1192 16127 1226 16149
rect 1192 16115 1226 16127
rect 1192 16059 1226 16077
rect 1192 16043 1226 16059
rect 1192 15991 1226 16005
rect 1192 15971 1226 15991
rect 1192 15923 1226 15933
rect 1192 15899 1226 15923
rect 1192 15855 1226 15861
rect 1192 15827 1226 15855
rect 1192 15787 1226 15789
rect 1192 15755 1226 15787
rect 1192 15685 1226 15717
rect 1192 15683 1226 15685
rect 1192 15617 1226 15645
rect 1192 15611 1226 15617
rect 1192 15549 1226 15573
rect 1192 15539 1226 15549
rect 1192 15481 1226 15501
rect 1192 15467 1226 15481
rect 1192 15413 1226 15429
rect 1192 15395 1226 15413
rect 1192 15345 1226 15357
rect 1192 15323 1226 15345
rect 1192 15277 1226 15285
rect 1192 15251 1226 15277
rect 1192 15209 1226 15213
rect 1192 15179 1226 15209
rect 1192 15107 1226 15141
rect 1192 15039 1226 15069
rect 1192 15035 1226 15039
rect 1192 14971 1226 14997
rect 1192 14963 1226 14971
rect 1192 14903 1226 14925
rect 1192 14891 1226 14903
rect 1192 14835 1226 14853
rect 1192 14819 1226 14835
rect 1192 14767 1226 14781
rect 1192 14747 1226 14767
rect 1192 14699 1226 14709
rect 1192 14675 1226 14699
rect 1192 14631 1226 14637
rect 1192 14603 1226 14631
rect 1192 14563 1226 14565
rect 1192 14531 1226 14563
rect 1192 14461 1226 14493
rect 1192 14459 1226 14461
rect 1192 14393 1226 14421
rect 1192 14387 1226 14393
rect 1192 14325 1226 14349
rect 1192 14315 1226 14325
rect 1192 14257 1226 14277
rect 1192 14243 1226 14257
rect 1192 14189 1226 14205
rect 1192 14171 1226 14189
rect 1192 14121 1226 14133
rect 1192 14099 1226 14121
rect 1192 14053 1226 14061
rect 1192 14027 1226 14053
rect 1192 13985 1226 13989
rect 1192 13955 1226 13985
rect 1192 13883 1226 13917
rect 1192 13815 1226 13845
rect 1192 13811 1226 13815
rect 1192 13747 1226 13773
rect 1192 13739 1226 13747
rect 1192 13679 1226 13701
rect 1192 13667 1226 13679
rect 1192 13611 1226 13629
rect 1192 13595 1226 13611
rect 1192 13543 1226 13557
rect 1192 13523 1226 13543
rect 1192 13475 1226 13485
rect 1192 13451 1226 13475
rect 1192 13407 1226 13413
rect 1192 13379 1226 13407
rect 1192 13339 1226 13341
rect 1192 13307 1226 13339
rect 1192 13237 1226 13269
rect 1192 13235 1226 13237
rect 1192 13169 1226 13197
rect 1192 13163 1226 13169
rect 1192 13101 1226 13125
rect 1192 13091 1226 13101
rect 1192 13033 1226 13053
rect 1192 13019 1226 13033
rect 1192 12965 1226 12981
rect 1192 12947 1226 12965
rect 1192 12897 1226 12909
rect 1192 12875 1226 12897
rect 1192 12829 1226 12837
rect 1192 12803 1226 12829
rect 1192 12761 1226 12765
rect 1192 12731 1226 12761
rect 1192 12659 1226 12693
rect 1192 12591 1226 12621
rect 1192 12587 1226 12591
rect 1192 12523 1226 12549
rect 1192 12515 1226 12523
rect 1192 12455 1226 12477
rect 1192 12443 1226 12455
rect 1192 12387 1226 12405
rect 1192 12371 1226 12387
rect 1192 12319 1226 12333
rect 1192 12299 1226 12319
rect 1192 12251 1226 12261
rect 1192 12227 1226 12251
rect 1192 12183 1226 12189
rect 1192 12155 1226 12183
rect 1192 12115 1226 12117
rect 1192 12083 1226 12115
rect 1192 12013 1226 12045
rect 1192 12011 1226 12013
rect 1192 11945 1226 11973
rect 1192 11939 1226 11945
rect 1192 11877 1226 11901
rect 1192 11867 1226 11877
rect 1192 11809 1226 11829
rect 1192 11795 1226 11809
rect 1192 11741 1226 11757
rect 1192 11723 1226 11741
rect 1192 11673 1226 11685
rect 1192 11651 1226 11673
rect 1192 11605 1226 11613
rect 1192 11579 1226 11605
rect 1192 11537 1226 11541
rect 1192 11507 1226 11537
rect 1192 11435 1226 11469
rect 1192 11367 1226 11397
rect 1192 11363 1226 11367
rect 1192 11299 1226 11325
rect 1192 11291 1226 11299
rect 1192 11231 1226 11253
rect 1192 11219 1226 11231
rect 1192 11163 1226 11181
rect 1192 11147 1226 11163
rect 1192 11095 1226 11109
rect 1192 11075 1226 11095
rect 1192 11027 1226 11037
rect 1192 11003 1226 11027
rect 1192 10959 1226 10965
rect 1192 10931 1226 10959
rect 1192 10891 1226 10893
rect 1192 10859 1226 10891
rect 1192 10789 1226 10821
rect 1192 10787 1226 10789
rect 1192 10721 1226 10749
rect 1192 10715 1226 10721
rect 1192 10653 1226 10677
rect 1192 10643 1226 10653
rect 1192 10585 1226 10605
rect 1192 10571 1226 10585
rect 1192 10517 1226 10533
rect 1192 10499 1226 10517
rect 1192 10449 1226 10461
rect 1192 10427 1226 10449
rect 13768 21206 13802 21219
rect 13768 21185 13802 21206
rect 13768 21138 13802 21147
rect 13768 21113 13802 21138
rect 13768 21070 13802 21075
rect 13768 21041 13802 21070
rect 13768 21002 13802 21003
rect 13768 20969 13802 21002
rect 13768 20900 13802 20931
rect 13768 20897 13802 20900
rect 13768 20832 13802 20859
rect 13768 20825 13802 20832
rect 13768 20764 13802 20787
rect 13768 20753 13802 20764
rect 13768 20696 13802 20715
rect 13768 20681 13802 20696
rect 13768 20628 13802 20643
rect 13768 20609 13802 20628
rect 13768 20560 13802 20571
rect 13768 20537 13802 20560
rect 13768 20492 13802 20499
rect 13768 20465 13802 20492
rect 13768 20424 13802 20427
rect 13768 20393 13802 20424
rect 13768 20322 13802 20355
rect 13768 20321 13802 20322
rect 13768 20254 13802 20283
rect 13768 20249 13802 20254
rect 13768 20186 13802 20211
rect 13768 20177 13802 20186
rect 13768 20118 13802 20139
rect 13768 20105 13802 20118
rect 13768 20050 13802 20067
rect 13768 20033 13802 20050
rect 13768 19982 13802 19995
rect 13768 19961 13802 19982
rect 13768 19914 13802 19923
rect 13768 19889 13802 19914
rect 13768 19846 13802 19851
rect 13768 19817 13802 19846
rect 13768 19778 13802 19779
rect 13768 19745 13802 19778
rect 13768 19676 13802 19707
rect 13768 19673 13802 19676
rect 13768 19608 13802 19635
rect 13768 19601 13802 19608
rect 13768 19540 13802 19563
rect 13768 19529 13802 19540
rect 13768 19472 13802 19491
rect 13768 19457 13802 19472
rect 13768 19404 13802 19419
rect 13768 19385 13802 19404
rect 13768 19336 13802 19347
rect 13768 19313 13802 19336
rect 13768 19268 13802 19275
rect 13768 19241 13802 19268
rect 13768 19200 13802 19203
rect 13768 19169 13802 19200
rect 13768 19098 13802 19131
rect 13768 19097 13802 19098
rect 13768 19030 13802 19059
rect 13768 19025 13802 19030
rect 13768 18962 13802 18987
rect 13768 18953 13802 18962
rect 13768 18894 13802 18915
rect 13768 18881 13802 18894
rect 13768 18826 13802 18843
rect 13768 18809 13802 18826
rect 13768 18758 13802 18771
rect 13768 18737 13802 18758
rect 13768 18690 13802 18699
rect 13768 18665 13802 18690
rect 13768 18622 13802 18627
rect 13768 18593 13802 18622
rect 13768 18554 13802 18555
rect 13768 18521 13802 18554
rect 13768 18452 13802 18483
rect 13768 18449 13802 18452
rect 13768 18384 13802 18411
rect 13768 18377 13802 18384
rect 13768 18316 13802 18339
rect 13768 18305 13802 18316
rect 13768 18248 13802 18267
rect 13768 18233 13802 18248
rect 13768 18180 13802 18195
rect 13768 18161 13802 18180
rect 13768 18112 13802 18123
rect 13768 18089 13802 18112
rect 13768 18044 13802 18051
rect 13768 18017 13802 18044
rect 13768 17976 13802 17979
rect 13768 17945 13802 17976
rect 13768 17874 13802 17907
rect 13768 17873 13802 17874
rect 13768 17806 13802 17835
rect 13768 17801 13802 17806
rect 13768 17738 13802 17763
rect 13768 17729 13802 17738
rect 13768 17670 13802 17691
rect 13768 17657 13802 17670
rect 13768 17602 13802 17619
rect 13768 17585 13802 17602
rect 13768 17534 13802 17547
rect 13768 17513 13802 17534
rect 13768 17466 13802 17475
rect 13768 17441 13802 17466
rect 13768 17398 13802 17403
rect 13768 17369 13802 17398
rect 13768 17330 13802 17331
rect 13768 17297 13802 17330
rect 13768 17228 13802 17259
rect 13768 17225 13802 17228
rect 13768 17160 13802 17187
rect 13768 17153 13802 17160
rect 13768 17092 13802 17115
rect 13768 17081 13802 17092
rect 13768 17024 13802 17043
rect 13768 17009 13802 17024
rect 13768 16956 13802 16971
rect 13768 16937 13802 16956
rect 13768 16888 13802 16899
rect 13768 16865 13802 16888
rect 13768 16820 13802 16827
rect 13768 16793 13802 16820
rect 13768 16752 13802 16755
rect 13768 16721 13802 16752
rect 13768 16650 13802 16683
rect 13768 16649 13802 16650
rect 13768 16582 13802 16611
rect 13768 16577 13802 16582
rect 13768 16514 13802 16539
rect 13768 16505 13802 16514
rect 13768 16446 13802 16467
rect 13768 16433 13802 16446
rect 13768 16378 13802 16395
rect 13768 16361 13802 16378
rect 13768 16310 13802 16323
rect 13768 16289 13802 16310
rect 13768 16242 13802 16251
rect 13768 16217 13802 16242
rect 13768 16174 13802 16179
rect 13768 16145 13802 16174
rect 13768 16106 13802 16107
rect 13768 16073 13802 16106
rect 13768 16004 13802 16035
rect 13768 16001 13802 16004
rect 13768 15936 13802 15963
rect 13768 15929 13802 15936
rect 13768 15868 13802 15891
rect 13768 15857 13802 15868
rect 13768 15800 13802 15819
rect 13768 15785 13802 15800
rect 13768 15732 13802 15747
rect 13768 15713 13802 15732
rect 13768 15664 13802 15675
rect 13768 15641 13802 15664
rect 13768 15596 13802 15603
rect 13768 15569 13802 15596
rect 13768 15528 13802 15531
rect 13768 15497 13802 15528
rect 13768 15426 13802 15459
rect 13768 15425 13802 15426
rect 13768 15358 13802 15387
rect 13768 15353 13802 15358
rect 13768 15290 13802 15315
rect 13768 15281 13802 15290
rect 13768 15222 13802 15243
rect 13768 15209 13802 15222
rect 13768 15154 13802 15171
rect 13768 15137 13802 15154
rect 13768 15086 13802 15099
rect 13768 15065 13802 15086
rect 13768 15018 13802 15027
rect 13768 14993 13802 15018
rect 13768 14950 13802 14955
rect 13768 14921 13802 14950
rect 13768 14882 13802 14883
rect 13768 14849 13802 14882
rect 13768 14780 13802 14811
rect 13768 14777 13802 14780
rect 13768 14712 13802 14739
rect 13768 14705 13802 14712
rect 13768 14644 13802 14667
rect 13768 14633 13802 14644
rect 13768 14576 13802 14595
rect 13768 14561 13802 14576
rect 13768 14508 13802 14523
rect 13768 14489 13802 14508
rect 13768 14440 13802 14451
rect 13768 14417 13802 14440
rect 13768 14372 13802 14379
rect 13768 14345 13802 14372
rect 13768 14304 13802 14307
rect 13768 14273 13802 14304
rect 13768 14202 13802 14235
rect 13768 14201 13802 14202
rect 13768 14134 13802 14163
rect 13768 14129 13802 14134
rect 13768 14066 13802 14091
rect 13768 14057 13802 14066
rect 13768 13998 13802 14019
rect 13768 13985 13802 13998
rect 13768 13930 13802 13947
rect 13768 13913 13802 13930
rect 13768 13862 13802 13875
rect 13768 13841 13802 13862
rect 13768 13794 13802 13803
rect 13768 13769 13802 13794
rect 13768 13726 13802 13731
rect 13768 13697 13802 13726
rect 13768 13658 13802 13659
rect 13768 13625 13802 13658
rect 13768 13556 13802 13587
rect 13768 13553 13802 13556
rect 13768 13488 13802 13515
rect 13768 13481 13802 13488
rect 13768 13420 13802 13443
rect 13768 13409 13802 13420
rect 13768 13352 13802 13371
rect 13768 13337 13802 13352
rect 13768 13284 13802 13299
rect 13768 13265 13802 13284
rect 13768 13216 13802 13227
rect 13768 13193 13802 13216
rect 13768 13148 13802 13155
rect 13768 13121 13802 13148
rect 13768 13080 13802 13083
rect 13768 13049 13802 13080
rect 13768 12978 13802 13011
rect 13768 12977 13802 12978
rect 13768 12910 13802 12939
rect 13768 12905 13802 12910
rect 13768 12842 13802 12867
rect 13768 12833 13802 12842
rect 13768 12774 13802 12795
rect 13768 12761 13802 12774
rect 13768 12706 13802 12723
rect 13768 12689 13802 12706
rect 13768 12638 13802 12651
rect 13768 12617 13802 12638
rect 13768 12570 13802 12579
rect 13768 12545 13802 12570
rect 13768 12502 13802 12507
rect 13768 12473 13802 12502
rect 13768 12434 13802 12435
rect 13768 12401 13802 12434
rect 13768 12332 13802 12363
rect 13768 12329 13802 12332
rect 13768 12264 13802 12291
rect 13768 12257 13802 12264
rect 13768 12196 13802 12219
rect 13768 12185 13802 12196
rect 13768 12128 13802 12147
rect 13768 12113 13802 12128
rect 13768 12060 13802 12075
rect 13768 12041 13802 12060
rect 13768 11992 13802 12003
rect 13768 11969 13802 11992
rect 13768 11924 13802 11931
rect 13768 11897 13802 11924
rect 13768 11856 13802 11859
rect 13768 11825 13802 11856
rect 13768 11754 13802 11787
rect 13768 11753 13802 11754
rect 13768 11686 13802 11715
rect 13768 11681 13802 11686
rect 13768 11618 13802 11643
rect 13768 11609 13802 11618
rect 13768 11550 13802 11571
rect 13768 11537 13802 11550
rect 13768 11482 13802 11499
rect 13768 11465 13802 11482
rect 13768 11414 13802 11427
rect 13768 11393 13802 11414
rect 13768 11346 13802 11355
rect 13768 11321 13802 11346
rect 13768 11278 13802 11283
rect 13768 11249 13802 11278
rect 13768 11210 13802 11211
rect 13768 11177 13802 11210
rect 13768 11108 13802 11139
rect 13768 11105 13802 11108
rect 13768 11040 13802 11067
rect 13768 11033 13802 11040
rect 13768 10972 13802 10995
rect 13768 10961 13802 10972
rect 13768 10904 13802 10923
rect 13768 10889 13802 10904
rect 13768 10836 13802 10851
rect 13768 10817 13802 10836
rect 13768 10768 13802 10779
rect 13768 10745 13802 10768
rect 13768 10700 13802 10707
rect 13768 10673 13802 10700
rect 13768 10632 13802 10635
rect 13768 10601 13802 10632
rect 13768 10530 13802 10563
rect 13768 10529 13802 10530
rect 13768 10462 13802 10491
rect 13768 10457 13802 10462
rect 13768 10394 13802 10419
rect 13768 10385 13802 10394
rect 1327 10284 1329 10318
rect 1329 10284 1361 10318
rect 1399 10284 1431 10318
rect 1431 10284 1433 10318
rect 1471 10284 1499 10318
rect 1499 10284 1505 10318
rect 1543 10284 1567 10318
rect 1567 10284 1577 10318
rect 1615 10284 1635 10318
rect 1635 10284 1649 10318
rect 1687 10284 1703 10318
rect 1703 10284 1721 10318
rect 1759 10284 1771 10318
rect 1771 10284 1793 10318
rect 1831 10284 1839 10318
rect 1839 10284 1865 10318
rect 1903 10284 1907 10318
rect 1907 10284 1937 10318
rect 1975 10284 2009 10318
rect 2047 10284 2077 10318
rect 2077 10284 2081 10318
rect 2119 10284 2145 10318
rect 2145 10284 2153 10318
rect 2191 10284 2213 10318
rect 2213 10284 2225 10318
rect 2263 10284 2281 10318
rect 2281 10284 2297 10318
rect 2335 10284 2349 10318
rect 2349 10284 2369 10318
rect 2407 10284 2417 10318
rect 2417 10284 2441 10318
rect 2479 10284 2485 10318
rect 2485 10284 2513 10318
rect 2551 10284 2553 10318
rect 2553 10284 2585 10318
rect 2623 10284 2655 10318
rect 2655 10284 2657 10318
rect 2695 10284 2723 10318
rect 2723 10284 2729 10318
rect 2767 10284 2791 10318
rect 2791 10284 2801 10318
rect 2839 10284 2859 10318
rect 2859 10284 2873 10318
rect 2911 10284 2927 10318
rect 2927 10284 2945 10318
rect 2983 10284 2995 10318
rect 2995 10284 3017 10318
rect 3055 10284 3063 10318
rect 3063 10284 3089 10318
rect 3127 10284 3131 10318
rect 3131 10284 3161 10318
rect 3199 10284 3233 10318
rect 3271 10284 3301 10318
rect 3301 10284 3305 10318
rect 3343 10284 3369 10318
rect 3369 10284 3377 10318
rect 3415 10284 3437 10318
rect 3437 10284 3449 10318
rect 3487 10284 3505 10318
rect 3505 10284 3521 10318
rect 3559 10284 3573 10318
rect 3573 10284 3593 10318
rect 3631 10284 3641 10318
rect 3641 10284 3665 10318
rect 3703 10284 3709 10318
rect 3709 10284 3737 10318
rect 3775 10284 3777 10318
rect 3777 10284 3809 10318
rect 3847 10284 3879 10318
rect 3879 10284 3881 10318
rect 3919 10284 3947 10318
rect 3947 10284 3953 10318
rect 3991 10284 4015 10318
rect 4015 10284 4025 10318
rect 4063 10284 4083 10318
rect 4083 10284 4097 10318
rect 4135 10284 4151 10318
rect 4151 10284 4169 10318
rect 4207 10284 4219 10318
rect 4219 10284 4241 10318
rect 4279 10284 4287 10318
rect 4287 10284 4313 10318
rect 4351 10284 4355 10318
rect 4355 10284 4385 10318
rect 4423 10284 4457 10318
rect 4495 10284 4525 10318
rect 4525 10284 4529 10318
rect 4567 10284 4593 10318
rect 4593 10284 4601 10318
rect 4639 10284 4661 10318
rect 4661 10284 4673 10318
rect 4711 10284 4729 10318
rect 4729 10284 4745 10318
rect 4783 10284 4797 10318
rect 4797 10284 4817 10318
rect 4855 10284 4865 10318
rect 4865 10284 4889 10318
rect 4927 10284 4933 10318
rect 4933 10284 4961 10318
rect 4999 10284 5001 10318
rect 5001 10284 5033 10318
rect 5071 10284 5103 10318
rect 5103 10284 5105 10318
rect 5143 10284 5171 10318
rect 5171 10284 5177 10318
rect 5215 10284 5239 10318
rect 5239 10284 5249 10318
rect 5287 10284 5307 10318
rect 5307 10284 5321 10318
rect 5359 10284 5375 10318
rect 5375 10284 5393 10318
rect 5431 10284 5443 10318
rect 5443 10284 5465 10318
rect 5503 10284 5511 10318
rect 5511 10284 5537 10318
rect 5575 10284 5579 10318
rect 5579 10284 5609 10318
rect 5647 10284 5681 10318
rect 5719 10284 5749 10318
rect 5749 10284 5753 10318
rect 5791 10284 5817 10318
rect 5817 10284 5825 10318
rect 5863 10284 5885 10318
rect 5885 10284 5897 10318
rect 5935 10284 5953 10318
rect 5953 10284 5969 10318
rect 6007 10284 6021 10318
rect 6021 10284 6041 10318
rect 6079 10284 6089 10318
rect 6089 10284 6113 10318
rect 6151 10284 6157 10318
rect 6157 10284 6185 10318
rect 6223 10284 6225 10318
rect 6225 10284 6257 10318
rect 6295 10284 6327 10318
rect 6327 10284 6329 10318
rect 6367 10284 6395 10318
rect 6395 10284 6401 10318
rect 6439 10284 6463 10318
rect 6463 10284 6473 10318
rect 6511 10284 6531 10318
rect 6531 10284 6545 10318
rect 6583 10284 6599 10318
rect 6599 10284 6617 10318
rect 6655 10284 6667 10318
rect 6667 10284 6689 10318
rect 6727 10284 6735 10318
rect 6735 10284 6761 10318
rect 6799 10284 6803 10318
rect 6803 10284 6833 10318
rect 6871 10284 6905 10318
rect 6943 10284 6973 10318
rect 6973 10284 6977 10318
rect 7015 10284 7041 10318
rect 7041 10284 7049 10318
rect 7087 10284 7109 10318
rect 7109 10284 7121 10318
rect 7159 10284 7177 10318
rect 7177 10284 7193 10318
rect 7231 10284 7245 10318
rect 7245 10284 7265 10318
rect 7303 10284 7313 10318
rect 7313 10284 7337 10318
rect 7375 10284 7381 10318
rect 7381 10284 7409 10318
rect 7447 10284 7449 10318
rect 7449 10284 7481 10318
rect 7519 10284 7551 10318
rect 7551 10284 7553 10318
rect 7591 10284 7619 10318
rect 7619 10284 7625 10318
rect 7663 10284 7687 10318
rect 7687 10284 7697 10318
rect 7735 10284 7755 10318
rect 7755 10284 7769 10318
rect 7807 10284 7823 10318
rect 7823 10284 7841 10318
rect 7879 10284 7891 10318
rect 7891 10284 7913 10318
rect 7951 10284 7959 10318
rect 7959 10284 7985 10318
rect 8023 10284 8027 10318
rect 8027 10284 8057 10318
rect 8095 10284 8129 10318
rect 8167 10284 8197 10318
rect 8197 10284 8201 10318
rect 8239 10284 8265 10318
rect 8265 10284 8273 10318
rect 8311 10284 8333 10318
rect 8333 10284 8345 10318
rect 8383 10284 8401 10318
rect 8401 10284 8417 10318
rect 8455 10284 8469 10318
rect 8469 10284 8489 10318
rect 8527 10284 8537 10318
rect 8537 10284 8561 10318
rect 8599 10284 8605 10318
rect 8605 10284 8633 10318
rect 8671 10284 8673 10318
rect 8673 10284 8705 10318
rect 8743 10284 8775 10318
rect 8775 10284 8777 10318
rect 8815 10284 8843 10318
rect 8843 10284 8849 10318
rect 8887 10284 8911 10318
rect 8911 10284 8921 10318
rect 8959 10284 8979 10318
rect 8979 10284 8993 10318
rect 9031 10284 9047 10318
rect 9047 10284 9065 10318
rect 9103 10284 9115 10318
rect 9115 10284 9137 10318
rect 9175 10284 9183 10318
rect 9183 10284 9209 10318
rect 9247 10284 9251 10318
rect 9251 10284 9281 10318
rect 9319 10284 9353 10318
rect 9391 10284 9421 10318
rect 9421 10284 9425 10318
rect 9463 10284 9489 10318
rect 9489 10284 9497 10318
rect 9535 10284 9557 10318
rect 9557 10284 9569 10318
rect 9607 10284 9625 10318
rect 9625 10284 9641 10318
rect 9679 10284 9693 10318
rect 9693 10284 9713 10318
rect 9751 10284 9761 10318
rect 9761 10284 9785 10318
rect 9823 10284 9829 10318
rect 9829 10284 9857 10318
rect 9895 10284 9897 10318
rect 9897 10284 9929 10318
rect 9967 10284 9999 10318
rect 9999 10284 10001 10318
rect 10039 10284 10067 10318
rect 10067 10284 10073 10318
rect 10111 10284 10135 10318
rect 10135 10284 10145 10318
rect 10183 10284 10203 10318
rect 10203 10284 10217 10318
rect 10255 10284 10271 10318
rect 10271 10284 10289 10318
rect 10327 10284 10339 10318
rect 10339 10284 10361 10318
rect 10399 10284 10407 10318
rect 10407 10284 10433 10318
rect 10471 10284 10475 10318
rect 10475 10284 10505 10318
rect 10543 10284 10577 10318
rect 10615 10284 10645 10318
rect 10645 10284 10649 10318
rect 10687 10284 10713 10318
rect 10713 10284 10721 10318
rect 10759 10284 10781 10318
rect 10781 10284 10793 10318
rect 10831 10284 10849 10318
rect 10849 10284 10865 10318
rect 10903 10284 10917 10318
rect 10917 10284 10937 10318
rect 10975 10284 10985 10318
rect 10985 10284 11009 10318
rect 11047 10284 11053 10318
rect 11053 10284 11081 10318
rect 11119 10284 11121 10318
rect 11121 10284 11153 10318
rect 11191 10284 11223 10318
rect 11223 10284 11225 10318
rect 11263 10284 11291 10318
rect 11291 10284 11297 10318
rect 11335 10284 11359 10318
rect 11359 10284 11369 10318
rect 11407 10284 11427 10318
rect 11427 10284 11441 10318
rect 11479 10284 11495 10318
rect 11495 10284 11513 10318
rect 11551 10284 11563 10318
rect 11563 10284 11585 10318
rect 11623 10284 11631 10318
rect 11631 10284 11657 10318
rect 11695 10284 11699 10318
rect 11699 10284 11729 10318
rect 11767 10284 11801 10318
rect 11839 10284 11869 10318
rect 11869 10284 11873 10318
rect 11911 10284 11937 10318
rect 11937 10284 11945 10318
rect 11983 10284 12005 10318
rect 12005 10284 12017 10318
rect 12055 10284 12073 10318
rect 12073 10284 12089 10318
rect 12127 10284 12141 10318
rect 12141 10284 12161 10318
rect 12199 10284 12209 10318
rect 12209 10284 12233 10318
rect 12271 10284 12277 10318
rect 12277 10284 12305 10318
rect 12343 10284 12345 10318
rect 12345 10284 12377 10318
rect 12415 10284 12447 10318
rect 12447 10284 12449 10318
rect 12487 10284 12515 10318
rect 12515 10284 12521 10318
rect 12559 10284 12583 10318
rect 12583 10284 12593 10318
rect 12631 10284 12651 10318
rect 12651 10284 12665 10318
rect 12703 10284 12719 10318
rect 12719 10284 12737 10318
rect 12775 10284 12787 10318
rect 12787 10284 12809 10318
rect 12847 10284 12855 10318
rect 12855 10284 12881 10318
rect 12919 10284 12923 10318
rect 12923 10284 12953 10318
rect 12991 10284 13025 10318
rect 13063 10284 13093 10318
rect 13093 10284 13097 10318
rect 13135 10284 13161 10318
rect 13161 10284 13169 10318
rect 13207 10284 13229 10318
rect 13229 10284 13241 10318
rect 13279 10284 13297 10318
rect 13297 10284 13313 10318
rect 13351 10284 13365 10318
rect 13365 10284 13385 10318
rect 13423 10284 13433 10318
rect 13433 10284 13457 10318
rect 13495 10284 13501 10318
rect 13501 10284 13529 10318
rect 13567 10284 13569 10318
rect 13569 10284 13601 10318
rect 13639 10284 13671 10318
rect 13671 10284 13673 10318
rect 14142 34691 14176 34725
rect 14142 34619 14176 34653
rect 14142 34547 14176 34581
rect 14142 34475 14176 34509
rect 14142 34403 14176 34437
rect 14142 34331 14176 34365
rect 14142 34259 14176 34293
rect 14142 34187 14176 34221
rect 14142 34115 14176 34149
rect 14142 34043 14176 34077
rect 14142 33971 14176 34005
rect 14142 33899 14176 33933
rect 14142 33827 14176 33861
rect 14142 33755 14176 33789
rect 14142 33683 14176 33717
rect 14142 33611 14176 33645
rect 14142 33539 14176 33573
rect 14142 33467 14176 33501
rect 14142 33395 14176 33429
rect 14142 33323 14176 33357
rect 14142 33251 14176 33285
rect 14142 33179 14176 33213
rect 14142 33107 14176 33141
rect 14142 33035 14176 33069
rect 14142 32963 14176 32997
rect 14142 32891 14176 32925
rect 14142 32819 14176 32853
rect 14142 32747 14176 32781
rect 14142 32675 14176 32709
rect 14142 32603 14176 32637
rect 14142 32531 14176 32565
rect 14142 32459 14176 32493
rect 14142 32387 14176 32421
rect 14142 32315 14176 32349
rect 14142 32243 14176 32277
rect 14142 32171 14176 32205
rect 14142 32099 14176 32133
rect 14142 32027 14176 32061
rect 14142 31955 14176 31989
rect 14142 31883 14176 31917
rect 14142 31811 14176 31845
rect 14142 31739 14176 31773
rect 14142 31667 14176 31701
rect 14142 31595 14176 31629
rect 14142 31523 14176 31557
rect 14142 31451 14176 31485
rect 14142 31379 14176 31413
rect 14142 31307 14176 31341
rect 14142 31235 14176 31269
rect 14142 31163 14176 31197
rect 14142 31091 14176 31125
rect 14142 31019 14176 31053
rect 14142 30947 14176 30981
rect 14142 30875 14176 30909
rect 14142 30803 14176 30837
rect 14142 30731 14176 30765
rect 14142 30659 14176 30693
rect 14142 30587 14176 30621
rect 14142 30515 14176 30549
rect 14142 30443 14176 30477
rect 14142 30371 14176 30405
rect 14142 30299 14176 30333
rect 14142 30227 14176 30261
rect 14142 30155 14176 30189
rect 14142 30083 14176 30117
rect 14142 30011 14176 30045
rect 14142 29939 14176 29973
rect 14142 29867 14176 29901
rect 14142 29795 14176 29829
rect 14142 29723 14176 29757
rect 14142 29651 14176 29685
rect 14142 29579 14176 29613
rect 14142 29507 14176 29541
rect 14142 29435 14176 29469
rect 14142 29363 14176 29397
rect 14142 29291 14176 29325
rect 14142 29219 14176 29253
rect 14142 29147 14176 29181
rect 14142 29075 14176 29109
rect 14142 29003 14176 29037
rect 14142 28931 14176 28965
rect 14142 28859 14176 28893
rect 14142 28787 14176 28821
rect 14142 28715 14176 28749
rect 14142 28643 14176 28677
rect 14142 28571 14176 28605
rect 14142 28499 14176 28533
rect 14142 28427 14176 28461
rect 14142 28355 14176 28389
rect 14142 28283 14176 28317
rect 14142 28211 14176 28245
rect 14142 28139 14176 28173
rect 14142 28067 14176 28101
rect 14142 27995 14176 28029
rect 14142 27923 14176 27957
rect 14142 27851 14176 27885
rect 14142 27779 14176 27813
rect 14142 27707 14176 27741
rect 14142 27635 14176 27669
rect 14142 27563 14176 27597
rect 14142 27491 14176 27525
rect 14142 27419 14176 27453
rect 14142 27347 14176 27381
rect 14142 27275 14176 27309
rect 14142 27203 14176 27237
rect 14142 27131 14176 27165
rect 14142 27059 14176 27093
rect 14142 26987 14176 27021
rect 14142 26915 14176 26949
rect 14142 26843 14176 26877
rect 14142 26771 14176 26805
rect 14142 26699 14176 26733
rect 14142 26627 14176 26661
rect 14142 26555 14176 26589
rect 14142 26483 14176 26517
rect 14142 26411 14176 26445
rect 14142 26339 14176 26373
rect 14142 26267 14176 26301
rect 14142 26195 14176 26229
rect 14142 26123 14176 26157
rect 14142 26051 14176 26085
rect 14142 25979 14176 26013
rect 14142 25907 14176 25941
rect 14142 25835 14176 25869
rect 14142 25763 14176 25797
rect 14142 25691 14176 25725
rect 14142 25619 14176 25653
rect 14142 25547 14176 25581
rect 14142 25475 14176 25509
rect 14142 25403 14176 25437
rect 14142 25331 14176 25365
rect 14142 25259 14176 25293
rect 14142 25187 14176 25221
rect 14142 25115 14176 25149
rect 14142 25043 14176 25077
rect 14142 24971 14176 25005
rect 14142 24899 14176 24933
rect 14142 24827 14176 24861
rect 14142 24755 14176 24789
rect 14142 24683 14176 24717
rect 14142 24611 14176 24645
rect 14142 24539 14176 24573
rect 14142 24467 14176 24501
rect 14142 24395 14176 24429
rect 14142 24323 14176 24357
rect 14142 24251 14176 24285
rect 14142 24179 14176 24213
rect 14142 24107 14176 24141
rect 14142 24035 14176 24069
rect 14142 23963 14176 23997
rect 14142 23891 14176 23925
rect 14142 23819 14176 23853
rect 14142 23747 14176 23781
rect 14142 23675 14176 23709
rect 14142 23603 14176 23637
rect 14142 23531 14176 23565
rect 14142 23459 14176 23493
rect 14142 23387 14176 23421
rect 14142 23315 14176 23349
rect 14142 23243 14176 23277
rect 14142 23171 14176 23205
rect 14142 23099 14176 23133
rect 14142 23027 14176 23061
rect 14142 22955 14176 22989
rect 14142 22883 14176 22917
rect 14142 22811 14176 22845
rect 14142 22739 14176 22773
rect 14142 22667 14176 22701
rect 14142 22595 14176 22629
rect 14142 22523 14176 22557
rect 14142 22451 14176 22485
rect 14142 22379 14176 22413
rect 14142 22307 14176 22341
rect 14142 22235 14176 22269
rect 14142 22163 14176 22197
rect 14142 22091 14176 22125
rect 14142 22019 14176 22053
rect 14142 21947 14176 21981
rect 14142 21875 14176 21909
rect 14142 21803 14176 21837
rect 14142 21731 14176 21765
rect 14142 21659 14176 21693
rect 14142 21587 14176 21621
rect 14142 21515 14176 21549
rect 14142 21443 14176 21477
rect 14142 21371 14176 21405
rect 14142 21299 14176 21333
rect 14142 21227 14176 21261
rect 14142 21155 14176 21189
rect 14142 21083 14176 21117
rect 14142 21011 14176 21045
rect 14142 20939 14176 20973
rect 14142 20867 14176 20901
rect 14142 20795 14176 20829
rect 14142 20723 14176 20757
rect 14142 20651 14176 20685
rect 14142 20579 14176 20613
rect 14142 20507 14176 20541
rect 14142 20435 14176 20469
rect 14142 20363 14176 20397
rect 14142 20291 14176 20325
rect 14142 20219 14176 20253
rect 14142 20147 14176 20181
rect 14142 20075 14176 20109
rect 14142 20003 14176 20037
rect 14142 19931 14176 19965
rect 14142 19859 14176 19893
rect 14142 19787 14176 19821
rect 14142 19715 14176 19749
rect 14142 19643 14176 19677
rect 14142 19571 14176 19605
rect 14142 19499 14176 19533
rect 14142 19427 14176 19461
rect 14142 19355 14176 19389
rect 14142 19283 14176 19317
rect 14142 19211 14176 19245
rect 14142 19139 14176 19173
rect 14142 19067 14176 19101
rect 14142 18995 14176 19029
rect 14142 18923 14176 18957
rect 14142 18851 14176 18885
rect 14142 18779 14176 18813
rect 14142 18707 14176 18741
rect 14142 18635 14176 18669
rect 14142 18563 14176 18597
rect 14142 18491 14176 18525
rect 14142 18419 14176 18453
rect 14142 18347 14176 18381
rect 14142 18275 14176 18309
rect 14142 18203 14176 18237
rect 14142 18131 14176 18165
rect 14142 18059 14176 18093
rect 14142 17987 14176 18021
rect 14142 17915 14176 17949
rect 14142 17843 14176 17877
rect 14142 17771 14176 17805
rect 14142 17699 14176 17733
rect 14142 17627 14176 17661
rect 14142 17555 14176 17589
rect 14142 17483 14176 17517
rect 14142 17411 14176 17445
rect 14142 17339 14176 17373
rect 14142 17267 14176 17301
rect 14142 17195 14176 17229
rect 14142 17123 14176 17157
rect 14142 17051 14176 17085
rect 14142 16979 14176 17013
rect 14142 16907 14176 16941
rect 14142 16835 14176 16869
rect 14142 16763 14176 16797
rect 14142 16691 14176 16725
rect 14142 16619 14176 16653
rect 14142 16547 14176 16581
rect 14142 16475 14176 16509
rect 14142 16403 14176 16437
rect 14142 16331 14176 16365
rect 14142 16259 14176 16293
rect 14142 16187 14176 16221
rect 14142 16115 14176 16149
rect 14142 16043 14176 16077
rect 14142 15971 14176 16005
rect 14142 15899 14176 15933
rect 14142 15827 14176 15861
rect 14142 15755 14176 15789
rect 14142 15683 14176 15717
rect 14142 15611 14176 15645
rect 14142 15539 14176 15573
rect 14142 15467 14176 15501
rect 14142 15395 14176 15429
rect 14142 15323 14176 15357
rect 14142 15251 14176 15285
rect 14142 15179 14176 15213
rect 14142 15107 14176 15141
rect 14142 15035 14176 15069
rect 14142 14963 14176 14997
rect 14142 14891 14176 14925
rect 14142 14819 14176 14853
rect 14142 14747 14176 14781
rect 14142 14675 14176 14709
rect 14142 14603 14176 14637
rect 14142 14531 14176 14565
rect 14142 14459 14176 14493
rect 14142 14387 14176 14421
rect 14142 14315 14176 14349
rect 14142 14243 14176 14277
rect 14142 14171 14176 14205
rect 14142 14099 14176 14133
rect 14142 14027 14176 14061
rect 14142 13955 14176 13989
rect 14142 13883 14176 13917
rect 14142 13811 14176 13845
rect 14142 13739 14176 13773
rect 14142 13667 14176 13701
rect 14142 13595 14176 13629
rect 14142 13523 14176 13557
rect 14142 13451 14176 13485
rect 14142 13379 14176 13413
rect 14142 13307 14176 13341
rect 14142 13235 14176 13269
rect 14142 13163 14176 13197
rect 14142 13091 14176 13125
rect 14142 13019 14176 13053
rect 14142 12947 14176 12981
rect 14142 12875 14176 12909
rect 14142 12803 14176 12837
rect 14142 12731 14176 12765
rect 14142 12659 14176 12693
rect 14142 12587 14176 12621
rect 14142 12515 14176 12549
rect 14142 12443 14176 12477
rect 14142 12371 14176 12405
rect 14142 12299 14176 12333
rect 14142 12227 14176 12261
rect 14142 12155 14176 12189
rect 14142 12083 14176 12117
rect 14142 12011 14176 12045
rect 14142 11939 14176 11973
rect 14142 11867 14176 11901
rect 14142 11795 14176 11829
rect 14142 11723 14176 11757
rect 14142 11651 14176 11685
rect 14142 11579 14176 11613
rect 14142 11507 14176 11541
rect 14142 11435 14176 11469
rect 14142 11363 14176 11397
rect 14142 11291 14176 11325
rect 14142 11219 14176 11253
rect 14142 11147 14176 11181
rect 14142 11075 14176 11109
rect 14142 11003 14176 11037
rect 14142 10931 14176 10965
rect 14142 10859 14176 10893
rect 14142 10787 14176 10821
rect 14142 10715 14176 10749
rect 14142 10643 14176 10677
rect 14142 10571 14176 10605
rect 14142 10499 14176 10533
rect 14142 10427 14176 10461
rect 14142 10355 14176 10389
rect 14142 10283 14176 10317
rect 807 10146 841 10180
rect 807 10074 841 10108
rect 14142 10211 14176 10245
rect 14142 10139 14176 10173
rect 14142 10067 14176 10101
rect 891 9908 925 9942
rect 963 9908 997 9942
rect 1035 9908 1069 9942
rect 1107 9908 1141 9942
rect 1179 9908 1213 9942
rect 1251 9908 1285 9942
rect 1323 9908 1357 9942
rect 1395 9908 1429 9942
rect 1467 9908 1501 9942
rect 1539 9908 1573 9942
rect 1611 9908 1645 9942
rect 1683 9908 1717 9942
rect 1755 9908 1789 9942
rect 1827 9908 1861 9942
rect 1899 9908 1933 9942
rect 1971 9908 2005 9942
rect 2043 9908 2077 9942
rect 2115 9908 2149 9942
rect 2187 9908 2221 9942
rect 2259 9908 2293 9942
rect 2331 9908 2365 9942
rect 2403 9908 2437 9942
rect 2475 9908 2509 9942
rect 2547 9908 2581 9942
rect 2619 9908 2653 9942
rect 2691 9908 2725 9942
rect 2763 9908 2797 9942
rect 2835 9908 2869 9942
rect 2907 9908 2941 9942
rect 2979 9908 3013 9942
rect 3051 9908 3085 9942
rect 3123 9908 3157 9942
rect 3195 9908 3229 9942
rect 3267 9908 3301 9942
rect 3339 9908 3373 9942
rect 3411 9908 3445 9942
rect 3483 9908 3517 9942
rect 3555 9908 3589 9942
rect 3627 9908 3661 9942
rect 3699 9908 3733 9942
rect 3771 9908 3805 9942
rect 3843 9908 3877 9942
rect 3915 9908 3949 9942
rect 3987 9908 4021 9942
rect 4059 9908 4093 9942
rect 4131 9908 4165 9942
rect 4203 9908 4237 9942
rect 4275 9908 4309 9942
rect 4347 9908 4381 9942
rect 4419 9908 4453 9942
rect 4491 9908 4525 9942
rect 4563 9908 4597 9942
rect 4635 9908 4669 9942
rect 4707 9908 4741 9942
rect 4779 9908 4813 9942
rect 4851 9908 4885 9942
rect 4923 9908 4957 9942
rect 4995 9908 5029 9942
rect 5067 9908 5101 9942
rect 5139 9908 5173 9942
rect 5211 9908 5245 9942
rect 5283 9908 5317 9942
rect 5355 9908 5389 9942
rect 5427 9908 5461 9942
rect 5499 9908 5533 9942
rect 5571 9908 5605 9942
rect 5643 9908 5677 9942
rect 5715 9908 5749 9942
rect 5787 9908 5821 9942
rect 5859 9908 5893 9942
rect 5931 9908 5965 9942
rect 6003 9908 6037 9942
rect 6075 9908 6109 9942
rect 6147 9908 6181 9942
rect 6219 9908 6253 9942
rect 6291 9908 6325 9942
rect 6363 9908 6397 9942
rect 6435 9908 6469 9942
rect 6507 9908 6541 9942
rect 6579 9908 6613 9942
rect 6651 9908 6685 9942
rect 6723 9908 6757 9942
rect 6795 9908 6829 9942
rect 6867 9908 6901 9942
rect 6939 9908 6973 9942
rect 7011 9908 7045 9942
rect 7083 9908 7117 9942
rect 7155 9908 7189 9942
rect 7227 9908 7261 9942
rect 7299 9908 7333 9942
rect 7371 9908 7405 9942
rect 7443 9908 7477 9942
rect 7515 9908 7549 9942
rect 7587 9908 7621 9942
rect 7659 9908 7693 9942
rect 7731 9908 7765 9942
rect 7803 9908 7837 9942
rect 7875 9908 7909 9942
rect 7947 9908 7981 9942
rect 8019 9908 8053 9942
rect 8091 9908 8125 9942
rect 8163 9908 8197 9942
rect 8235 9908 8269 9942
rect 8307 9908 8341 9942
rect 8379 9908 8413 9942
rect 8451 9908 8485 9942
rect 8523 9908 8557 9942
rect 8595 9908 8629 9942
rect 8667 9908 8701 9942
rect 8739 9908 8773 9942
rect 8811 9908 8845 9942
rect 8883 9908 8917 9942
rect 8955 9908 8989 9942
rect 9027 9908 9061 9942
rect 9099 9908 9133 9942
rect 9171 9908 9205 9942
rect 9243 9908 9277 9942
rect 9315 9908 9349 9942
rect 9387 9908 9421 9942
rect 9459 9908 9493 9942
rect 9531 9908 9565 9942
rect 9603 9908 9637 9942
rect 9675 9908 9709 9942
rect 9747 9908 9781 9942
rect 9819 9908 9853 9942
rect 9891 9908 9925 9942
rect 9963 9908 9997 9942
rect 10035 9908 10069 9942
rect 10107 9908 10141 9942
rect 10179 9908 10213 9942
rect 10251 9908 10285 9942
rect 10323 9908 10357 9942
rect 10395 9908 10429 9942
rect 10467 9908 10501 9942
rect 10539 9908 10573 9942
rect 10611 9908 10645 9942
rect 10683 9908 10717 9942
rect 10755 9908 10789 9942
rect 10827 9908 10861 9942
rect 10899 9908 10933 9942
rect 10971 9908 11005 9942
rect 11043 9908 11077 9942
rect 11115 9908 11149 9942
rect 11187 9908 11221 9942
rect 11259 9908 11293 9942
rect 11331 9908 11365 9942
rect 11403 9908 11437 9942
rect 11475 9908 11509 9942
rect 11547 9908 11581 9942
rect 11619 9908 11653 9942
rect 11691 9908 11725 9942
rect 11763 9908 11797 9942
rect 11835 9908 11869 9942
rect 11907 9908 11941 9942
rect 11979 9908 12013 9942
rect 12051 9908 12085 9942
rect 12123 9908 12157 9942
rect 12195 9908 12229 9942
rect 12267 9908 12301 9942
rect 12339 9908 12373 9942
rect 12411 9908 12445 9942
rect 12483 9908 12517 9942
rect 12555 9908 12589 9942
rect 12627 9908 12661 9942
rect 12699 9908 12733 9942
rect 12771 9908 12805 9942
rect 12843 9908 12877 9942
rect 12915 9908 12949 9942
rect 12987 9908 13021 9942
rect 13059 9908 13093 9942
rect 13131 9908 13165 9942
rect 13203 9908 13237 9942
rect 13275 9908 13309 9942
rect 13347 9908 13381 9942
rect 13419 9908 13453 9942
rect 13491 9908 13525 9942
rect 13563 9908 13597 9942
rect 13635 9908 13669 9942
rect 13707 9908 13741 9942
rect 13779 9908 13813 9942
rect 13851 9908 13885 9942
rect 13923 9908 13957 9942
rect 13995 9908 14029 9942
rect 883 9741 915 9775
rect 915 9741 917 9775
rect 955 9741 983 9775
rect 983 9741 989 9775
rect 1027 9741 1051 9775
rect 1051 9741 1061 9775
rect 1099 9741 1119 9775
rect 1119 9741 1133 9775
rect 1171 9741 1187 9775
rect 1187 9741 1205 9775
rect 1243 9741 1255 9775
rect 1255 9741 1277 9775
rect 1315 9741 1323 9775
rect 1323 9741 1349 9775
rect 1387 9741 1391 9775
rect 1391 9741 1421 9775
rect 1459 9741 1493 9775
rect 1531 9741 1561 9775
rect 1561 9741 1565 9775
rect 1603 9741 1629 9775
rect 1629 9741 1637 9775
rect 1675 9741 1697 9775
rect 1697 9741 1709 9775
rect 1747 9741 1765 9775
rect 1765 9741 1781 9775
rect 1819 9741 1833 9775
rect 1833 9741 1853 9775
rect 1891 9741 1901 9775
rect 1901 9741 1925 9775
rect 1963 9741 1969 9775
rect 1969 9741 1997 9775
rect 2035 9741 2037 9775
rect 2037 9741 2069 9775
rect 12883 9740 12915 9774
rect 12915 9740 12917 9774
rect 12955 9740 12983 9774
rect 12983 9740 12989 9774
rect 13027 9740 13051 9774
rect 13051 9740 13061 9774
rect 13099 9740 13119 9774
rect 13119 9740 13133 9774
rect 13171 9740 13187 9774
rect 13187 9740 13205 9774
rect 13243 9740 13255 9774
rect 13255 9740 13277 9774
rect 13315 9740 13323 9774
rect 13323 9740 13349 9774
rect 13387 9740 13391 9774
rect 13391 9740 13421 9774
rect 13459 9740 13493 9774
rect 13531 9740 13561 9774
rect 13561 9740 13565 9774
rect 13603 9740 13629 9774
rect 13629 9740 13637 9774
rect 13675 9740 13697 9774
rect 13697 9740 13709 9774
rect 13747 9740 13765 9774
rect 13765 9740 13781 9774
rect 13819 9740 13833 9774
rect 13833 9740 13853 9774
rect 13891 9740 13901 9774
rect 13901 9740 13925 9774
rect 13963 9740 13969 9774
rect 13969 9740 13997 9774
rect 14035 9740 14037 9774
rect 14037 9740 14069 9774
rect 14614 36173 14648 36190
rect 14614 36156 14645 36173
rect 14645 36156 14648 36173
rect 14614 36105 14648 36118
rect 14614 36084 14645 36105
rect 14645 36084 14648 36105
rect 14614 36037 14648 36046
rect 14614 36012 14645 36037
rect 14645 36012 14648 36037
rect 14614 35969 14648 35974
rect 14614 35940 14645 35969
rect 14645 35940 14648 35969
rect 14614 35901 14648 35902
rect 14614 35868 14645 35901
rect 14645 35868 14648 35901
rect 14614 35799 14645 35830
rect 14645 35799 14648 35830
rect 14614 35796 14648 35799
rect 14614 35731 14645 35758
rect 14645 35731 14648 35758
rect 14614 35724 14648 35731
rect 14614 35663 14645 35686
rect 14645 35663 14648 35686
rect 14614 35652 14648 35663
rect 14614 35595 14645 35614
rect 14645 35595 14648 35614
rect 14614 35580 14648 35595
rect 14614 35527 14645 35542
rect 14645 35527 14648 35542
rect 14614 35508 14648 35527
rect 14614 35459 14645 35470
rect 14645 35459 14648 35470
rect 14614 35436 14648 35459
rect 14614 35391 14645 35398
rect 14645 35391 14648 35398
rect 14614 35364 14648 35391
rect 14614 35323 14645 35326
rect 14645 35323 14648 35326
rect 14614 35292 14648 35323
rect 14614 35221 14648 35254
rect 14614 35220 14645 35221
rect 14645 35220 14648 35221
rect 14614 35153 14648 35182
rect 14614 35148 14645 35153
rect 14645 35148 14648 35153
rect 14614 35085 14648 35110
rect 14614 35076 14645 35085
rect 14645 35076 14648 35085
rect 14614 35017 14648 35038
rect 14614 35004 14645 35017
rect 14645 35004 14648 35017
rect 14614 34949 14648 34966
rect 14614 34932 14645 34949
rect 14645 34932 14648 34949
rect 14614 34881 14648 34894
rect 14614 34860 14645 34881
rect 14645 34860 14648 34881
rect 14614 34813 14648 34822
rect 14614 34788 14645 34813
rect 14645 34788 14648 34813
rect 14614 34745 14648 34750
rect 14614 34716 14645 34745
rect 14645 34716 14648 34745
rect 14614 34677 14648 34678
rect 14614 34644 14645 34677
rect 14645 34644 14648 34677
rect 14614 34575 14645 34606
rect 14645 34575 14648 34606
rect 14614 34572 14648 34575
rect 14614 34507 14645 34534
rect 14645 34507 14648 34534
rect 14614 34500 14648 34507
rect 14614 34439 14645 34462
rect 14645 34439 14648 34462
rect 14614 34428 14648 34439
rect 14614 34371 14645 34390
rect 14645 34371 14648 34390
rect 14614 34356 14648 34371
rect 14614 34303 14645 34318
rect 14645 34303 14648 34318
rect 14614 34284 14648 34303
rect 14614 34235 14645 34246
rect 14645 34235 14648 34246
rect 14614 34212 14648 34235
rect 14614 34167 14645 34174
rect 14645 34167 14648 34174
rect 14614 34140 14648 34167
rect 14614 34099 14645 34102
rect 14645 34099 14648 34102
rect 14614 34068 14648 34099
rect 14614 33997 14648 34030
rect 14614 33996 14645 33997
rect 14645 33996 14648 33997
rect 14614 33929 14648 33958
rect 14614 33924 14645 33929
rect 14645 33924 14648 33929
rect 14614 33861 14648 33886
rect 14614 33852 14645 33861
rect 14645 33852 14648 33861
rect 14614 33793 14648 33814
rect 14614 33780 14645 33793
rect 14645 33780 14648 33793
rect 14614 33725 14648 33742
rect 14614 33708 14645 33725
rect 14645 33708 14648 33725
rect 14614 33657 14648 33670
rect 14614 33636 14645 33657
rect 14645 33636 14648 33657
rect 14614 33589 14648 33598
rect 14614 33564 14645 33589
rect 14645 33564 14648 33589
rect 14614 33521 14648 33526
rect 14614 33492 14645 33521
rect 14645 33492 14648 33521
rect 14614 33453 14648 33454
rect 14614 33420 14645 33453
rect 14645 33420 14648 33453
rect 14614 33351 14645 33382
rect 14645 33351 14648 33382
rect 14614 33348 14648 33351
rect 14614 33283 14645 33310
rect 14645 33283 14648 33310
rect 14614 33276 14648 33283
rect 14614 33215 14645 33238
rect 14645 33215 14648 33238
rect 14614 33204 14648 33215
rect 14614 33147 14645 33166
rect 14645 33147 14648 33166
rect 14614 33132 14648 33147
rect 14614 33079 14645 33094
rect 14645 33079 14648 33094
rect 14614 33060 14648 33079
rect 14614 33011 14645 33022
rect 14645 33011 14648 33022
rect 14614 32988 14648 33011
rect 14614 32943 14645 32950
rect 14645 32943 14648 32950
rect 14614 32916 14648 32943
rect 14614 32875 14645 32878
rect 14645 32875 14648 32878
rect 14614 32844 14648 32875
rect 14614 32773 14648 32806
rect 14614 32772 14645 32773
rect 14645 32772 14648 32773
rect 14614 32705 14648 32734
rect 14614 32700 14645 32705
rect 14645 32700 14648 32705
rect 14614 32637 14648 32662
rect 14614 32628 14645 32637
rect 14645 32628 14648 32637
rect 14614 32569 14648 32590
rect 14614 32556 14645 32569
rect 14645 32556 14648 32569
rect 14614 32501 14648 32518
rect 14614 32484 14645 32501
rect 14645 32484 14648 32501
rect 14614 32433 14648 32446
rect 14614 32412 14645 32433
rect 14645 32412 14648 32433
rect 14614 32365 14648 32374
rect 14614 32340 14645 32365
rect 14645 32340 14648 32365
rect 14614 32297 14648 32302
rect 14614 32268 14645 32297
rect 14645 32268 14648 32297
rect 14614 32229 14648 32230
rect 14614 32196 14645 32229
rect 14645 32196 14648 32229
rect 14614 32127 14645 32158
rect 14645 32127 14648 32158
rect 14614 32124 14648 32127
rect 14614 32059 14645 32086
rect 14645 32059 14648 32086
rect 14614 32052 14648 32059
rect 14614 31991 14645 32014
rect 14645 31991 14648 32014
rect 14614 31980 14648 31991
rect 14614 31923 14645 31942
rect 14645 31923 14648 31942
rect 14614 31908 14648 31923
rect 14614 31855 14645 31870
rect 14645 31855 14648 31870
rect 14614 31836 14648 31855
rect 14614 31787 14645 31798
rect 14645 31787 14648 31798
rect 14614 31764 14648 31787
rect 14614 31719 14645 31726
rect 14645 31719 14648 31726
rect 14614 31692 14648 31719
rect 14614 31651 14645 31654
rect 14645 31651 14648 31654
rect 14614 31620 14648 31651
rect 14614 31549 14648 31582
rect 14614 31548 14645 31549
rect 14645 31548 14648 31549
rect 14614 31481 14648 31510
rect 14614 31476 14645 31481
rect 14645 31476 14648 31481
rect 14614 31413 14648 31438
rect 14614 31404 14645 31413
rect 14645 31404 14648 31413
rect 14614 31345 14648 31366
rect 14614 31332 14645 31345
rect 14645 31332 14648 31345
rect 14614 31277 14648 31294
rect 14614 31260 14645 31277
rect 14645 31260 14648 31277
rect 14614 31209 14648 31222
rect 14614 31188 14645 31209
rect 14645 31188 14648 31209
rect 14614 31141 14648 31150
rect 14614 31116 14645 31141
rect 14645 31116 14648 31141
rect 14614 31073 14648 31078
rect 14614 31044 14645 31073
rect 14645 31044 14648 31073
rect 14614 31005 14648 31006
rect 14614 30972 14645 31005
rect 14645 30972 14648 31005
rect 14614 30903 14645 30934
rect 14645 30903 14648 30934
rect 14614 30900 14648 30903
rect 14614 30835 14645 30862
rect 14645 30835 14648 30862
rect 14614 30828 14648 30835
rect 14614 30767 14645 30790
rect 14645 30767 14648 30790
rect 14614 30756 14648 30767
rect 14614 30699 14645 30718
rect 14645 30699 14648 30718
rect 14614 30684 14648 30699
rect 14614 30631 14645 30646
rect 14645 30631 14648 30646
rect 14614 30612 14648 30631
rect 14614 30563 14645 30574
rect 14645 30563 14648 30574
rect 14614 30540 14648 30563
rect 14614 30495 14645 30502
rect 14645 30495 14648 30502
rect 14614 30468 14648 30495
rect 14614 30427 14645 30430
rect 14645 30427 14648 30430
rect 14614 30396 14648 30427
rect 14614 30325 14648 30358
rect 14614 30324 14645 30325
rect 14645 30324 14648 30325
rect 14614 30257 14648 30286
rect 14614 30252 14645 30257
rect 14645 30252 14648 30257
rect 14614 30189 14648 30214
rect 14614 30180 14645 30189
rect 14645 30180 14648 30189
rect 14614 30121 14648 30142
rect 14614 30108 14645 30121
rect 14645 30108 14648 30121
rect 14614 30053 14648 30070
rect 14614 30036 14645 30053
rect 14645 30036 14648 30053
rect 14614 29985 14648 29998
rect 14614 29964 14645 29985
rect 14645 29964 14648 29985
rect 14614 29917 14648 29926
rect 14614 29892 14645 29917
rect 14645 29892 14648 29917
rect 14614 29849 14648 29854
rect 14614 29820 14645 29849
rect 14645 29820 14648 29849
rect 14614 29781 14648 29782
rect 14614 29748 14645 29781
rect 14645 29748 14648 29781
rect 14614 29679 14645 29710
rect 14645 29679 14648 29710
rect 14614 29676 14648 29679
rect 14614 29611 14645 29638
rect 14645 29611 14648 29638
rect 14614 29604 14648 29611
rect 14614 29543 14645 29566
rect 14645 29543 14648 29566
rect 14614 29532 14648 29543
rect 14614 29475 14645 29494
rect 14645 29475 14648 29494
rect 14614 29460 14648 29475
rect 14614 29407 14645 29422
rect 14645 29407 14648 29422
rect 14614 29388 14648 29407
rect 14614 29339 14645 29350
rect 14645 29339 14648 29350
rect 14614 29316 14648 29339
rect 14614 29271 14645 29278
rect 14645 29271 14648 29278
rect 14614 29244 14648 29271
rect 14614 29203 14645 29206
rect 14645 29203 14648 29206
rect 14614 29172 14648 29203
rect 14614 29101 14648 29134
rect 14614 29100 14645 29101
rect 14645 29100 14648 29101
rect 14614 29033 14648 29062
rect 14614 29028 14645 29033
rect 14645 29028 14648 29033
rect 14614 28965 14648 28990
rect 14614 28956 14645 28965
rect 14645 28956 14648 28965
rect 14614 28897 14648 28918
rect 14614 28884 14645 28897
rect 14645 28884 14648 28897
rect 14614 28829 14648 28846
rect 14614 28812 14645 28829
rect 14645 28812 14648 28829
rect 14614 28761 14648 28774
rect 14614 28740 14645 28761
rect 14645 28740 14648 28761
rect 14614 28693 14648 28702
rect 14614 28668 14645 28693
rect 14645 28668 14648 28693
rect 14614 28625 14648 28630
rect 14614 28596 14645 28625
rect 14645 28596 14648 28625
rect 14614 28557 14648 28558
rect 14614 28524 14645 28557
rect 14645 28524 14648 28557
rect 14614 28455 14645 28486
rect 14645 28455 14648 28486
rect 14614 28452 14648 28455
rect 14614 28387 14645 28414
rect 14645 28387 14648 28414
rect 14614 28380 14648 28387
rect 14614 28319 14645 28342
rect 14645 28319 14648 28342
rect 14614 28308 14648 28319
rect 14614 28251 14645 28270
rect 14645 28251 14648 28270
rect 14614 28236 14648 28251
rect 14614 28183 14645 28198
rect 14645 28183 14648 28198
rect 14614 28164 14648 28183
rect 14614 28115 14645 28126
rect 14645 28115 14648 28126
rect 14614 28092 14648 28115
rect 14614 28047 14645 28054
rect 14645 28047 14648 28054
rect 14614 28020 14648 28047
rect 14614 27979 14645 27982
rect 14645 27979 14648 27982
rect 14614 27948 14648 27979
rect 14614 27877 14648 27910
rect 14614 27876 14645 27877
rect 14645 27876 14648 27877
rect 14614 27809 14648 27838
rect 14614 27804 14645 27809
rect 14645 27804 14648 27809
rect 14614 27741 14648 27766
rect 14614 27732 14645 27741
rect 14645 27732 14648 27741
rect 14614 27673 14648 27694
rect 14614 27660 14645 27673
rect 14645 27660 14648 27673
rect 14614 27605 14648 27622
rect 14614 27588 14645 27605
rect 14645 27588 14648 27605
rect 14614 27537 14648 27550
rect 14614 27516 14645 27537
rect 14645 27516 14648 27537
rect 14614 27469 14648 27478
rect 14614 27444 14645 27469
rect 14645 27444 14648 27469
rect 14614 27401 14648 27406
rect 14614 27372 14645 27401
rect 14645 27372 14648 27401
rect 14614 27333 14648 27334
rect 14614 27300 14645 27333
rect 14645 27300 14648 27333
rect 14614 27231 14645 27262
rect 14645 27231 14648 27262
rect 14614 27228 14648 27231
rect 14614 27163 14645 27190
rect 14645 27163 14648 27190
rect 14614 27156 14648 27163
rect 14614 27095 14645 27118
rect 14645 27095 14648 27118
rect 14614 27084 14648 27095
rect 14614 27027 14645 27046
rect 14645 27027 14648 27046
rect 14614 27012 14648 27027
rect 14614 26959 14645 26974
rect 14645 26959 14648 26974
rect 14614 26940 14648 26959
rect 14614 26891 14645 26902
rect 14645 26891 14648 26902
rect 14614 26868 14648 26891
rect 14614 26823 14645 26830
rect 14645 26823 14648 26830
rect 14614 26796 14648 26823
rect 14614 26755 14645 26758
rect 14645 26755 14648 26758
rect 14614 26724 14648 26755
rect 14614 26653 14648 26686
rect 14614 26652 14645 26653
rect 14645 26652 14648 26653
rect 14614 26585 14648 26614
rect 14614 26580 14645 26585
rect 14645 26580 14648 26585
rect 14614 26517 14648 26542
rect 14614 26508 14645 26517
rect 14645 26508 14648 26517
rect 14614 26449 14648 26470
rect 14614 26436 14645 26449
rect 14645 26436 14648 26449
rect 14614 26381 14648 26398
rect 14614 26364 14645 26381
rect 14645 26364 14648 26381
rect 14614 26313 14648 26326
rect 14614 26292 14645 26313
rect 14645 26292 14648 26313
rect 14614 26245 14648 26254
rect 14614 26220 14645 26245
rect 14645 26220 14648 26245
rect 14614 26177 14648 26182
rect 14614 26148 14645 26177
rect 14645 26148 14648 26177
rect 14614 26109 14648 26110
rect 14614 26076 14645 26109
rect 14645 26076 14648 26109
rect 14614 26007 14645 26038
rect 14645 26007 14648 26038
rect 14614 26004 14648 26007
rect 14614 25939 14645 25966
rect 14645 25939 14648 25966
rect 14614 25932 14648 25939
rect 14614 25871 14645 25894
rect 14645 25871 14648 25894
rect 14614 25860 14648 25871
rect 14614 25803 14645 25822
rect 14645 25803 14648 25822
rect 14614 25788 14648 25803
rect 14614 25735 14645 25750
rect 14645 25735 14648 25750
rect 14614 25716 14648 25735
rect 14614 25667 14645 25678
rect 14645 25667 14648 25678
rect 14614 25644 14648 25667
rect 14614 25599 14645 25606
rect 14645 25599 14648 25606
rect 14614 25572 14648 25599
rect 14614 25531 14645 25534
rect 14645 25531 14648 25534
rect 14614 25500 14648 25531
rect 14614 25429 14648 25462
rect 14614 25428 14645 25429
rect 14645 25428 14648 25429
rect 14614 25361 14648 25390
rect 14614 25356 14645 25361
rect 14645 25356 14648 25361
rect 14614 25293 14648 25318
rect 14614 25284 14645 25293
rect 14645 25284 14648 25293
rect 14614 25225 14648 25246
rect 14614 25212 14645 25225
rect 14645 25212 14648 25225
rect 14614 25157 14648 25174
rect 14614 25140 14645 25157
rect 14645 25140 14648 25157
rect 14614 25089 14648 25102
rect 14614 25068 14645 25089
rect 14645 25068 14648 25089
rect 14614 25021 14648 25030
rect 14614 24996 14645 25021
rect 14645 24996 14648 25021
rect 14614 24953 14648 24958
rect 14614 24924 14645 24953
rect 14645 24924 14648 24953
rect 14614 24885 14648 24886
rect 14614 24852 14645 24885
rect 14645 24852 14648 24885
rect 14614 24783 14645 24814
rect 14645 24783 14648 24814
rect 14614 24780 14648 24783
rect 14614 24715 14645 24742
rect 14645 24715 14648 24742
rect 14614 24708 14648 24715
rect 14614 24647 14645 24670
rect 14645 24647 14648 24670
rect 14614 24636 14648 24647
rect 14614 24579 14645 24598
rect 14645 24579 14648 24598
rect 14614 24564 14648 24579
rect 14614 24511 14645 24526
rect 14645 24511 14648 24526
rect 14614 24492 14648 24511
rect 14614 24443 14645 24454
rect 14645 24443 14648 24454
rect 14614 24420 14648 24443
rect 14614 24375 14645 24382
rect 14645 24375 14648 24382
rect 14614 24348 14648 24375
rect 14614 24307 14645 24310
rect 14645 24307 14648 24310
rect 14614 24276 14648 24307
rect 14614 24205 14648 24238
rect 14614 24204 14645 24205
rect 14645 24204 14648 24205
rect 14614 24137 14648 24166
rect 14614 24132 14645 24137
rect 14645 24132 14648 24137
rect 14614 24069 14648 24094
rect 14614 24060 14645 24069
rect 14645 24060 14648 24069
rect 14614 24001 14648 24022
rect 14614 23988 14645 24001
rect 14645 23988 14648 24001
rect 14614 23933 14648 23950
rect 14614 23916 14645 23933
rect 14645 23916 14648 23933
rect 14614 23865 14648 23878
rect 14614 23844 14645 23865
rect 14645 23844 14648 23865
rect 14614 23797 14648 23806
rect 14614 23772 14645 23797
rect 14645 23772 14648 23797
rect 14614 23729 14648 23734
rect 14614 23700 14645 23729
rect 14645 23700 14648 23729
rect 14614 23661 14648 23662
rect 14614 23628 14645 23661
rect 14645 23628 14648 23661
rect 14614 23559 14645 23590
rect 14645 23559 14648 23590
rect 14614 23556 14648 23559
rect 14614 23491 14645 23518
rect 14645 23491 14648 23518
rect 14614 23484 14648 23491
rect 14614 23423 14645 23446
rect 14645 23423 14648 23446
rect 14614 23412 14648 23423
rect 14614 23355 14645 23374
rect 14645 23355 14648 23374
rect 14614 23340 14648 23355
rect 14614 23287 14645 23302
rect 14645 23287 14648 23302
rect 14614 23268 14648 23287
rect 14614 23219 14645 23230
rect 14645 23219 14648 23230
rect 14614 23196 14648 23219
rect 14614 23151 14645 23158
rect 14645 23151 14648 23158
rect 14614 23124 14648 23151
rect 14614 23083 14645 23086
rect 14645 23083 14648 23086
rect 14614 23052 14648 23083
rect 14614 22981 14648 23014
rect 14614 22980 14645 22981
rect 14645 22980 14648 22981
rect 14614 22913 14648 22942
rect 14614 22908 14645 22913
rect 14645 22908 14648 22913
rect 14614 22845 14648 22870
rect 14614 22836 14645 22845
rect 14645 22836 14648 22845
rect 14614 22777 14648 22798
rect 14614 22764 14645 22777
rect 14645 22764 14648 22777
rect 14614 22709 14648 22726
rect 14614 22692 14645 22709
rect 14645 22692 14648 22709
rect 14614 22641 14648 22654
rect 14614 22620 14645 22641
rect 14645 22620 14648 22641
rect 14614 22573 14648 22582
rect 14614 22548 14645 22573
rect 14645 22548 14648 22573
rect 14614 22505 14648 22510
rect 14614 22476 14645 22505
rect 14645 22476 14648 22505
rect 14614 22437 14648 22438
rect 14614 22404 14645 22437
rect 14645 22404 14648 22437
rect 14614 22335 14645 22366
rect 14645 22335 14648 22366
rect 14614 22332 14648 22335
rect 14614 22267 14645 22294
rect 14645 22267 14648 22294
rect 14614 22260 14648 22267
rect 14614 22199 14645 22222
rect 14645 22199 14648 22222
rect 14614 22188 14648 22199
rect 14614 22131 14645 22150
rect 14645 22131 14648 22150
rect 14614 22116 14648 22131
rect 14614 22063 14645 22078
rect 14645 22063 14648 22078
rect 14614 22044 14648 22063
rect 14614 21995 14645 22006
rect 14645 21995 14648 22006
rect 14614 21972 14648 21995
rect 14614 21927 14645 21934
rect 14645 21927 14648 21934
rect 14614 21900 14648 21927
rect 14614 21859 14645 21862
rect 14645 21859 14648 21862
rect 14614 21828 14648 21859
rect 14614 21757 14648 21790
rect 14614 21756 14645 21757
rect 14645 21756 14648 21757
rect 14614 21689 14648 21718
rect 14614 21684 14645 21689
rect 14645 21684 14648 21689
rect 14614 21621 14648 21646
rect 14614 21612 14645 21621
rect 14645 21612 14648 21621
rect 14614 21553 14648 21574
rect 14614 21540 14645 21553
rect 14645 21540 14648 21553
rect 14614 21485 14648 21502
rect 14614 21468 14645 21485
rect 14645 21468 14648 21485
rect 14614 21417 14648 21430
rect 14614 21396 14645 21417
rect 14645 21396 14648 21417
rect 14614 21349 14648 21358
rect 14614 21324 14645 21349
rect 14645 21324 14648 21349
rect 14614 21281 14648 21286
rect 14614 21252 14645 21281
rect 14645 21252 14648 21281
rect 14614 21213 14648 21214
rect 14614 21180 14645 21213
rect 14645 21180 14648 21213
rect 14614 21111 14645 21142
rect 14645 21111 14648 21142
rect 14614 21108 14648 21111
rect 14614 21043 14645 21070
rect 14645 21043 14648 21070
rect 14614 21036 14648 21043
rect 14614 20975 14645 20998
rect 14645 20975 14648 20998
rect 14614 20964 14648 20975
rect 14614 20907 14645 20926
rect 14645 20907 14648 20926
rect 14614 20892 14648 20907
rect 14614 20839 14645 20854
rect 14645 20839 14648 20854
rect 14614 20820 14648 20839
rect 14614 20771 14645 20782
rect 14645 20771 14648 20782
rect 14614 20748 14648 20771
rect 14614 20703 14645 20710
rect 14645 20703 14648 20710
rect 14614 20676 14648 20703
rect 14614 20635 14645 20638
rect 14645 20635 14648 20638
rect 14614 20604 14648 20635
rect 14614 20533 14648 20566
rect 14614 20532 14645 20533
rect 14645 20532 14648 20533
rect 14614 20465 14648 20494
rect 14614 20460 14645 20465
rect 14645 20460 14648 20465
rect 14614 20397 14648 20422
rect 14614 20388 14645 20397
rect 14645 20388 14648 20397
rect 14614 20329 14648 20350
rect 14614 20316 14645 20329
rect 14645 20316 14648 20329
rect 14614 20261 14648 20278
rect 14614 20244 14645 20261
rect 14645 20244 14648 20261
rect 14614 20193 14648 20206
rect 14614 20172 14645 20193
rect 14645 20172 14648 20193
rect 14614 20125 14648 20134
rect 14614 20100 14645 20125
rect 14645 20100 14648 20125
rect 14614 20057 14648 20062
rect 14614 20028 14645 20057
rect 14645 20028 14648 20057
rect 14614 19989 14648 19990
rect 14614 19956 14645 19989
rect 14645 19956 14648 19989
rect 14614 19887 14645 19918
rect 14645 19887 14648 19918
rect 14614 19884 14648 19887
rect 14614 19819 14645 19846
rect 14645 19819 14648 19846
rect 14614 19812 14648 19819
rect 14614 19751 14645 19774
rect 14645 19751 14648 19774
rect 14614 19740 14648 19751
rect 14614 19683 14645 19702
rect 14645 19683 14648 19702
rect 14614 19668 14648 19683
rect 14614 19615 14645 19630
rect 14645 19615 14648 19630
rect 14614 19596 14648 19615
rect 14614 19547 14645 19558
rect 14645 19547 14648 19558
rect 14614 19524 14648 19547
rect 14614 19479 14645 19486
rect 14645 19479 14648 19486
rect 14614 19452 14648 19479
rect 14614 19411 14645 19414
rect 14645 19411 14648 19414
rect 14614 19380 14648 19411
rect 14614 19309 14648 19342
rect 14614 19308 14645 19309
rect 14645 19308 14648 19309
rect 14614 19241 14648 19270
rect 14614 19236 14645 19241
rect 14645 19236 14648 19241
rect 14614 19173 14648 19198
rect 14614 19164 14645 19173
rect 14645 19164 14648 19173
rect 14614 19105 14648 19126
rect 14614 19092 14645 19105
rect 14645 19092 14648 19105
rect 14614 19037 14648 19054
rect 14614 19020 14645 19037
rect 14645 19020 14648 19037
rect 14614 18969 14648 18982
rect 14614 18948 14645 18969
rect 14645 18948 14648 18969
rect 14614 18901 14648 18910
rect 14614 18876 14645 18901
rect 14645 18876 14648 18901
rect 14614 18833 14648 18838
rect 14614 18804 14645 18833
rect 14645 18804 14648 18833
rect 14614 18765 14648 18766
rect 14614 18732 14645 18765
rect 14645 18732 14648 18765
rect 14614 18663 14645 18694
rect 14645 18663 14648 18694
rect 14614 18660 14648 18663
rect 14614 18595 14645 18622
rect 14645 18595 14648 18622
rect 14614 18588 14648 18595
rect 14614 18527 14645 18550
rect 14645 18527 14648 18550
rect 14614 18516 14648 18527
rect 14614 18459 14645 18478
rect 14645 18459 14648 18478
rect 14614 18444 14648 18459
rect 14614 18391 14645 18406
rect 14645 18391 14648 18406
rect 14614 18372 14648 18391
rect 14614 18323 14645 18334
rect 14645 18323 14648 18334
rect 14614 18300 14648 18323
rect 14614 18255 14645 18262
rect 14645 18255 14648 18262
rect 14614 18228 14648 18255
rect 14614 18187 14645 18190
rect 14645 18187 14648 18190
rect 14614 18156 14648 18187
rect 14614 18085 14648 18118
rect 14614 18084 14645 18085
rect 14645 18084 14648 18085
rect 14614 18017 14648 18046
rect 14614 18012 14645 18017
rect 14645 18012 14648 18017
rect 14614 17949 14648 17974
rect 14614 17940 14645 17949
rect 14645 17940 14648 17949
rect 14614 17881 14648 17902
rect 14614 17868 14645 17881
rect 14645 17868 14648 17881
rect 14614 17813 14648 17830
rect 14614 17796 14645 17813
rect 14645 17796 14648 17813
rect 14614 17745 14648 17758
rect 14614 17724 14645 17745
rect 14645 17724 14648 17745
rect 14614 17677 14648 17686
rect 14614 17652 14645 17677
rect 14645 17652 14648 17677
rect 14614 17609 14648 17614
rect 14614 17580 14645 17609
rect 14645 17580 14648 17609
rect 14614 17541 14648 17542
rect 14614 17508 14645 17541
rect 14645 17508 14648 17541
rect 14614 17439 14645 17470
rect 14645 17439 14648 17470
rect 14614 17436 14648 17439
rect 14614 17371 14645 17398
rect 14645 17371 14648 17398
rect 14614 17364 14648 17371
rect 14614 17303 14645 17326
rect 14645 17303 14648 17326
rect 14614 17292 14648 17303
rect 14614 17235 14645 17254
rect 14645 17235 14648 17254
rect 14614 17220 14648 17235
rect 14614 17167 14645 17182
rect 14645 17167 14648 17182
rect 14614 17148 14648 17167
rect 14614 17099 14645 17110
rect 14645 17099 14648 17110
rect 14614 17076 14648 17099
rect 14614 17031 14645 17038
rect 14645 17031 14648 17038
rect 14614 17004 14648 17031
rect 14614 16963 14645 16966
rect 14645 16963 14648 16966
rect 14614 16932 14648 16963
rect 14614 16861 14648 16894
rect 14614 16860 14645 16861
rect 14645 16860 14648 16861
rect 14614 16793 14648 16822
rect 14614 16788 14645 16793
rect 14645 16788 14648 16793
rect 14614 16725 14648 16750
rect 14614 16716 14645 16725
rect 14645 16716 14648 16725
rect 14614 16657 14648 16678
rect 14614 16644 14645 16657
rect 14645 16644 14648 16657
rect 14614 16589 14648 16606
rect 14614 16572 14645 16589
rect 14645 16572 14648 16589
rect 14614 16521 14648 16534
rect 14614 16500 14645 16521
rect 14645 16500 14648 16521
rect 14614 16453 14648 16462
rect 14614 16428 14645 16453
rect 14645 16428 14648 16453
rect 14614 16385 14648 16390
rect 14614 16356 14645 16385
rect 14645 16356 14648 16385
rect 14614 16317 14648 16318
rect 14614 16284 14645 16317
rect 14645 16284 14648 16317
rect 14614 16215 14645 16246
rect 14645 16215 14648 16246
rect 14614 16212 14648 16215
rect 14614 16147 14645 16174
rect 14645 16147 14648 16174
rect 14614 16140 14648 16147
rect 14614 16079 14645 16102
rect 14645 16079 14648 16102
rect 14614 16068 14648 16079
rect 14614 16011 14645 16030
rect 14645 16011 14648 16030
rect 14614 15996 14648 16011
rect 14614 15943 14645 15958
rect 14645 15943 14648 15958
rect 14614 15924 14648 15943
rect 14614 15875 14645 15886
rect 14645 15875 14648 15886
rect 14614 15852 14648 15875
rect 14614 15807 14645 15814
rect 14645 15807 14648 15814
rect 14614 15780 14648 15807
rect 14614 15739 14645 15742
rect 14645 15739 14648 15742
rect 14614 15708 14648 15739
rect 14614 15637 14648 15670
rect 14614 15636 14645 15637
rect 14645 15636 14648 15637
rect 14614 15569 14648 15598
rect 14614 15564 14645 15569
rect 14645 15564 14648 15569
rect 14614 15501 14648 15526
rect 14614 15492 14645 15501
rect 14645 15492 14648 15501
rect 14614 15433 14648 15454
rect 14614 15420 14645 15433
rect 14645 15420 14648 15433
rect 14614 15365 14648 15382
rect 14614 15348 14645 15365
rect 14645 15348 14648 15365
rect 14614 15297 14648 15310
rect 14614 15276 14645 15297
rect 14645 15276 14648 15297
rect 14614 15229 14648 15238
rect 14614 15204 14645 15229
rect 14645 15204 14648 15229
rect 14614 15161 14648 15166
rect 14614 15132 14645 15161
rect 14645 15132 14648 15161
rect 14614 15093 14648 15094
rect 14614 15060 14645 15093
rect 14645 15060 14648 15093
rect 14614 14991 14645 15022
rect 14645 14991 14648 15022
rect 14614 14988 14648 14991
rect 14614 14923 14645 14950
rect 14645 14923 14648 14950
rect 14614 14916 14648 14923
rect 14614 14855 14645 14878
rect 14645 14855 14648 14878
rect 14614 14844 14648 14855
rect 14614 14787 14645 14806
rect 14645 14787 14648 14806
rect 14614 14772 14648 14787
rect 14614 14719 14645 14734
rect 14645 14719 14648 14734
rect 14614 14700 14648 14719
rect 14614 14651 14645 14662
rect 14645 14651 14648 14662
rect 14614 14628 14648 14651
rect 14614 14583 14645 14590
rect 14645 14583 14648 14590
rect 14614 14556 14648 14583
rect 14614 14515 14645 14518
rect 14645 14515 14648 14518
rect 14614 14484 14648 14515
rect 14614 14413 14648 14446
rect 14614 14412 14645 14413
rect 14645 14412 14648 14413
rect 14614 14345 14648 14374
rect 14614 14340 14645 14345
rect 14645 14340 14648 14345
rect 14614 14277 14648 14302
rect 14614 14268 14645 14277
rect 14645 14268 14648 14277
rect 14614 14209 14648 14230
rect 14614 14196 14645 14209
rect 14645 14196 14648 14209
rect 14614 14141 14648 14158
rect 14614 14124 14645 14141
rect 14645 14124 14648 14141
rect 14614 14073 14648 14086
rect 14614 14052 14645 14073
rect 14645 14052 14648 14073
rect 14614 14005 14648 14014
rect 14614 13980 14645 14005
rect 14645 13980 14648 14005
rect 14614 13937 14648 13942
rect 14614 13908 14645 13937
rect 14645 13908 14648 13937
rect 14614 13869 14648 13870
rect 14614 13836 14645 13869
rect 14645 13836 14648 13869
rect 14614 13767 14645 13798
rect 14645 13767 14648 13798
rect 14614 13764 14648 13767
rect 14614 13699 14645 13726
rect 14645 13699 14648 13726
rect 14614 13692 14648 13699
rect 14614 13631 14645 13654
rect 14645 13631 14648 13654
rect 14614 13620 14648 13631
rect 14614 13563 14645 13582
rect 14645 13563 14648 13582
rect 14614 13548 14648 13563
rect 14614 13495 14645 13510
rect 14645 13495 14648 13510
rect 14614 13476 14648 13495
rect 14614 13427 14645 13438
rect 14645 13427 14648 13438
rect 14614 13404 14648 13427
rect 14614 13359 14645 13366
rect 14645 13359 14648 13366
rect 14614 13332 14648 13359
rect 14614 13291 14645 13294
rect 14645 13291 14648 13294
rect 14614 13260 14648 13291
rect 14614 13189 14648 13222
rect 14614 13188 14645 13189
rect 14645 13188 14648 13189
rect 14614 13121 14648 13150
rect 14614 13116 14645 13121
rect 14645 13116 14648 13121
rect 14614 13053 14648 13078
rect 14614 13044 14645 13053
rect 14645 13044 14648 13053
rect 14614 12985 14648 13006
rect 14614 12972 14645 12985
rect 14645 12972 14648 12985
rect 14614 12917 14648 12934
rect 14614 12900 14645 12917
rect 14645 12900 14648 12917
rect 14614 12849 14648 12862
rect 14614 12828 14645 12849
rect 14645 12828 14648 12849
rect 14614 12781 14648 12790
rect 14614 12756 14645 12781
rect 14645 12756 14648 12781
rect 14614 12713 14648 12718
rect 14614 12684 14645 12713
rect 14645 12684 14648 12713
rect 14614 12645 14648 12646
rect 14614 12612 14645 12645
rect 14645 12612 14648 12645
rect 14614 12543 14645 12574
rect 14645 12543 14648 12574
rect 14614 12540 14648 12543
rect 14614 12475 14645 12502
rect 14645 12475 14648 12502
rect 14614 12468 14648 12475
rect 14614 12407 14645 12430
rect 14645 12407 14648 12430
rect 14614 12396 14648 12407
rect 14614 12339 14645 12358
rect 14645 12339 14648 12358
rect 14614 12324 14648 12339
rect 14614 12271 14645 12286
rect 14645 12271 14648 12286
rect 14614 12252 14648 12271
rect 14614 12203 14645 12214
rect 14645 12203 14648 12214
rect 14614 12180 14648 12203
rect 14614 12135 14645 12142
rect 14645 12135 14648 12142
rect 14614 12108 14648 12135
rect 14614 12067 14645 12070
rect 14645 12067 14648 12070
rect 14614 12036 14648 12067
rect 14614 11965 14648 11998
rect 14614 11964 14645 11965
rect 14645 11964 14648 11965
rect 14614 11897 14648 11926
rect 14614 11892 14645 11897
rect 14645 11892 14648 11897
rect 14614 11829 14648 11854
rect 14614 11820 14645 11829
rect 14645 11820 14648 11829
rect 14614 11761 14648 11782
rect 14614 11748 14645 11761
rect 14645 11748 14648 11761
rect 14614 11693 14648 11710
rect 14614 11676 14645 11693
rect 14645 11676 14648 11693
rect 14614 11625 14648 11638
rect 14614 11604 14645 11625
rect 14645 11604 14648 11625
rect 14614 11557 14648 11566
rect 14614 11532 14645 11557
rect 14645 11532 14648 11557
rect 14614 11489 14648 11494
rect 14614 11460 14645 11489
rect 14645 11460 14648 11489
rect 14614 11421 14648 11422
rect 14614 11388 14645 11421
rect 14645 11388 14648 11421
rect 14614 11319 14645 11350
rect 14645 11319 14648 11350
rect 14614 11316 14648 11319
rect 14614 11251 14645 11278
rect 14645 11251 14648 11278
rect 14614 11244 14648 11251
rect 14614 11183 14645 11206
rect 14645 11183 14648 11206
rect 14614 11172 14648 11183
rect 14614 11115 14645 11134
rect 14645 11115 14648 11134
rect 14614 11100 14648 11115
rect 14614 11047 14645 11062
rect 14645 11047 14648 11062
rect 14614 11028 14648 11047
rect 14614 10979 14645 10990
rect 14645 10979 14648 10990
rect 14614 10956 14648 10979
rect 14614 10911 14645 10918
rect 14645 10911 14648 10918
rect 14614 10884 14648 10911
rect 14614 10843 14645 10846
rect 14645 10843 14648 10846
rect 14614 10812 14648 10843
rect 14614 10741 14648 10774
rect 14614 10740 14645 10741
rect 14645 10740 14648 10741
rect 14614 10673 14648 10702
rect 14614 10668 14645 10673
rect 14645 10668 14648 10673
rect 14614 10605 14648 10630
rect 14614 10596 14645 10605
rect 14645 10596 14648 10605
rect 14614 10537 14648 10558
rect 14614 10524 14645 10537
rect 14645 10524 14648 10537
rect 14614 10469 14648 10486
rect 14614 10452 14645 10469
rect 14645 10452 14648 10469
rect 14614 10401 14648 10414
rect 14614 10380 14645 10401
rect 14645 10380 14648 10401
rect 14614 10333 14648 10342
rect 14614 10308 14645 10333
rect 14645 10308 14648 10333
rect 14614 10265 14648 10270
rect 14614 10236 14645 10265
rect 14645 10236 14648 10265
rect 14614 10197 14648 10198
rect 14614 10164 14645 10197
rect 14645 10164 14648 10197
rect 14614 10095 14645 10126
rect 14645 10095 14648 10126
rect 14614 10092 14648 10095
rect 14614 10027 14645 10054
rect 14645 10027 14648 10054
rect 14614 10020 14648 10027
rect 14614 9959 14645 9982
rect 14645 9959 14648 9982
rect 14614 9948 14648 9959
rect 14614 9891 14645 9910
rect 14645 9891 14648 9910
rect 14614 9876 14648 9891
rect 14614 9823 14645 9838
rect 14645 9823 14648 9838
rect 14614 9804 14648 9823
rect 14614 9755 14645 9766
rect 14645 9755 14648 9766
rect 14614 9732 14648 9755
rect 320 9689 351 9697
rect 351 9689 354 9697
rect 320 9663 354 9689
rect 14614 9687 14645 9694
rect 14645 9687 14648 9694
rect 14614 9660 14648 9687
rect 320 9418 354 9452
rect 610 9450 644 9452
rect 2311 9450 2345 9452
rect 2383 9450 2417 9452
rect 2455 9450 2489 9452
rect 2527 9450 2561 9452
rect 2599 9450 2633 9452
rect 2671 9450 2705 9452
rect 2743 9450 2777 9452
rect 2815 9450 2849 9452
rect 2887 9450 2921 9452
rect 2959 9450 2993 9452
rect 3031 9450 3065 9452
rect 3103 9450 3137 9452
rect 3175 9450 3209 9452
rect 3247 9450 3281 9452
rect 3319 9450 3353 9452
rect 3391 9450 3425 9452
rect 3463 9450 3497 9452
rect 3535 9450 3569 9452
rect 3607 9450 3641 9452
rect 3679 9450 3713 9452
rect 3751 9450 3785 9452
rect 3823 9450 3857 9452
rect 3895 9450 3929 9452
rect 3967 9450 4001 9452
rect 4039 9450 4073 9452
rect 4111 9450 4145 9452
rect 4183 9450 4217 9452
rect 4255 9450 4289 9452
rect 4327 9450 4361 9452
rect 4399 9450 4433 9452
rect 4471 9450 4505 9452
rect 4543 9450 4577 9452
rect 4615 9450 4649 9452
rect 4687 9450 4721 9452
rect 4759 9450 4793 9452
rect 4831 9450 4865 9452
rect 4903 9450 4937 9452
rect 4975 9450 5009 9452
rect 5047 9450 5081 9452
rect 5119 9450 5153 9452
rect 5191 9450 5225 9452
rect 5263 9450 5297 9452
rect 5335 9450 5369 9452
rect 5407 9450 5441 9452
rect 5479 9450 5513 9452
rect 5551 9450 5585 9452
rect 5623 9450 5657 9452
rect 5695 9450 5729 9452
rect 5767 9450 5801 9452
rect 5839 9450 5873 9452
rect 5911 9450 5945 9452
rect 5983 9450 6017 9452
rect 6055 9450 6089 9452
rect 6127 9450 6161 9452
rect 6199 9450 6233 9452
rect 6271 9450 6305 9452
rect 6343 9450 6377 9452
rect 6415 9450 6449 9452
rect 6487 9450 6521 9452
rect 6559 9450 6593 9452
rect 6631 9450 6665 9452
rect 6703 9450 6737 9452
rect 6775 9450 6809 9452
rect 6847 9450 6881 9452
rect 6919 9450 6953 9452
rect 6991 9450 7025 9452
rect 7063 9450 7097 9452
rect 7135 9450 7169 9452
rect 7207 9450 7241 9452
rect 7279 9450 7313 9452
rect 7351 9450 7385 9452
rect 7423 9450 7457 9452
rect 7495 9450 7529 9452
rect 7567 9450 7601 9452
rect 7639 9450 7673 9452
rect 7711 9450 7745 9452
rect 7783 9450 7817 9452
rect 7855 9450 7889 9452
rect 7927 9450 7961 9452
rect 7999 9450 8033 9452
rect 8071 9450 8105 9452
rect 8143 9450 8177 9452
rect 8215 9450 8249 9452
rect 8287 9450 8321 9452
rect 8359 9450 8393 9452
rect 8431 9450 8465 9452
rect 8503 9450 8537 9452
rect 8575 9450 8609 9452
rect 8647 9450 8681 9452
rect 8719 9450 8753 9452
rect 8791 9450 8825 9452
rect 8863 9450 8897 9452
rect 8935 9450 8969 9452
rect 9007 9450 9041 9452
rect 9079 9450 9113 9452
rect 9151 9450 9185 9452
rect 9223 9450 9257 9452
rect 9295 9450 9329 9452
rect 9367 9450 9401 9452
rect 9439 9450 9473 9452
rect 9511 9450 9545 9452
rect 9583 9450 9617 9452
rect 9655 9450 9689 9452
rect 9727 9450 9761 9452
rect 9799 9450 9833 9452
rect 9871 9450 9905 9452
rect 9943 9450 9977 9452
rect 10015 9450 10049 9452
rect 10087 9450 10121 9452
rect 10159 9450 10193 9452
rect 10231 9450 10265 9452
rect 10303 9450 10337 9452
rect 10375 9450 10409 9452
rect 10447 9450 10481 9452
rect 10519 9450 10553 9452
rect 10591 9450 10625 9452
rect 10663 9450 10697 9452
rect 10735 9450 10769 9452
rect 10807 9450 10841 9452
rect 10879 9450 10913 9452
rect 10951 9450 10985 9452
rect 11023 9450 11057 9452
rect 11095 9450 11129 9452
rect 11167 9450 11201 9452
rect 11239 9450 11273 9452
rect 11311 9450 11345 9452
rect 11383 9450 11417 9452
rect 11455 9450 11489 9452
rect 11527 9450 11561 9452
rect 11599 9450 11633 9452
rect 11671 9450 11705 9452
rect 11743 9450 11777 9452
rect 11815 9450 11849 9452
rect 11887 9450 11921 9452
rect 11959 9450 11993 9452
rect 12031 9450 12065 9452
rect 12103 9450 12137 9452
rect 12175 9450 12209 9452
rect 12247 9450 12281 9452
rect 12319 9450 12353 9452
rect 12391 9450 12425 9452
rect 12463 9450 12497 9452
rect 12535 9450 12569 9452
rect 12607 9450 12641 9452
rect 14314 9450 14348 9452
rect 610 9418 642 9450
rect 642 9418 644 9450
rect 2311 9418 2342 9450
rect 2342 9418 2345 9450
rect 2383 9418 2410 9450
rect 2410 9418 2417 9450
rect 2455 9418 2478 9450
rect 2478 9418 2489 9450
rect 2527 9418 2546 9450
rect 2546 9418 2561 9450
rect 2599 9418 2614 9450
rect 2614 9418 2633 9450
rect 2671 9418 2682 9450
rect 2682 9418 2705 9450
rect 2743 9418 2750 9450
rect 2750 9418 2777 9450
rect 2815 9418 2818 9450
rect 2818 9418 2849 9450
rect 2887 9418 2920 9450
rect 2920 9418 2921 9450
rect 2959 9418 2988 9450
rect 2988 9418 2993 9450
rect 3031 9418 3056 9450
rect 3056 9418 3065 9450
rect 3103 9418 3124 9450
rect 3124 9418 3137 9450
rect 3175 9418 3192 9450
rect 3192 9418 3209 9450
rect 3247 9418 3260 9450
rect 3260 9418 3281 9450
rect 3319 9418 3328 9450
rect 3328 9418 3353 9450
rect 3391 9418 3396 9450
rect 3396 9418 3425 9450
rect 3463 9418 3464 9450
rect 3464 9418 3497 9450
rect 3535 9418 3566 9450
rect 3566 9418 3569 9450
rect 3607 9418 3634 9450
rect 3634 9418 3641 9450
rect 3679 9418 3702 9450
rect 3702 9418 3713 9450
rect 3751 9418 3770 9450
rect 3770 9418 3785 9450
rect 3823 9418 3838 9450
rect 3838 9418 3857 9450
rect 3895 9418 3906 9450
rect 3906 9418 3929 9450
rect 3967 9418 3974 9450
rect 3974 9418 4001 9450
rect 4039 9418 4042 9450
rect 4042 9418 4073 9450
rect 4111 9418 4144 9450
rect 4144 9418 4145 9450
rect 4183 9418 4212 9450
rect 4212 9418 4217 9450
rect 4255 9418 4280 9450
rect 4280 9418 4289 9450
rect 4327 9418 4348 9450
rect 4348 9418 4361 9450
rect 4399 9418 4416 9450
rect 4416 9418 4433 9450
rect 4471 9418 4484 9450
rect 4484 9418 4505 9450
rect 4543 9418 4552 9450
rect 4552 9418 4577 9450
rect 4615 9418 4620 9450
rect 4620 9418 4649 9450
rect 4687 9418 4688 9450
rect 4688 9418 4721 9450
rect 4759 9418 4790 9450
rect 4790 9418 4793 9450
rect 4831 9418 4858 9450
rect 4858 9418 4865 9450
rect 4903 9418 4926 9450
rect 4926 9418 4937 9450
rect 4975 9418 4994 9450
rect 4994 9418 5009 9450
rect 5047 9418 5062 9450
rect 5062 9418 5081 9450
rect 5119 9418 5130 9450
rect 5130 9418 5153 9450
rect 5191 9418 5198 9450
rect 5198 9418 5225 9450
rect 5263 9418 5266 9450
rect 5266 9418 5297 9450
rect 5335 9418 5368 9450
rect 5368 9418 5369 9450
rect 5407 9418 5436 9450
rect 5436 9418 5441 9450
rect 5479 9418 5504 9450
rect 5504 9418 5513 9450
rect 5551 9418 5572 9450
rect 5572 9418 5585 9450
rect 5623 9418 5640 9450
rect 5640 9418 5657 9450
rect 5695 9418 5708 9450
rect 5708 9418 5729 9450
rect 5767 9418 5776 9450
rect 5776 9418 5801 9450
rect 5839 9418 5844 9450
rect 5844 9418 5873 9450
rect 5911 9418 5912 9450
rect 5912 9418 5945 9450
rect 5983 9418 6014 9450
rect 6014 9418 6017 9450
rect 6055 9418 6082 9450
rect 6082 9418 6089 9450
rect 6127 9418 6150 9450
rect 6150 9418 6161 9450
rect 6199 9418 6218 9450
rect 6218 9418 6233 9450
rect 6271 9418 6286 9450
rect 6286 9418 6305 9450
rect 6343 9418 6354 9450
rect 6354 9418 6377 9450
rect 6415 9418 6422 9450
rect 6422 9418 6449 9450
rect 6487 9418 6490 9450
rect 6490 9418 6521 9450
rect 6559 9418 6592 9450
rect 6592 9418 6593 9450
rect 6631 9418 6660 9450
rect 6660 9418 6665 9450
rect 6703 9418 6728 9450
rect 6728 9418 6737 9450
rect 6775 9418 6796 9450
rect 6796 9418 6809 9450
rect 6847 9418 6864 9450
rect 6864 9418 6881 9450
rect 6919 9418 6932 9450
rect 6932 9418 6953 9450
rect 6991 9418 7000 9450
rect 7000 9418 7025 9450
rect 7063 9418 7068 9450
rect 7068 9418 7097 9450
rect 7135 9418 7136 9450
rect 7136 9418 7169 9450
rect 7207 9418 7238 9450
rect 7238 9418 7241 9450
rect 7279 9418 7306 9450
rect 7306 9418 7313 9450
rect 7351 9418 7374 9450
rect 7374 9418 7385 9450
rect 7423 9418 7442 9450
rect 7442 9418 7457 9450
rect 7495 9418 7510 9450
rect 7510 9418 7529 9450
rect 7567 9418 7578 9450
rect 7578 9418 7601 9450
rect 7639 9418 7646 9450
rect 7646 9418 7673 9450
rect 7711 9418 7714 9450
rect 7714 9418 7745 9450
rect 7783 9418 7816 9450
rect 7816 9418 7817 9450
rect 7855 9418 7884 9450
rect 7884 9418 7889 9450
rect 7927 9418 7952 9450
rect 7952 9418 7961 9450
rect 7999 9418 8020 9450
rect 8020 9418 8033 9450
rect 8071 9418 8088 9450
rect 8088 9418 8105 9450
rect 8143 9418 8156 9450
rect 8156 9418 8177 9450
rect 8215 9418 8224 9450
rect 8224 9418 8249 9450
rect 8287 9418 8292 9450
rect 8292 9418 8321 9450
rect 8359 9418 8360 9450
rect 8360 9418 8393 9450
rect 8431 9418 8462 9450
rect 8462 9418 8465 9450
rect 8503 9418 8530 9450
rect 8530 9418 8537 9450
rect 8575 9418 8598 9450
rect 8598 9418 8609 9450
rect 8647 9418 8666 9450
rect 8666 9418 8681 9450
rect 8719 9418 8734 9450
rect 8734 9418 8753 9450
rect 8791 9418 8802 9450
rect 8802 9418 8825 9450
rect 8863 9418 8870 9450
rect 8870 9418 8897 9450
rect 8935 9418 8938 9450
rect 8938 9418 8969 9450
rect 9007 9418 9040 9450
rect 9040 9418 9041 9450
rect 9079 9418 9108 9450
rect 9108 9418 9113 9450
rect 9151 9418 9176 9450
rect 9176 9418 9185 9450
rect 9223 9418 9244 9450
rect 9244 9418 9257 9450
rect 9295 9418 9312 9450
rect 9312 9418 9329 9450
rect 9367 9418 9380 9450
rect 9380 9418 9401 9450
rect 9439 9418 9448 9450
rect 9448 9418 9473 9450
rect 9511 9418 9516 9450
rect 9516 9418 9545 9450
rect 9583 9418 9584 9450
rect 9584 9418 9617 9450
rect 9655 9418 9686 9450
rect 9686 9418 9689 9450
rect 9727 9418 9754 9450
rect 9754 9418 9761 9450
rect 9799 9418 9822 9450
rect 9822 9418 9833 9450
rect 9871 9418 9890 9450
rect 9890 9418 9905 9450
rect 9943 9418 9958 9450
rect 9958 9418 9977 9450
rect 10015 9418 10026 9450
rect 10026 9418 10049 9450
rect 10087 9418 10094 9450
rect 10094 9418 10121 9450
rect 10159 9418 10162 9450
rect 10162 9418 10193 9450
rect 10231 9418 10264 9450
rect 10264 9418 10265 9450
rect 10303 9418 10332 9450
rect 10332 9418 10337 9450
rect 10375 9418 10400 9450
rect 10400 9418 10409 9450
rect 10447 9418 10468 9450
rect 10468 9418 10481 9450
rect 10519 9418 10536 9450
rect 10536 9418 10553 9450
rect 10591 9418 10604 9450
rect 10604 9418 10625 9450
rect 10663 9418 10672 9450
rect 10672 9418 10697 9450
rect 10735 9418 10740 9450
rect 10740 9418 10769 9450
rect 10807 9418 10808 9450
rect 10808 9418 10841 9450
rect 10879 9418 10910 9450
rect 10910 9418 10913 9450
rect 10951 9418 10978 9450
rect 10978 9418 10985 9450
rect 11023 9418 11046 9450
rect 11046 9418 11057 9450
rect 11095 9418 11114 9450
rect 11114 9418 11129 9450
rect 11167 9418 11182 9450
rect 11182 9418 11201 9450
rect 11239 9418 11250 9450
rect 11250 9418 11273 9450
rect 11311 9418 11318 9450
rect 11318 9418 11345 9450
rect 11383 9418 11386 9450
rect 11386 9418 11417 9450
rect 11455 9418 11488 9450
rect 11488 9418 11489 9450
rect 11527 9418 11556 9450
rect 11556 9418 11561 9450
rect 11599 9418 11624 9450
rect 11624 9418 11633 9450
rect 11671 9418 11692 9450
rect 11692 9418 11705 9450
rect 11743 9418 11760 9450
rect 11760 9418 11777 9450
rect 11815 9418 11828 9450
rect 11828 9418 11849 9450
rect 11887 9418 11896 9450
rect 11896 9418 11921 9450
rect 11959 9418 11964 9450
rect 11964 9418 11993 9450
rect 12031 9418 12032 9450
rect 12032 9418 12065 9450
rect 12103 9418 12134 9450
rect 12134 9418 12137 9450
rect 12175 9418 12202 9450
rect 12202 9418 12209 9450
rect 12247 9418 12270 9450
rect 12270 9418 12281 9450
rect 12319 9418 12338 9450
rect 12338 9418 12353 9450
rect 12391 9418 12406 9450
rect 12406 9418 12425 9450
rect 12463 9418 12474 9450
rect 12474 9418 12497 9450
rect 12535 9418 12542 9450
rect 12542 9418 12569 9450
rect 12607 9418 12610 9450
rect 12610 9418 12641 9450
rect 14314 9418 14344 9450
rect 14344 9418 14348 9450
rect 14614 9418 14648 9452
<< metal1 >>
rect 245 36534 14724 36574
rect 245 36500 320 36534
rect 354 36533 14724 36534
rect 354 36500 14614 36533
rect 245 36499 14614 36500
rect 14648 36499 14724 36533
rect 245 36498 14724 36499
rect 245 36464 556 36498
rect 590 36464 628 36498
rect 662 36464 700 36498
rect 734 36464 772 36498
rect 806 36464 844 36498
rect 878 36464 916 36498
rect 950 36464 988 36498
rect 1022 36464 1060 36498
rect 1094 36464 1132 36498
rect 1166 36464 1204 36498
rect 1238 36464 1276 36498
rect 1310 36464 1348 36498
rect 1382 36464 1420 36498
rect 1454 36464 1492 36498
rect 1526 36464 1564 36498
rect 1598 36464 1636 36498
rect 1670 36464 1708 36498
rect 1742 36464 1780 36498
rect 1814 36464 1852 36498
rect 1886 36464 1924 36498
rect 1958 36464 1996 36498
rect 2030 36464 2068 36498
rect 2102 36464 2140 36498
rect 2174 36464 2212 36498
rect 2246 36464 2284 36498
rect 2318 36464 2356 36498
rect 2390 36464 2428 36498
rect 2462 36464 2500 36498
rect 2534 36464 2572 36498
rect 2606 36464 2644 36498
rect 2678 36464 2716 36498
rect 2750 36464 2788 36498
rect 2822 36464 2860 36498
rect 2894 36464 2932 36498
rect 2966 36464 3004 36498
rect 3038 36464 3076 36498
rect 3110 36464 3148 36498
rect 3182 36464 3220 36498
rect 3254 36464 3292 36498
rect 3326 36464 3364 36498
rect 3398 36464 3436 36498
rect 3470 36464 3508 36498
rect 3542 36464 3580 36498
rect 3614 36464 3652 36498
rect 3686 36464 3724 36498
rect 3758 36464 3796 36498
rect 3830 36464 3868 36498
rect 3902 36464 3940 36498
rect 3974 36464 4012 36498
rect 4046 36464 4084 36498
rect 4118 36464 4156 36498
rect 4190 36464 4228 36498
rect 4262 36464 4300 36498
rect 4334 36464 4372 36498
rect 4406 36464 4444 36498
rect 4478 36464 4516 36498
rect 4550 36464 4588 36498
rect 4622 36464 4660 36498
rect 4694 36464 4732 36498
rect 4766 36464 4804 36498
rect 4838 36464 4876 36498
rect 4910 36464 4948 36498
rect 4982 36464 5020 36498
rect 5054 36464 5092 36498
rect 5126 36464 5164 36498
rect 5198 36464 5236 36498
rect 5270 36464 5308 36498
rect 5342 36464 5380 36498
rect 5414 36464 5452 36498
rect 5486 36464 5524 36498
rect 5558 36464 5596 36498
rect 5630 36464 5668 36498
rect 5702 36464 5740 36498
rect 5774 36464 5812 36498
rect 5846 36464 5884 36498
rect 5918 36464 5956 36498
rect 5990 36464 6028 36498
rect 6062 36464 6100 36498
rect 6134 36464 6172 36498
rect 6206 36464 6244 36498
rect 6278 36464 6316 36498
rect 6350 36464 6388 36498
rect 6422 36464 6460 36498
rect 6494 36464 6532 36498
rect 6566 36464 6604 36498
rect 6638 36464 6676 36498
rect 6710 36464 6748 36498
rect 6782 36464 6820 36498
rect 6854 36464 6892 36498
rect 6926 36464 6964 36498
rect 6998 36464 7036 36498
rect 7070 36464 7108 36498
rect 7142 36464 7180 36498
rect 7214 36464 7252 36498
rect 7286 36464 7324 36498
rect 7358 36464 7396 36498
rect 7430 36464 7468 36498
rect 7502 36464 7540 36498
rect 7574 36464 7612 36498
rect 7646 36464 7684 36498
rect 7718 36464 7756 36498
rect 7790 36464 7828 36498
rect 7862 36464 7900 36498
rect 7934 36464 7972 36498
rect 8006 36464 8044 36498
rect 8078 36464 8116 36498
rect 8150 36464 8188 36498
rect 8222 36464 8260 36498
rect 8294 36464 8332 36498
rect 8366 36464 8404 36498
rect 8438 36464 8476 36498
rect 8510 36464 8548 36498
rect 8582 36464 8620 36498
rect 8654 36464 8692 36498
rect 8726 36464 8764 36498
rect 8798 36464 8836 36498
rect 8870 36464 8908 36498
rect 8942 36464 8980 36498
rect 9014 36464 9052 36498
rect 9086 36464 9124 36498
rect 9158 36464 9196 36498
rect 9230 36464 9268 36498
rect 9302 36464 9340 36498
rect 9374 36464 9412 36498
rect 9446 36464 9484 36498
rect 9518 36464 9556 36498
rect 9590 36464 9628 36498
rect 9662 36464 9700 36498
rect 9734 36464 9772 36498
rect 9806 36464 9844 36498
rect 9878 36464 9916 36498
rect 9950 36464 9988 36498
rect 10022 36464 10060 36498
rect 10094 36464 10132 36498
rect 10166 36464 10204 36498
rect 10238 36464 10276 36498
rect 10310 36464 10348 36498
rect 10382 36464 10420 36498
rect 10454 36464 10492 36498
rect 10526 36464 10564 36498
rect 10598 36464 10636 36498
rect 10670 36464 10708 36498
rect 10742 36464 10780 36498
rect 10814 36464 10852 36498
rect 10886 36464 10924 36498
rect 10958 36464 10996 36498
rect 11030 36464 11068 36498
rect 11102 36464 11140 36498
rect 11174 36464 11212 36498
rect 11246 36464 11284 36498
rect 11318 36464 11356 36498
rect 11390 36464 11428 36498
rect 11462 36464 11500 36498
rect 11534 36464 11572 36498
rect 11606 36464 11644 36498
rect 11678 36464 11716 36498
rect 11750 36464 11788 36498
rect 11822 36464 11860 36498
rect 11894 36464 11932 36498
rect 11966 36464 12004 36498
rect 12038 36464 12076 36498
rect 12110 36464 12148 36498
rect 12182 36464 12220 36498
rect 12254 36464 12292 36498
rect 12326 36464 12364 36498
rect 12398 36464 12436 36498
rect 12470 36464 12508 36498
rect 12542 36464 12580 36498
rect 12614 36464 12652 36498
rect 12686 36464 12724 36498
rect 12758 36464 12796 36498
rect 12830 36464 12868 36498
rect 12902 36464 12940 36498
rect 12974 36464 13012 36498
rect 13046 36464 13084 36498
rect 13118 36464 13156 36498
rect 13190 36464 13228 36498
rect 13262 36464 13300 36498
rect 13334 36464 13372 36498
rect 13406 36464 13444 36498
rect 13478 36464 13516 36498
rect 13550 36464 13588 36498
rect 13622 36464 13660 36498
rect 13694 36464 13732 36498
rect 13766 36464 13804 36498
rect 13838 36464 13876 36498
rect 13910 36464 13948 36498
rect 13982 36464 14020 36498
rect 14054 36464 14092 36498
rect 14126 36464 14164 36498
rect 14198 36464 14236 36498
rect 14270 36464 14308 36498
rect 14342 36464 14380 36498
rect 14414 36464 14724 36498
rect 245 36462 14724 36464
rect 245 36428 320 36462
rect 354 36461 14724 36462
rect 354 36428 14614 36461
rect 245 36427 14614 36428
rect 14648 36427 14724 36461
rect 245 36389 14724 36427
rect 245 36265 430 36389
rect 245 36231 320 36265
rect 354 36231 430 36265
rect 245 36193 430 36231
rect 245 36159 320 36193
rect 354 36159 430 36193
rect 245 36121 430 36159
rect 245 36087 320 36121
rect 354 36087 430 36121
rect 245 36049 430 36087
rect 14539 36262 14724 36389
rect 14539 36228 14614 36262
rect 14648 36228 14724 36262
rect 14539 36190 14724 36228
rect 14539 36156 14614 36190
rect 14648 36156 14724 36190
rect 14539 36118 14724 36156
rect 14539 36084 14614 36118
rect 14648 36084 14724 36118
rect 245 36015 320 36049
rect 354 36015 430 36049
tri 850 36046 857 36053 se
rect 857 36046 14119 36053
tri 14119 36046 14126 36053 sw
rect 14539 36046 14724 36084
tri 823 36019 850 36046 se
rect 850 36019 14126 36046
rect 245 35977 430 36015
tri 816 36012 823 36019 se
rect 823 36012 14126 36019
tri 14126 36012 14160 36046 sw
rect 14539 36012 14614 36046
rect 14648 36012 14724 36046
tri 807 36003 816 36012 se
rect 816 36003 14160 36012
rect 245 35943 320 35977
rect 354 35943 430 35977
tri 773 35969 807 36003 se
rect 807 35969 1007 36003
rect 1041 35969 1079 36003
rect 1113 35969 1151 36003
rect 1185 35969 1223 36003
rect 1257 35969 1295 36003
rect 1329 35969 1367 36003
rect 1401 35969 1439 36003
rect 1473 35969 1511 36003
rect 1545 35969 1583 36003
rect 1617 35969 1655 36003
rect 1689 35969 1727 36003
rect 1761 35969 1799 36003
rect 1833 35969 1871 36003
rect 1905 35969 1943 36003
rect 1977 35969 2015 36003
rect 2049 35969 2087 36003
rect 2121 35969 2159 36003
rect 2193 35969 2231 36003
rect 2265 35969 2303 36003
rect 2337 35969 2375 36003
rect 2409 35969 2447 36003
rect 2481 35969 2519 36003
rect 2553 35969 2591 36003
rect 2625 35969 2663 36003
rect 2697 35969 2735 36003
rect 2769 35969 2807 36003
rect 2841 35969 2879 36003
rect 2913 35969 2951 36003
rect 2985 35969 3023 36003
rect 3057 35969 3095 36003
rect 3129 35969 3167 36003
rect 3201 35969 3239 36003
rect 3273 35969 3311 36003
rect 3345 35969 3383 36003
rect 3417 35969 3455 36003
rect 3489 35969 3527 36003
rect 3561 35969 3599 36003
rect 3633 35969 3671 36003
rect 3705 35969 3743 36003
rect 3777 35969 3815 36003
rect 3849 35969 3887 36003
rect 3921 35969 3959 36003
rect 3993 35969 4031 36003
rect 4065 35969 4103 36003
rect 4137 35969 4175 36003
rect 4209 35969 4247 36003
rect 4281 35969 4319 36003
rect 4353 35969 4391 36003
rect 4425 35969 4463 36003
rect 4497 35969 4535 36003
rect 4569 35969 4607 36003
rect 4641 35969 4679 36003
rect 4713 35969 4751 36003
rect 4785 35969 4823 36003
rect 4857 35969 4895 36003
rect 4929 35969 4967 36003
rect 5001 35969 5039 36003
rect 5073 35969 5111 36003
rect 5145 35969 5183 36003
rect 5217 35969 5255 36003
rect 5289 35969 5327 36003
rect 5361 35969 5399 36003
rect 5433 35969 5471 36003
rect 5505 35969 5543 36003
rect 5577 35969 5615 36003
rect 5649 35969 5687 36003
rect 5721 35969 5759 36003
rect 5793 35969 5831 36003
rect 5865 35969 5903 36003
rect 5937 35969 5975 36003
rect 6009 35969 6047 36003
rect 6081 35969 6119 36003
rect 6153 35969 6191 36003
rect 6225 35969 6263 36003
rect 6297 35969 6335 36003
rect 6369 35969 6407 36003
rect 6441 35969 6479 36003
rect 6513 35969 6551 36003
rect 6585 35969 6623 36003
rect 6657 35969 6695 36003
rect 6729 35969 6767 36003
rect 6801 35969 6839 36003
rect 6873 35969 6911 36003
rect 6945 35969 6983 36003
rect 7017 35969 7055 36003
rect 7089 35969 7127 36003
rect 7161 35969 7199 36003
rect 7233 35969 7271 36003
rect 7305 35969 7343 36003
rect 7377 35969 7415 36003
rect 7449 35969 7487 36003
rect 7521 35969 7559 36003
rect 7593 35969 7631 36003
rect 7665 35969 7703 36003
rect 7737 35969 7775 36003
rect 7809 35969 7847 36003
rect 7881 35969 7919 36003
rect 7953 35969 7991 36003
rect 8025 35969 8063 36003
rect 8097 35969 8135 36003
rect 8169 35969 8207 36003
rect 8241 35969 8279 36003
rect 8313 35969 8351 36003
rect 8385 35969 8423 36003
rect 8457 35969 8495 36003
rect 8529 35969 8567 36003
rect 8601 35969 8639 36003
rect 8673 35969 8711 36003
rect 8745 35969 8783 36003
rect 8817 35969 8855 36003
rect 8889 35969 8927 36003
rect 8961 35969 8999 36003
rect 9033 35969 9071 36003
rect 9105 35969 9143 36003
rect 9177 35969 9215 36003
rect 9249 35969 9287 36003
rect 9321 35969 9359 36003
rect 9393 35969 9431 36003
rect 9465 35969 9503 36003
rect 9537 35969 9575 36003
rect 9609 35969 9647 36003
rect 9681 35969 9719 36003
rect 9753 35969 9791 36003
rect 9825 35969 9863 36003
rect 9897 35969 9935 36003
rect 9969 35969 10007 36003
rect 10041 35969 10079 36003
rect 10113 35969 10151 36003
rect 10185 35969 10223 36003
rect 10257 35969 10295 36003
rect 10329 35969 10367 36003
rect 10401 35969 10439 36003
rect 10473 35969 10511 36003
rect 10545 35969 10583 36003
rect 10617 35969 10655 36003
rect 10689 35969 10727 36003
rect 10761 35969 10799 36003
rect 10833 35969 10871 36003
rect 10905 35969 10943 36003
rect 10977 35969 11015 36003
rect 11049 35969 11087 36003
rect 11121 35969 11159 36003
rect 11193 35969 11231 36003
rect 11265 35969 11303 36003
rect 11337 35969 11375 36003
rect 11409 35969 11447 36003
rect 11481 35969 11519 36003
rect 11553 35969 11591 36003
rect 11625 35969 11663 36003
rect 11697 35969 11735 36003
rect 11769 35969 11807 36003
rect 11841 35969 11879 36003
rect 11913 35969 11951 36003
rect 11985 35969 12023 36003
rect 12057 35969 12095 36003
rect 12129 35969 12167 36003
rect 12201 35969 12239 36003
rect 12273 35969 12311 36003
rect 12345 35969 12383 36003
rect 12417 35969 12455 36003
rect 12489 35969 12527 36003
rect 12561 35969 12599 36003
rect 12633 35969 12671 36003
rect 12705 35969 12743 36003
rect 12777 35969 12815 36003
rect 12849 35969 12887 36003
rect 12921 35969 12959 36003
rect 12993 35969 13031 36003
rect 13065 35969 13103 36003
rect 13137 35969 13175 36003
rect 13209 35969 13247 36003
rect 13281 35969 13319 36003
rect 13353 35969 13391 36003
rect 13425 35969 13463 36003
rect 13497 35969 13535 36003
rect 13569 35969 13607 36003
rect 13641 35969 13679 36003
rect 13713 35969 13751 36003
rect 13785 35969 13823 36003
rect 13857 35969 13895 36003
rect 13929 35969 13967 36003
rect 14001 35974 14160 36003
tri 14160 35974 14198 36012 sw
rect 14539 35974 14724 36012
rect 14001 35969 14198 35974
rect 245 35905 430 35943
rect 245 35871 320 35905
rect 354 35871 430 35905
rect 245 35833 430 35871
rect 245 35799 320 35833
rect 354 35799 430 35833
rect 245 35761 430 35799
rect 245 35727 320 35761
rect 354 35727 430 35761
rect 245 35689 430 35727
rect 245 35655 320 35689
rect 354 35655 430 35689
rect 245 35617 430 35655
rect 245 35583 320 35617
rect 354 35583 430 35617
rect 245 35545 430 35583
rect 245 35511 320 35545
rect 354 35511 430 35545
rect 245 35473 430 35511
rect 245 35439 320 35473
rect 354 35439 430 35473
rect 245 35401 430 35439
rect 245 35367 320 35401
rect 354 35367 430 35401
rect 245 35329 430 35367
rect 245 35295 320 35329
rect 354 35295 430 35329
rect 245 35257 430 35295
rect 245 35223 320 35257
rect 354 35223 430 35257
rect 245 35185 430 35223
rect 245 35151 320 35185
rect 354 35151 430 35185
rect 245 35113 430 35151
rect 245 35079 320 35113
rect 354 35079 430 35113
rect 245 35041 430 35079
rect 245 35007 320 35041
rect 354 35007 430 35041
rect 245 34969 430 35007
rect 245 34935 320 34969
rect 354 34935 430 34969
rect 245 34897 430 34935
rect 245 34863 320 34897
rect 354 34863 430 34897
rect 245 34825 430 34863
rect 245 34791 320 34825
rect 354 34791 430 34825
rect 245 34753 430 34791
rect 245 34719 320 34753
rect 354 34719 430 34753
rect 245 34681 430 34719
rect 245 34647 320 34681
rect 354 34647 430 34681
rect 245 34609 430 34647
rect 245 34575 320 34609
rect 354 34575 430 34609
rect 245 34537 430 34575
rect 245 34503 320 34537
rect 354 34503 430 34537
rect 245 34465 430 34503
rect 245 34431 320 34465
rect 354 34431 430 34465
rect 245 34393 430 34431
rect 245 34359 320 34393
rect 354 34359 430 34393
rect 245 34321 430 34359
rect 245 34287 320 34321
rect 354 34287 430 34321
rect 245 34249 430 34287
rect 245 34215 320 34249
rect 354 34215 430 34249
rect 245 34177 430 34215
rect 245 34143 320 34177
rect 354 34143 430 34177
rect 245 34105 430 34143
rect 245 34071 320 34105
rect 354 34071 430 34105
rect 245 34033 430 34071
rect 245 33999 320 34033
rect 354 33999 430 34033
rect 245 33961 430 33999
rect 245 33927 320 33961
rect 354 33927 430 33961
rect 245 33889 430 33927
rect 245 33855 320 33889
rect 354 33855 430 33889
rect 245 33817 430 33855
rect 245 33783 320 33817
rect 354 33783 430 33817
rect 245 33745 430 33783
rect 245 33711 320 33745
rect 354 33711 430 33745
rect 245 33673 430 33711
rect 245 33639 320 33673
rect 354 33639 430 33673
rect 245 33601 430 33639
rect 245 33567 320 33601
rect 354 33567 430 33601
rect 245 33529 430 33567
rect 245 33495 320 33529
rect 354 33495 430 33529
rect 245 33457 430 33495
rect 245 33423 320 33457
rect 354 33423 430 33457
rect 245 33385 430 33423
rect 245 33351 320 33385
rect 354 33351 430 33385
rect 245 33313 430 33351
rect 245 33279 320 33313
rect 354 33279 430 33313
rect 245 33241 430 33279
rect 245 33207 320 33241
rect 354 33207 430 33241
rect 245 33169 430 33207
rect 245 33135 320 33169
rect 354 33135 430 33169
rect 245 33097 430 33135
rect 245 33063 320 33097
rect 354 33063 430 33097
rect 245 33025 430 33063
rect 245 32991 320 33025
rect 354 32991 430 33025
rect 245 32953 430 32991
rect 245 32919 320 32953
rect 354 32919 430 32953
rect 245 32881 430 32919
rect 245 32847 320 32881
rect 354 32847 430 32881
rect 245 32809 430 32847
rect 245 32775 320 32809
rect 354 32775 430 32809
rect 245 32737 430 32775
rect 245 32703 320 32737
rect 354 32703 430 32737
rect 245 32665 430 32703
rect 245 32631 320 32665
rect 354 32631 430 32665
rect 245 32593 430 32631
rect 245 32559 320 32593
rect 354 32559 430 32593
rect 245 32521 430 32559
rect 245 32487 320 32521
rect 354 32487 430 32521
rect 245 32449 430 32487
rect 245 32415 320 32449
rect 354 32415 430 32449
rect 245 32377 430 32415
rect 245 32343 320 32377
rect 354 32343 430 32377
rect 245 32305 430 32343
rect 245 32271 320 32305
rect 354 32271 430 32305
rect 245 32233 430 32271
rect 245 32199 320 32233
rect 354 32199 430 32233
rect 245 32161 430 32199
rect 245 32127 320 32161
rect 354 32127 430 32161
rect 245 32089 430 32127
rect 245 32055 320 32089
rect 354 32055 430 32089
rect 245 32017 430 32055
rect 245 31983 320 32017
rect 354 31983 430 32017
rect 245 31945 430 31983
rect 245 31911 320 31945
rect 354 31911 430 31945
rect 245 31873 430 31911
rect 245 31839 320 31873
rect 354 31839 430 31873
rect 245 31801 430 31839
rect 245 31767 320 31801
rect 354 31767 430 31801
rect 245 31729 430 31767
rect 245 31695 320 31729
rect 354 31695 430 31729
rect 245 31657 430 31695
rect 245 31623 320 31657
rect 354 31623 430 31657
rect 245 31585 430 31623
rect 245 31551 320 31585
rect 354 31551 430 31585
rect 245 31513 430 31551
rect 245 31479 320 31513
rect 354 31479 430 31513
rect 245 31441 430 31479
rect 245 31407 320 31441
rect 354 31407 430 31441
rect 245 31369 430 31407
rect 245 31335 320 31369
rect 354 31335 430 31369
rect 245 31297 430 31335
rect 245 31263 320 31297
rect 354 31263 430 31297
rect 245 31225 430 31263
rect 245 31191 320 31225
rect 354 31191 430 31225
rect 245 31153 430 31191
rect 245 31119 320 31153
rect 354 31119 430 31153
rect 245 31081 430 31119
rect 245 31047 320 31081
rect 354 31047 430 31081
rect 245 31009 430 31047
rect 245 30975 320 31009
rect 354 30975 430 31009
rect 245 30937 430 30975
rect 245 30903 320 30937
rect 354 30903 430 30937
rect 245 30865 430 30903
rect 245 30831 320 30865
rect 354 30831 430 30865
rect 245 30793 430 30831
rect 245 30759 320 30793
rect 354 30759 430 30793
rect 245 30721 430 30759
rect 245 30687 320 30721
rect 354 30687 430 30721
rect 245 30649 430 30687
rect 245 30615 320 30649
rect 354 30615 430 30649
rect 245 30577 430 30615
rect 245 30543 320 30577
rect 354 30543 430 30577
rect 245 30505 430 30543
rect 245 30471 320 30505
rect 354 30471 430 30505
rect 245 30433 430 30471
rect 245 30399 320 30433
rect 354 30399 430 30433
rect 245 30361 430 30399
rect 245 30327 320 30361
rect 354 30327 430 30361
rect 245 30289 430 30327
rect 245 30255 320 30289
rect 354 30255 430 30289
rect 245 30217 430 30255
rect 245 30183 320 30217
rect 354 30183 430 30217
rect 245 30145 430 30183
rect 245 30111 320 30145
rect 354 30111 430 30145
rect 245 30073 430 30111
rect 245 30039 320 30073
rect 354 30039 430 30073
rect 245 30001 430 30039
rect 245 29967 320 30001
rect 354 29967 430 30001
rect 245 29929 430 29967
rect 245 29895 320 29929
rect 354 29895 430 29929
rect 245 29857 430 29895
rect 245 29823 320 29857
rect 354 29823 430 29857
rect 245 29785 430 29823
rect 245 29751 320 29785
rect 354 29751 430 29785
rect 245 29713 430 29751
rect 245 29679 320 29713
rect 354 29679 430 29713
rect 245 29641 430 29679
rect 245 29607 320 29641
rect 354 29607 430 29641
rect 245 29569 430 29607
rect 245 29535 320 29569
rect 354 29535 430 29569
rect 245 29497 430 29535
rect 245 29463 320 29497
rect 354 29463 430 29497
rect 245 29425 430 29463
rect 245 29391 320 29425
rect 354 29391 430 29425
rect 245 29353 430 29391
rect 245 29319 320 29353
rect 354 29319 430 29353
rect 245 29281 430 29319
rect 245 29247 320 29281
rect 354 29247 430 29281
rect 245 29209 430 29247
rect 245 29175 320 29209
rect 354 29175 430 29209
rect 245 29137 430 29175
rect 245 29103 320 29137
rect 354 29103 430 29137
rect 245 29065 430 29103
rect 245 29031 320 29065
rect 354 29031 430 29065
rect 245 28993 430 29031
rect 245 28959 320 28993
rect 354 28959 430 28993
rect 245 28921 430 28959
rect 245 28887 320 28921
rect 354 28887 430 28921
rect 245 28849 430 28887
rect 245 28815 320 28849
rect 354 28815 430 28849
rect 245 28777 430 28815
rect 245 28743 320 28777
rect 354 28743 430 28777
rect 245 28705 430 28743
rect 245 28671 320 28705
rect 354 28671 430 28705
rect 245 28633 430 28671
rect 245 28599 320 28633
rect 354 28599 430 28633
rect 245 28561 430 28599
rect 245 28527 320 28561
rect 354 28527 430 28561
rect 245 28489 430 28527
rect 245 28455 320 28489
rect 354 28455 430 28489
rect 245 28417 430 28455
rect 245 28383 320 28417
rect 354 28383 430 28417
rect 245 28345 430 28383
rect 245 28311 320 28345
rect 354 28311 430 28345
rect 245 28273 430 28311
rect 245 28239 320 28273
rect 354 28239 430 28273
rect 245 28201 430 28239
rect 245 28167 320 28201
rect 354 28167 430 28201
rect 245 28129 430 28167
rect 245 28095 320 28129
rect 354 28095 430 28129
rect 245 28057 430 28095
rect 245 28023 320 28057
rect 354 28023 430 28057
rect 245 27985 430 28023
rect 245 27951 320 27985
rect 354 27951 430 27985
rect 245 27913 430 27951
rect 245 27879 320 27913
rect 354 27879 430 27913
rect 245 27841 430 27879
rect 245 27807 320 27841
rect 354 27807 430 27841
rect 245 27769 430 27807
rect 245 27735 320 27769
rect 354 27735 430 27769
rect 245 27697 430 27735
rect 245 27663 320 27697
rect 354 27663 430 27697
rect 245 27625 430 27663
rect 245 27591 320 27625
rect 354 27591 430 27625
rect 245 27553 430 27591
rect 245 27519 320 27553
rect 354 27519 430 27553
rect 245 27481 430 27519
rect 245 27447 320 27481
rect 354 27447 430 27481
rect 245 27409 430 27447
rect 245 27375 320 27409
rect 354 27375 430 27409
rect 245 27337 430 27375
rect 245 27303 320 27337
rect 354 27303 430 27337
rect 245 27265 430 27303
rect 245 27231 320 27265
rect 354 27231 430 27265
rect 245 27193 430 27231
rect 245 27159 320 27193
rect 354 27159 430 27193
rect 245 27121 430 27159
rect 245 27087 320 27121
rect 354 27087 430 27121
rect 245 27049 430 27087
rect 245 27015 320 27049
rect 354 27015 430 27049
rect 245 26977 430 27015
rect 245 26943 320 26977
rect 354 26943 430 26977
rect 245 26905 430 26943
rect 245 26871 320 26905
rect 354 26871 430 26905
rect 245 26833 430 26871
rect 245 26799 320 26833
rect 354 26799 430 26833
rect 245 26761 430 26799
rect 245 26727 320 26761
rect 354 26727 430 26761
rect 245 26689 430 26727
rect 245 26655 320 26689
rect 354 26655 430 26689
rect 245 26617 430 26655
rect 245 26583 320 26617
rect 354 26583 430 26617
rect 245 26545 430 26583
rect 245 26511 320 26545
rect 354 26511 430 26545
rect 245 26473 430 26511
rect 245 26439 320 26473
rect 354 26439 430 26473
rect 245 26401 430 26439
rect 245 26367 320 26401
rect 354 26367 430 26401
rect 245 26329 430 26367
rect 245 26295 320 26329
rect 354 26295 430 26329
rect 245 26257 430 26295
rect 245 26223 320 26257
rect 354 26223 430 26257
rect 245 26185 430 26223
rect 245 26151 320 26185
rect 354 26151 430 26185
rect 245 26113 430 26151
rect 245 26079 320 26113
rect 354 26079 430 26113
rect 245 26041 430 26079
rect 245 26007 320 26041
rect 354 26007 430 26041
rect 245 25969 430 26007
rect 245 25935 320 25969
rect 354 25935 430 25969
rect 245 25897 430 25935
rect 245 25863 320 25897
rect 354 25863 430 25897
rect 245 25825 430 25863
rect 245 25791 320 25825
rect 354 25791 430 25825
rect 245 25753 430 25791
rect 245 25719 320 25753
rect 354 25719 430 25753
rect 245 25681 430 25719
rect 245 25647 320 25681
rect 354 25647 430 25681
rect 245 25609 430 25647
rect 245 25575 320 25609
rect 354 25575 430 25609
rect 245 25537 430 25575
rect 245 25503 320 25537
rect 354 25503 430 25537
rect 245 25465 430 25503
rect 245 25431 320 25465
rect 354 25431 430 25465
rect 245 25393 430 25431
rect 245 25359 320 25393
rect 354 25359 430 25393
rect 245 25321 430 25359
rect 245 25287 320 25321
rect 354 25287 430 25321
rect 245 25249 430 25287
rect 245 25215 320 25249
rect 354 25215 430 25249
rect 245 25177 430 25215
rect 245 25143 320 25177
rect 354 25143 430 25177
rect 245 25105 430 25143
rect 245 25071 320 25105
rect 354 25071 430 25105
rect 245 25033 430 25071
rect 245 24999 320 25033
rect 354 24999 430 25033
rect 245 24961 430 24999
rect 245 24927 320 24961
rect 354 24927 430 24961
rect 245 24889 430 24927
rect 245 24855 320 24889
rect 354 24855 430 24889
rect 245 24817 430 24855
rect 245 24783 320 24817
rect 354 24783 430 24817
rect 245 24745 430 24783
rect 245 24711 320 24745
rect 354 24711 430 24745
rect 245 24673 430 24711
rect 245 24639 320 24673
rect 354 24639 430 24673
rect 245 24601 430 24639
rect 245 24567 320 24601
rect 354 24567 430 24601
rect 245 24529 430 24567
rect 245 24495 320 24529
rect 354 24495 430 24529
rect 245 24457 430 24495
rect 245 24423 320 24457
rect 354 24423 430 24457
rect 245 24385 430 24423
rect 245 24351 320 24385
rect 354 24351 430 24385
rect 245 24313 430 24351
rect 245 24279 320 24313
rect 354 24279 430 24313
rect 245 24241 430 24279
rect 245 24207 320 24241
rect 354 24207 430 24241
rect 245 24169 430 24207
rect 245 24135 320 24169
rect 354 24135 430 24169
rect 245 24097 430 24135
rect 245 24063 320 24097
rect 354 24063 430 24097
rect 245 24025 430 24063
rect 245 23991 320 24025
rect 354 23991 430 24025
rect 245 23953 430 23991
rect 245 23919 320 23953
rect 354 23919 430 23953
rect 245 23881 430 23919
rect 245 23847 320 23881
rect 354 23847 430 23881
rect 245 23809 430 23847
rect 245 23775 320 23809
rect 354 23775 430 23809
rect 245 23737 430 23775
rect 245 23703 320 23737
rect 354 23703 430 23737
rect 245 23665 430 23703
rect 245 23631 320 23665
rect 354 23631 430 23665
rect 245 23593 430 23631
rect 245 23559 320 23593
rect 354 23559 430 23593
rect 245 23521 430 23559
rect 245 23487 320 23521
rect 354 23487 430 23521
rect 245 23449 430 23487
rect 245 23415 320 23449
rect 354 23415 430 23449
rect 245 23377 430 23415
rect 245 23343 320 23377
rect 354 23343 430 23377
rect 245 23305 430 23343
rect 245 23271 320 23305
rect 354 23271 430 23305
rect 245 23233 430 23271
rect 245 23199 320 23233
rect 354 23199 430 23233
rect 245 23161 430 23199
rect 245 23127 320 23161
rect 354 23127 430 23161
rect 245 23089 430 23127
rect 245 23055 320 23089
rect 354 23055 430 23089
rect 245 23017 430 23055
rect 245 22983 320 23017
rect 354 22983 430 23017
rect 245 22945 430 22983
rect 245 22911 320 22945
rect 354 22911 430 22945
rect 245 22873 430 22911
rect 245 22839 320 22873
rect 354 22839 430 22873
rect 245 22801 430 22839
rect 245 22767 320 22801
rect 354 22767 430 22801
rect 245 22729 430 22767
rect 245 22695 320 22729
rect 354 22695 430 22729
rect 245 22657 430 22695
rect 245 22623 320 22657
rect 354 22623 430 22657
rect 245 22585 430 22623
rect 245 22551 320 22585
rect 354 22551 430 22585
rect 245 22513 430 22551
rect 245 22479 320 22513
rect 354 22479 430 22513
rect 245 22441 430 22479
rect 245 22407 320 22441
rect 354 22407 430 22441
rect 245 22369 430 22407
rect 245 22335 320 22369
rect 354 22335 430 22369
rect 245 22297 430 22335
rect 245 22263 320 22297
rect 354 22263 430 22297
rect 245 22225 430 22263
rect 245 22191 320 22225
rect 354 22191 430 22225
rect 245 22153 430 22191
rect 245 22119 320 22153
rect 354 22119 430 22153
rect 245 22081 430 22119
rect 245 22047 320 22081
rect 354 22047 430 22081
rect 245 22009 430 22047
rect 245 21975 320 22009
rect 354 21975 430 22009
rect 245 21937 430 21975
rect 245 21903 320 21937
rect 354 21903 430 21937
rect 245 21865 430 21903
rect 245 21831 320 21865
rect 354 21831 430 21865
rect 245 21793 430 21831
rect 245 21759 320 21793
rect 354 21759 430 21793
rect 245 21721 430 21759
rect 245 21687 320 21721
rect 354 21687 430 21721
rect 245 21649 430 21687
rect 245 21615 320 21649
rect 354 21615 430 21649
rect 245 21577 430 21615
rect 245 21543 320 21577
rect 354 21543 430 21577
rect 245 21505 430 21543
rect 245 21471 320 21505
rect 354 21471 430 21505
rect 245 21433 430 21471
rect 245 21399 320 21433
rect 354 21399 430 21433
rect 245 21361 430 21399
rect 245 21327 320 21361
rect 354 21327 430 21361
rect 245 21289 430 21327
rect 245 21255 320 21289
rect 354 21255 430 21289
rect 245 21217 430 21255
rect 245 21183 320 21217
rect 354 21183 430 21217
rect 245 21145 430 21183
rect 245 21111 320 21145
rect 354 21111 430 21145
rect 245 21073 430 21111
rect 245 21039 320 21073
rect 354 21039 430 21073
rect 245 21001 430 21039
rect 245 20967 320 21001
rect 354 20967 430 21001
rect 245 20929 430 20967
rect 245 20895 320 20929
rect 354 20895 430 20929
rect 245 20857 430 20895
rect 245 20823 320 20857
rect 354 20823 430 20857
rect 245 20785 430 20823
rect 245 20751 320 20785
rect 354 20751 430 20785
rect 245 20713 430 20751
rect 245 20679 320 20713
rect 354 20679 430 20713
rect 245 20641 430 20679
rect 245 20607 320 20641
rect 354 20607 430 20641
rect 245 20569 430 20607
rect 245 20535 320 20569
rect 354 20535 430 20569
rect 245 20497 430 20535
rect 245 20463 320 20497
rect 354 20463 430 20497
rect 245 20425 430 20463
rect 245 20391 320 20425
rect 354 20391 430 20425
rect 245 20353 430 20391
rect 245 20319 320 20353
rect 354 20319 430 20353
rect 245 20281 430 20319
rect 245 20247 320 20281
rect 354 20247 430 20281
rect 245 20209 430 20247
rect 245 20175 320 20209
rect 354 20175 430 20209
rect 245 20137 430 20175
rect 245 20103 320 20137
rect 354 20103 430 20137
rect 245 20065 430 20103
rect 245 20031 320 20065
rect 354 20031 430 20065
rect 245 19993 430 20031
rect 245 19959 320 19993
rect 354 19959 430 19993
rect 245 19921 430 19959
rect 245 19887 320 19921
rect 354 19887 430 19921
rect 245 19849 430 19887
rect 245 19815 320 19849
rect 354 19815 430 19849
rect 245 19777 430 19815
rect 245 19743 320 19777
rect 354 19743 430 19777
rect 245 19705 430 19743
rect 245 19671 320 19705
rect 354 19671 430 19705
rect 245 19633 430 19671
rect 245 19599 320 19633
rect 354 19599 430 19633
rect 245 19561 430 19599
rect 245 19527 320 19561
rect 354 19527 430 19561
rect 245 19489 430 19527
rect 245 19455 320 19489
rect 354 19455 430 19489
rect 245 19417 430 19455
rect 245 19383 320 19417
rect 354 19383 430 19417
rect 245 19345 430 19383
rect 245 19311 320 19345
rect 354 19311 430 19345
rect 245 19273 430 19311
rect 245 19239 320 19273
rect 354 19239 430 19273
rect 245 19201 430 19239
rect 245 19167 320 19201
rect 354 19167 430 19201
rect 245 19129 430 19167
rect 245 19095 320 19129
rect 354 19095 430 19129
rect 245 19057 430 19095
rect 245 19023 320 19057
rect 354 19023 430 19057
rect 245 18985 430 19023
rect 245 18951 320 18985
rect 354 18951 430 18985
rect 245 18913 430 18951
rect 245 18879 320 18913
rect 354 18879 430 18913
rect 245 18841 430 18879
rect 245 18807 320 18841
rect 354 18807 430 18841
rect 245 18769 430 18807
rect 245 18735 320 18769
rect 354 18735 430 18769
rect 245 18697 430 18735
rect 245 18663 320 18697
rect 354 18663 430 18697
rect 245 18625 430 18663
rect 245 18591 320 18625
rect 354 18591 430 18625
rect 245 18553 430 18591
rect 245 18519 320 18553
rect 354 18519 430 18553
rect 245 18481 430 18519
rect 245 18447 320 18481
rect 354 18447 430 18481
rect 245 18409 430 18447
rect 245 18375 320 18409
rect 354 18375 430 18409
rect 245 18337 430 18375
rect 245 18303 320 18337
rect 354 18303 430 18337
rect 245 18265 430 18303
rect 245 18231 320 18265
rect 354 18231 430 18265
rect 245 18193 430 18231
rect 245 18159 320 18193
rect 354 18159 430 18193
rect 245 18121 430 18159
rect 245 18087 320 18121
rect 354 18087 430 18121
rect 245 18049 430 18087
rect 245 18015 320 18049
rect 354 18015 430 18049
rect 245 17977 430 18015
rect 245 17943 320 17977
rect 354 17943 430 17977
rect 245 17905 430 17943
rect 245 17871 320 17905
rect 354 17871 430 17905
rect 245 17833 430 17871
rect 245 17799 320 17833
rect 354 17799 430 17833
rect 245 17761 430 17799
rect 245 17727 320 17761
rect 354 17727 430 17761
rect 245 17689 430 17727
rect 245 17655 320 17689
rect 354 17655 430 17689
rect 245 17617 430 17655
rect 245 17583 320 17617
rect 354 17583 430 17617
rect 245 17545 430 17583
rect 245 17511 320 17545
rect 354 17511 430 17545
rect 245 17473 430 17511
rect 245 17439 320 17473
rect 354 17439 430 17473
rect 245 17401 430 17439
rect 245 17367 320 17401
rect 354 17367 430 17401
rect 245 17329 430 17367
rect 245 17295 320 17329
rect 354 17295 430 17329
rect 245 17257 430 17295
rect 245 17223 320 17257
rect 354 17223 430 17257
rect 245 17185 430 17223
rect 245 17151 320 17185
rect 354 17151 430 17185
rect 245 17113 430 17151
rect 245 17079 320 17113
rect 354 17079 430 17113
rect 245 17041 430 17079
rect 245 17007 320 17041
rect 354 17007 430 17041
rect 245 16969 430 17007
rect 245 16935 320 16969
rect 354 16935 430 16969
rect 245 16897 430 16935
rect 245 16863 320 16897
rect 354 16863 430 16897
rect 245 16825 430 16863
rect 245 16791 320 16825
rect 354 16791 430 16825
rect 245 16753 430 16791
rect 245 16719 320 16753
rect 354 16719 430 16753
rect 245 16681 430 16719
rect 245 16647 320 16681
rect 354 16647 430 16681
rect 245 16609 430 16647
rect 245 16575 320 16609
rect 354 16575 430 16609
rect 245 16537 430 16575
rect 245 16503 320 16537
rect 354 16503 430 16537
rect 245 16465 430 16503
rect 245 16431 320 16465
rect 354 16431 430 16465
rect 245 16393 430 16431
rect 245 16359 320 16393
rect 354 16359 430 16393
rect 245 16321 430 16359
rect 245 16287 320 16321
rect 354 16287 430 16321
rect 245 16249 430 16287
rect 245 16215 320 16249
rect 354 16215 430 16249
rect 245 16177 430 16215
rect 245 16143 320 16177
rect 354 16143 430 16177
rect 245 16105 430 16143
rect 245 16071 320 16105
rect 354 16071 430 16105
rect 245 16033 430 16071
rect 245 15999 320 16033
rect 354 15999 430 16033
rect 245 15961 430 15999
rect 245 15927 320 15961
rect 354 15927 430 15961
rect 245 15889 430 15927
rect 245 15855 320 15889
rect 354 15855 430 15889
rect 245 15817 430 15855
rect 245 15783 320 15817
rect 354 15783 430 15817
rect 245 15745 430 15783
rect 245 15711 320 15745
rect 354 15711 430 15745
rect 245 15673 430 15711
rect 245 15639 320 15673
rect 354 15639 430 15673
rect 245 15601 430 15639
rect 245 15567 320 15601
rect 354 15567 430 15601
rect 245 15529 430 15567
rect 245 15495 320 15529
rect 354 15495 430 15529
rect 245 15457 430 15495
rect 245 15423 320 15457
rect 354 15423 430 15457
rect 245 15385 430 15423
rect 245 15351 320 15385
rect 354 15351 430 15385
rect 245 15313 430 15351
rect 245 15279 320 15313
rect 354 15279 430 15313
rect 245 15241 430 15279
rect 245 15207 320 15241
rect 354 15207 430 15241
rect 245 15169 430 15207
rect 245 15135 320 15169
rect 354 15135 430 15169
rect 245 15097 430 15135
rect 245 15063 320 15097
rect 354 15063 430 15097
rect 245 15025 430 15063
rect 245 14991 320 15025
rect 354 14991 430 15025
rect 245 14953 430 14991
rect 245 14919 320 14953
rect 354 14919 430 14953
rect 245 14881 430 14919
rect 245 14847 320 14881
rect 354 14847 430 14881
rect 245 14809 430 14847
rect 245 14775 320 14809
rect 354 14775 430 14809
rect 245 14737 430 14775
rect 245 14703 320 14737
rect 354 14703 430 14737
rect 245 14665 430 14703
rect 245 14631 320 14665
rect 354 14631 430 14665
rect 245 14593 430 14631
rect 245 14559 320 14593
rect 354 14559 430 14593
rect 245 14521 430 14559
rect 245 14487 320 14521
rect 354 14487 430 14521
rect 245 14449 430 14487
rect 245 14415 320 14449
rect 354 14415 430 14449
rect 245 14377 430 14415
rect 245 14343 320 14377
rect 354 14343 430 14377
rect 245 14305 430 14343
rect 245 14271 320 14305
rect 354 14271 430 14305
rect 245 14233 430 14271
rect 245 14199 320 14233
rect 354 14199 430 14233
rect 245 14161 430 14199
rect 245 14127 320 14161
rect 354 14127 430 14161
rect 245 14089 430 14127
rect 245 14055 320 14089
rect 354 14055 430 14089
rect 245 14017 430 14055
rect 245 13983 320 14017
rect 354 13983 430 14017
rect 245 13945 430 13983
rect 245 13911 320 13945
rect 354 13911 430 13945
rect 245 13873 430 13911
rect 245 13839 320 13873
rect 354 13839 430 13873
rect 245 13801 430 13839
rect 245 13767 320 13801
rect 354 13767 430 13801
rect 245 13729 430 13767
rect 245 13695 320 13729
rect 354 13695 430 13729
rect 245 13657 430 13695
rect 245 13623 320 13657
rect 354 13623 430 13657
rect 245 13585 430 13623
rect 245 13551 320 13585
rect 354 13551 430 13585
rect 245 13513 430 13551
rect 245 13479 320 13513
rect 354 13479 430 13513
rect 245 13441 430 13479
rect 245 13407 320 13441
rect 354 13407 430 13441
rect 245 13369 430 13407
rect 245 13335 320 13369
rect 354 13335 430 13369
rect 245 13297 430 13335
rect 245 13263 320 13297
rect 354 13263 430 13297
rect 245 13225 430 13263
rect 245 13191 320 13225
rect 354 13191 430 13225
rect 245 13153 430 13191
rect 245 13119 320 13153
rect 354 13119 430 13153
rect 245 13081 430 13119
rect 245 13047 320 13081
rect 354 13047 430 13081
rect 245 13009 430 13047
rect 245 12975 320 13009
rect 354 12975 430 13009
rect 245 12937 430 12975
rect 245 12903 320 12937
rect 354 12903 430 12937
rect 245 12865 430 12903
rect 245 12831 320 12865
rect 354 12831 430 12865
rect 245 12793 430 12831
rect 245 12759 320 12793
rect 354 12759 430 12793
rect 245 12721 430 12759
rect 245 12687 320 12721
rect 354 12687 430 12721
rect 245 12649 430 12687
rect 245 12615 320 12649
rect 354 12615 430 12649
rect 245 12577 430 12615
rect 245 12543 320 12577
rect 354 12543 430 12577
rect 245 12505 430 12543
rect 245 12471 320 12505
rect 354 12471 430 12505
rect 245 12433 430 12471
rect 245 12399 320 12433
rect 354 12399 430 12433
rect 245 12361 430 12399
rect 245 12327 320 12361
rect 354 12327 430 12361
rect 245 12289 430 12327
rect 245 12255 320 12289
rect 354 12255 430 12289
rect 245 12217 430 12255
rect 245 12183 320 12217
rect 354 12183 430 12217
rect 245 12145 430 12183
rect 245 12111 320 12145
rect 354 12111 430 12145
rect 245 12073 430 12111
rect 245 12039 320 12073
rect 354 12039 430 12073
rect 245 12001 430 12039
rect 245 11967 320 12001
rect 354 11967 430 12001
rect 245 11929 430 11967
rect 245 11895 320 11929
rect 354 11895 430 11929
rect 245 11857 430 11895
rect 245 11823 320 11857
rect 354 11823 430 11857
rect 245 11785 430 11823
rect 245 11751 320 11785
rect 354 11751 430 11785
rect 245 11713 430 11751
rect 245 11679 320 11713
rect 354 11679 430 11713
rect 245 11641 430 11679
rect 245 11607 320 11641
rect 354 11607 430 11641
rect 245 11569 430 11607
rect 245 11535 320 11569
rect 354 11535 430 11569
rect 245 11497 430 11535
rect 245 11463 320 11497
rect 354 11463 430 11497
rect 245 11425 430 11463
rect 245 11391 320 11425
rect 354 11391 430 11425
rect 245 11353 430 11391
rect 245 11319 320 11353
rect 354 11319 430 11353
rect 245 11281 430 11319
rect 245 11247 320 11281
rect 354 11247 430 11281
rect 245 11209 430 11247
rect 245 11175 320 11209
rect 354 11175 430 11209
rect 245 11137 430 11175
rect 245 11103 320 11137
rect 354 11103 430 11137
rect 245 11065 430 11103
rect 245 11031 320 11065
rect 354 11031 430 11065
rect 245 10993 430 11031
rect 245 10959 320 10993
rect 354 10959 430 10993
rect 245 10921 430 10959
rect 245 10887 320 10921
rect 354 10887 430 10921
rect 245 10849 430 10887
rect 245 10815 320 10849
rect 354 10815 430 10849
rect 245 10777 430 10815
rect 245 10743 320 10777
rect 354 10743 430 10777
rect 245 10705 430 10743
rect 245 10671 320 10705
rect 354 10671 430 10705
rect 245 10633 430 10671
rect 245 10599 320 10633
rect 354 10599 430 10633
rect 245 10561 430 10599
rect 245 10527 320 10561
rect 354 10527 430 10561
rect 245 10489 430 10527
rect 245 10455 320 10489
rect 354 10455 430 10489
rect 245 10417 430 10455
rect 245 10383 320 10417
rect 354 10383 430 10417
rect 245 10345 430 10383
rect 245 10311 320 10345
rect 354 10311 430 10345
rect 245 10273 430 10311
rect 245 10239 320 10273
rect 354 10239 430 10273
rect 245 10201 430 10239
rect 245 10167 320 10201
rect 354 10167 430 10201
rect 245 10129 430 10167
rect 245 10095 320 10129
rect 354 10095 430 10129
rect 245 10057 430 10095
rect 245 10023 320 10057
rect 354 10023 430 10057
rect 245 9985 430 10023
rect 245 9951 320 9985
rect 354 9951 430 9985
rect 245 9913 430 9951
tri 757 35953 773 35969 se
rect 773 35953 14198 35969
tri 14198 35953 14219 35974 sw
rect 757 35933 14219 35953
rect 757 35902 886 35933
tri 886 35902 917 35933 nw
tri 14059 35902 14090 35933 ne
rect 14090 35902 14219 35933
rect 757 35884 877 35902
tri 877 35893 886 35902 nw
tri 14090 35893 14099 35902 ne
rect 757 35850 807 35884
rect 841 35850 877 35884
rect 757 35812 877 35850
rect 757 35778 807 35812
rect 841 35778 877 35812
rect 757 35740 877 35778
rect 757 35706 807 35740
rect 841 35706 877 35740
rect 757 35668 877 35706
rect 757 35634 807 35668
rect 841 35634 877 35668
rect 757 35596 877 35634
rect 757 35562 807 35596
rect 841 35562 877 35596
rect 757 35524 877 35562
rect 757 35490 807 35524
rect 841 35490 877 35524
rect 757 35452 877 35490
rect 757 35418 807 35452
rect 841 35418 877 35452
rect 757 35380 877 35418
rect 757 35346 807 35380
rect 841 35346 877 35380
rect 757 35308 877 35346
rect 757 35274 807 35308
rect 841 35274 877 35308
rect 757 35236 877 35274
rect 757 35202 807 35236
rect 841 35202 877 35236
rect 757 35164 877 35202
rect 757 35130 807 35164
rect 841 35130 877 35164
rect 757 35092 877 35130
rect 757 35058 807 35092
rect 841 35058 877 35092
rect 757 35020 877 35058
rect 757 34986 807 35020
rect 841 34986 877 35020
rect 757 34948 877 34986
rect 757 34914 807 34948
rect 841 34914 877 34948
rect 757 34876 877 34914
rect 757 34842 807 34876
rect 841 34842 877 34876
rect 757 34804 877 34842
rect 757 34770 807 34804
rect 841 34770 877 34804
rect 757 34732 877 34770
rect 757 34698 807 34732
rect 841 34698 877 34732
rect 757 34660 877 34698
rect 14099 35805 14219 35902
rect 14099 35771 14142 35805
rect 14176 35771 14219 35805
rect 14099 35733 14219 35771
rect 14099 35699 14142 35733
rect 14176 35699 14219 35733
rect 14099 35661 14219 35699
rect 14099 35627 14142 35661
rect 14176 35627 14219 35661
rect 14099 35589 14219 35627
rect 14099 35555 14142 35589
rect 14176 35555 14219 35589
rect 14099 35517 14219 35555
rect 14099 35483 14142 35517
rect 14176 35483 14219 35517
rect 14099 35445 14219 35483
rect 14099 35411 14142 35445
rect 14176 35411 14219 35445
rect 14099 35373 14219 35411
rect 14099 35339 14142 35373
rect 14176 35339 14219 35373
rect 14099 35301 14219 35339
rect 14099 35267 14142 35301
rect 14176 35267 14219 35301
rect 14099 35229 14219 35267
rect 14099 35195 14142 35229
rect 14176 35195 14219 35229
rect 14099 35157 14219 35195
rect 14099 35123 14142 35157
rect 14176 35123 14219 35157
rect 14099 35085 14219 35123
rect 14099 35051 14142 35085
rect 14176 35051 14219 35085
rect 14099 35013 14219 35051
rect 14099 34979 14142 35013
rect 14176 34979 14219 35013
rect 14099 34941 14219 34979
rect 14099 34907 14142 34941
rect 14176 34907 14219 34941
rect 14099 34869 14219 34907
rect 14099 34835 14142 34869
rect 14176 34835 14219 34869
rect 14099 34797 14219 34835
rect 14099 34763 14142 34797
rect 14176 34763 14219 34797
rect 14099 34725 14219 34763
rect 757 34626 807 34660
rect 841 34626 877 34660
rect 757 34588 877 34626
rect 757 34554 807 34588
rect 841 34554 877 34588
rect 757 34516 877 34554
rect 757 34482 807 34516
rect 841 34482 877 34516
rect 757 34444 877 34482
rect 757 34410 807 34444
rect 841 34410 877 34444
rect 757 34372 877 34410
rect 757 34338 807 34372
rect 841 34338 877 34372
rect 757 34300 877 34338
rect 757 34266 807 34300
rect 841 34266 877 34300
rect 757 34228 877 34266
rect 757 34194 807 34228
rect 841 34194 877 34228
rect 757 34156 877 34194
rect 757 34122 807 34156
rect 841 34122 877 34156
rect 757 34084 877 34122
rect 757 34050 807 34084
rect 841 34050 877 34084
rect 757 34012 877 34050
rect 757 33978 807 34012
rect 841 33978 877 34012
rect 757 33940 877 33978
rect 757 33906 807 33940
rect 841 33906 877 33940
rect 757 33868 877 33906
rect 757 33834 807 33868
rect 841 33834 877 33868
rect 757 33796 877 33834
rect 757 33762 807 33796
rect 841 33762 877 33796
rect 757 33724 877 33762
rect 757 33690 807 33724
rect 841 33690 877 33724
rect 757 33652 877 33690
rect 757 33618 807 33652
rect 841 33618 877 33652
rect 757 33580 877 33618
rect 757 33546 807 33580
rect 841 33546 877 33580
rect 757 33508 877 33546
rect 757 33474 807 33508
rect 841 33474 877 33508
rect 757 33436 877 33474
rect 757 33402 807 33436
rect 841 33402 877 33436
rect 757 33364 877 33402
rect 757 33330 807 33364
rect 841 33330 877 33364
rect 757 33292 877 33330
rect 757 33258 807 33292
rect 841 33258 877 33292
rect 757 33220 877 33258
rect 757 33186 807 33220
rect 841 33186 877 33220
rect 757 33148 877 33186
rect 757 33114 807 33148
rect 841 33114 877 33148
rect 757 33076 877 33114
rect 757 33042 807 33076
rect 841 33042 877 33076
rect 757 33004 877 33042
rect 757 32970 807 33004
rect 841 32970 877 33004
rect 757 32932 877 32970
rect 757 32898 807 32932
rect 841 32898 877 32932
rect 757 32860 877 32898
rect 757 32826 807 32860
rect 841 32826 877 32860
rect 757 32788 877 32826
rect 757 32754 807 32788
rect 841 32754 877 32788
rect 757 32716 877 32754
rect 757 32682 807 32716
rect 841 32682 877 32716
rect 757 32644 877 32682
rect 757 32610 807 32644
rect 841 32610 877 32644
rect 757 32572 877 32610
rect 757 32538 807 32572
rect 841 32538 877 32572
rect 757 32500 877 32538
rect 757 32466 807 32500
rect 841 32466 877 32500
rect 757 32428 877 32466
rect 757 32394 807 32428
rect 841 32394 877 32428
rect 757 32356 877 32394
rect 757 32322 807 32356
rect 841 32322 877 32356
rect 757 32284 877 32322
rect 757 32250 807 32284
rect 841 32250 877 32284
rect 757 32212 877 32250
rect 757 32178 807 32212
rect 841 32178 877 32212
rect 757 32140 877 32178
rect 757 32106 807 32140
rect 841 32106 877 32140
rect 757 32068 877 32106
rect 757 32034 807 32068
rect 841 32034 877 32068
rect 757 31996 877 32034
rect 757 31962 807 31996
rect 841 31962 877 31996
rect 757 31924 877 31962
rect 757 31890 807 31924
rect 841 31890 877 31924
rect 757 31852 877 31890
rect 757 31818 807 31852
rect 841 31818 877 31852
rect 757 31780 877 31818
rect 757 31746 807 31780
rect 841 31746 877 31780
rect 757 31708 877 31746
rect 757 31674 807 31708
rect 841 31674 877 31708
rect 757 31636 877 31674
rect 757 31602 807 31636
rect 841 31602 877 31636
rect 757 31564 877 31602
rect 757 31530 807 31564
rect 841 31530 877 31564
rect 757 31492 877 31530
rect 757 31458 807 31492
rect 841 31458 877 31492
rect 757 31420 877 31458
rect 757 31386 807 31420
rect 841 31386 877 31420
rect 757 31348 877 31386
rect 757 31314 807 31348
rect 841 31314 877 31348
rect 757 31276 877 31314
rect 757 31242 807 31276
rect 841 31242 877 31276
rect 757 31204 877 31242
rect 757 31170 807 31204
rect 841 31170 877 31204
rect 757 31132 877 31170
rect 757 31098 807 31132
rect 841 31098 877 31132
rect 757 31060 877 31098
rect 757 31026 807 31060
rect 841 31026 877 31060
rect 757 30988 877 31026
rect 757 30954 807 30988
rect 841 30954 877 30988
rect 757 30916 877 30954
rect 757 30882 807 30916
rect 841 30882 877 30916
rect 757 30844 877 30882
rect 757 30810 807 30844
rect 841 30810 877 30844
rect 757 30772 877 30810
rect 757 30738 807 30772
rect 841 30738 877 30772
rect 757 30700 877 30738
rect 757 30666 807 30700
rect 841 30666 877 30700
rect 757 30628 877 30666
rect 757 30594 807 30628
rect 841 30594 877 30628
rect 757 30556 877 30594
rect 757 30522 807 30556
rect 841 30522 877 30556
rect 757 30484 877 30522
rect 757 30450 807 30484
rect 841 30450 877 30484
rect 757 30412 877 30450
rect 757 30378 807 30412
rect 841 30378 877 30412
rect 757 30340 877 30378
rect 757 30306 807 30340
rect 841 30306 877 30340
rect 757 30268 877 30306
rect 757 30234 807 30268
rect 841 30234 877 30268
rect 757 30196 877 30234
rect 757 30162 807 30196
rect 841 30162 877 30196
rect 757 30124 877 30162
rect 757 30090 807 30124
rect 841 30090 877 30124
rect 757 30052 877 30090
rect 757 30018 807 30052
rect 841 30018 877 30052
rect 757 29980 877 30018
rect 757 29946 807 29980
rect 841 29946 877 29980
rect 757 29908 877 29946
rect 757 29874 807 29908
rect 841 29874 877 29908
rect 757 29836 877 29874
rect 757 29802 807 29836
rect 841 29802 877 29836
rect 757 29764 877 29802
rect 757 29730 807 29764
rect 841 29730 877 29764
rect 757 29692 877 29730
rect 757 29658 807 29692
rect 841 29658 877 29692
rect 757 29620 877 29658
rect 757 29586 807 29620
rect 841 29586 877 29620
rect 757 29548 877 29586
rect 757 29514 807 29548
rect 841 29514 877 29548
rect 757 29476 877 29514
rect 757 29442 807 29476
rect 841 29442 877 29476
rect 757 29404 877 29442
rect 757 29370 807 29404
rect 841 29370 877 29404
rect 757 29332 877 29370
rect 757 29298 807 29332
rect 841 29298 877 29332
rect 757 29260 877 29298
rect 757 29226 807 29260
rect 841 29226 877 29260
rect 757 29188 877 29226
rect 757 29154 807 29188
rect 841 29154 877 29188
rect 757 29116 877 29154
rect 757 29082 807 29116
rect 841 29082 877 29116
rect 757 29044 877 29082
rect 757 29010 807 29044
rect 841 29010 877 29044
rect 757 28972 877 29010
rect 757 28938 807 28972
rect 841 28938 877 28972
rect 757 28900 877 28938
rect 757 28866 807 28900
rect 841 28866 877 28900
rect 757 28828 877 28866
rect 757 28794 807 28828
rect 841 28794 877 28828
rect 757 28756 877 28794
rect 757 28722 807 28756
rect 841 28722 877 28756
rect 757 28684 877 28722
rect 757 28650 807 28684
rect 841 28650 877 28684
rect 757 28612 877 28650
rect 757 28578 807 28612
rect 841 28578 877 28612
rect 757 28540 877 28578
rect 757 28506 807 28540
rect 841 28506 877 28540
rect 757 28468 877 28506
rect 757 28434 807 28468
rect 841 28434 877 28468
rect 757 28396 877 28434
rect 757 28362 807 28396
rect 841 28362 877 28396
rect 757 28324 877 28362
rect 757 28290 807 28324
rect 841 28290 877 28324
rect 757 28252 877 28290
rect 757 28218 807 28252
rect 841 28218 877 28252
rect 757 28180 877 28218
rect 757 28146 807 28180
rect 841 28146 877 28180
rect 757 28108 877 28146
rect 757 28074 807 28108
rect 841 28074 877 28108
rect 757 28036 877 28074
rect 757 28002 807 28036
rect 841 28002 877 28036
rect 757 27964 877 28002
rect 757 27930 807 27964
rect 841 27930 877 27964
rect 757 27892 877 27930
rect 757 27858 807 27892
rect 841 27858 877 27892
rect 757 27820 877 27858
rect 757 27786 807 27820
rect 841 27786 877 27820
rect 757 27748 877 27786
rect 757 27714 807 27748
rect 841 27714 877 27748
rect 757 27676 877 27714
rect 757 27642 807 27676
rect 841 27642 877 27676
rect 757 27604 877 27642
rect 757 27570 807 27604
rect 841 27570 877 27604
rect 757 27532 877 27570
rect 757 27498 807 27532
rect 841 27498 877 27532
rect 757 27460 877 27498
rect 757 27426 807 27460
rect 841 27426 877 27460
rect 757 27388 877 27426
rect 757 27354 807 27388
rect 841 27354 877 27388
rect 757 27316 877 27354
rect 757 27282 807 27316
rect 841 27282 877 27316
rect 757 27244 877 27282
rect 757 27210 807 27244
rect 841 27210 877 27244
rect 757 27172 877 27210
rect 757 27138 807 27172
rect 841 27138 877 27172
rect 757 27100 877 27138
rect 757 27066 807 27100
rect 841 27066 877 27100
rect 757 27028 877 27066
rect 757 26994 807 27028
rect 841 26994 877 27028
rect 757 26956 877 26994
rect 757 26922 807 26956
rect 841 26922 877 26956
rect 757 26884 877 26922
rect 757 26850 807 26884
rect 841 26850 877 26884
rect 757 26812 877 26850
rect 757 26778 807 26812
rect 841 26778 877 26812
rect 757 26740 877 26778
rect 757 26706 807 26740
rect 841 26706 877 26740
rect 757 26668 877 26706
rect 757 26634 807 26668
rect 841 26634 877 26668
rect 757 26596 877 26634
rect 757 26562 807 26596
rect 841 26562 877 26596
rect 757 26524 877 26562
rect 757 26490 807 26524
rect 841 26490 877 26524
rect 757 26452 877 26490
rect 757 26418 807 26452
rect 841 26418 877 26452
rect 757 26380 877 26418
rect 757 26346 807 26380
rect 841 26346 877 26380
rect 757 26308 877 26346
rect 757 26274 807 26308
rect 841 26274 877 26308
rect 757 26236 877 26274
rect 757 26202 807 26236
rect 841 26202 877 26236
rect 757 26164 877 26202
rect 757 26130 807 26164
rect 841 26130 877 26164
rect 757 26092 877 26130
rect 757 26058 807 26092
rect 841 26058 877 26092
rect 757 26020 877 26058
rect 757 25986 807 26020
rect 841 25986 877 26020
rect 757 25948 877 25986
rect 757 25914 807 25948
rect 841 25914 877 25948
rect 757 25876 877 25914
rect 757 25842 807 25876
rect 841 25842 877 25876
rect 757 25804 877 25842
rect 757 25770 807 25804
rect 841 25770 877 25804
rect 757 25732 877 25770
rect 757 25698 807 25732
rect 841 25698 877 25732
rect 757 25660 877 25698
rect 757 25626 807 25660
rect 841 25626 877 25660
rect 757 25588 877 25626
rect 757 25554 807 25588
rect 841 25554 877 25588
rect 757 25516 877 25554
rect 757 25482 807 25516
rect 841 25482 877 25516
rect 757 25444 877 25482
rect 757 25410 807 25444
rect 841 25410 877 25444
rect 757 25372 877 25410
rect 757 25338 807 25372
rect 841 25338 877 25372
rect 757 25300 877 25338
rect 757 25266 807 25300
rect 841 25266 877 25300
rect 757 25228 877 25266
rect 757 25194 807 25228
rect 841 25194 877 25228
rect 757 25156 877 25194
rect 757 25122 807 25156
rect 841 25122 877 25156
rect 757 25084 877 25122
rect 757 25050 807 25084
rect 841 25050 877 25084
rect 757 25012 877 25050
rect 757 24978 807 25012
rect 841 24978 877 25012
rect 757 24940 877 24978
rect 757 24906 807 24940
rect 841 24906 877 24940
rect 757 24868 877 24906
rect 757 24834 807 24868
rect 841 24834 877 24868
rect 757 24796 877 24834
rect 757 24762 807 24796
rect 841 24762 877 24796
rect 757 24724 877 24762
rect 757 24690 807 24724
rect 841 24690 877 24724
rect 757 24652 877 24690
rect 757 24618 807 24652
rect 841 24618 877 24652
rect 757 24580 877 24618
rect 757 24546 807 24580
rect 841 24546 877 24580
rect 757 24508 877 24546
rect 757 24474 807 24508
rect 841 24474 877 24508
rect 757 24436 877 24474
rect 757 24402 807 24436
rect 841 24402 877 24436
rect 757 24364 877 24402
rect 757 24330 807 24364
rect 841 24330 877 24364
rect 757 24292 877 24330
rect 757 24258 807 24292
rect 841 24258 877 24292
rect 757 24220 877 24258
rect 757 24186 807 24220
rect 841 24186 877 24220
rect 757 24148 877 24186
rect 757 24114 807 24148
rect 841 24114 877 24148
rect 757 24076 877 24114
rect 757 24042 807 24076
rect 841 24042 877 24076
rect 757 24004 877 24042
rect 757 23970 807 24004
rect 841 23970 877 24004
rect 757 23932 877 23970
rect 757 23898 807 23932
rect 841 23898 877 23932
rect 757 23860 877 23898
rect 757 23826 807 23860
rect 841 23826 877 23860
rect 757 23788 877 23826
rect 757 23754 807 23788
rect 841 23754 877 23788
rect 757 23716 877 23754
rect 757 23682 807 23716
rect 841 23682 877 23716
rect 757 23644 877 23682
rect 757 23610 807 23644
rect 841 23610 877 23644
rect 757 23572 877 23610
rect 757 23538 807 23572
rect 841 23538 877 23572
rect 757 23500 877 23538
rect 757 23466 807 23500
rect 841 23466 877 23500
rect 757 23428 877 23466
rect 757 23394 807 23428
rect 841 23394 877 23428
rect 757 23356 877 23394
rect 757 23322 807 23356
rect 841 23322 877 23356
rect 757 23284 877 23322
rect 757 23250 807 23284
rect 841 23250 877 23284
rect 757 23212 877 23250
rect 757 23178 807 23212
rect 841 23178 877 23212
rect 757 23140 877 23178
rect 757 23106 807 23140
rect 841 23106 877 23140
rect 757 23068 877 23106
rect 757 23034 807 23068
rect 841 23034 877 23068
rect 757 22996 877 23034
rect 757 22962 807 22996
rect 841 22962 877 22996
rect 757 22924 877 22962
rect 757 22890 807 22924
rect 841 22890 877 22924
rect 757 22852 877 22890
rect 757 22818 807 22852
rect 841 22818 877 22852
rect 757 22780 877 22818
rect 757 22746 807 22780
rect 841 22746 877 22780
rect 757 22708 877 22746
rect 757 22674 807 22708
rect 841 22674 877 22708
rect 757 22636 877 22674
rect 757 22602 807 22636
rect 841 22602 877 22636
rect 757 22564 877 22602
rect 757 22530 807 22564
rect 841 22530 877 22564
rect 757 22492 877 22530
rect 757 22458 807 22492
rect 841 22458 877 22492
rect 757 22420 877 22458
rect 757 22386 807 22420
rect 841 22386 877 22420
rect 757 22348 877 22386
rect 757 22314 807 22348
rect 841 22314 877 22348
rect 757 22276 877 22314
rect 757 22242 807 22276
rect 841 22242 877 22276
rect 757 22204 877 22242
rect 757 22170 807 22204
rect 841 22170 877 22204
rect 757 22132 877 22170
rect 757 22098 807 22132
rect 841 22098 877 22132
rect 757 22060 877 22098
rect 757 22026 807 22060
rect 841 22026 877 22060
rect 757 21988 877 22026
rect 757 21954 807 21988
rect 841 21954 877 21988
rect 757 21916 877 21954
rect 757 21882 807 21916
rect 841 21882 877 21916
rect 757 21844 877 21882
rect 757 21810 807 21844
rect 841 21810 877 21844
rect 757 21772 877 21810
rect 757 21738 807 21772
rect 841 21738 877 21772
rect 757 21700 877 21738
rect 757 21666 807 21700
rect 841 21666 877 21700
rect 757 21628 877 21666
rect 757 21594 807 21628
rect 841 21594 877 21628
rect 757 21556 877 21594
rect 757 21522 807 21556
rect 841 21522 877 21556
rect 757 21484 877 21522
rect 757 21450 807 21484
rect 841 21450 877 21484
rect 757 21412 877 21450
rect 757 21378 807 21412
rect 841 21378 877 21412
rect 757 21340 877 21378
rect 757 21306 807 21340
rect 841 21306 877 21340
rect 757 21268 877 21306
rect 757 21234 807 21268
rect 841 21234 877 21268
rect 757 21196 877 21234
rect 757 21162 807 21196
rect 841 21162 877 21196
rect 757 21124 877 21162
rect 757 21090 807 21124
rect 841 21090 877 21124
rect 757 21052 877 21090
rect 757 21018 807 21052
rect 841 21018 877 21052
rect 757 20980 877 21018
rect 757 20946 807 20980
rect 841 20946 877 20980
rect 757 20908 877 20946
rect 757 20874 807 20908
rect 841 20874 877 20908
rect 757 20836 877 20874
rect 757 20802 807 20836
rect 841 20802 877 20836
rect 757 20764 877 20802
rect 757 20730 807 20764
rect 841 20730 877 20764
rect 757 20692 877 20730
rect 757 20658 807 20692
rect 841 20658 877 20692
rect 757 20620 877 20658
rect 757 20586 807 20620
rect 841 20586 877 20620
rect 757 20548 877 20586
rect 757 20514 807 20548
rect 841 20514 877 20548
rect 757 20476 877 20514
rect 757 20442 807 20476
rect 841 20442 877 20476
rect 757 20404 877 20442
rect 757 20370 807 20404
rect 841 20370 877 20404
rect 757 20332 877 20370
rect 757 20298 807 20332
rect 841 20298 877 20332
rect 757 20260 877 20298
rect 757 20226 807 20260
rect 841 20226 877 20260
rect 757 20188 877 20226
rect 757 20154 807 20188
rect 841 20154 877 20188
rect 757 20116 877 20154
rect 757 20082 807 20116
rect 841 20082 877 20116
rect 757 20044 877 20082
rect 757 20010 807 20044
rect 841 20010 877 20044
rect 757 19972 877 20010
rect 757 19938 807 19972
rect 841 19938 877 19972
rect 757 19900 877 19938
rect 757 19866 807 19900
rect 841 19866 877 19900
rect 757 19828 877 19866
rect 757 19794 807 19828
rect 841 19794 877 19828
rect 757 19756 877 19794
rect 757 19722 807 19756
rect 841 19722 877 19756
rect 757 19684 877 19722
rect 757 19650 807 19684
rect 841 19650 877 19684
rect 757 19612 877 19650
rect 757 19578 807 19612
rect 841 19578 877 19612
rect 757 19540 877 19578
rect 757 19506 807 19540
rect 841 19506 877 19540
rect 757 19468 877 19506
rect 757 19434 807 19468
rect 841 19434 877 19468
rect 757 19396 877 19434
rect 757 19362 807 19396
rect 841 19362 877 19396
rect 757 19324 877 19362
rect 757 19290 807 19324
rect 841 19290 877 19324
rect 757 19252 877 19290
rect 757 19218 807 19252
rect 841 19218 877 19252
rect 757 19180 877 19218
rect 757 19146 807 19180
rect 841 19146 877 19180
rect 757 19108 877 19146
rect 757 19074 807 19108
rect 841 19074 877 19108
rect 757 19036 877 19074
rect 757 19002 807 19036
rect 841 19002 877 19036
rect 757 18964 877 19002
rect 757 18930 807 18964
rect 841 18930 877 18964
rect 757 18892 877 18930
rect 757 18858 807 18892
rect 841 18858 877 18892
rect 757 18820 877 18858
rect 757 18786 807 18820
rect 841 18786 877 18820
rect 757 18748 877 18786
rect 757 18714 807 18748
rect 841 18714 877 18748
rect 757 18676 877 18714
rect 757 18642 807 18676
rect 841 18642 877 18676
rect 757 18604 877 18642
rect 757 18570 807 18604
rect 841 18570 877 18604
rect 757 18532 877 18570
rect 757 18498 807 18532
rect 841 18498 877 18532
rect 757 18460 877 18498
rect 757 18426 807 18460
rect 841 18426 877 18460
rect 757 18388 877 18426
rect 757 18354 807 18388
rect 841 18354 877 18388
rect 757 18316 877 18354
rect 757 18282 807 18316
rect 841 18282 877 18316
rect 757 18244 877 18282
rect 757 18210 807 18244
rect 841 18210 877 18244
rect 757 18172 877 18210
rect 757 18138 807 18172
rect 841 18138 877 18172
rect 757 18100 877 18138
rect 757 18066 807 18100
rect 841 18066 877 18100
rect 757 18028 877 18066
rect 757 17994 807 18028
rect 841 17994 877 18028
rect 757 17956 877 17994
rect 757 17922 807 17956
rect 841 17922 877 17956
rect 757 17884 877 17922
rect 757 17850 807 17884
rect 841 17850 877 17884
rect 757 17812 877 17850
rect 757 17778 807 17812
rect 841 17778 877 17812
rect 757 17740 877 17778
rect 757 17706 807 17740
rect 841 17706 877 17740
rect 757 17668 877 17706
rect 757 17634 807 17668
rect 841 17634 877 17668
rect 757 17596 877 17634
rect 757 17562 807 17596
rect 841 17562 877 17596
rect 757 17524 877 17562
rect 757 17490 807 17524
rect 841 17490 877 17524
rect 757 17452 877 17490
rect 757 17418 807 17452
rect 841 17418 877 17452
rect 757 17380 877 17418
rect 757 17346 807 17380
rect 841 17346 877 17380
rect 757 17308 877 17346
rect 757 17274 807 17308
rect 841 17274 877 17308
rect 757 17236 877 17274
rect 757 17202 807 17236
rect 841 17202 877 17236
rect 757 17164 877 17202
rect 757 17130 807 17164
rect 841 17130 877 17164
rect 757 17092 877 17130
rect 757 17058 807 17092
rect 841 17058 877 17092
rect 757 17020 877 17058
rect 757 16986 807 17020
rect 841 16986 877 17020
rect 757 16948 877 16986
rect 757 16914 807 16948
rect 841 16914 877 16948
rect 757 16876 877 16914
rect 757 16842 807 16876
rect 841 16842 877 16876
rect 757 16804 877 16842
rect 757 16770 807 16804
rect 841 16770 877 16804
rect 757 16732 877 16770
rect 757 16698 807 16732
rect 841 16698 877 16732
rect 757 16660 877 16698
rect 757 16626 807 16660
rect 841 16626 877 16660
rect 757 16588 877 16626
rect 757 16554 807 16588
rect 841 16554 877 16588
rect 757 16516 877 16554
rect 757 16482 807 16516
rect 841 16482 877 16516
rect 757 16444 877 16482
rect 757 16410 807 16444
rect 841 16410 877 16444
rect 757 16372 877 16410
rect 757 16338 807 16372
rect 841 16338 877 16372
rect 757 16300 877 16338
rect 757 16266 807 16300
rect 841 16266 877 16300
rect 757 16228 877 16266
rect 757 16194 807 16228
rect 841 16194 877 16228
rect 757 16156 877 16194
rect 757 16122 807 16156
rect 841 16122 877 16156
rect 757 16084 877 16122
rect 757 16050 807 16084
rect 841 16050 877 16084
rect 757 16012 877 16050
rect 757 15978 807 16012
rect 841 15978 877 16012
rect 757 15940 877 15978
rect 757 15906 807 15940
rect 841 15906 877 15940
rect 757 15868 877 15906
rect 757 15834 807 15868
rect 841 15834 877 15868
rect 757 15796 877 15834
rect 757 15762 807 15796
rect 841 15762 877 15796
rect 757 15724 877 15762
rect 757 15690 807 15724
rect 841 15690 877 15724
rect 757 15652 877 15690
rect 757 15618 807 15652
rect 841 15618 877 15652
rect 757 15580 877 15618
rect 757 15546 807 15580
rect 841 15546 877 15580
rect 757 15508 877 15546
rect 757 15474 807 15508
rect 841 15474 877 15508
rect 757 15436 877 15474
rect 757 15402 807 15436
rect 841 15402 877 15436
rect 757 15364 877 15402
rect 757 15330 807 15364
rect 841 15330 877 15364
rect 757 15292 877 15330
rect 757 15258 807 15292
rect 841 15258 877 15292
rect 757 15220 877 15258
rect 757 15186 807 15220
rect 841 15186 877 15220
rect 757 15148 877 15186
rect 757 15114 807 15148
rect 841 15114 877 15148
rect 757 15076 877 15114
rect 757 15042 807 15076
rect 841 15042 877 15076
rect 757 15004 877 15042
rect 757 14970 807 15004
rect 841 14970 877 15004
rect 757 14932 877 14970
rect 757 14898 807 14932
rect 841 14898 877 14932
rect 757 14860 877 14898
rect 757 14826 807 14860
rect 841 14826 877 14860
rect 757 14788 877 14826
rect 757 14754 807 14788
rect 841 14754 877 14788
rect 757 14716 877 14754
rect 757 14682 807 14716
rect 841 14682 877 14716
rect 757 14644 877 14682
rect 757 14610 807 14644
rect 841 14610 877 14644
rect 757 14572 877 14610
rect 757 14538 807 14572
rect 841 14538 877 14572
rect 757 14500 877 14538
rect 757 14466 807 14500
rect 841 14466 877 14500
rect 757 14428 877 14466
rect 757 14394 807 14428
rect 841 14394 877 14428
rect 757 14356 877 14394
rect 757 14322 807 14356
rect 841 14322 877 14356
rect 757 14284 877 14322
rect 757 14250 807 14284
rect 841 14250 877 14284
rect 757 14212 877 14250
rect 757 14178 807 14212
rect 841 14178 877 14212
rect 757 14140 877 14178
rect 757 14106 807 14140
rect 841 14106 877 14140
rect 757 14068 877 14106
rect 757 14034 807 14068
rect 841 14034 877 14068
rect 757 13996 877 14034
rect 757 13962 807 13996
rect 841 13962 877 13996
rect 757 13924 877 13962
rect 757 13890 807 13924
rect 841 13890 877 13924
rect 757 13852 877 13890
rect 757 13818 807 13852
rect 841 13818 877 13852
rect 757 13780 877 13818
rect 757 13746 807 13780
rect 841 13746 877 13780
rect 757 13708 877 13746
rect 757 13674 807 13708
rect 841 13674 877 13708
rect 757 13636 877 13674
rect 757 13602 807 13636
rect 841 13602 877 13636
rect 757 13564 877 13602
rect 757 13530 807 13564
rect 841 13530 877 13564
rect 757 13492 877 13530
rect 757 13458 807 13492
rect 841 13458 877 13492
rect 757 13420 877 13458
rect 757 13386 807 13420
rect 841 13386 877 13420
rect 757 13348 877 13386
rect 757 13314 807 13348
rect 841 13314 877 13348
rect 757 13276 877 13314
rect 757 13242 807 13276
rect 841 13242 877 13276
rect 757 13204 877 13242
rect 757 13170 807 13204
rect 841 13170 877 13204
rect 757 13132 877 13170
rect 757 13098 807 13132
rect 841 13098 877 13132
rect 757 13060 877 13098
rect 757 13026 807 13060
rect 841 13026 877 13060
rect 757 12988 877 13026
rect 757 12954 807 12988
rect 841 12954 877 12988
rect 757 12916 877 12954
rect 757 12882 807 12916
rect 841 12882 877 12916
rect 757 12844 877 12882
rect 757 12810 807 12844
rect 841 12810 877 12844
rect 757 12772 877 12810
rect 757 12738 807 12772
rect 841 12738 877 12772
rect 757 12700 877 12738
rect 757 12666 807 12700
rect 841 12666 877 12700
rect 757 12628 877 12666
rect 757 12594 807 12628
rect 841 12594 877 12628
rect 757 12556 877 12594
rect 757 12522 807 12556
rect 841 12522 877 12556
rect 757 12484 877 12522
rect 757 12450 807 12484
rect 841 12450 877 12484
rect 757 12412 877 12450
rect 757 12378 807 12412
rect 841 12378 877 12412
rect 757 12340 877 12378
rect 757 12306 807 12340
rect 841 12306 877 12340
rect 757 12268 877 12306
rect 757 12234 807 12268
rect 841 12234 877 12268
rect 757 12196 877 12234
rect 757 12162 807 12196
rect 841 12162 877 12196
rect 757 12124 877 12162
rect 757 12090 807 12124
rect 841 12090 877 12124
rect 757 12052 877 12090
rect 757 12018 807 12052
rect 841 12018 877 12052
rect 757 11980 877 12018
rect 757 11946 807 11980
rect 841 11946 877 11980
rect 757 11908 877 11946
rect 757 11874 807 11908
rect 841 11874 877 11908
rect 757 11836 877 11874
rect 757 11802 807 11836
rect 841 11802 877 11836
rect 757 11764 877 11802
rect 757 11730 807 11764
rect 841 11730 877 11764
rect 757 11692 877 11730
rect 757 11658 807 11692
rect 841 11658 877 11692
rect 757 11620 877 11658
rect 757 11586 807 11620
rect 841 11586 877 11620
rect 757 11548 877 11586
rect 757 11514 807 11548
rect 841 11514 877 11548
rect 757 11476 877 11514
rect 757 11442 807 11476
rect 841 11442 877 11476
rect 757 11404 877 11442
rect 757 11370 807 11404
rect 841 11370 877 11404
rect 757 11332 877 11370
rect 757 11298 807 11332
rect 841 11298 877 11332
rect 757 11260 877 11298
rect 757 11226 807 11260
rect 841 11226 877 11260
rect 757 11188 877 11226
rect 757 11154 807 11188
rect 841 11154 877 11188
rect 757 11116 877 11154
rect 757 11082 807 11116
rect 841 11082 877 11116
rect 757 11044 877 11082
rect 757 11010 807 11044
rect 841 11010 877 11044
rect 757 10972 877 11010
rect 757 10938 807 10972
rect 841 10938 877 10972
rect 757 10900 877 10938
rect 757 10866 807 10900
rect 841 10866 877 10900
rect 757 10828 877 10866
rect 757 10794 807 10828
rect 841 10794 877 10828
rect 757 10756 877 10794
rect 757 10722 807 10756
rect 841 10722 877 10756
rect 757 10684 877 10722
rect 757 10650 807 10684
rect 841 10650 877 10684
rect 757 10612 877 10650
rect 757 10578 807 10612
rect 841 10578 877 10612
rect 757 10540 877 10578
rect 757 10506 807 10540
rect 841 10506 877 10540
rect 757 10468 877 10506
rect 757 10434 807 10468
rect 841 10434 877 10468
rect 757 10396 877 10434
rect 757 10362 807 10396
rect 841 10362 877 10396
rect 757 10324 877 10362
rect 757 10290 807 10324
rect 841 10290 877 10324
rect 757 10252 877 10290
rect 757 10218 807 10252
rect 841 10218 877 10252
rect 1148 34650 13844 34694
rect 1148 34616 1325 34650
rect 1359 34616 1397 34650
rect 1431 34616 1469 34650
rect 1503 34616 1541 34650
rect 1575 34616 1613 34650
rect 1647 34616 1685 34650
rect 1719 34616 1757 34650
rect 1791 34616 1829 34650
rect 1863 34616 1901 34650
rect 1935 34616 1973 34650
rect 2007 34616 2045 34650
rect 2079 34616 2117 34650
rect 2151 34616 2189 34650
rect 2223 34616 2261 34650
rect 2295 34616 2333 34650
rect 2367 34616 2405 34650
rect 2439 34616 2477 34650
rect 2511 34616 2549 34650
rect 2583 34616 2621 34650
rect 2655 34616 2693 34650
rect 2727 34616 2765 34650
rect 2799 34616 2837 34650
rect 2871 34616 2909 34650
rect 2943 34616 2981 34650
rect 3015 34616 3053 34650
rect 3087 34616 3125 34650
rect 3159 34616 3197 34650
rect 3231 34616 3269 34650
rect 3303 34616 3341 34650
rect 3375 34616 3413 34650
rect 3447 34616 3485 34650
rect 3519 34616 3557 34650
rect 3591 34616 3629 34650
rect 3663 34616 3701 34650
rect 3735 34616 3773 34650
rect 3807 34616 3845 34650
rect 3879 34616 3917 34650
rect 3951 34616 3989 34650
rect 4023 34616 4061 34650
rect 4095 34616 4133 34650
rect 4167 34616 4205 34650
rect 4239 34616 4277 34650
rect 4311 34616 4349 34650
rect 4383 34616 4421 34650
rect 4455 34616 4493 34650
rect 4527 34616 4565 34650
rect 4599 34616 4637 34650
rect 4671 34616 4709 34650
rect 4743 34616 4781 34650
rect 4815 34616 4853 34650
rect 4887 34616 4925 34650
rect 4959 34616 4997 34650
rect 5031 34616 5069 34650
rect 5103 34616 5141 34650
rect 5175 34616 5213 34650
rect 5247 34616 5285 34650
rect 5319 34616 5357 34650
rect 5391 34616 5429 34650
rect 5463 34616 5501 34650
rect 5535 34616 5573 34650
rect 5607 34616 5645 34650
rect 5679 34616 5717 34650
rect 5751 34616 5789 34650
rect 5823 34616 5861 34650
rect 5895 34616 5933 34650
rect 5967 34616 6005 34650
rect 6039 34616 6077 34650
rect 6111 34616 6149 34650
rect 6183 34616 6221 34650
rect 6255 34616 6293 34650
rect 6327 34616 6365 34650
rect 6399 34616 6437 34650
rect 6471 34616 6509 34650
rect 6543 34616 6581 34650
rect 6615 34616 6653 34650
rect 6687 34616 6725 34650
rect 6759 34616 6797 34650
rect 6831 34616 6869 34650
rect 6903 34616 6941 34650
rect 6975 34616 7013 34650
rect 7047 34616 7085 34650
rect 7119 34616 7157 34650
rect 7191 34616 7229 34650
rect 7263 34616 7301 34650
rect 7335 34616 7373 34650
rect 7407 34616 7445 34650
rect 7479 34616 7517 34650
rect 7551 34616 7589 34650
rect 7623 34616 7661 34650
rect 7695 34616 7733 34650
rect 7767 34616 7805 34650
rect 7839 34616 7877 34650
rect 7911 34616 7949 34650
rect 7983 34616 8021 34650
rect 8055 34616 8093 34650
rect 8127 34616 8165 34650
rect 8199 34616 8237 34650
rect 8271 34616 8309 34650
rect 8343 34616 8381 34650
rect 8415 34616 8453 34650
rect 8487 34616 8525 34650
rect 8559 34616 8597 34650
rect 8631 34616 8669 34650
rect 8703 34616 8741 34650
rect 8775 34616 8813 34650
rect 8847 34616 8885 34650
rect 8919 34616 8957 34650
rect 8991 34616 9029 34650
rect 9063 34616 9101 34650
rect 9135 34616 9173 34650
rect 9207 34616 9245 34650
rect 9279 34616 9317 34650
rect 9351 34616 9389 34650
rect 9423 34616 9461 34650
rect 9495 34616 9533 34650
rect 9567 34616 9605 34650
rect 9639 34616 9677 34650
rect 9711 34616 9749 34650
rect 9783 34616 9821 34650
rect 9855 34616 9893 34650
rect 9927 34616 9965 34650
rect 9999 34616 10037 34650
rect 10071 34616 10109 34650
rect 10143 34616 10181 34650
rect 10215 34616 10253 34650
rect 10287 34616 10325 34650
rect 10359 34616 10397 34650
rect 10431 34616 10469 34650
rect 10503 34616 10541 34650
rect 10575 34616 10613 34650
rect 10647 34616 10685 34650
rect 10719 34616 10757 34650
rect 10791 34616 10829 34650
rect 10863 34616 10901 34650
rect 10935 34616 10973 34650
rect 11007 34616 11045 34650
rect 11079 34616 11117 34650
rect 11151 34616 11189 34650
rect 11223 34616 11261 34650
rect 11295 34616 11333 34650
rect 11367 34616 11405 34650
rect 11439 34616 11477 34650
rect 11511 34616 11549 34650
rect 11583 34616 11621 34650
rect 11655 34616 11693 34650
rect 11727 34616 11765 34650
rect 11799 34616 11837 34650
rect 11871 34616 11909 34650
rect 11943 34616 11981 34650
rect 12015 34616 12053 34650
rect 12087 34616 12125 34650
rect 12159 34616 12197 34650
rect 12231 34616 12269 34650
rect 12303 34616 12341 34650
rect 12375 34616 12413 34650
rect 12447 34616 12485 34650
rect 12519 34616 12557 34650
rect 12591 34616 12629 34650
rect 12663 34616 12701 34650
rect 12735 34616 12773 34650
rect 12807 34616 12845 34650
rect 12879 34616 12917 34650
rect 12951 34616 12989 34650
rect 13023 34616 13061 34650
rect 13095 34616 13133 34650
rect 13167 34616 13205 34650
rect 13239 34616 13277 34650
rect 13311 34616 13349 34650
rect 13383 34616 13421 34650
rect 13455 34616 13493 34650
rect 13527 34616 13565 34650
rect 13599 34616 13637 34650
rect 13671 34616 13844 34650
rect 1148 34574 13844 34616
rect 1148 34509 1268 34574
rect 1148 34475 1192 34509
rect 1226 34475 1268 34509
rect 1148 34437 1268 34475
rect 1148 34403 1192 34437
rect 1226 34403 1268 34437
rect 1148 34365 1268 34403
rect 1148 34331 1192 34365
rect 1226 34331 1268 34365
rect 1148 34293 1268 34331
rect 1148 34259 1192 34293
rect 1226 34259 1268 34293
rect 1148 34221 1268 34259
rect 1148 34187 1192 34221
rect 1226 34187 1268 34221
rect 1148 34149 1268 34187
rect 1148 34115 1192 34149
rect 1226 34115 1268 34149
rect 1148 34077 1268 34115
rect 1148 34043 1192 34077
rect 1226 34043 1268 34077
rect 1148 34005 1268 34043
rect 1148 33971 1192 34005
rect 1226 33971 1268 34005
rect 1148 33933 1268 33971
rect 1148 33899 1192 33933
rect 1226 33899 1268 33933
rect 1148 33861 1268 33899
rect 1148 33827 1192 33861
rect 1226 33827 1268 33861
rect 1148 33789 1268 33827
rect 1148 33755 1192 33789
rect 1226 33755 1268 33789
rect 1148 33717 1268 33755
rect 1148 33683 1192 33717
rect 1226 33683 1268 33717
rect 1148 33645 1268 33683
rect 1148 33611 1192 33645
rect 1226 33611 1268 33645
rect 1148 33573 1268 33611
rect 1148 33539 1192 33573
rect 1226 33539 1268 33573
rect 1148 33501 1268 33539
rect 1148 33467 1192 33501
rect 1226 33467 1268 33501
rect 1148 33429 1268 33467
rect 1148 33395 1192 33429
rect 1226 33395 1268 33429
rect 1148 33357 1268 33395
rect 1148 33323 1192 33357
rect 1226 33323 1268 33357
rect 1148 33285 1268 33323
rect 1148 33251 1192 33285
rect 1226 33251 1268 33285
rect 1148 33213 1268 33251
rect 1148 33179 1192 33213
rect 1226 33179 1268 33213
rect 1148 33141 1268 33179
rect 1148 33107 1192 33141
rect 1226 33107 1268 33141
rect 1148 33069 1268 33107
rect 1148 33035 1192 33069
rect 1226 33035 1268 33069
rect 1148 32997 1268 33035
rect 1148 32963 1192 32997
rect 1226 32963 1268 32997
rect 1148 32925 1268 32963
rect 1148 32891 1192 32925
rect 1226 32891 1268 32925
rect 1148 32853 1268 32891
rect 1148 32819 1192 32853
rect 1226 32819 1268 32853
rect 1148 32781 1268 32819
rect 1148 32747 1192 32781
rect 1226 32751 1268 32781
rect 13724 34508 13844 34574
rect 13724 34474 13768 34508
rect 13802 34474 13844 34508
rect 13724 34436 13844 34474
rect 13724 34402 13768 34436
rect 13802 34402 13844 34436
rect 13724 34364 13844 34402
rect 13724 34330 13768 34364
rect 13802 34330 13844 34364
rect 13724 34292 13844 34330
rect 13724 34258 13768 34292
rect 13802 34258 13844 34292
rect 13724 34220 13844 34258
rect 13724 34186 13768 34220
rect 13802 34186 13844 34220
rect 13724 34148 13844 34186
rect 13724 34114 13768 34148
rect 13802 34114 13844 34148
rect 13724 34076 13844 34114
rect 13724 34042 13768 34076
rect 13802 34042 13844 34076
rect 13724 34004 13844 34042
rect 13724 33970 13768 34004
rect 13802 33970 13844 34004
rect 13724 33932 13844 33970
rect 13724 33898 13768 33932
rect 13802 33898 13844 33932
rect 13724 33860 13844 33898
rect 13724 33826 13768 33860
rect 13802 33826 13844 33860
rect 13724 33788 13844 33826
rect 13724 33754 13768 33788
rect 13802 33754 13844 33788
rect 13724 33716 13844 33754
rect 13724 33682 13768 33716
rect 13802 33682 13844 33716
rect 13724 33644 13844 33682
rect 13724 33610 13768 33644
rect 13802 33610 13844 33644
rect 13724 33572 13844 33610
rect 13724 33538 13768 33572
rect 13802 33538 13844 33572
rect 13724 33500 13844 33538
rect 13724 33466 13768 33500
rect 13802 33466 13844 33500
rect 13724 33428 13844 33466
rect 13724 33394 13768 33428
rect 13802 33394 13844 33428
rect 13724 33356 13844 33394
rect 13724 33322 13768 33356
rect 13802 33322 13844 33356
rect 13724 33284 13844 33322
rect 13724 33250 13768 33284
rect 13802 33250 13844 33284
rect 13724 33212 13844 33250
rect 13724 33178 13768 33212
rect 13802 33178 13844 33212
rect 13724 33140 13844 33178
rect 13724 33106 13768 33140
rect 13802 33106 13844 33140
rect 13724 33068 13844 33106
rect 13724 33034 13768 33068
rect 13802 33034 13844 33068
rect 13724 32996 13844 33034
rect 13724 32962 13768 32996
rect 13802 32962 13844 32996
rect 13724 32924 13844 32962
rect 13724 32890 13768 32924
rect 13802 32890 13844 32924
rect 13724 32852 13844 32890
rect 13724 32818 13768 32852
rect 13802 32818 13844 32852
rect 13724 32780 13844 32818
rect 1226 32747 10091 32751
rect 1148 32746 10091 32747
tri 10091 32746 10096 32751 sw
rect 13724 32746 13768 32780
rect 13802 32746 13844 32780
rect 1148 32734 10096 32746
tri 10096 32734 10108 32746 sw
rect 1148 32709 10108 32734
tri 10108 32709 10133 32734 sw
rect 1148 32675 1192 32709
rect 1226 32708 10133 32709
tri 10133 32708 10134 32709 sw
rect 13724 32708 13844 32746
rect 1226 32697 10134 32708
rect 1226 32675 4944 32697
rect 1148 32637 4944 32675
rect 1148 32603 1192 32637
rect 1226 32603 4944 32637
rect 1148 32565 4944 32603
rect 1148 32531 1192 32565
rect 1226 32531 4944 32565
rect 1148 32493 4944 32531
rect 1148 32459 1192 32493
rect 1226 32459 4944 32493
rect 1148 32421 4944 32459
rect 1148 32387 1192 32421
rect 1226 32387 4944 32421
rect 1148 32349 4944 32387
rect 1148 32315 1192 32349
rect 1226 32315 4944 32349
rect 1148 32277 4944 32315
rect 1148 32243 1192 32277
rect 1226 32243 4944 32277
rect 1148 32205 4944 32243
rect 1148 32171 1192 32205
rect 1226 32171 4944 32205
rect 1148 32133 4944 32171
rect 1148 32099 1192 32133
rect 1226 32099 4944 32133
rect 1148 32061 4944 32099
rect 1148 32027 1192 32061
rect 1226 32027 4944 32061
rect 1148 31989 4944 32027
rect 1148 31955 1192 31989
rect 1226 31955 4944 31989
rect 1148 31917 4944 31955
rect 1148 31883 1192 31917
rect 1226 31883 4944 31917
rect 1148 31877 4944 31883
rect 7236 31877 7745 32697
rect 10037 32674 10134 32697
tri 10134 32674 10168 32708 sw
rect 13724 32674 13768 32708
rect 13802 32674 13844 32708
rect 10037 32662 10168 32674
tri 10168 32662 10180 32674 sw
rect 10037 32637 10180 32662
tri 10180 32637 10205 32662 sw
rect 10037 32636 10205 32637
tri 10205 32636 10206 32637 sw
rect 13724 32636 13844 32674
rect 10037 32602 10206 32636
tri 10206 32602 10240 32636 sw
rect 13724 32602 13768 32636
rect 13802 32602 13844 32636
rect 10037 32590 10240 32602
tri 10240 32590 10252 32602 sw
rect 10037 32565 10252 32590
tri 10252 32565 10277 32590 sw
rect 10037 32564 10277 32565
tri 10277 32564 10278 32565 sw
rect 13724 32564 13844 32602
rect 10037 32551 10278 32564
tri 10278 32551 10291 32564 sw
rect 10037 32023 10291 32551
rect 10037 32014 10282 32023
tri 10282 32014 10291 32023 nw
rect 13724 32530 13768 32564
rect 13802 32530 13844 32564
rect 13724 32492 13844 32530
rect 13724 32458 13768 32492
rect 13802 32458 13844 32492
rect 13724 32420 13844 32458
rect 13724 32386 13768 32420
rect 13802 32386 13844 32420
rect 13724 32348 13844 32386
rect 13724 32314 13768 32348
rect 13802 32314 13844 32348
rect 13724 32276 13844 32314
rect 13724 32242 13768 32276
rect 13802 32242 13844 32276
rect 13724 32204 13844 32242
rect 13724 32170 13768 32204
rect 13802 32170 13844 32204
rect 13724 32132 13844 32170
rect 13724 32098 13768 32132
rect 13802 32098 13844 32132
rect 13724 32060 13844 32098
rect 13724 32026 13768 32060
rect 13802 32026 13844 32060
rect 10037 31989 10257 32014
tri 10257 31989 10282 32014 nw
rect 10037 31988 10256 31989
tri 10256 31988 10257 31989 nw
rect 13724 31988 13844 32026
rect 10037 31954 10222 31988
tri 10222 31954 10256 31988 nw
rect 13724 31954 13768 31988
rect 13802 31954 13844 31988
rect 10037 31942 10210 31954
tri 10210 31942 10222 31954 nw
rect 10037 31917 10185 31942
tri 10185 31917 10210 31942 nw
rect 10037 31916 10184 31917
tri 10184 31916 10185 31917 nw
rect 13724 31916 13844 31954
rect 10037 31882 10150 31916
tri 10150 31882 10184 31916 nw
rect 13724 31882 13768 31916
rect 13802 31882 13844 31916
rect 10037 31877 10138 31882
rect 1148 31870 10138 31877
tri 10138 31870 10150 31882 nw
rect 1148 31845 10113 31870
tri 10113 31845 10138 31870 nw
rect 1148 31811 1192 31845
rect 1226 31844 10112 31845
tri 10112 31844 10113 31845 nw
rect 13724 31844 13844 31882
rect 1226 31823 10091 31844
tri 10091 31823 10112 31844 nw
rect 1226 31811 1442 31823
rect 1148 31773 1442 31811
rect 1148 31739 1192 31773
rect 1226 31739 1442 31773
rect 1148 31701 1442 31739
rect 1148 31667 1192 31701
rect 1226 31667 1442 31701
rect 1148 31629 1442 31667
rect 1148 31595 1192 31629
rect 1226 31595 1442 31629
rect 1148 31557 1442 31595
rect 1148 31523 1192 31557
rect 1226 31523 1442 31557
rect 1148 31485 1442 31523
rect 1148 31451 1192 31485
rect 1226 31451 1442 31485
rect 1148 31413 1442 31451
rect 1148 31379 1192 31413
rect 1226 31379 1442 31413
rect 13724 31810 13768 31844
rect 13802 31810 13844 31844
rect 13724 31772 13844 31810
rect 13724 31738 13768 31772
rect 13802 31738 13844 31772
rect 13724 31700 13844 31738
rect 13724 31666 13768 31700
rect 13802 31666 13844 31700
rect 13724 31628 13844 31666
rect 13724 31594 13768 31628
rect 13802 31594 13844 31628
rect 13724 31556 13844 31594
rect 13724 31522 13768 31556
rect 13802 31522 13844 31556
rect 13724 31484 13844 31522
rect 13724 31450 13768 31484
rect 13802 31450 13844 31484
rect 13724 31412 13844 31450
rect 1148 31341 1442 31379
tri 1858 31378 1859 31379 se
rect 1859 31378 13157 31379
tri 13157 31378 13158 31379 sw
rect 13724 31378 13768 31412
rect 13802 31378 13844 31412
tri 1846 31366 1858 31378 se
rect 1858 31366 13158 31378
tri 13158 31366 13170 31378 sw
tri 1832 31352 1846 31366 se
rect 1846 31352 13170 31366
tri 13170 31352 13184 31366 sw
tri 1831 31351 1832 31352 se
rect 1832 31351 13184 31352
tri 1825 31345 1831 31351 se
rect 1831 31345 13184 31351
rect 1148 31307 1192 31341
rect 1226 31307 1442 31341
rect 1148 31269 1442 31307
rect 1148 31235 1192 31269
rect 1226 31235 1442 31269
rect 1148 31197 1442 31235
rect 1148 31163 1192 31197
rect 1226 31163 1442 31197
rect 1148 31125 1442 31163
rect 1148 31091 1192 31125
rect 1226 31091 1442 31125
rect 1148 31053 1442 31091
rect 1148 31019 1192 31053
rect 1226 31019 1442 31053
rect 1148 30981 1442 31019
rect 1148 30947 1192 30981
rect 1226 30947 1442 30981
rect 1148 30909 1442 30947
rect 1148 30875 1192 30909
rect 1226 30875 1442 30909
rect 1148 30837 1442 30875
rect 1148 30803 1192 30837
rect 1226 30803 1442 30837
rect 1148 30765 1442 30803
rect 1148 30731 1192 30765
rect 1226 30731 1442 30765
rect 1148 30693 1442 30731
rect 1148 30659 1192 30693
rect 1226 30659 1442 30693
rect 1148 30621 1442 30659
rect 1148 30587 1192 30621
rect 1226 30587 1442 30621
rect 1148 30549 1442 30587
rect 1148 30515 1192 30549
rect 1226 30515 1442 30549
rect 1148 30477 1442 30515
rect 1148 30443 1192 30477
rect 1226 30443 1442 30477
rect 1148 30405 1442 30443
rect 1148 30371 1192 30405
rect 1226 30371 1442 30405
rect 1148 30333 1442 30371
rect 1148 30299 1192 30333
rect 1226 30299 1442 30333
rect 1148 30261 1442 30299
rect 1148 30227 1192 30261
rect 1226 30227 1442 30261
rect 1148 30189 1442 30227
rect 1148 30155 1192 30189
rect 1226 30155 1442 30189
rect 1148 30117 1442 30155
rect 1148 30083 1192 30117
rect 1226 30083 1442 30117
rect 1148 30045 1442 30083
rect 1148 30011 1192 30045
rect 1226 30011 1442 30045
rect 1148 29973 1442 30011
rect 1148 29939 1192 29973
rect 1226 29939 1442 29973
rect 1148 29901 1442 29939
rect 1148 29867 1192 29901
rect 1226 29867 1442 29901
rect 1148 29829 1442 29867
rect 1148 29795 1192 29829
rect 1226 29795 1442 29829
rect 1148 29757 1442 29795
rect 1148 29723 1192 29757
rect 1226 29723 1442 29757
rect 1148 29685 1442 29723
rect 1148 29651 1192 29685
rect 1226 29651 1442 29685
rect 1148 29613 1442 29651
rect 1148 29579 1192 29613
rect 1226 29579 1442 29613
rect 1148 29541 1442 29579
rect 1148 29507 1192 29541
rect 1226 29507 1442 29541
rect 1148 29469 1442 29507
rect 1148 29435 1192 29469
rect 1226 29435 1442 29469
rect 1148 29397 1442 29435
rect 1148 29363 1192 29397
rect 1226 29363 1442 29397
rect 1148 29325 1442 29363
rect 1148 29291 1192 29325
rect 1226 29291 1442 29325
rect 1148 29253 1442 29291
rect 1148 29219 1192 29253
rect 1226 29219 1442 29253
rect 1148 29181 1442 29219
rect 1148 29147 1192 29181
rect 1226 29147 1442 29181
rect 1148 29109 1442 29147
rect 1148 29075 1192 29109
rect 1226 29075 1442 29109
rect 1148 29037 1442 29075
rect 1148 29003 1192 29037
rect 1226 29003 1442 29037
rect 1148 28965 1442 29003
rect 1148 28931 1192 28965
rect 1226 28931 1442 28965
rect 1148 28893 1442 28931
rect 1148 28859 1192 28893
rect 1226 28859 1442 28893
rect 1148 28821 1442 28859
rect 1148 28787 1192 28821
rect 1226 28787 1442 28821
rect 1148 28749 1442 28787
rect 1148 28715 1192 28749
rect 1226 28715 1442 28749
rect 1148 28677 1442 28715
rect 1148 28643 1192 28677
rect 1226 28643 1442 28677
rect 1148 28605 1442 28643
rect 1148 28571 1192 28605
rect 1226 28571 1442 28605
rect 1148 28533 1442 28571
rect 1148 28499 1192 28533
rect 1226 28499 1442 28533
rect 1148 28461 1442 28499
rect 1148 28427 1192 28461
rect 1226 28427 1442 28461
rect 1148 28389 1442 28427
rect 1148 28355 1192 28389
rect 1226 28355 1442 28389
rect 1148 28317 1442 28355
rect 1148 28283 1192 28317
rect 1226 28283 1442 28317
rect 1148 28245 1442 28283
rect 1148 28211 1192 28245
rect 1226 28211 1442 28245
rect 1148 28173 1442 28211
rect 1148 28139 1192 28173
rect 1226 28139 1442 28173
rect 1148 28101 1442 28139
rect 1148 28067 1192 28101
rect 1226 28067 1442 28101
rect 1148 28029 1442 28067
rect 1148 27995 1192 28029
rect 1226 27995 1442 28029
rect 1148 27957 1442 27995
rect 1148 27923 1192 27957
rect 1226 27923 1442 27957
rect 1148 27885 1442 27923
rect 1148 27851 1192 27885
rect 1226 27851 1442 27885
rect 1148 27813 1442 27851
rect 1148 27779 1192 27813
rect 1226 27779 1442 27813
rect 1148 27741 1442 27779
rect 1148 27707 1192 27741
rect 1226 27707 1442 27741
rect 1148 27669 1442 27707
rect 1148 27635 1192 27669
rect 1226 27635 1442 27669
rect 1148 27597 1442 27635
rect 1148 27563 1192 27597
rect 1226 27563 1442 27597
rect 1148 27525 1442 27563
rect 1148 27491 1192 27525
rect 1226 27491 1442 27525
rect 1148 27453 1442 27491
rect 1148 27419 1192 27453
rect 1226 27419 1442 27453
rect 1148 27381 1442 27419
rect 1148 27347 1192 27381
rect 1226 27347 1442 27381
rect 1148 27309 1442 27347
rect 1148 27275 1192 27309
rect 1226 27275 1442 27309
rect 1148 27237 1442 27275
rect 1148 27203 1192 27237
rect 1226 27203 1442 27237
rect 1148 27165 1442 27203
rect 1148 27131 1192 27165
rect 1226 27131 1442 27165
rect 1148 27093 1442 27131
rect 1148 27059 1192 27093
rect 1226 27059 1442 27093
tri 1659 31179 1825 31345 se
rect 1825 31179 1982 31345
rect 1659 31023 1982 31179
rect 13032 31341 13184 31345
tri 13184 31341 13195 31352 sw
rect 13032 31307 13195 31341
tri 13195 31307 13229 31341 sw
rect 13724 31332 13844 31378
rect 14099 34691 14142 34725
rect 14176 34691 14219 34725
rect 14099 34653 14219 34691
rect 14099 34619 14142 34653
rect 14176 34619 14219 34653
rect 14099 34581 14219 34619
rect 14099 34547 14142 34581
rect 14176 34547 14219 34581
rect 14099 34509 14219 34547
rect 14099 34475 14142 34509
rect 14176 34475 14219 34509
rect 14099 34437 14219 34475
rect 14099 34403 14142 34437
rect 14176 34403 14219 34437
rect 14099 34365 14219 34403
rect 14099 34331 14142 34365
rect 14176 34331 14219 34365
rect 14099 34293 14219 34331
rect 14099 34259 14142 34293
rect 14176 34259 14219 34293
rect 14099 34221 14219 34259
rect 14099 34187 14142 34221
rect 14176 34187 14219 34221
rect 14099 34149 14219 34187
rect 14099 34115 14142 34149
rect 14176 34115 14219 34149
rect 14099 34077 14219 34115
rect 14099 34043 14142 34077
rect 14176 34043 14219 34077
rect 14099 34005 14219 34043
rect 14099 33971 14142 34005
rect 14176 33971 14219 34005
rect 14099 33933 14219 33971
rect 14099 33899 14142 33933
rect 14176 33899 14219 33933
rect 14099 33861 14219 33899
rect 14099 33827 14142 33861
rect 14176 33827 14219 33861
rect 14099 33789 14219 33827
rect 14099 33755 14142 33789
rect 14176 33755 14219 33789
rect 14099 33717 14219 33755
rect 14099 33683 14142 33717
rect 14176 33683 14219 33717
rect 14099 33645 14219 33683
rect 14099 33611 14142 33645
rect 14176 33611 14219 33645
rect 14099 33573 14219 33611
rect 14099 33539 14142 33573
rect 14176 33539 14219 33573
rect 14099 33501 14219 33539
rect 14099 33467 14142 33501
rect 14176 33467 14219 33501
rect 14099 33429 14219 33467
rect 14099 33395 14142 33429
rect 14176 33395 14219 33429
rect 14099 33357 14219 33395
rect 14099 33323 14142 33357
rect 14176 33323 14219 33357
rect 14099 33285 14219 33323
rect 14099 33251 14142 33285
rect 14176 33251 14219 33285
rect 14099 33213 14219 33251
rect 14099 33179 14142 33213
rect 14176 33179 14219 33213
rect 14099 33141 14219 33179
rect 14099 33107 14142 33141
rect 14176 33107 14219 33141
rect 14099 33069 14219 33107
rect 14099 33035 14142 33069
rect 14176 33035 14219 33069
rect 14099 32997 14219 33035
rect 14099 32963 14142 32997
rect 14176 32963 14219 32997
rect 14099 32925 14219 32963
rect 14099 32891 14142 32925
rect 14176 32891 14219 32925
rect 14099 32853 14219 32891
rect 14099 32819 14142 32853
rect 14176 32819 14219 32853
rect 14099 32781 14219 32819
rect 14099 32747 14142 32781
rect 14176 32747 14219 32781
rect 14099 32709 14219 32747
rect 14099 32675 14142 32709
rect 14176 32675 14219 32709
rect 14099 32637 14219 32675
rect 14099 32603 14142 32637
rect 14176 32603 14219 32637
rect 14099 32565 14219 32603
rect 14099 32531 14142 32565
rect 14176 32531 14219 32565
rect 14099 32493 14219 32531
rect 14099 32459 14142 32493
rect 14176 32459 14219 32493
rect 14099 32421 14219 32459
rect 14099 32387 14142 32421
rect 14176 32387 14219 32421
rect 14099 32349 14219 32387
rect 14099 32315 14142 32349
rect 14176 32315 14219 32349
rect 14099 32277 14219 32315
rect 14099 32243 14142 32277
rect 14176 32243 14219 32277
rect 14099 32205 14219 32243
rect 14099 32171 14142 32205
rect 14176 32171 14219 32205
rect 14099 32133 14219 32171
rect 14099 32099 14142 32133
rect 14176 32099 14219 32133
rect 14099 32061 14219 32099
rect 14099 32027 14142 32061
rect 14176 32027 14219 32061
rect 14099 31989 14219 32027
rect 14099 31955 14142 31989
rect 14176 31955 14219 31989
rect 14099 31917 14219 31955
rect 14099 31883 14142 31917
rect 14176 31883 14219 31917
rect 14099 31845 14219 31883
rect 14099 31811 14142 31845
rect 14176 31811 14219 31845
rect 14099 31773 14219 31811
rect 14099 31739 14142 31773
rect 14176 31739 14219 31773
rect 14099 31701 14219 31739
rect 14099 31667 14142 31701
rect 14176 31667 14219 31701
rect 14099 31629 14219 31667
rect 14099 31595 14142 31629
rect 14176 31595 14219 31629
rect 14099 31557 14219 31595
rect 14099 31523 14142 31557
rect 14176 31523 14219 31557
rect 14099 31485 14219 31523
rect 14099 31451 14142 31485
rect 14176 31451 14219 31485
rect 14099 31413 14219 31451
rect 14099 31379 14142 31413
rect 14176 31379 14219 31413
rect 14099 31341 14219 31379
rect 14099 31307 14142 31341
rect 14176 31307 14219 31341
rect 13032 31294 13229 31307
tri 13229 31294 13242 31307 sw
rect 13032 31269 13242 31294
tri 13242 31269 13267 31294 sw
rect 14099 31269 14219 31307
rect 13032 31235 13267 31269
tri 13267 31235 13301 31269 sw
rect 14099 31235 14142 31269
rect 14176 31235 14219 31269
rect 13032 31222 13301 31235
tri 13301 31222 13314 31235 sw
rect 13032 31197 13314 31222
tri 13314 31197 13339 31222 sw
rect 14099 31197 14219 31235
rect 13032 31163 13339 31197
tri 13339 31163 13373 31197 sw
rect 14099 31163 14142 31197
rect 14176 31163 14219 31197
rect 13032 31150 13373 31163
tri 13373 31150 13386 31163 sw
rect 13032 31125 13386 31150
tri 13386 31125 13411 31150 sw
rect 14099 31125 14219 31163
rect 13032 31091 13411 31125
tri 13411 31091 13445 31125 sw
rect 14099 31091 14142 31125
rect 14176 31091 14219 31125
rect 13032 31078 13445 31091
tri 13445 31078 13458 31091 sw
rect 13032 31053 13458 31078
tri 13458 31053 13483 31078 sw
rect 14099 31053 14219 31091
rect 13032 31023 13483 31053
rect 1659 31019 13483 31023
tri 13483 31019 13517 31053 sw
rect 14099 31019 14142 31053
rect 14176 31019 14219 31053
rect 1659 31006 13517 31019
tri 13517 31006 13530 31019 sw
rect 1659 30985 13530 31006
rect 1659 30981 2129 30985
tri 2129 30981 2133 30985 nw
tri 12883 30981 12887 30985 ne
rect 12887 30981 13530 30985
tri 13530 30981 13555 31006 sw
rect 14099 30981 14219 31019
rect 1659 30955 2103 30981
tri 2103 30955 2129 30981 nw
tri 12887 30955 12913 30981 ne
rect 12913 30955 13555 30981
tri 13555 30955 13581 30981 sw
rect 1659 30948 2095 30955
rect 1659 27458 1726 30948
rect 1976 30947 2095 30948
tri 2095 30947 2103 30955 nw
tri 12913 30947 12921 30955 ne
rect 12921 30947 13581 30955
tri 13581 30947 13589 30955 sw
rect 14099 30947 14142 30981
rect 14176 30947 14219 30981
rect 1976 27458 2093 30947
tri 2093 30945 2095 30947 nw
tri 12921 30945 12923 30947 ne
rect 12923 30941 13589 30947
tri 2320 30744 2420 30844 se
rect 2420 30799 12596 30844
rect 2420 30744 4939 30799
rect 2320 30683 4939 30744
rect 7231 30683 7750 30799
rect 10042 30744 12596 30799
tri 12596 30744 12696 30844 sw
rect 10042 30683 12696 30744
rect 2320 30632 12696 30683
rect 2509 30486 4482 30512
rect 4481 30370 4482 30486
rect 2509 30344 4482 30370
rect 10500 30486 12473 30512
rect 12472 30370 12473 30486
rect 10500 30344 12473 30370
rect 2422 30183 12572 30228
rect 2422 30067 4939 30183
rect 7231 30067 7750 30183
rect 10042 30067 12572 30183
rect 2422 30016 12572 30067
rect 2509 29870 4482 29896
rect 4481 29754 4482 29870
rect 2509 29728 4482 29754
rect 10500 29870 12473 29896
rect 12472 29754 12473 29870
rect 10500 29728 12473 29754
rect 2422 29567 12572 29612
rect 2422 29451 4939 29567
rect 7231 29451 7750 29567
rect 10042 29451 12572 29567
rect 2422 29400 12572 29451
rect 2509 29254 4482 29280
rect 4481 29138 4482 29254
rect 2509 29112 4482 29138
rect 10500 29254 12473 29280
rect 12472 29138 12473 29254
rect 10500 29112 12473 29138
rect 2422 28951 12572 28996
rect 2422 28835 4939 28951
rect 7231 28835 7750 28951
rect 10042 28835 12572 28951
rect 2422 28784 12572 28835
rect 2509 28638 4482 28664
rect 4481 28522 4482 28638
rect 2509 28496 4482 28522
rect 10500 28638 12473 28664
rect 12472 28522 12473 28638
rect 10500 28496 12473 28522
rect 2422 28335 12572 28380
rect 2422 28219 4939 28335
rect 7231 28219 7750 28335
rect 10042 28219 12572 28335
rect 2422 28168 12572 28219
rect 2509 28022 4482 28048
rect 4481 27906 4482 28022
rect 2509 27880 4482 27906
rect 10500 28022 12473 28048
rect 12472 27906 12473 28022
rect 10500 27880 12473 27906
rect 2320 27719 12696 27764
rect 2320 27652 4939 27719
tri 2320 27552 2420 27652 ne
rect 2420 27603 4939 27652
rect 7231 27603 7750 27719
rect 10042 27652 12696 27719
rect 10042 27603 12596 27652
rect 2420 27552 12596 27603
tri 12596 27552 12696 27652 nw
rect 1659 27437 2093 27458
rect 12923 27451 13031 30941
rect 13281 30934 13589 30941
tri 13589 30934 13602 30947 sw
rect 13281 30909 13602 30934
tri 13602 30909 13627 30934 sw
rect 14099 30909 14219 30947
rect 13281 30875 13627 30909
tri 13627 30875 13661 30909 sw
rect 14099 30875 14142 30909
rect 14176 30875 14219 30909
rect 13281 30862 13661 30875
tri 13661 30862 13674 30875 sw
rect 13281 30837 13674 30862
tri 13674 30837 13699 30862 sw
rect 14099 30837 14219 30875
rect 13281 30803 13699 30837
tri 13699 30803 13733 30837 sw
rect 14099 30803 14142 30837
rect 14176 30803 14219 30837
rect 13281 30790 13733 30803
tri 13733 30790 13746 30803 sw
rect 13281 30765 13746 30790
tri 13746 30765 13771 30790 sw
rect 14099 30765 14219 30803
rect 13281 30753 13771 30765
tri 13771 30753 13783 30765 sw
rect 13281 27451 13783 30753
tri 2093 27437 2107 27451 sw
tri 12909 27437 12923 27451 se
rect 12923 27437 13783 27451
rect 1659 27419 2107 27437
tri 2107 27419 2125 27437 sw
tri 12891 27419 12909 27437 se
rect 12909 27419 13783 27437
rect 1659 27411 2125 27419
tri 2125 27411 2133 27419 sw
tri 12883 27411 12891 27419 se
rect 12891 27411 13783 27419
rect 1659 27334 13783 27411
rect 1659 27217 1985 27334
tri 1659 27084 1792 27217 ne
rect 1792 27084 1985 27217
rect 13035 27217 13783 27334
rect 13035 27203 13343 27217
tri 13343 27203 13357 27217 nw
rect 13035 27190 13330 27203
tri 13330 27190 13343 27203 nw
rect 13035 27165 13305 27190
tri 13305 27165 13330 27190 nw
rect 13035 27131 13271 27165
tri 13271 27131 13305 27165 nw
rect 13035 27118 13258 27131
tri 13258 27118 13271 27131 nw
rect 13035 27093 13233 27118
tri 13233 27093 13258 27118 nw
rect 13035 27084 13199 27093
tri 1792 27059 1817 27084 ne
rect 1817 27059 13199 27084
tri 13199 27059 13233 27093 nw
rect 1148 27021 1442 27059
tri 1817 27053 1823 27059 ne
rect 1823 27053 13186 27059
tri 1823 27046 1830 27053 ne
rect 1830 27046 13186 27053
tri 13186 27046 13199 27059 nw
tri 1830 27021 1855 27046 ne
rect 1855 27021 13161 27046
tri 13161 27021 13186 27046 nw
rect 1148 26987 1192 27021
rect 1226 26987 1442 27021
tri 1855 27017 1859 27021 ne
rect 1859 27017 13157 27021
tri 13157 27017 13161 27021 nw
rect 1148 26949 1442 26987
rect 1148 26915 1192 26949
rect 1226 26915 1442 26949
rect 1148 26877 1442 26915
rect 1148 26843 1192 26877
rect 1226 26843 1442 26877
rect 1148 26805 1442 26843
rect 1148 26771 1192 26805
rect 1226 26771 1442 26805
rect 1148 26733 1442 26771
rect 1148 26699 1192 26733
rect 1226 26699 1442 26733
rect 1148 26661 1442 26699
rect 1148 26627 1192 26661
rect 1226 26627 1442 26661
rect 1148 26589 1442 26627
rect 1148 26555 1192 26589
rect 1226 26555 1442 26589
rect 1148 26517 1442 26555
rect 1148 26483 1192 26517
rect 1226 26483 1442 26517
rect 1148 26445 1442 26483
rect 1148 26411 1192 26445
rect 1226 26411 1442 26445
rect 1148 26373 1442 26411
rect 1148 26339 1192 26373
rect 1226 26339 1442 26373
rect 1148 26320 1442 26339
rect 1148 26301 1734 26320
rect 1148 26267 1192 26301
rect 1226 26267 1734 26301
rect 1148 26229 1734 26267
rect 1148 26195 1192 26229
rect 1226 26195 1734 26229
rect 1148 26157 1734 26195
tri 2383 26157 2406 26180 se
rect 2406 26157 12582 26180
tri 12582 26157 12605 26180 sw
rect 1148 26123 1192 26157
rect 1226 26123 1734 26157
tri 2349 26123 2383 26157 se
rect 2383 26153 12605 26157
rect 2383 26123 4933 26153
rect 1148 26085 1734 26123
tri 2336 26110 2349 26123 se
rect 2349 26110 4933 26123
rect 1148 26051 1192 26085
rect 1226 26051 1734 26085
rect 1148 26013 1734 26051
rect 1148 25979 1192 26013
rect 1226 25979 1734 26013
tri 2326 26100 2336 26110 se
rect 2336 26100 4933 26110
rect 2326 26037 4933 26100
rect 7225 26037 7757 26153
rect 10049 26123 12605 26153
tri 12605 26123 12639 26157 sw
rect 10049 26110 12639 26123
tri 12639 26110 12652 26123 sw
rect 10049 26100 12652 26110
tri 12652 26100 12662 26110 sw
rect 10049 26037 12662 26100
rect 2326 26008 12662 26037
rect 1148 25941 1734 25979
rect 1148 25907 1192 25941
rect 1226 25907 1734 25941
rect 1148 25869 1734 25907
rect 1148 25835 1192 25869
rect 1226 25835 1734 25869
rect 1148 25797 1734 25835
rect 1148 25763 1192 25797
rect 1226 25763 1734 25797
rect 1148 25725 1734 25763
rect 2528 25887 4472 25909
rect 2528 25771 2546 25887
rect 4454 25771 4472 25887
rect 2528 25749 4472 25771
rect 10510 25887 12454 25909
rect 10510 25771 10528 25887
rect 12436 25771 12454 25887
rect 10510 25749 12454 25771
rect 1148 25691 1192 25725
rect 1226 25691 1734 25725
rect 1148 25653 1734 25691
rect 1148 25619 1192 25653
rect 1226 25619 1734 25653
rect 1148 25581 1734 25619
rect 1148 25547 1192 25581
rect 1226 25547 1734 25581
rect 1148 25509 1734 25547
rect 1148 25475 1192 25509
rect 1226 25475 1734 25509
rect 2456 25621 12536 25648
rect 2456 25505 4933 25621
rect 7225 25505 7757 25621
rect 10049 25505 12536 25621
rect 2456 25476 12536 25505
rect 1148 25437 1734 25475
rect 1148 25403 1192 25437
rect 1226 25403 1734 25437
rect 1148 25365 1734 25403
rect 1148 25331 1192 25365
rect 1226 25331 1734 25365
rect 1148 25293 1734 25331
rect 1148 25259 1192 25293
rect 1226 25259 1734 25293
rect 1148 25221 1734 25259
rect 1148 25187 1192 25221
rect 1226 25187 1734 25221
rect 2528 25355 4472 25377
rect 2528 25239 2546 25355
rect 4454 25239 4472 25355
rect 2528 25217 4472 25239
rect 10510 25355 12454 25377
rect 10510 25239 10528 25355
rect 12436 25239 12454 25355
rect 10510 25217 12454 25239
rect 1148 25149 1734 25187
rect 1148 25115 1192 25149
rect 1226 25115 1734 25149
rect 1148 25077 1734 25115
rect 1148 25043 1192 25077
rect 1226 25043 1734 25077
rect 1148 25005 1734 25043
rect 1148 24971 1192 25005
rect 1226 24971 1734 25005
rect 1148 24933 1734 24971
rect 2456 25112 4826 25116
rect 7344 25112 12536 25116
rect 2456 25089 12536 25112
rect 2456 24973 4933 25089
rect 7225 24973 7757 25089
rect 10049 24973 12536 25089
rect 2456 24944 12536 24973
rect 1148 24899 1192 24933
rect 1226 24899 1734 24933
rect 1148 24861 1734 24899
rect 1148 24827 1192 24861
rect 1226 24827 1734 24861
rect 1148 24789 1734 24827
rect 1148 24755 1192 24789
rect 1226 24755 1734 24789
rect 1148 24717 1734 24755
rect 1148 24683 1192 24717
rect 1226 24683 1734 24717
rect 2528 24823 4472 24845
rect 2528 24707 2546 24823
rect 4454 24707 4472 24823
rect 2528 24685 4472 24707
rect 10510 24823 12454 24845
rect 10510 24707 10528 24823
rect 12436 24707 12454 24823
rect 10510 24685 12454 24707
rect 1148 24645 1734 24683
rect 1148 24611 1192 24645
rect 1226 24611 1734 24645
rect 1148 24573 1734 24611
rect 1148 24539 1192 24573
rect 1226 24539 1734 24573
rect 1148 24501 1734 24539
rect 1148 24467 1192 24501
rect 1226 24467 1734 24501
rect 1148 24429 1734 24467
rect 1148 24395 1192 24429
rect 1226 24395 1734 24429
rect 2456 24557 12536 24584
rect 2456 24441 4933 24557
rect 7225 24441 7757 24557
rect 10049 24441 12536 24557
rect 2456 24412 12536 24441
rect 1148 24357 1734 24395
rect 1148 24323 1192 24357
rect 1226 24323 1734 24357
rect 1148 24285 1734 24323
rect 1148 24251 1192 24285
rect 1226 24251 1734 24285
rect 1148 24213 1734 24251
rect 1148 24179 1192 24213
rect 1226 24179 1734 24213
rect 1148 24141 1734 24179
rect 2528 24291 4472 24313
rect 2528 24175 2546 24291
rect 4454 24175 4472 24291
rect 2528 24153 4472 24175
rect 10510 24291 12454 24313
rect 10510 24175 10528 24291
rect 12436 24175 12454 24291
rect 10510 24153 12454 24175
rect 1148 24107 1192 24141
rect 1226 24107 1734 24141
rect 1148 24069 1734 24107
rect 1148 24035 1192 24069
rect 1226 24035 1734 24069
rect 1148 23997 1734 24035
rect 1148 23963 1192 23997
rect 1226 23963 1734 23997
rect 1148 23925 1734 23963
rect 1148 23891 1192 23925
rect 1226 23891 1734 23925
rect 1148 23853 1734 23891
rect 2456 24025 12536 24052
rect 2456 23909 4933 24025
rect 7225 23909 7757 24025
rect 10049 23909 12536 24025
rect 2456 23880 12536 23909
rect 1148 23819 1192 23853
rect 1226 23819 1734 23853
rect 1148 23781 1734 23819
rect 1148 23747 1192 23781
rect 1226 23747 1734 23781
rect 1148 23709 1734 23747
rect 1148 23675 1192 23709
rect 1226 23675 1734 23709
rect 1148 23637 1734 23675
rect 1148 23603 1192 23637
rect 1226 23603 1734 23637
rect 2528 23759 4472 23781
rect 2528 23643 2546 23759
rect 4454 23643 4472 23759
rect 2528 23621 4472 23643
rect 10510 23759 12454 23781
rect 10510 23643 10528 23759
rect 12436 23643 12454 23759
rect 10510 23621 12454 23643
rect 1148 23565 1734 23603
rect 1148 23531 1192 23565
rect 1226 23531 1734 23565
rect 1148 23493 1734 23531
rect 1148 23459 1192 23493
rect 1226 23459 1734 23493
rect 1148 23421 1734 23459
rect 2326 23493 12662 23520
rect 2326 23428 4933 23493
tri 2326 23421 2333 23428 ne
rect 2333 23421 4933 23428
rect 1148 23387 1192 23421
rect 1226 23387 1734 23421
tri 2333 23387 2367 23421 ne
rect 2367 23387 4933 23421
rect 1148 23349 1734 23387
tri 2367 23374 2380 23387 ne
rect 2380 23377 4933 23387
rect 7225 23377 7757 23493
rect 10049 23428 12662 23493
rect 10049 23421 12655 23428
tri 12655 23421 12662 23428 nw
rect 10049 23387 12621 23421
tri 12621 23387 12655 23421 nw
rect 10049 23377 12608 23387
rect 2380 23374 12608 23377
tri 12608 23374 12621 23387 nw
tri 2380 23349 2405 23374 ne
rect 2405 23349 12583 23374
tri 12583 23349 12608 23374 nw
rect 1148 23315 1192 23349
rect 1226 23315 1734 23349
tri 2405 23348 2406 23349 ne
rect 2406 23348 12582 23349
tri 12582 23348 12583 23349 nw
rect 1148 23277 1734 23315
rect 1148 23243 1192 23277
rect 1226 23243 1734 23277
rect 1148 23208 1734 23243
rect 1148 23205 1268 23208
rect 1148 23171 1192 23205
rect 1226 23171 1268 23205
rect 1148 23133 1268 23171
rect 1148 23099 1192 23133
rect 1226 23099 1268 23133
rect 1148 23061 1268 23099
rect 1148 23027 1192 23061
rect 1226 23027 1268 23061
rect 1148 22989 1268 23027
rect 1148 22955 1192 22989
rect 1226 22955 1268 22989
rect 1148 22917 1268 22955
rect 1148 22883 1192 22917
rect 1226 22883 1268 22917
rect 1148 22845 1268 22883
rect 1148 22811 1192 22845
rect 1226 22811 1268 22845
rect 1148 22773 1268 22811
rect 1148 22739 1192 22773
rect 1226 22739 1268 22773
rect 1148 22701 1268 22739
rect 1148 22667 1192 22701
rect 1226 22667 1268 22701
rect 1148 22629 1268 22667
rect 1148 22595 1192 22629
rect 1226 22595 1268 22629
rect 1148 22557 1268 22595
rect 1148 22523 1192 22557
rect 1226 22523 1268 22557
rect 13527 22543 13783 27217
tri 4871 22523 4891 22543 se
rect 4891 22523 13783 22543
rect 1148 22485 1268 22523
tri 4858 22510 4871 22523 se
rect 4871 22510 13783 22523
tri 4833 22485 4858 22510 se
rect 4858 22489 13783 22510
rect 4858 22485 4945 22489
rect 1148 22451 1192 22485
rect 1226 22451 1268 22485
tri 4799 22451 4833 22485 se
rect 4833 22451 4945 22485
rect 1148 22413 1268 22451
tri 4786 22438 4799 22451 se
rect 4799 22438 4945 22451
tri 4761 22413 4786 22438 se
rect 4786 22413 4945 22438
rect 1148 22379 1192 22413
rect 1226 22379 1268 22413
tri 4727 22379 4761 22413 se
rect 4761 22379 4945 22413
rect 1148 22341 1268 22379
tri 4714 22366 4727 22379 se
rect 4727 22366 4945 22379
rect 1148 22307 1192 22341
rect 1226 22307 1268 22341
rect 1148 22269 1268 22307
rect 1148 22235 1192 22269
rect 1226 22235 1268 22269
rect 1148 22197 1268 22235
rect 1148 22163 1192 22197
rect 1226 22163 1268 22197
rect 1148 22125 1268 22163
rect 1148 22091 1192 22125
rect 1226 22091 1268 22125
rect 1148 22053 1268 22091
rect 1148 22019 1192 22053
rect 1226 22019 1268 22053
rect 1148 21981 1268 22019
rect 1148 21947 1192 21981
rect 1226 21947 1268 21981
rect 1148 21909 1268 21947
rect 1148 21875 1192 21909
rect 1226 21875 1268 21909
rect 1148 21837 1268 21875
rect 1148 21803 1192 21837
rect 1226 21803 1268 21837
tri 4691 22343 4714 22366 se
rect 4714 22343 4945 22366
rect 4691 21815 4945 22343
tri 4691 21803 4703 21815 ne
rect 4703 21803 4945 21815
rect 1148 21765 1268 21803
tri 4703 21790 4716 21803 ne
rect 4716 21790 4945 21803
tri 4716 21765 4741 21790 ne
rect 4741 21765 4945 21790
rect 1148 21731 1192 21765
rect 1226 21731 1268 21765
tri 4741 21731 4775 21765 ne
rect 4775 21731 4945 21765
rect 1148 21693 1268 21731
tri 4775 21718 4788 21731 ne
rect 4788 21718 4945 21731
tri 4788 21693 4813 21718 ne
rect 4813 21693 4945 21718
rect 1148 21659 1192 21693
rect 1226 21659 1268 21693
tri 4813 21659 4847 21693 ne
rect 4847 21669 4945 21693
rect 7237 21669 7744 22489
rect 10036 22041 13783 22489
rect 10036 22019 13761 22041
tri 13761 22019 13783 22041 nw
rect 14099 30731 14142 30765
rect 14176 30731 14219 30765
rect 14099 30693 14219 30731
rect 14099 30659 14142 30693
rect 14176 30659 14219 30693
rect 14099 30621 14219 30659
rect 14099 30587 14142 30621
rect 14176 30587 14219 30621
rect 14099 30549 14219 30587
rect 14099 30515 14142 30549
rect 14176 30515 14219 30549
rect 14099 30477 14219 30515
rect 14099 30443 14142 30477
rect 14176 30443 14219 30477
rect 14099 30405 14219 30443
rect 14099 30371 14142 30405
rect 14176 30371 14219 30405
rect 14099 30333 14219 30371
rect 14099 30299 14142 30333
rect 14176 30299 14219 30333
rect 14099 30261 14219 30299
rect 14099 30227 14142 30261
rect 14176 30227 14219 30261
rect 14099 30189 14219 30227
rect 14099 30155 14142 30189
rect 14176 30155 14219 30189
rect 14099 30117 14219 30155
rect 14099 30083 14142 30117
rect 14176 30083 14219 30117
rect 14099 30045 14219 30083
rect 14099 30011 14142 30045
rect 14176 30011 14219 30045
rect 14099 29973 14219 30011
rect 14099 29939 14142 29973
rect 14176 29939 14219 29973
rect 14099 29901 14219 29939
rect 14099 29867 14142 29901
rect 14176 29867 14219 29901
rect 14099 29829 14219 29867
rect 14099 29795 14142 29829
rect 14176 29795 14219 29829
rect 14099 29757 14219 29795
rect 14099 29723 14142 29757
rect 14176 29723 14219 29757
rect 14099 29685 14219 29723
rect 14099 29651 14142 29685
rect 14176 29651 14219 29685
rect 14099 29613 14219 29651
rect 14099 29579 14142 29613
rect 14176 29579 14219 29613
rect 14099 29541 14219 29579
rect 14099 29507 14142 29541
rect 14176 29507 14219 29541
rect 14099 29469 14219 29507
rect 14099 29435 14142 29469
rect 14176 29435 14219 29469
rect 14099 29397 14219 29435
rect 14099 29363 14142 29397
rect 14176 29363 14219 29397
rect 14099 29325 14219 29363
rect 14099 29291 14142 29325
rect 14176 29291 14219 29325
rect 14099 29253 14219 29291
rect 14099 29219 14142 29253
rect 14176 29219 14219 29253
rect 14099 29181 14219 29219
rect 14099 29147 14142 29181
rect 14176 29147 14219 29181
rect 14099 29109 14219 29147
rect 14099 29075 14142 29109
rect 14176 29075 14219 29109
rect 14099 29037 14219 29075
rect 14099 29003 14142 29037
rect 14176 29003 14219 29037
rect 14099 28965 14219 29003
rect 14099 28931 14142 28965
rect 14176 28931 14219 28965
rect 14099 28893 14219 28931
rect 14099 28859 14142 28893
rect 14176 28859 14219 28893
rect 14099 28821 14219 28859
rect 14099 28787 14142 28821
rect 14176 28787 14219 28821
rect 14099 28749 14219 28787
rect 14099 28715 14142 28749
rect 14176 28715 14219 28749
rect 14099 28677 14219 28715
rect 14099 28643 14142 28677
rect 14176 28643 14219 28677
rect 14099 28605 14219 28643
rect 14099 28571 14142 28605
rect 14176 28571 14219 28605
rect 14099 28533 14219 28571
rect 14099 28499 14142 28533
rect 14176 28499 14219 28533
rect 14099 28461 14219 28499
rect 14099 28427 14142 28461
rect 14176 28427 14219 28461
rect 14099 28389 14219 28427
rect 14099 28355 14142 28389
rect 14176 28355 14219 28389
rect 14099 28317 14219 28355
rect 14099 28283 14142 28317
rect 14176 28283 14219 28317
rect 14099 28245 14219 28283
rect 14099 28211 14142 28245
rect 14176 28211 14219 28245
rect 14099 28173 14219 28211
rect 14099 28139 14142 28173
rect 14176 28139 14219 28173
rect 14099 28101 14219 28139
rect 14099 28067 14142 28101
rect 14176 28067 14219 28101
rect 14099 28029 14219 28067
rect 14099 27995 14142 28029
rect 14176 27995 14219 28029
rect 14099 27957 14219 27995
rect 14099 27923 14142 27957
rect 14176 27923 14219 27957
rect 14099 27885 14219 27923
rect 14099 27851 14142 27885
rect 14176 27851 14219 27885
rect 14099 27813 14219 27851
rect 14099 27779 14142 27813
rect 14176 27779 14219 27813
rect 14099 27741 14219 27779
rect 14099 27707 14142 27741
rect 14176 27707 14219 27741
rect 14099 27669 14219 27707
rect 14099 27635 14142 27669
rect 14176 27635 14219 27669
rect 14099 27597 14219 27635
rect 14099 27563 14142 27597
rect 14176 27563 14219 27597
rect 14099 27525 14219 27563
rect 14099 27491 14142 27525
rect 14176 27491 14219 27525
rect 14099 27453 14219 27491
rect 14099 27419 14142 27453
rect 14176 27419 14219 27453
rect 14099 27381 14219 27419
rect 14099 27347 14142 27381
rect 14176 27347 14219 27381
rect 14099 27309 14219 27347
rect 14099 27275 14142 27309
rect 14176 27275 14219 27309
rect 14099 27237 14219 27275
rect 14099 27203 14142 27237
rect 14176 27203 14219 27237
rect 14099 27165 14219 27203
rect 14099 27131 14142 27165
rect 14176 27131 14219 27165
rect 14099 27093 14219 27131
rect 14099 27059 14142 27093
rect 14176 27059 14219 27093
rect 14099 27021 14219 27059
rect 14099 26987 14142 27021
rect 14176 26987 14219 27021
rect 14099 26949 14219 26987
rect 14099 26915 14142 26949
rect 14176 26915 14219 26949
rect 14099 26877 14219 26915
rect 14099 26843 14142 26877
rect 14176 26843 14219 26877
rect 14099 26805 14219 26843
rect 14099 26771 14142 26805
rect 14176 26771 14219 26805
rect 14099 26733 14219 26771
rect 14099 26699 14142 26733
rect 14176 26699 14219 26733
rect 14099 26661 14219 26699
rect 14099 26627 14142 26661
rect 14176 26627 14219 26661
rect 14099 26589 14219 26627
rect 14099 26555 14142 26589
rect 14176 26555 14219 26589
rect 14099 26517 14219 26555
rect 14099 26483 14142 26517
rect 14176 26483 14219 26517
rect 14099 26445 14219 26483
rect 14099 26411 14142 26445
rect 14176 26411 14219 26445
rect 14099 26373 14219 26411
rect 14099 26339 14142 26373
rect 14176 26339 14219 26373
rect 14099 26301 14219 26339
rect 14099 26267 14142 26301
rect 14176 26267 14219 26301
rect 14099 26229 14219 26267
rect 14099 26195 14142 26229
rect 14176 26195 14219 26229
rect 14099 26157 14219 26195
rect 14099 26123 14142 26157
rect 14176 26123 14219 26157
rect 14099 26085 14219 26123
rect 14099 26051 14142 26085
rect 14176 26051 14219 26085
rect 14099 26013 14219 26051
rect 14099 25979 14142 26013
rect 14176 25979 14219 26013
rect 14099 25941 14219 25979
rect 14099 25907 14142 25941
rect 14176 25907 14219 25941
rect 14099 25869 14219 25907
rect 14099 25835 14142 25869
rect 14176 25835 14219 25869
rect 14099 25797 14219 25835
rect 14099 25763 14142 25797
rect 14176 25763 14219 25797
rect 14099 25725 14219 25763
rect 14099 25691 14142 25725
rect 14176 25691 14219 25725
rect 14099 25653 14219 25691
rect 14099 25619 14142 25653
rect 14176 25619 14219 25653
rect 14099 25581 14219 25619
rect 14099 25547 14142 25581
rect 14176 25547 14219 25581
rect 14099 25509 14219 25547
rect 14099 25475 14142 25509
rect 14176 25475 14219 25509
rect 14099 25437 14219 25475
rect 14099 25403 14142 25437
rect 14176 25403 14219 25437
rect 14099 25365 14219 25403
rect 14099 25331 14142 25365
rect 14176 25331 14219 25365
rect 14099 25293 14219 25331
rect 14099 25259 14142 25293
rect 14176 25259 14219 25293
rect 14099 25221 14219 25259
rect 14099 25187 14142 25221
rect 14176 25187 14219 25221
rect 14099 25149 14219 25187
rect 14099 25115 14142 25149
rect 14176 25115 14219 25149
rect 14099 25077 14219 25115
rect 14099 25043 14142 25077
rect 14176 25043 14219 25077
rect 14099 25005 14219 25043
rect 14099 24971 14142 25005
rect 14176 24971 14219 25005
rect 14099 24933 14219 24971
rect 14099 24899 14142 24933
rect 14176 24899 14219 24933
rect 14099 24861 14219 24899
rect 14099 24827 14142 24861
rect 14176 24827 14219 24861
rect 14099 24789 14219 24827
rect 14099 24755 14142 24789
rect 14176 24755 14219 24789
rect 14099 24717 14219 24755
rect 14099 24683 14142 24717
rect 14176 24683 14219 24717
rect 14099 24645 14219 24683
rect 14099 24611 14142 24645
rect 14176 24611 14219 24645
rect 14099 24573 14219 24611
rect 14099 24539 14142 24573
rect 14176 24539 14219 24573
rect 14099 24501 14219 24539
rect 14099 24467 14142 24501
rect 14176 24467 14219 24501
rect 14099 24429 14219 24467
rect 14099 24395 14142 24429
rect 14176 24395 14219 24429
rect 14099 24357 14219 24395
rect 14099 24323 14142 24357
rect 14176 24323 14219 24357
rect 14099 24285 14219 24323
rect 14099 24251 14142 24285
rect 14176 24251 14219 24285
rect 14099 24213 14219 24251
rect 14099 24179 14142 24213
rect 14176 24179 14219 24213
rect 14099 24141 14219 24179
rect 14099 24107 14142 24141
rect 14176 24107 14219 24141
rect 14099 24069 14219 24107
rect 14099 24035 14142 24069
rect 14176 24035 14219 24069
rect 14099 23997 14219 24035
rect 14099 23963 14142 23997
rect 14176 23963 14219 23997
rect 14099 23925 14219 23963
rect 14099 23891 14142 23925
rect 14176 23891 14219 23925
rect 14099 23853 14219 23891
rect 14099 23819 14142 23853
rect 14176 23819 14219 23853
rect 14099 23781 14219 23819
rect 14099 23747 14142 23781
rect 14176 23747 14219 23781
rect 14099 23709 14219 23747
rect 14099 23675 14142 23709
rect 14176 23675 14219 23709
rect 14099 23637 14219 23675
rect 14099 23603 14142 23637
rect 14176 23603 14219 23637
rect 14099 23565 14219 23603
rect 14099 23531 14142 23565
rect 14176 23531 14219 23565
rect 14099 23493 14219 23531
rect 14099 23459 14142 23493
rect 14176 23459 14219 23493
rect 14099 23421 14219 23459
rect 14099 23387 14142 23421
rect 14176 23387 14219 23421
rect 14099 23349 14219 23387
rect 14099 23315 14142 23349
rect 14176 23315 14219 23349
rect 14099 23277 14219 23315
rect 14099 23243 14142 23277
rect 14176 23243 14219 23277
rect 14099 23205 14219 23243
rect 14099 23171 14142 23205
rect 14176 23171 14219 23205
rect 14099 23133 14219 23171
rect 14099 23099 14142 23133
rect 14176 23099 14219 23133
rect 14099 23061 14219 23099
rect 14099 23027 14142 23061
rect 14176 23027 14219 23061
rect 14099 22989 14219 23027
rect 14099 22955 14142 22989
rect 14176 22955 14219 22989
rect 14099 22917 14219 22955
rect 14099 22883 14142 22917
rect 14176 22883 14219 22917
rect 14099 22845 14219 22883
rect 14099 22811 14142 22845
rect 14176 22811 14219 22845
rect 14099 22773 14219 22811
rect 14099 22739 14142 22773
rect 14176 22739 14219 22773
rect 14099 22701 14219 22739
rect 14099 22667 14142 22701
rect 14176 22667 14219 22701
rect 14099 22629 14219 22667
rect 14099 22595 14142 22629
rect 14176 22595 14219 22629
rect 14099 22557 14219 22595
rect 14099 22523 14142 22557
rect 14176 22523 14219 22557
rect 14099 22485 14219 22523
rect 14099 22451 14142 22485
rect 14176 22451 14219 22485
rect 14099 22413 14219 22451
rect 14099 22379 14142 22413
rect 14176 22379 14219 22413
rect 14099 22341 14219 22379
rect 14099 22307 14142 22341
rect 14176 22307 14219 22341
rect 14099 22269 14219 22307
rect 14099 22235 14142 22269
rect 14176 22235 14219 22269
rect 14099 22197 14219 22235
rect 14099 22163 14142 22197
rect 14176 22163 14219 22197
rect 14099 22125 14219 22163
rect 14099 22091 14142 22125
rect 14176 22091 14219 22125
rect 14099 22053 14219 22091
rect 14099 22019 14142 22053
rect 14176 22019 14219 22053
rect 10036 22006 13748 22019
tri 13748 22006 13761 22019 nw
rect 10036 21981 13723 22006
tri 13723 21981 13748 22006 nw
rect 14099 21981 14219 22019
rect 10036 21947 13689 21981
tri 13689 21947 13723 21981 nw
rect 14099 21947 14142 21981
rect 14176 21947 14219 21981
rect 10036 21934 13676 21947
tri 13676 21934 13689 21947 nw
rect 10036 21909 13651 21934
tri 13651 21909 13676 21934 nw
rect 14099 21909 14219 21947
rect 10036 21875 13617 21909
tri 13617 21875 13651 21909 nw
rect 14099 21875 14142 21909
rect 14176 21875 14219 21909
rect 10036 21862 13604 21875
tri 13604 21862 13617 21875 nw
rect 10036 21837 13579 21862
tri 13579 21837 13604 21862 nw
rect 14099 21837 14219 21875
rect 10036 21803 13545 21837
tri 13545 21803 13579 21837 nw
rect 14099 21803 14142 21837
rect 14176 21803 14219 21837
rect 10036 21790 13532 21803
tri 13532 21790 13545 21803 nw
rect 10036 21765 13507 21790
tri 13507 21765 13532 21790 nw
rect 14099 21765 14219 21803
rect 10036 21731 13473 21765
tri 13473 21731 13507 21765 nw
rect 14099 21731 14142 21765
rect 14176 21731 14219 21765
rect 10036 21718 13460 21731
tri 13460 21718 13473 21731 nw
rect 10036 21693 13435 21718
tri 13435 21693 13460 21718 nw
rect 14099 21693 14219 21731
rect 10036 21669 13401 21693
rect 4847 21659 13401 21669
tri 13401 21659 13435 21693 nw
rect 14099 21659 14142 21693
rect 14176 21659 14219 21693
rect 1148 21621 1268 21659
tri 4847 21646 4860 21659 ne
rect 4860 21646 13388 21659
tri 13388 21646 13401 21659 nw
tri 4860 21621 4885 21646 ne
rect 4885 21621 13363 21646
tri 13363 21621 13388 21646 nw
rect 14099 21621 14219 21659
rect 1148 21587 1192 21621
rect 1226 21587 1268 21621
tri 4885 21615 4891 21621 ne
rect 4891 21615 13357 21621
tri 13357 21615 13363 21621 nw
rect 1148 21549 1268 21587
rect 1148 21515 1192 21549
rect 1226 21515 1268 21549
rect 1148 21477 1268 21515
rect 1148 21443 1192 21477
rect 1226 21443 1268 21477
rect 1148 21405 1268 21443
rect 1148 21371 1192 21405
rect 1226 21371 1268 21405
rect 1148 21333 1268 21371
rect 1148 21299 1192 21333
rect 1226 21299 1268 21333
rect 1148 21261 1268 21299
rect 14099 21587 14142 21621
rect 14176 21587 14219 21621
rect 14099 21549 14219 21587
rect 14099 21515 14142 21549
rect 14176 21515 14219 21549
rect 14099 21477 14219 21515
rect 14099 21443 14142 21477
rect 14176 21443 14219 21477
rect 14099 21405 14219 21443
rect 14099 21371 14142 21405
rect 14176 21371 14219 21405
rect 14099 21333 14219 21371
rect 14099 21299 14142 21333
rect 14176 21299 14219 21333
rect 1148 21227 1192 21261
rect 1226 21227 1268 21261
rect 1148 21189 1268 21227
rect 1148 21155 1192 21189
rect 1226 21155 1268 21189
rect 1148 21117 1268 21155
rect 1148 21083 1192 21117
rect 1226 21083 1268 21117
rect 1148 21045 1268 21083
rect 1148 21011 1192 21045
rect 1226 21011 1268 21045
rect 1148 20973 1268 21011
rect 1148 20939 1192 20973
rect 1226 20939 1268 20973
rect 1148 20901 1268 20939
rect 1148 20867 1192 20901
rect 1226 20867 1268 20901
rect 1148 20829 1268 20867
rect 1148 20795 1192 20829
rect 1226 20795 1268 20829
rect 1148 20757 1268 20795
rect 1148 20723 1192 20757
rect 1226 20723 1268 20757
rect 1148 20685 1268 20723
rect 1148 20651 1192 20685
rect 1226 20651 1268 20685
rect 1148 20613 1268 20651
rect 1148 20579 1192 20613
rect 1226 20579 1268 20613
rect 1148 20541 1268 20579
rect 1148 20507 1192 20541
rect 1226 20507 1268 20541
rect 1148 20469 1268 20507
rect 1148 20435 1192 20469
rect 1226 20435 1268 20469
rect 1148 20397 1268 20435
rect 1148 20363 1192 20397
rect 1226 20363 1268 20397
rect 1148 20325 1268 20363
rect 1148 20291 1192 20325
rect 1226 20291 1268 20325
rect 1148 20253 1268 20291
rect 1148 20219 1192 20253
rect 1226 20219 1268 20253
rect 1148 20181 1268 20219
rect 1148 20147 1192 20181
rect 1226 20147 1268 20181
rect 1148 20109 1268 20147
rect 1148 20075 1192 20109
rect 1226 20075 1268 20109
rect 1148 20037 1268 20075
rect 1148 20003 1192 20037
rect 1226 20003 1268 20037
rect 1148 19965 1268 20003
rect 1148 19931 1192 19965
rect 1226 19931 1268 19965
rect 1148 19893 1268 19931
rect 1148 19859 1192 19893
rect 1226 19859 1268 19893
rect 1148 19821 1268 19859
rect 1148 19787 1192 19821
rect 1226 19787 1268 19821
rect 1148 19749 1268 19787
rect 1148 19715 1192 19749
rect 1226 19715 1268 19749
rect 1148 19677 1268 19715
rect 1148 19643 1192 19677
rect 1226 19643 1268 19677
rect 1148 19605 1268 19643
rect 1148 19571 1192 19605
rect 1226 19571 1268 19605
rect 1148 19533 1268 19571
rect 1148 19499 1192 19533
rect 1226 19499 1268 19533
rect 1148 19461 1268 19499
rect 1148 19427 1192 19461
rect 1226 19427 1268 19461
rect 1148 19389 1268 19427
rect 1148 19355 1192 19389
rect 1226 19355 1268 19389
rect 1148 19317 1268 19355
rect 1148 19283 1192 19317
rect 1226 19283 1268 19317
rect 1148 19245 1268 19283
rect 1148 19211 1192 19245
rect 1226 19211 1268 19245
rect 1148 19173 1268 19211
rect 1148 19139 1192 19173
rect 1226 19139 1268 19173
rect 1148 19101 1268 19139
rect 1148 19067 1192 19101
rect 1226 19067 1268 19101
rect 1148 19029 1268 19067
rect 1148 18995 1192 19029
rect 1226 18995 1268 19029
rect 1148 18957 1268 18995
rect 1148 18923 1192 18957
rect 1226 18923 1268 18957
rect 1148 18885 1268 18923
rect 1148 18851 1192 18885
rect 1226 18851 1268 18885
rect 1148 18813 1268 18851
rect 1148 18779 1192 18813
rect 1226 18779 1268 18813
rect 1148 18741 1268 18779
rect 1148 18707 1192 18741
rect 1226 18707 1268 18741
rect 1148 18669 1268 18707
rect 1148 18635 1192 18669
rect 1226 18635 1268 18669
rect 1148 18597 1268 18635
rect 1148 18563 1192 18597
rect 1226 18563 1268 18597
rect 1148 18525 1268 18563
rect 1148 18491 1192 18525
rect 1226 18491 1268 18525
rect 1148 18453 1268 18491
rect 1148 18419 1192 18453
rect 1226 18419 1268 18453
rect 1148 18381 1268 18419
rect 1148 18347 1192 18381
rect 1226 18347 1268 18381
rect 1148 18309 1268 18347
rect 1148 18275 1192 18309
rect 1226 18275 1268 18309
rect 1148 18237 1268 18275
rect 1148 18203 1192 18237
rect 1226 18203 1268 18237
rect 1148 18165 1268 18203
rect 1148 18131 1192 18165
rect 1226 18131 1268 18165
rect 1148 18093 1268 18131
rect 1148 18059 1192 18093
rect 1226 18059 1268 18093
rect 1148 18021 1268 18059
rect 1148 17987 1192 18021
rect 1226 17987 1268 18021
rect 1148 17949 1268 17987
rect 1148 17915 1192 17949
rect 1226 17915 1268 17949
rect 1148 17877 1268 17915
rect 1148 17843 1192 17877
rect 1226 17843 1268 17877
rect 1148 17805 1268 17843
rect 1148 17771 1192 17805
rect 1226 17771 1268 17805
rect 1148 17733 1268 17771
rect 1148 17699 1192 17733
rect 1226 17699 1268 17733
rect 1148 17661 1268 17699
rect 1148 17627 1192 17661
rect 1226 17627 1268 17661
rect 1148 17589 1268 17627
rect 1148 17555 1192 17589
rect 1226 17555 1268 17589
rect 1148 17517 1268 17555
rect 1148 17483 1192 17517
rect 1226 17483 1268 17517
rect 1148 17445 1268 17483
rect 1148 17411 1192 17445
rect 1226 17411 1268 17445
rect 1148 17373 1268 17411
rect 1148 17339 1192 17373
rect 1226 17339 1268 17373
rect 1148 17301 1268 17339
rect 1148 17267 1192 17301
rect 1226 17267 1268 17301
rect 1148 17229 1268 17267
rect 1148 17195 1192 17229
rect 1226 17195 1268 17229
rect 1148 17157 1268 17195
rect 1148 17123 1192 17157
rect 1226 17123 1268 17157
rect 1148 17085 1268 17123
rect 1148 17051 1192 17085
rect 1226 17051 1268 17085
rect 1148 17013 1268 17051
rect 1148 16979 1192 17013
rect 1226 16979 1268 17013
rect 1148 16941 1268 16979
rect 1148 16907 1192 16941
rect 1226 16907 1268 16941
rect 1148 16869 1268 16907
rect 1148 16835 1192 16869
rect 1226 16835 1268 16869
rect 1148 16797 1268 16835
rect 1148 16763 1192 16797
rect 1226 16763 1268 16797
rect 1148 16725 1268 16763
rect 1148 16691 1192 16725
rect 1226 16691 1268 16725
rect 1148 16653 1268 16691
rect 1148 16619 1192 16653
rect 1226 16619 1268 16653
rect 1148 16581 1268 16619
rect 1148 16547 1192 16581
rect 1226 16547 1268 16581
rect 1148 16509 1268 16547
rect 1148 16475 1192 16509
rect 1226 16475 1268 16509
rect 1148 16437 1268 16475
rect 1148 16403 1192 16437
rect 1226 16403 1268 16437
rect 1148 16365 1268 16403
rect 1148 16331 1192 16365
rect 1226 16331 1268 16365
rect 1148 16293 1268 16331
rect 1148 16259 1192 16293
rect 1226 16259 1268 16293
rect 1148 16221 1268 16259
rect 1148 16187 1192 16221
rect 1226 16187 1268 16221
rect 1148 16149 1268 16187
rect 1148 16115 1192 16149
rect 1226 16115 1268 16149
rect 1148 16077 1268 16115
rect 1148 16043 1192 16077
rect 1226 16043 1268 16077
rect 1148 16005 1268 16043
rect 1148 15971 1192 16005
rect 1226 15971 1268 16005
rect 1148 15933 1268 15971
rect 1148 15899 1192 15933
rect 1226 15899 1268 15933
rect 1148 15861 1268 15899
rect 1148 15827 1192 15861
rect 1226 15827 1268 15861
rect 1148 15789 1268 15827
rect 1148 15755 1192 15789
rect 1226 15755 1268 15789
rect 1148 15717 1268 15755
rect 1148 15683 1192 15717
rect 1226 15683 1268 15717
rect 1148 15645 1268 15683
rect 1148 15611 1192 15645
rect 1226 15611 1268 15645
rect 1148 15573 1268 15611
rect 1148 15539 1192 15573
rect 1226 15539 1268 15573
rect 1148 15501 1268 15539
rect 1148 15467 1192 15501
rect 1226 15467 1268 15501
rect 1148 15429 1268 15467
rect 1148 15395 1192 15429
rect 1226 15395 1268 15429
rect 1148 15357 1268 15395
rect 1148 15323 1192 15357
rect 1226 15323 1268 15357
rect 1148 15285 1268 15323
rect 1148 15251 1192 15285
rect 1226 15251 1268 15285
rect 1148 15213 1268 15251
rect 1148 15179 1192 15213
rect 1226 15179 1268 15213
rect 1148 15141 1268 15179
rect 1148 15107 1192 15141
rect 1226 15107 1268 15141
rect 1148 15069 1268 15107
rect 1148 15035 1192 15069
rect 1226 15035 1268 15069
rect 1148 14997 1268 15035
rect 1148 14963 1192 14997
rect 1226 14963 1268 14997
rect 1148 14925 1268 14963
rect 1148 14891 1192 14925
rect 1226 14891 1268 14925
rect 1148 14853 1268 14891
rect 1148 14819 1192 14853
rect 1226 14819 1268 14853
rect 1148 14781 1268 14819
rect 1148 14747 1192 14781
rect 1226 14747 1268 14781
rect 1148 14709 1268 14747
rect 1148 14675 1192 14709
rect 1226 14675 1268 14709
rect 1148 14637 1268 14675
rect 1148 14603 1192 14637
rect 1226 14603 1268 14637
rect 1148 14565 1268 14603
rect 1148 14531 1192 14565
rect 1226 14531 1268 14565
rect 1148 14493 1268 14531
rect 1148 14459 1192 14493
rect 1226 14459 1268 14493
rect 1148 14421 1268 14459
rect 1148 14387 1192 14421
rect 1226 14387 1268 14421
rect 1148 14349 1268 14387
rect 1148 14315 1192 14349
rect 1226 14315 1268 14349
rect 1148 14277 1268 14315
rect 1148 14243 1192 14277
rect 1226 14243 1268 14277
rect 1148 14205 1268 14243
rect 1148 14171 1192 14205
rect 1226 14171 1268 14205
rect 1148 14133 1268 14171
rect 1148 14099 1192 14133
rect 1226 14099 1268 14133
rect 1148 14061 1268 14099
rect 1148 14027 1192 14061
rect 1226 14027 1268 14061
rect 1148 13989 1268 14027
rect 1148 13955 1192 13989
rect 1226 13955 1268 13989
rect 1148 13917 1268 13955
rect 1148 13883 1192 13917
rect 1226 13883 1268 13917
rect 1148 13845 1268 13883
rect 1148 13811 1192 13845
rect 1226 13811 1268 13845
rect 1148 13773 1268 13811
rect 1148 13739 1192 13773
rect 1226 13739 1268 13773
rect 1148 13701 1268 13739
rect 1148 13667 1192 13701
rect 1226 13667 1268 13701
rect 1148 13629 1268 13667
rect 1148 13595 1192 13629
rect 1226 13595 1268 13629
rect 1148 13557 1268 13595
rect 1148 13523 1192 13557
rect 1226 13523 1268 13557
rect 1148 13485 1268 13523
rect 1148 13451 1192 13485
rect 1226 13451 1268 13485
rect 1148 13413 1268 13451
rect 1148 13379 1192 13413
rect 1226 13379 1268 13413
rect 1148 13341 1268 13379
rect 1148 13307 1192 13341
rect 1226 13307 1268 13341
rect 1148 13269 1268 13307
rect 1148 13235 1192 13269
rect 1226 13235 1268 13269
rect 1148 13197 1268 13235
rect 1148 13163 1192 13197
rect 1226 13163 1268 13197
rect 1148 13125 1268 13163
rect 1148 13091 1192 13125
rect 1226 13091 1268 13125
rect 1148 13053 1268 13091
rect 1148 13019 1192 13053
rect 1226 13019 1268 13053
rect 1148 12981 1268 13019
rect 1148 12947 1192 12981
rect 1226 12947 1268 12981
rect 1148 12909 1268 12947
rect 1148 12875 1192 12909
rect 1226 12875 1268 12909
rect 1148 12837 1268 12875
rect 1148 12803 1192 12837
rect 1226 12803 1268 12837
rect 1148 12765 1268 12803
rect 1148 12731 1192 12765
rect 1226 12731 1268 12765
rect 1148 12693 1268 12731
rect 1148 12659 1192 12693
rect 1226 12659 1268 12693
rect 1148 12621 1268 12659
rect 1148 12587 1192 12621
rect 1226 12587 1268 12621
rect 1148 12549 1268 12587
rect 1148 12515 1192 12549
rect 1226 12515 1268 12549
rect 1148 12477 1268 12515
rect 1148 12443 1192 12477
rect 1226 12443 1268 12477
rect 1148 12405 1268 12443
rect 1148 12371 1192 12405
rect 1226 12371 1268 12405
rect 1148 12333 1268 12371
rect 1148 12299 1192 12333
rect 1226 12299 1268 12333
rect 1148 12261 1268 12299
rect 1148 12227 1192 12261
rect 1226 12227 1268 12261
rect 1148 12189 1268 12227
rect 1148 12155 1192 12189
rect 1226 12155 1268 12189
rect 1148 12117 1268 12155
rect 1148 12083 1192 12117
rect 1226 12083 1268 12117
rect 1148 12045 1268 12083
rect 1148 12011 1192 12045
rect 1226 12011 1268 12045
rect 1148 11973 1268 12011
rect 1148 11939 1192 11973
rect 1226 11939 1268 11973
rect 1148 11901 1268 11939
rect 1148 11867 1192 11901
rect 1226 11867 1268 11901
rect 1148 11829 1268 11867
rect 1148 11795 1192 11829
rect 1226 11795 1268 11829
rect 1148 11757 1268 11795
rect 1148 11723 1192 11757
rect 1226 11723 1268 11757
rect 1148 11685 1268 11723
rect 1148 11651 1192 11685
rect 1226 11651 1268 11685
rect 1148 11613 1268 11651
rect 1148 11579 1192 11613
rect 1226 11579 1268 11613
rect 1148 11541 1268 11579
rect 1148 11507 1192 11541
rect 1226 11507 1268 11541
rect 1148 11469 1268 11507
rect 1148 11435 1192 11469
rect 1226 11435 1268 11469
rect 1148 11397 1268 11435
rect 1148 11363 1192 11397
rect 1226 11363 1268 11397
rect 1148 11325 1268 11363
rect 1148 11291 1192 11325
rect 1226 11291 1268 11325
rect 1148 11253 1268 11291
rect 1148 11219 1192 11253
rect 1226 11219 1268 11253
rect 1148 11181 1268 11219
rect 1148 11147 1192 11181
rect 1226 11147 1268 11181
rect 1148 11109 1268 11147
rect 1148 11075 1192 11109
rect 1226 11075 1268 11109
rect 1148 11037 1268 11075
rect 1148 11003 1192 11037
rect 1226 11003 1268 11037
rect 1148 10965 1268 11003
rect 1148 10931 1192 10965
rect 1226 10931 1268 10965
rect 1148 10893 1268 10931
rect 1148 10859 1192 10893
rect 1226 10859 1268 10893
rect 1148 10821 1268 10859
rect 1148 10787 1192 10821
rect 1226 10787 1268 10821
rect 1148 10749 1268 10787
rect 1148 10715 1192 10749
rect 1226 10715 1268 10749
rect 1148 10677 1268 10715
rect 1148 10643 1192 10677
rect 1226 10643 1268 10677
rect 1148 10605 1268 10643
rect 1148 10571 1192 10605
rect 1226 10571 1268 10605
rect 1148 10533 1268 10571
rect 1148 10499 1192 10533
rect 1226 10499 1268 10533
rect 1148 10461 1268 10499
rect 1148 10427 1192 10461
rect 1226 10427 1268 10461
rect 1148 10362 1268 10427
rect 13724 21219 13844 21262
rect 13724 21185 13768 21219
rect 13802 21185 13844 21219
rect 13724 21147 13844 21185
rect 13724 21113 13768 21147
rect 13802 21113 13844 21147
rect 13724 21075 13844 21113
rect 13724 21041 13768 21075
rect 13802 21041 13844 21075
rect 13724 21003 13844 21041
rect 13724 20969 13768 21003
rect 13802 20969 13844 21003
rect 13724 20931 13844 20969
rect 13724 20897 13768 20931
rect 13802 20897 13844 20931
rect 13724 20859 13844 20897
rect 13724 20825 13768 20859
rect 13802 20825 13844 20859
rect 13724 20787 13844 20825
rect 13724 20753 13768 20787
rect 13802 20753 13844 20787
rect 13724 20715 13844 20753
rect 13724 20681 13768 20715
rect 13802 20681 13844 20715
rect 13724 20643 13844 20681
rect 13724 20609 13768 20643
rect 13802 20609 13844 20643
rect 13724 20571 13844 20609
rect 13724 20537 13768 20571
rect 13802 20537 13844 20571
rect 13724 20499 13844 20537
rect 13724 20465 13768 20499
rect 13802 20465 13844 20499
rect 13724 20427 13844 20465
rect 13724 20393 13768 20427
rect 13802 20393 13844 20427
rect 13724 20355 13844 20393
rect 13724 20321 13768 20355
rect 13802 20321 13844 20355
rect 13724 20283 13844 20321
rect 13724 20249 13768 20283
rect 13802 20249 13844 20283
rect 13724 20211 13844 20249
rect 13724 20177 13768 20211
rect 13802 20177 13844 20211
rect 13724 20139 13844 20177
rect 13724 20105 13768 20139
rect 13802 20105 13844 20139
rect 13724 20067 13844 20105
rect 13724 20033 13768 20067
rect 13802 20033 13844 20067
rect 13724 19995 13844 20033
rect 13724 19961 13768 19995
rect 13802 19961 13844 19995
rect 13724 19923 13844 19961
rect 13724 19889 13768 19923
rect 13802 19889 13844 19923
rect 13724 19851 13844 19889
rect 13724 19817 13768 19851
rect 13802 19817 13844 19851
rect 13724 19779 13844 19817
rect 13724 19745 13768 19779
rect 13802 19745 13844 19779
rect 13724 19707 13844 19745
rect 13724 19673 13768 19707
rect 13802 19673 13844 19707
rect 13724 19635 13844 19673
rect 13724 19601 13768 19635
rect 13802 19601 13844 19635
rect 13724 19563 13844 19601
rect 13724 19529 13768 19563
rect 13802 19529 13844 19563
rect 13724 19491 13844 19529
rect 13724 19457 13768 19491
rect 13802 19457 13844 19491
rect 13724 19419 13844 19457
rect 13724 19385 13768 19419
rect 13802 19385 13844 19419
rect 13724 19347 13844 19385
rect 13724 19313 13768 19347
rect 13802 19313 13844 19347
rect 13724 19275 13844 19313
rect 13724 19241 13768 19275
rect 13802 19241 13844 19275
rect 13724 19203 13844 19241
rect 13724 19169 13768 19203
rect 13802 19169 13844 19203
rect 13724 19131 13844 19169
rect 13724 19097 13768 19131
rect 13802 19097 13844 19131
rect 13724 19059 13844 19097
rect 13724 19025 13768 19059
rect 13802 19025 13844 19059
rect 13724 18987 13844 19025
rect 13724 18953 13768 18987
rect 13802 18953 13844 18987
rect 13724 18915 13844 18953
rect 13724 18881 13768 18915
rect 13802 18881 13844 18915
rect 13724 18843 13844 18881
rect 13724 18809 13768 18843
rect 13802 18809 13844 18843
rect 13724 18771 13844 18809
rect 13724 18737 13768 18771
rect 13802 18737 13844 18771
rect 13724 18699 13844 18737
rect 13724 18665 13768 18699
rect 13802 18665 13844 18699
rect 13724 18627 13844 18665
rect 13724 18593 13768 18627
rect 13802 18593 13844 18627
rect 13724 18555 13844 18593
rect 13724 18521 13768 18555
rect 13802 18521 13844 18555
rect 13724 18483 13844 18521
rect 13724 18449 13768 18483
rect 13802 18449 13844 18483
rect 13724 18411 13844 18449
rect 13724 18377 13768 18411
rect 13802 18377 13844 18411
rect 13724 18339 13844 18377
rect 13724 18305 13768 18339
rect 13802 18305 13844 18339
rect 13724 18267 13844 18305
rect 13724 18233 13768 18267
rect 13802 18233 13844 18267
rect 13724 18195 13844 18233
rect 13724 18161 13768 18195
rect 13802 18161 13844 18195
rect 13724 18123 13844 18161
rect 13724 18089 13768 18123
rect 13802 18089 13844 18123
rect 13724 18051 13844 18089
rect 13724 18017 13768 18051
rect 13802 18017 13844 18051
rect 13724 17979 13844 18017
rect 13724 17945 13768 17979
rect 13802 17945 13844 17979
rect 13724 17907 13844 17945
rect 13724 17873 13768 17907
rect 13802 17873 13844 17907
rect 13724 17835 13844 17873
rect 13724 17801 13768 17835
rect 13802 17801 13844 17835
rect 13724 17763 13844 17801
rect 13724 17729 13768 17763
rect 13802 17729 13844 17763
rect 13724 17691 13844 17729
rect 13724 17657 13768 17691
rect 13802 17657 13844 17691
rect 13724 17619 13844 17657
rect 13724 17585 13768 17619
rect 13802 17585 13844 17619
rect 13724 17547 13844 17585
rect 13724 17513 13768 17547
rect 13802 17513 13844 17547
rect 13724 17475 13844 17513
rect 13724 17441 13768 17475
rect 13802 17441 13844 17475
rect 13724 17403 13844 17441
rect 13724 17369 13768 17403
rect 13802 17369 13844 17403
rect 13724 17331 13844 17369
rect 13724 17297 13768 17331
rect 13802 17297 13844 17331
rect 13724 17259 13844 17297
rect 13724 17225 13768 17259
rect 13802 17225 13844 17259
rect 13724 17187 13844 17225
rect 13724 17153 13768 17187
rect 13802 17153 13844 17187
rect 13724 17115 13844 17153
rect 13724 17081 13768 17115
rect 13802 17081 13844 17115
rect 13724 17043 13844 17081
rect 13724 17009 13768 17043
rect 13802 17009 13844 17043
rect 13724 16971 13844 17009
rect 13724 16937 13768 16971
rect 13802 16937 13844 16971
rect 13724 16899 13844 16937
rect 13724 16865 13768 16899
rect 13802 16865 13844 16899
rect 13724 16827 13844 16865
rect 13724 16793 13768 16827
rect 13802 16793 13844 16827
rect 13724 16755 13844 16793
rect 13724 16721 13768 16755
rect 13802 16721 13844 16755
rect 13724 16683 13844 16721
rect 13724 16649 13768 16683
rect 13802 16649 13844 16683
rect 13724 16611 13844 16649
rect 13724 16577 13768 16611
rect 13802 16577 13844 16611
rect 13724 16539 13844 16577
rect 13724 16505 13768 16539
rect 13802 16505 13844 16539
rect 13724 16467 13844 16505
rect 13724 16433 13768 16467
rect 13802 16433 13844 16467
rect 13724 16395 13844 16433
rect 13724 16361 13768 16395
rect 13802 16361 13844 16395
rect 13724 16323 13844 16361
rect 13724 16289 13768 16323
rect 13802 16289 13844 16323
rect 13724 16251 13844 16289
rect 13724 16217 13768 16251
rect 13802 16217 13844 16251
rect 13724 16179 13844 16217
rect 13724 16145 13768 16179
rect 13802 16145 13844 16179
rect 13724 16107 13844 16145
rect 13724 16073 13768 16107
rect 13802 16073 13844 16107
rect 13724 16035 13844 16073
rect 13724 16001 13768 16035
rect 13802 16001 13844 16035
rect 13724 15963 13844 16001
rect 13724 15929 13768 15963
rect 13802 15929 13844 15963
rect 13724 15891 13844 15929
rect 13724 15857 13768 15891
rect 13802 15857 13844 15891
rect 13724 15819 13844 15857
rect 13724 15785 13768 15819
rect 13802 15785 13844 15819
rect 13724 15747 13844 15785
rect 13724 15713 13768 15747
rect 13802 15713 13844 15747
rect 13724 15675 13844 15713
rect 13724 15641 13768 15675
rect 13802 15641 13844 15675
rect 13724 15603 13844 15641
rect 13724 15569 13768 15603
rect 13802 15569 13844 15603
rect 13724 15531 13844 15569
rect 13724 15497 13768 15531
rect 13802 15497 13844 15531
rect 13724 15459 13844 15497
rect 13724 15425 13768 15459
rect 13802 15425 13844 15459
rect 13724 15387 13844 15425
rect 13724 15353 13768 15387
rect 13802 15353 13844 15387
rect 13724 15315 13844 15353
rect 13724 15281 13768 15315
rect 13802 15281 13844 15315
rect 13724 15243 13844 15281
rect 13724 15209 13768 15243
rect 13802 15209 13844 15243
rect 13724 15171 13844 15209
rect 13724 15137 13768 15171
rect 13802 15137 13844 15171
rect 13724 15099 13844 15137
rect 13724 15065 13768 15099
rect 13802 15065 13844 15099
rect 13724 15027 13844 15065
rect 13724 14993 13768 15027
rect 13802 14993 13844 15027
rect 13724 14955 13844 14993
rect 13724 14921 13768 14955
rect 13802 14921 13844 14955
rect 13724 14883 13844 14921
rect 13724 14849 13768 14883
rect 13802 14849 13844 14883
rect 13724 14811 13844 14849
rect 13724 14777 13768 14811
rect 13802 14777 13844 14811
rect 13724 14739 13844 14777
rect 13724 14705 13768 14739
rect 13802 14705 13844 14739
rect 13724 14667 13844 14705
rect 13724 14633 13768 14667
rect 13802 14633 13844 14667
rect 13724 14595 13844 14633
rect 13724 14561 13768 14595
rect 13802 14561 13844 14595
rect 13724 14523 13844 14561
rect 13724 14489 13768 14523
rect 13802 14489 13844 14523
rect 13724 14451 13844 14489
rect 13724 14417 13768 14451
rect 13802 14417 13844 14451
rect 13724 14379 13844 14417
rect 13724 14345 13768 14379
rect 13802 14345 13844 14379
rect 13724 14307 13844 14345
rect 13724 14273 13768 14307
rect 13802 14273 13844 14307
rect 13724 14235 13844 14273
rect 13724 14201 13768 14235
rect 13802 14201 13844 14235
rect 13724 14163 13844 14201
rect 13724 14129 13768 14163
rect 13802 14129 13844 14163
rect 13724 14091 13844 14129
rect 13724 14057 13768 14091
rect 13802 14057 13844 14091
rect 13724 14019 13844 14057
rect 13724 13985 13768 14019
rect 13802 13985 13844 14019
rect 13724 13947 13844 13985
rect 13724 13913 13768 13947
rect 13802 13913 13844 13947
rect 13724 13875 13844 13913
rect 13724 13841 13768 13875
rect 13802 13841 13844 13875
rect 13724 13803 13844 13841
rect 13724 13769 13768 13803
rect 13802 13769 13844 13803
rect 13724 13731 13844 13769
rect 13724 13697 13768 13731
rect 13802 13697 13844 13731
rect 13724 13659 13844 13697
rect 13724 13625 13768 13659
rect 13802 13625 13844 13659
rect 13724 13587 13844 13625
rect 13724 13553 13768 13587
rect 13802 13553 13844 13587
rect 13724 13515 13844 13553
rect 13724 13481 13768 13515
rect 13802 13481 13844 13515
rect 13724 13443 13844 13481
rect 13724 13409 13768 13443
rect 13802 13409 13844 13443
rect 13724 13371 13844 13409
rect 13724 13337 13768 13371
rect 13802 13337 13844 13371
rect 13724 13299 13844 13337
rect 13724 13265 13768 13299
rect 13802 13265 13844 13299
rect 13724 13227 13844 13265
rect 13724 13193 13768 13227
rect 13802 13193 13844 13227
rect 13724 13155 13844 13193
rect 13724 13121 13768 13155
rect 13802 13121 13844 13155
rect 13724 13083 13844 13121
rect 13724 13049 13768 13083
rect 13802 13049 13844 13083
rect 13724 13011 13844 13049
rect 13724 12977 13768 13011
rect 13802 12977 13844 13011
rect 13724 12939 13844 12977
rect 13724 12905 13768 12939
rect 13802 12905 13844 12939
rect 13724 12867 13844 12905
rect 13724 12833 13768 12867
rect 13802 12833 13844 12867
rect 13724 12795 13844 12833
rect 13724 12761 13768 12795
rect 13802 12761 13844 12795
rect 13724 12723 13844 12761
rect 13724 12689 13768 12723
rect 13802 12689 13844 12723
rect 13724 12651 13844 12689
rect 13724 12617 13768 12651
rect 13802 12617 13844 12651
rect 13724 12579 13844 12617
rect 13724 12545 13768 12579
rect 13802 12545 13844 12579
rect 13724 12507 13844 12545
rect 13724 12473 13768 12507
rect 13802 12473 13844 12507
rect 13724 12435 13844 12473
rect 13724 12401 13768 12435
rect 13802 12401 13844 12435
rect 13724 12363 13844 12401
rect 13724 12329 13768 12363
rect 13802 12329 13844 12363
rect 13724 12291 13844 12329
rect 13724 12257 13768 12291
rect 13802 12257 13844 12291
rect 13724 12219 13844 12257
rect 13724 12185 13768 12219
rect 13802 12185 13844 12219
rect 13724 12147 13844 12185
rect 13724 12113 13768 12147
rect 13802 12113 13844 12147
rect 13724 12075 13844 12113
rect 13724 12041 13768 12075
rect 13802 12041 13844 12075
rect 13724 12003 13844 12041
rect 13724 11969 13768 12003
rect 13802 11969 13844 12003
rect 13724 11931 13844 11969
rect 13724 11897 13768 11931
rect 13802 11897 13844 11931
rect 13724 11859 13844 11897
rect 13724 11825 13768 11859
rect 13802 11825 13844 11859
rect 13724 11787 13844 11825
rect 13724 11753 13768 11787
rect 13802 11753 13844 11787
rect 13724 11715 13844 11753
rect 13724 11681 13768 11715
rect 13802 11681 13844 11715
rect 13724 11643 13844 11681
rect 13724 11609 13768 11643
rect 13802 11609 13844 11643
rect 13724 11571 13844 11609
rect 13724 11537 13768 11571
rect 13802 11537 13844 11571
rect 13724 11499 13844 11537
rect 13724 11465 13768 11499
rect 13802 11465 13844 11499
rect 13724 11427 13844 11465
rect 13724 11393 13768 11427
rect 13802 11393 13844 11427
rect 13724 11355 13844 11393
rect 13724 11321 13768 11355
rect 13802 11321 13844 11355
rect 13724 11283 13844 11321
rect 13724 11249 13768 11283
rect 13802 11249 13844 11283
rect 13724 11211 13844 11249
rect 13724 11177 13768 11211
rect 13802 11177 13844 11211
rect 13724 11139 13844 11177
rect 13724 11105 13768 11139
rect 13802 11105 13844 11139
rect 13724 11067 13844 11105
rect 13724 11033 13768 11067
rect 13802 11033 13844 11067
rect 13724 10995 13844 11033
rect 13724 10961 13768 10995
rect 13802 10961 13844 10995
rect 13724 10923 13844 10961
rect 13724 10889 13768 10923
rect 13802 10889 13844 10923
rect 13724 10851 13844 10889
rect 13724 10817 13768 10851
rect 13802 10817 13844 10851
rect 13724 10779 13844 10817
rect 13724 10745 13768 10779
rect 13802 10745 13844 10779
rect 13724 10707 13844 10745
rect 13724 10673 13768 10707
rect 13802 10673 13844 10707
rect 13724 10635 13844 10673
rect 13724 10601 13768 10635
rect 13802 10601 13844 10635
rect 13724 10563 13844 10601
rect 13724 10529 13768 10563
rect 13802 10529 13844 10563
rect 13724 10491 13844 10529
rect 13724 10457 13768 10491
rect 13802 10457 13844 10491
rect 13724 10419 13844 10457
rect 13724 10385 13768 10419
rect 13802 10385 13844 10419
rect 13724 10362 13844 10385
rect 1148 10318 13844 10362
rect 1148 10284 1327 10318
rect 1361 10284 1399 10318
rect 1433 10284 1471 10318
rect 1505 10284 1543 10318
rect 1577 10284 1615 10318
rect 1649 10284 1687 10318
rect 1721 10284 1759 10318
rect 1793 10284 1831 10318
rect 1865 10284 1903 10318
rect 1937 10284 1975 10318
rect 2009 10284 2047 10318
rect 2081 10284 2119 10318
rect 2153 10284 2191 10318
rect 2225 10284 2263 10318
rect 2297 10284 2335 10318
rect 2369 10284 2407 10318
rect 2441 10284 2479 10318
rect 2513 10284 2551 10318
rect 2585 10284 2623 10318
rect 2657 10284 2695 10318
rect 2729 10284 2767 10318
rect 2801 10284 2839 10318
rect 2873 10284 2911 10318
rect 2945 10284 2983 10318
rect 3017 10284 3055 10318
rect 3089 10284 3127 10318
rect 3161 10284 3199 10318
rect 3233 10284 3271 10318
rect 3305 10284 3343 10318
rect 3377 10284 3415 10318
rect 3449 10284 3487 10318
rect 3521 10284 3559 10318
rect 3593 10284 3631 10318
rect 3665 10284 3703 10318
rect 3737 10284 3775 10318
rect 3809 10284 3847 10318
rect 3881 10284 3919 10318
rect 3953 10284 3991 10318
rect 4025 10284 4063 10318
rect 4097 10284 4135 10318
rect 4169 10284 4207 10318
rect 4241 10284 4279 10318
rect 4313 10284 4351 10318
rect 4385 10284 4423 10318
rect 4457 10284 4495 10318
rect 4529 10284 4567 10318
rect 4601 10284 4639 10318
rect 4673 10284 4711 10318
rect 4745 10284 4783 10318
rect 4817 10284 4855 10318
rect 4889 10284 4927 10318
rect 4961 10284 4999 10318
rect 5033 10284 5071 10318
rect 5105 10284 5143 10318
rect 5177 10284 5215 10318
rect 5249 10284 5287 10318
rect 5321 10284 5359 10318
rect 5393 10284 5431 10318
rect 5465 10284 5503 10318
rect 5537 10284 5575 10318
rect 5609 10284 5647 10318
rect 5681 10284 5719 10318
rect 5753 10284 5791 10318
rect 5825 10284 5863 10318
rect 5897 10284 5935 10318
rect 5969 10284 6007 10318
rect 6041 10284 6079 10318
rect 6113 10284 6151 10318
rect 6185 10284 6223 10318
rect 6257 10284 6295 10318
rect 6329 10284 6367 10318
rect 6401 10284 6439 10318
rect 6473 10284 6511 10318
rect 6545 10284 6583 10318
rect 6617 10284 6655 10318
rect 6689 10284 6727 10318
rect 6761 10284 6799 10318
rect 6833 10284 6871 10318
rect 6905 10284 6943 10318
rect 6977 10284 7015 10318
rect 7049 10284 7087 10318
rect 7121 10284 7159 10318
rect 7193 10284 7231 10318
rect 7265 10284 7303 10318
rect 7337 10284 7375 10318
rect 7409 10284 7447 10318
rect 7481 10284 7519 10318
rect 7553 10284 7591 10318
rect 7625 10284 7663 10318
rect 7697 10284 7735 10318
rect 7769 10284 7807 10318
rect 7841 10284 7879 10318
rect 7913 10284 7951 10318
rect 7985 10284 8023 10318
rect 8057 10284 8095 10318
rect 8129 10284 8167 10318
rect 8201 10284 8239 10318
rect 8273 10284 8311 10318
rect 8345 10284 8383 10318
rect 8417 10284 8455 10318
rect 8489 10284 8527 10318
rect 8561 10284 8599 10318
rect 8633 10284 8671 10318
rect 8705 10284 8743 10318
rect 8777 10284 8815 10318
rect 8849 10284 8887 10318
rect 8921 10284 8959 10318
rect 8993 10284 9031 10318
rect 9065 10284 9103 10318
rect 9137 10284 9175 10318
rect 9209 10284 9247 10318
rect 9281 10284 9319 10318
rect 9353 10284 9391 10318
rect 9425 10284 9463 10318
rect 9497 10284 9535 10318
rect 9569 10284 9607 10318
rect 9641 10284 9679 10318
rect 9713 10284 9751 10318
rect 9785 10284 9823 10318
rect 9857 10284 9895 10318
rect 9929 10284 9967 10318
rect 10001 10284 10039 10318
rect 10073 10284 10111 10318
rect 10145 10284 10183 10318
rect 10217 10284 10255 10318
rect 10289 10284 10327 10318
rect 10361 10284 10399 10318
rect 10433 10284 10471 10318
rect 10505 10284 10543 10318
rect 10577 10284 10615 10318
rect 10649 10284 10687 10318
rect 10721 10284 10759 10318
rect 10793 10284 10831 10318
rect 10865 10284 10903 10318
rect 10937 10284 10975 10318
rect 11009 10284 11047 10318
rect 11081 10284 11119 10318
rect 11153 10284 11191 10318
rect 11225 10284 11263 10318
rect 11297 10284 11335 10318
rect 11369 10284 11407 10318
rect 11441 10284 11479 10318
rect 11513 10284 11551 10318
rect 11585 10284 11623 10318
rect 11657 10284 11695 10318
rect 11729 10284 11767 10318
rect 11801 10284 11839 10318
rect 11873 10284 11911 10318
rect 11945 10284 11983 10318
rect 12017 10284 12055 10318
rect 12089 10284 12127 10318
rect 12161 10284 12199 10318
rect 12233 10284 12271 10318
rect 12305 10284 12343 10318
rect 12377 10284 12415 10318
rect 12449 10284 12487 10318
rect 12521 10284 12559 10318
rect 12593 10284 12631 10318
rect 12665 10284 12703 10318
rect 12737 10284 12775 10318
rect 12809 10284 12847 10318
rect 12881 10284 12919 10318
rect 12953 10284 12991 10318
rect 13025 10284 13063 10318
rect 13097 10284 13135 10318
rect 13169 10284 13207 10318
rect 13241 10284 13279 10318
rect 13313 10284 13351 10318
rect 13385 10284 13423 10318
rect 13457 10284 13495 10318
rect 13529 10284 13567 10318
rect 13601 10284 13639 10318
rect 13673 10284 13844 10318
rect 1148 10242 13844 10284
rect 14099 21261 14219 21299
rect 14099 21227 14142 21261
rect 14176 21227 14219 21261
rect 14099 21189 14219 21227
rect 14099 21155 14142 21189
rect 14176 21155 14219 21189
rect 14099 21117 14219 21155
rect 14099 21083 14142 21117
rect 14176 21083 14219 21117
rect 14099 21045 14219 21083
rect 14099 21011 14142 21045
rect 14176 21011 14219 21045
rect 14099 20973 14219 21011
rect 14099 20939 14142 20973
rect 14176 20939 14219 20973
rect 14099 20901 14219 20939
rect 14099 20867 14142 20901
rect 14176 20867 14219 20901
rect 14099 20829 14219 20867
rect 14099 20795 14142 20829
rect 14176 20795 14219 20829
rect 14099 20757 14219 20795
rect 14099 20723 14142 20757
rect 14176 20723 14219 20757
rect 14099 20685 14219 20723
rect 14099 20651 14142 20685
rect 14176 20651 14219 20685
rect 14099 20613 14219 20651
rect 14099 20579 14142 20613
rect 14176 20579 14219 20613
rect 14099 20541 14219 20579
rect 14099 20507 14142 20541
rect 14176 20507 14219 20541
rect 14099 20469 14219 20507
rect 14099 20435 14142 20469
rect 14176 20435 14219 20469
rect 14099 20397 14219 20435
rect 14099 20363 14142 20397
rect 14176 20363 14219 20397
rect 14099 20325 14219 20363
rect 14099 20291 14142 20325
rect 14176 20291 14219 20325
rect 14099 20253 14219 20291
rect 14099 20219 14142 20253
rect 14176 20219 14219 20253
rect 14099 20181 14219 20219
rect 14099 20147 14142 20181
rect 14176 20147 14219 20181
rect 14099 20109 14219 20147
rect 14099 20075 14142 20109
rect 14176 20075 14219 20109
rect 14099 20037 14219 20075
rect 14099 20003 14142 20037
rect 14176 20003 14219 20037
rect 14099 19965 14219 20003
rect 14099 19931 14142 19965
rect 14176 19931 14219 19965
rect 14099 19893 14219 19931
rect 14099 19859 14142 19893
rect 14176 19859 14219 19893
rect 14099 19821 14219 19859
rect 14099 19787 14142 19821
rect 14176 19787 14219 19821
rect 14099 19749 14219 19787
rect 14099 19715 14142 19749
rect 14176 19715 14219 19749
rect 14099 19677 14219 19715
rect 14099 19643 14142 19677
rect 14176 19643 14219 19677
rect 14099 19605 14219 19643
rect 14099 19571 14142 19605
rect 14176 19571 14219 19605
rect 14099 19533 14219 19571
rect 14099 19499 14142 19533
rect 14176 19499 14219 19533
rect 14099 19461 14219 19499
rect 14099 19427 14142 19461
rect 14176 19427 14219 19461
rect 14099 19389 14219 19427
rect 14099 19355 14142 19389
rect 14176 19355 14219 19389
rect 14099 19317 14219 19355
rect 14099 19283 14142 19317
rect 14176 19283 14219 19317
rect 14099 19245 14219 19283
rect 14099 19211 14142 19245
rect 14176 19211 14219 19245
rect 14099 19173 14219 19211
rect 14099 19139 14142 19173
rect 14176 19139 14219 19173
rect 14099 19101 14219 19139
rect 14099 19067 14142 19101
rect 14176 19067 14219 19101
rect 14099 19029 14219 19067
rect 14099 18995 14142 19029
rect 14176 18995 14219 19029
rect 14099 18957 14219 18995
rect 14099 18923 14142 18957
rect 14176 18923 14219 18957
rect 14099 18885 14219 18923
rect 14099 18851 14142 18885
rect 14176 18851 14219 18885
rect 14099 18813 14219 18851
rect 14099 18779 14142 18813
rect 14176 18779 14219 18813
rect 14099 18741 14219 18779
rect 14099 18707 14142 18741
rect 14176 18707 14219 18741
rect 14099 18669 14219 18707
rect 14099 18635 14142 18669
rect 14176 18635 14219 18669
rect 14099 18597 14219 18635
rect 14099 18563 14142 18597
rect 14176 18563 14219 18597
rect 14099 18525 14219 18563
rect 14099 18491 14142 18525
rect 14176 18491 14219 18525
rect 14099 18453 14219 18491
rect 14099 18419 14142 18453
rect 14176 18419 14219 18453
rect 14099 18381 14219 18419
rect 14099 18347 14142 18381
rect 14176 18347 14219 18381
rect 14099 18309 14219 18347
rect 14099 18275 14142 18309
rect 14176 18275 14219 18309
rect 14099 18237 14219 18275
rect 14099 18203 14142 18237
rect 14176 18203 14219 18237
rect 14099 18165 14219 18203
rect 14099 18131 14142 18165
rect 14176 18131 14219 18165
rect 14099 18093 14219 18131
rect 14099 18059 14142 18093
rect 14176 18059 14219 18093
rect 14099 18021 14219 18059
rect 14099 17987 14142 18021
rect 14176 17987 14219 18021
rect 14099 17949 14219 17987
rect 14099 17915 14142 17949
rect 14176 17915 14219 17949
rect 14099 17877 14219 17915
rect 14099 17843 14142 17877
rect 14176 17843 14219 17877
rect 14099 17805 14219 17843
rect 14099 17771 14142 17805
rect 14176 17771 14219 17805
rect 14099 17733 14219 17771
rect 14099 17699 14142 17733
rect 14176 17699 14219 17733
rect 14099 17661 14219 17699
rect 14099 17627 14142 17661
rect 14176 17627 14219 17661
rect 14099 17589 14219 17627
rect 14099 17555 14142 17589
rect 14176 17555 14219 17589
rect 14099 17517 14219 17555
rect 14099 17483 14142 17517
rect 14176 17483 14219 17517
rect 14099 17445 14219 17483
rect 14099 17411 14142 17445
rect 14176 17411 14219 17445
rect 14099 17373 14219 17411
rect 14099 17339 14142 17373
rect 14176 17339 14219 17373
rect 14099 17301 14219 17339
rect 14099 17267 14142 17301
rect 14176 17267 14219 17301
rect 14099 17229 14219 17267
rect 14099 17195 14142 17229
rect 14176 17195 14219 17229
rect 14099 17157 14219 17195
rect 14099 17123 14142 17157
rect 14176 17123 14219 17157
rect 14099 17085 14219 17123
rect 14099 17051 14142 17085
rect 14176 17051 14219 17085
rect 14099 17013 14219 17051
rect 14099 16979 14142 17013
rect 14176 16979 14219 17013
rect 14099 16941 14219 16979
rect 14099 16907 14142 16941
rect 14176 16907 14219 16941
rect 14099 16869 14219 16907
rect 14099 16835 14142 16869
rect 14176 16835 14219 16869
rect 14099 16797 14219 16835
rect 14099 16763 14142 16797
rect 14176 16763 14219 16797
rect 14099 16725 14219 16763
rect 14099 16691 14142 16725
rect 14176 16691 14219 16725
rect 14099 16653 14219 16691
rect 14099 16619 14142 16653
rect 14176 16619 14219 16653
rect 14099 16581 14219 16619
rect 14099 16547 14142 16581
rect 14176 16547 14219 16581
rect 14099 16509 14219 16547
rect 14099 16475 14142 16509
rect 14176 16475 14219 16509
rect 14099 16437 14219 16475
rect 14099 16403 14142 16437
rect 14176 16403 14219 16437
rect 14099 16365 14219 16403
rect 14099 16331 14142 16365
rect 14176 16331 14219 16365
rect 14099 16293 14219 16331
rect 14099 16259 14142 16293
rect 14176 16259 14219 16293
rect 14099 16221 14219 16259
rect 14099 16187 14142 16221
rect 14176 16187 14219 16221
rect 14099 16149 14219 16187
rect 14099 16115 14142 16149
rect 14176 16115 14219 16149
rect 14099 16077 14219 16115
rect 14099 16043 14142 16077
rect 14176 16043 14219 16077
rect 14099 16005 14219 16043
rect 14099 15971 14142 16005
rect 14176 15971 14219 16005
rect 14099 15933 14219 15971
rect 14099 15899 14142 15933
rect 14176 15899 14219 15933
rect 14099 15861 14219 15899
rect 14099 15827 14142 15861
rect 14176 15827 14219 15861
rect 14099 15789 14219 15827
rect 14099 15755 14142 15789
rect 14176 15755 14219 15789
rect 14099 15717 14219 15755
rect 14099 15683 14142 15717
rect 14176 15683 14219 15717
rect 14099 15645 14219 15683
rect 14099 15611 14142 15645
rect 14176 15611 14219 15645
rect 14099 15573 14219 15611
rect 14099 15539 14142 15573
rect 14176 15539 14219 15573
rect 14099 15501 14219 15539
rect 14099 15467 14142 15501
rect 14176 15467 14219 15501
rect 14099 15429 14219 15467
rect 14099 15395 14142 15429
rect 14176 15395 14219 15429
rect 14099 15357 14219 15395
rect 14099 15323 14142 15357
rect 14176 15323 14219 15357
rect 14099 15285 14219 15323
rect 14099 15251 14142 15285
rect 14176 15251 14219 15285
rect 14099 15213 14219 15251
rect 14099 15179 14142 15213
rect 14176 15179 14219 15213
rect 14099 15141 14219 15179
rect 14099 15107 14142 15141
rect 14176 15107 14219 15141
rect 14099 15069 14219 15107
rect 14099 15035 14142 15069
rect 14176 15035 14219 15069
rect 14099 14997 14219 15035
rect 14099 14963 14142 14997
rect 14176 14963 14219 14997
rect 14099 14925 14219 14963
rect 14099 14891 14142 14925
rect 14176 14891 14219 14925
rect 14099 14853 14219 14891
rect 14099 14819 14142 14853
rect 14176 14819 14219 14853
rect 14099 14781 14219 14819
rect 14099 14747 14142 14781
rect 14176 14747 14219 14781
rect 14099 14709 14219 14747
rect 14099 14675 14142 14709
rect 14176 14675 14219 14709
rect 14099 14637 14219 14675
rect 14099 14603 14142 14637
rect 14176 14603 14219 14637
rect 14099 14565 14219 14603
rect 14099 14531 14142 14565
rect 14176 14531 14219 14565
rect 14099 14493 14219 14531
rect 14099 14459 14142 14493
rect 14176 14459 14219 14493
rect 14099 14421 14219 14459
rect 14099 14387 14142 14421
rect 14176 14387 14219 14421
rect 14099 14349 14219 14387
rect 14099 14315 14142 14349
rect 14176 14315 14219 14349
rect 14099 14277 14219 14315
rect 14099 14243 14142 14277
rect 14176 14243 14219 14277
rect 14099 14205 14219 14243
rect 14099 14171 14142 14205
rect 14176 14171 14219 14205
rect 14099 14133 14219 14171
rect 14099 14099 14142 14133
rect 14176 14099 14219 14133
rect 14099 14061 14219 14099
rect 14099 14027 14142 14061
rect 14176 14027 14219 14061
rect 14099 13989 14219 14027
rect 14099 13955 14142 13989
rect 14176 13955 14219 13989
rect 14099 13917 14219 13955
rect 14099 13883 14142 13917
rect 14176 13883 14219 13917
rect 14099 13845 14219 13883
rect 14099 13811 14142 13845
rect 14176 13811 14219 13845
rect 14099 13773 14219 13811
rect 14099 13739 14142 13773
rect 14176 13739 14219 13773
rect 14099 13701 14219 13739
rect 14099 13667 14142 13701
rect 14176 13667 14219 13701
rect 14099 13629 14219 13667
rect 14099 13595 14142 13629
rect 14176 13595 14219 13629
rect 14099 13557 14219 13595
rect 14099 13523 14142 13557
rect 14176 13523 14219 13557
rect 14099 13485 14219 13523
rect 14099 13451 14142 13485
rect 14176 13451 14219 13485
rect 14099 13413 14219 13451
rect 14099 13379 14142 13413
rect 14176 13379 14219 13413
rect 14099 13341 14219 13379
rect 14099 13307 14142 13341
rect 14176 13307 14219 13341
rect 14099 13269 14219 13307
rect 14099 13235 14142 13269
rect 14176 13235 14219 13269
rect 14099 13197 14219 13235
rect 14099 13163 14142 13197
rect 14176 13163 14219 13197
rect 14099 13125 14219 13163
rect 14099 13091 14142 13125
rect 14176 13091 14219 13125
rect 14099 13053 14219 13091
rect 14099 13019 14142 13053
rect 14176 13019 14219 13053
rect 14099 12981 14219 13019
rect 14099 12947 14142 12981
rect 14176 12947 14219 12981
rect 14099 12909 14219 12947
rect 14099 12875 14142 12909
rect 14176 12875 14219 12909
rect 14099 12837 14219 12875
rect 14099 12803 14142 12837
rect 14176 12803 14219 12837
rect 14099 12765 14219 12803
rect 14099 12731 14142 12765
rect 14176 12731 14219 12765
rect 14099 12693 14219 12731
rect 14099 12659 14142 12693
rect 14176 12659 14219 12693
rect 14099 12621 14219 12659
rect 14099 12587 14142 12621
rect 14176 12587 14219 12621
rect 14099 12549 14219 12587
rect 14099 12515 14142 12549
rect 14176 12515 14219 12549
rect 14099 12477 14219 12515
rect 14099 12443 14142 12477
rect 14176 12443 14219 12477
rect 14099 12405 14219 12443
rect 14099 12371 14142 12405
rect 14176 12371 14219 12405
rect 14099 12333 14219 12371
rect 14099 12299 14142 12333
rect 14176 12299 14219 12333
rect 14099 12261 14219 12299
rect 14099 12227 14142 12261
rect 14176 12227 14219 12261
rect 14099 12189 14219 12227
rect 14099 12155 14142 12189
rect 14176 12155 14219 12189
rect 14099 12117 14219 12155
rect 14099 12083 14142 12117
rect 14176 12083 14219 12117
rect 14099 12045 14219 12083
rect 14099 12011 14142 12045
rect 14176 12011 14219 12045
rect 14099 11973 14219 12011
rect 14099 11939 14142 11973
rect 14176 11939 14219 11973
rect 14099 11901 14219 11939
rect 14099 11867 14142 11901
rect 14176 11867 14219 11901
rect 14099 11829 14219 11867
rect 14099 11795 14142 11829
rect 14176 11795 14219 11829
rect 14099 11757 14219 11795
rect 14099 11723 14142 11757
rect 14176 11723 14219 11757
rect 14099 11685 14219 11723
rect 14099 11651 14142 11685
rect 14176 11651 14219 11685
rect 14099 11613 14219 11651
rect 14099 11579 14142 11613
rect 14176 11579 14219 11613
rect 14099 11541 14219 11579
rect 14099 11507 14142 11541
rect 14176 11507 14219 11541
rect 14099 11469 14219 11507
rect 14099 11435 14142 11469
rect 14176 11435 14219 11469
rect 14099 11397 14219 11435
rect 14099 11363 14142 11397
rect 14176 11363 14219 11397
rect 14099 11325 14219 11363
rect 14099 11291 14142 11325
rect 14176 11291 14219 11325
rect 14099 11253 14219 11291
rect 14099 11219 14142 11253
rect 14176 11219 14219 11253
rect 14099 11181 14219 11219
rect 14099 11147 14142 11181
rect 14176 11147 14219 11181
rect 14099 11109 14219 11147
rect 14099 11075 14142 11109
rect 14176 11075 14219 11109
rect 14099 11037 14219 11075
rect 14099 11003 14142 11037
rect 14176 11003 14219 11037
rect 14099 10965 14219 11003
rect 14099 10931 14142 10965
rect 14176 10931 14219 10965
rect 14099 10893 14219 10931
rect 14099 10859 14142 10893
rect 14176 10859 14219 10893
rect 14099 10821 14219 10859
rect 14099 10787 14142 10821
rect 14176 10787 14219 10821
rect 14099 10749 14219 10787
rect 14099 10715 14142 10749
rect 14176 10715 14219 10749
rect 14099 10677 14219 10715
rect 14099 10643 14142 10677
rect 14176 10643 14219 10677
rect 14099 10605 14219 10643
rect 14099 10571 14142 10605
rect 14176 10571 14219 10605
rect 14099 10533 14219 10571
rect 14099 10499 14142 10533
rect 14176 10499 14219 10533
rect 14099 10461 14219 10499
rect 14099 10427 14142 10461
rect 14176 10427 14219 10461
rect 14099 10389 14219 10427
rect 14099 10355 14142 10389
rect 14176 10355 14219 10389
rect 14099 10317 14219 10355
rect 14099 10283 14142 10317
rect 14176 10283 14219 10317
rect 14099 10245 14219 10283
rect 757 10180 877 10218
rect 757 10146 807 10180
rect 841 10146 877 10180
rect 757 10108 877 10146
rect 757 10074 807 10108
rect 841 10074 877 10108
rect 757 9982 877 10074
rect 14099 10211 14142 10245
rect 14176 10211 14219 10245
rect 14099 10173 14219 10211
rect 14099 10139 14142 10173
rect 14176 10139 14219 10173
rect 14099 10101 14219 10139
rect 14099 10067 14142 10101
rect 14176 10067 14219 10101
tri 877 9982 898 10003 sw
tri 14078 9982 14099 10003 se
rect 14099 9982 14219 10067
rect 757 9963 898 9982
tri 898 9963 917 9982 sw
tri 14059 9963 14078 9982 se
rect 14078 9963 14219 9982
rect 757 9943 14219 9963
tri 757 9942 758 9943 ne
rect 758 9942 14186 9943
rect 245 9879 320 9913
rect 354 9879 430 9913
tri 758 9908 792 9942 ne
rect 792 9908 891 9942
rect 925 9908 963 9942
rect 997 9908 1035 9942
rect 1069 9908 1107 9942
rect 1141 9908 1179 9942
rect 1213 9908 1251 9942
rect 1285 9908 1323 9942
rect 1357 9908 1395 9942
rect 1429 9908 1467 9942
rect 1501 9908 1539 9942
rect 1573 9908 1611 9942
rect 1645 9908 1683 9942
rect 1717 9908 1755 9942
rect 1789 9908 1827 9942
rect 1861 9908 1899 9942
rect 1933 9908 1971 9942
rect 2005 9908 2043 9942
rect 2077 9908 2115 9942
rect 2149 9908 2187 9942
rect 2221 9908 2259 9942
rect 2293 9908 2331 9942
rect 2365 9908 2403 9942
rect 2437 9908 2475 9942
rect 2509 9908 2547 9942
rect 2581 9908 2619 9942
rect 2653 9908 2691 9942
rect 2725 9908 2763 9942
rect 2797 9908 2835 9942
rect 2869 9908 2907 9942
rect 2941 9908 2979 9942
rect 3013 9908 3051 9942
rect 3085 9908 3123 9942
rect 3157 9908 3195 9942
rect 3229 9908 3267 9942
rect 3301 9908 3339 9942
rect 3373 9908 3411 9942
rect 3445 9908 3483 9942
rect 3517 9908 3555 9942
rect 3589 9908 3627 9942
rect 3661 9908 3699 9942
rect 3733 9908 3771 9942
rect 3805 9908 3843 9942
rect 3877 9908 3915 9942
rect 3949 9908 3987 9942
rect 4021 9908 4059 9942
rect 4093 9908 4131 9942
rect 4165 9908 4203 9942
rect 4237 9908 4275 9942
rect 4309 9908 4347 9942
rect 4381 9908 4419 9942
rect 4453 9908 4491 9942
rect 4525 9908 4563 9942
rect 4597 9908 4635 9942
rect 4669 9908 4707 9942
rect 4741 9908 4779 9942
rect 4813 9908 4851 9942
rect 4885 9908 4923 9942
rect 4957 9908 4995 9942
rect 5029 9908 5067 9942
rect 5101 9908 5139 9942
rect 5173 9908 5211 9942
rect 5245 9908 5283 9942
rect 5317 9908 5355 9942
rect 5389 9908 5427 9942
rect 5461 9908 5499 9942
rect 5533 9908 5571 9942
rect 5605 9908 5643 9942
rect 5677 9908 5715 9942
rect 5749 9908 5787 9942
rect 5821 9908 5859 9942
rect 5893 9908 5931 9942
rect 5965 9908 6003 9942
rect 6037 9908 6075 9942
rect 6109 9908 6147 9942
rect 6181 9908 6219 9942
rect 6253 9908 6291 9942
rect 6325 9908 6363 9942
rect 6397 9908 6435 9942
rect 6469 9908 6507 9942
rect 6541 9908 6579 9942
rect 6613 9908 6651 9942
rect 6685 9908 6723 9942
rect 6757 9908 6795 9942
rect 6829 9908 6867 9942
rect 6901 9908 6939 9942
rect 6973 9908 7011 9942
rect 7045 9908 7083 9942
rect 7117 9908 7155 9942
rect 7189 9908 7227 9942
rect 7261 9908 7299 9942
rect 7333 9908 7371 9942
rect 7405 9908 7443 9942
rect 7477 9908 7515 9942
rect 7549 9908 7587 9942
rect 7621 9908 7659 9942
rect 7693 9908 7731 9942
rect 7765 9908 7803 9942
rect 7837 9908 7875 9942
rect 7909 9908 7947 9942
rect 7981 9908 8019 9942
rect 8053 9908 8091 9942
rect 8125 9908 8163 9942
rect 8197 9908 8235 9942
rect 8269 9908 8307 9942
rect 8341 9908 8379 9942
rect 8413 9908 8451 9942
rect 8485 9908 8523 9942
rect 8557 9908 8595 9942
rect 8629 9908 8667 9942
rect 8701 9908 8739 9942
rect 8773 9908 8811 9942
rect 8845 9908 8883 9942
rect 8917 9908 8955 9942
rect 8989 9908 9027 9942
rect 9061 9908 9099 9942
rect 9133 9908 9171 9942
rect 9205 9908 9243 9942
rect 9277 9908 9315 9942
rect 9349 9908 9387 9942
rect 9421 9908 9459 9942
rect 9493 9908 9531 9942
rect 9565 9908 9603 9942
rect 9637 9908 9675 9942
rect 9709 9908 9747 9942
rect 9781 9908 9819 9942
rect 9853 9908 9891 9942
rect 9925 9908 9963 9942
rect 9997 9908 10035 9942
rect 10069 9908 10107 9942
rect 10141 9908 10179 9942
rect 10213 9908 10251 9942
rect 10285 9908 10323 9942
rect 10357 9908 10395 9942
rect 10429 9908 10467 9942
rect 10501 9908 10539 9942
rect 10573 9908 10611 9942
rect 10645 9908 10683 9942
rect 10717 9908 10755 9942
rect 10789 9908 10827 9942
rect 10861 9908 10899 9942
rect 10933 9908 10971 9942
rect 11005 9908 11043 9942
rect 11077 9908 11115 9942
rect 11149 9908 11187 9942
rect 11221 9908 11259 9942
rect 11293 9908 11331 9942
rect 11365 9908 11403 9942
rect 11437 9908 11475 9942
rect 11509 9908 11547 9942
rect 11581 9908 11619 9942
rect 11653 9908 11691 9942
rect 11725 9908 11763 9942
rect 11797 9908 11835 9942
rect 11869 9908 11907 9942
rect 11941 9908 11979 9942
rect 12013 9908 12051 9942
rect 12085 9908 12123 9942
rect 12157 9908 12195 9942
rect 12229 9908 12267 9942
rect 12301 9908 12339 9942
rect 12373 9908 12411 9942
rect 12445 9908 12483 9942
rect 12517 9908 12555 9942
rect 12589 9908 12627 9942
rect 12661 9908 12699 9942
rect 12733 9908 12771 9942
rect 12805 9908 12843 9942
rect 12877 9908 12915 9942
rect 12949 9908 12987 9942
rect 13021 9908 13059 9942
rect 13093 9908 13131 9942
rect 13165 9908 13203 9942
rect 13237 9908 13275 9942
rect 13309 9908 13347 9942
rect 13381 9908 13419 9942
rect 13453 9908 13491 9942
rect 13525 9908 13563 9942
rect 13597 9908 13635 9942
rect 13669 9908 13707 9942
rect 13741 9908 13779 9942
rect 13813 9908 13851 9942
rect 13885 9908 13923 9942
rect 13957 9908 13995 9942
rect 14029 9910 14186 9942
tri 14186 9910 14219 9943 nw
rect 14539 35940 14614 35974
rect 14648 35940 14724 35974
rect 14539 35902 14724 35940
rect 14539 35868 14614 35902
rect 14648 35868 14724 35902
rect 14539 35830 14724 35868
rect 14539 35796 14614 35830
rect 14648 35796 14724 35830
rect 14539 35758 14724 35796
rect 14539 35724 14614 35758
rect 14648 35724 14724 35758
rect 14539 35686 14724 35724
rect 14539 35652 14614 35686
rect 14648 35652 14724 35686
rect 14539 35614 14724 35652
rect 14539 35580 14614 35614
rect 14648 35580 14724 35614
rect 14539 35542 14724 35580
rect 14539 35508 14614 35542
rect 14648 35508 14724 35542
rect 14539 35470 14724 35508
rect 14539 35436 14614 35470
rect 14648 35436 14724 35470
rect 14539 35398 14724 35436
rect 14539 35364 14614 35398
rect 14648 35364 14724 35398
rect 14539 35326 14724 35364
rect 14539 35292 14614 35326
rect 14648 35292 14724 35326
rect 14539 35254 14724 35292
rect 14539 35220 14614 35254
rect 14648 35220 14724 35254
rect 14539 35182 14724 35220
rect 14539 35148 14614 35182
rect 14648 35148 14724 35182
rect 14539 35110 14724 35148
rect 14539 35076 14614 35110
rect 14648 35076 14724 35110
rect 14539 35038 14724 35076
rect 14539 35004 14614 35038
rect 14648 35004 14724 35038
rect 14539 34966 14724 35004
rect 14539 34932 14614 34966
rect 14648 34932 14724 34966
rect 14539 34894 14724 34932
rect 14539 34860 14614 34894
rect 14648 34860 14724 34894
rect 14539 34822 14724 34860
rect 14539 34788 14614 34822
rect 14648 34788 14724 34822
rect 14539 34750 14724 34788
rect 14539 34716 14614 34750
rect 14648 34716 14724 34750
rect 14539 34678 14724 34716
rect 14539 34644 14614 34678
rect 14648 34644 14724 34678
rect 14539 34606 14724 34644
rect 14539 34572 14614 34606
rect 14648 34572 14724 34606
rect 14539 34534 14724 34572
rect 14539 34500 14614 34534
rect 14648 34500 14724 34534
rect 14539 34462 14724 34500
rect 14539 34428 14614 34462
rect 14648 34428 14724 34462
rect 14539 34390 14724 34428
rect 14539 34356 14614 34390
rect 14648 34356 14724 34390
rect 14539 34318 14724 34356
rect 14539 34284 14614 34318
rect 14648 34284 14724 34318
rect 14539 34246 14724 34284
rect 14539 34212 14614 34246
rect 14648 34212 14724 34246
rect 14539 34174 14724 34212
rect 14539 34140 14614 34174
rect 14648 34140 14724 34174
rect 14539 34102 14724 34140
rect 14539 34068 14614 34102
rect 14648 34068 14724 34102
rect 14539 34030 14724 34068
rect 14539 33996 14614 34030
rect 14648 33996 14724 34030
rect 14539 33958 14724 33996
rect 14539 33924 14614 33958
rect 14648 33924 14724 33958
rect 14539 33886 14724 33924
rect 14539 33852 14614 33886
rect 14648 33852 14724 33886
rect 14539 33814 14724 33852
rect 14539 33780 14614 33814
rect 14648 33780 14724 33814
rect 14539 33742 14724 33780
rect 14539 33708 14614 33742
rect 14648 33708 14724 33742
rect 14539 33670 14724 33708
rect 14539 33636 14614 33670
rect 14648 33636 14724 33670
rect 14539 33598 14724 33636
rect 14539 33564 14614 33598
rect 14648 33564 14724 33598
rect 14539 33526 14724 33564
rect 14539 33492 14614 33526
rect 14648 33492 14724 33526
rect 14539 33454 14724 33492
rect 14539 33420 14614 33454
rect 14648 33420 14724 33454
rect 14539 33382 14724 33420
rect 14539 33348 14614 33382
rect 14648 33348 14724 33382
rect 14539 33310 14724 33348
rect 14539 33276 14614 33310
rect 14648 33276 14724 33310
rect 14539 33238 14724 33276
rect 14539 33204 14614 33238
rect 14648 33204 14724 33238
rect 14539 33166 14724 33204
rect 14539 33132 14614 33166
rect 14648 33132 14724 33166
rect 14539 33094 14724 33132
rect 14539 33060 14614 33094
rect 14648 33060 14724 33094
rect 14539 33022 14724 33060
rect 14539 32988 14614 33022
rect 14648 32988 14724 33022
rect 14539 32950 14724 32988
rect 14539 32916 14614 32950
rect 14648 32916 14724 32950
rect 14539 32878 14724 32916
rect 14539 32844 14614 32878
rect 14648 32844 14724 32878
rect 14539 32806 14724 32844
rect 14539 32772 14614 32806
rect 14648 32772 14724 32806
rect 14539 32734 14724 32772
rect 14539 32700 14614 32734
rect 14648 32700 14724 32734
rect 14539 32662 14724 32700
rect 14539 32628 14614 32662
rect 14648 32628 14724 32662
rect 14539 32590 14724 32628
rect 14539 32556 14614 32590
rect 14648 32556 14724 32590
rect 14539 32518 14724 32556
rect 14539 32484 14614 32518
rect 14648 32484 14724 32518
rect 14539 32446 14724 32484
rect 14539 32412 14614 32446
rect 14648 32412 14724 32446
rect 14539 32374 14724 32412
rect 14539 32340 14614 32374
rect 14648 32340 14724 32374
rect 14539 32302 14724 32340
rect 14539 32268 14614 32302
rect 14648 32268 14724 32302
rect 14539 32230 14724 32268
rect 14539 32196 14614 32230
rect 14648 32196 14724 32230
rect 14539 32158 14724 32196
rect 14539 32124 14614 32158
rect 14648 32124 14724 32158
rect 14539 32086 14724 32124
rect 14539 32052 14614 32086
rect 14648 32052 14724 32086
rect 14539 32014 14724 32052
rect 14539 31980 14614 32014
rect 14648 31980 14724 32014
rect 14539 31942 14724 31980
rect 14539 31908 14614 31942
rect 14648 31908 14724 31942
rect 14539 31870 14724 31908
rect 14539 31836 14614 31870
rect 14648 31836 14724 31870
rect 14539 31798 14724 31836
rect 14539 31764 14614 31798
rect 14648 31764 14724 31798
rect 14539 31726 14724 31764
rect 14539 31692 14614 31726
rect 14648 31692 14724 31726
rect 14539 31654 14724 31692
rect 14539 31620 14614 31654
rect 14648 31620 14724 31654
rect 14539 31582 14724 31620
rect 14539 31548 14614 31582
rect 14648 31548 14724 31582
rect 14539 31510 14724 31548
rect 14539 31476 14614 31510
rect 14648 31476 14724 31510
rect 14539 31438 14724 31476
rect 14539 31404 14614 31438
rect 14648 31404 14724 31438
rect 14539 31366 14724 31404
rect 14539 31332 14614 31366
rect 14648 31332 14724 31366
rect 14539 31294 14724 31332
rect 14539 31260 14614 31294
rect 14648 31260 14724 31294
rect 14539 31222 14724 31260
rect 14539 31188 14614 31222
rect 14648 31188 14724 31222
rect 14539 31150 14724 31188
rect 14539 31116 14614 31150
rect 14648 31116 14724 31150
rect 14539 31078 14724 31116
rect 14539 31044 14614 31078
rect 14648 31044 14724 31078
rect 14539 31006 14724 31044
rect 14539 30972 14614 31006
rect 14648 30972 14724 31006
rect 14539 30934 14724 30972
rect 14539 30900 14614 30934
rect 14648 30900 14724 30934
rect 14539 30862 14724 30900
rect 14539 30828 14614 30862
rect 14648 30828 14724 30862
rect 14539 30790 14724 30828
rect 14539 30756 14614 30790
rect 14648 30756 14724 30790
rect 14539 30718 14724 30756
rect 14539 30684 14614 30718
rect 14648 30684 14724 30718
rect 14539 30646 14724 30684
rect 14539 30612 14614 30646
rect 14648 30612 14724 30646
rect 14539 30574 14724 30612
rect 14539 30540 14614 30574
rect 14648 30540 14724 30574
rect 14539 30502 14724 30540
rect 14539 30468 14614 30502
rect 14648 30468 14724 30502
rect 14539 30430 14724 30468
rect 14539 30396 14614 30430
rect 14648 30396 14724 30430
rect 14539 30358 14724 30396
rect 14539 30324 14614 30358
rect 14648 30324 14724 30358
rect 14539 30286 14724 30324
rect 14539 30252 14614 30286
rect 14648 30252 14724 30286
rect 14539 30214 14724 30252
rect 14539 30180 14614 30214
rect 14648 30180 14724 30214
rect 14539 30142 14724 30180
rect 14539 30108 14614 30142
rect 14648 30108 14724 30142
rect 14539 30070 14724 30108
rect 14539 30036 14614 30070
rect 14648 30036 14724 30070
rect 14539 29998 14724 30036
rect 14539 29964 14614 29998
rect 14648 29964 14724 29998
rect 14539 29926 14724 29964
rect 14539 29892 14614 29926
rect 14648 29892 14724 29926
rect 14539 29854 14724 29892
rect 14539 29820 14614 29854
rect 14648 29820 14724 29854
rect 14539 29782 14724 29820
rect 14539 29748 14614 29782
rect 14648 29748 14724 29782
rect 14539 29710 14724 29748
rect 14539 29676 14614 29710
rect 14648 29676 14724 29710
rect 14539 29638 14724 29676
rect 14539 29604 14614 29638
rect 14648 29604 14724 29638
rect 14539 29566 14724 29604
rect 14539 29532 14614 29566
rect 14648 29532 14724 29566
rect 14539 29494 14724 29532
rect 14539 29460 14614 29494
rect 14648 29460 14724 29494
rect 14539 29422 14724 29460
rect 14539 29388 14614 29422
rect 14648 29388 14724 29422
rect 14539 29350 14724 29388
rect 14539 29316 14614 29350
rect 14648 29316 14724 29350
rect 14539 29278 14724 29316
rect 14539 29244 14614 29278
rect 14648 29244 14724 29278
rect 14539 29206 14724 29244
rect 14539 29172 14614 29206
rect 14648 29172 14724 29206
rect 14539 29134 14724 29172
rect 14539 29100 14614 29134
rect 14648 29100 14724 29134
rect 14539 29062 14724 29100
rect 14539 29028 14614 29062
rect 14648 29028 14724 29062
rect 14539 28990 14724 29028
rect 14539 28956 14614 28990
rect 14648 28956 14724 28990
rect 14539 28918 14724 28956
rect 14539 28884 14614 28918
rect 14648 28884 14724 28918
rect 14539 28846 14724 28884
rect 14539 28812 14614 28846
rect 14648 28812 14724 28846
rect 14539 28774 14724 28812
rect 14539 28740 14614 28774
rect 14648 28740 14724 28774
rect 14539 28702 14724 28740
rect 14539 28668 14614 28702
rect 14648 28668 14724 28702
rect 14539 28630 14724 28668
rect 14539 28596 14614 28630
rect 14648 28596 14724 28630
rect 14539 28558 14724 28596
rect 14539 28524 14614 28558
rect 14648 28524 14724 28558
rect 14539 28486 14724 28524
rect 14539 28452 14614 28486
rect 14648 28452 14724 28486
rect 14539 28414 14724 28452
rect 14539 28380 14614 28414
rect 14648 28380 14724 28414
rect 14539 28342 14724 28380
rect 14539 28308 14614 28342
rect 14648 28308 14724 28342
rect 14539 28270 14724 28308
rect 14539 28236 14614 28270
rect 14648 28236 14724 28270
rect 14539 28198 14724 28236
rect 14539 28164 14614 28198
rect 14648 28164 14724 28198
rect 14539 28126 14724 28164
rect 14539 28092 14614 28126
rect 14648 28092 14724 28126
rect 14539 28054 14724 28092
rect 14539 28020 14614 28054
rect 14648 28020 14724 28054
rect 14539 27982 14724 28020
rect 14539 27948 14614 27982
rect 14648 27948 14724 27982
rect 14539 27910 14724 27948
rect 14539 27876 14614 27910
rect 14648 27876 14724 27910
rect 14539 27838 14724 27876
rect 14539 27804 14614 27838
rect 14648 27804 14724 27838
rect 14539 27766 14724 27804
rect 14539 27732 14614 27766
rect 14648 27732 14724 27766
rect 14539 27694 14724 27732
rect 14539 27660 14614 27694
rect 14648 27660 14724 27694
rect 14539 27622 14724 27660
rect 14539 27588 14614 27622
rect 14648 27588 14724 27622
rect 14539 27550 14724 27588
rect 14539 27516 14614 27550
rect 14648 27516 14724 27550
rect 14539 27478 14724 27516
rect 14539 27444 14614 27478
rect 14648 27444 14724 27478
rect 14539 27406 14724 27444
rect 14539 27372 14614 27406
rect 14648 27372 14724 27406
rect 14539 27334 14724 27372
rect 14539 27300 14614 27334
rect 14648 27300 14724 27334
rect 14539 27262 14724 27300
rect 14539 27228 14614 27262
rect 14648 27228 14724 27262
rect 14539 27190 14724 27228
rect 14539 27156 14614 27190
rect 14648 27156 14724 27190
rect 14539 27118 14724 27156
rect 14539 27084 14614 27118
rect 14648 27084 14724 27118
rect 14539 27046 14724 27084
rect 14539 27012 14614 27046
rect 14648 27012 14724 27046
rect 14539 26974 14724 27012
rect 14539 26940 14614 26974
rect 14648 26940 14724 26974
rect 14539 26902 14724 26940
rect 14539 26868 14614 26902
rect 14648 26868 14724 26902
rect 14539 26830 14724 26868
rect 14539 26796 14614 26830
rect 14648 26796 14724 26830
rect 14539 26758 14724 26796
rect 14539 26724 14614 26758
rect 14648 26724 14724 26758
rect 14539 26686 14724 26724
rect 14539 26652 14614 26686
rect 14648 26652 14724 26686
rect 14539 26614 14724 26652
rect 14539 26580 14614 26614
rect 14648 26580 14724 26614
rect 14539 26542 14724 26580
rect 14539 26508 14614 26542
rect 14648 26508 14724 26542
rect 14539 26470 14724 26508
rect 14539 26436 14614 26470
rect 14648 26436 14724 26470
rect 14539 26398 14724 26436
rect 14539 26364 14614 26398
rect 14648 26364 14724 26398
rect 14539 26326 14724 26364
rect 14539 26292 14614 26326
rect 14648 26292 14724 26326
rect 14539 26254 14724 26292
rect 14539 26220 14614 26254
rect 14648 26220 14724 26254
rect 14539 26182 14724 26220
rect 14539 26148 14614 26182
rect 14648 26148 14724 26182
rect 14539 26110 14724 26148
rect 14539 26076 14614 26110
rect 14648 26076 14724 26110
rect 14539 26038 14724 26076
rect 14539 26004 14614 26038
rect 14648 26004 14724 26038
rect 14539 25966 14724 26004
rect 14539 25932 14614 25966
rect 14648 25932 14724 25966
rect 14539 25894 14724 25932
rect 14539 25860 14614 25894
rect 14648 25860 14724 25894
rect 14539 25822 14724 25860
rect 14539 25788 14614 25822
rect 14648 25788 14724 25822
rect 14539 25750 14724 25788
rect 14539 25716 14614 25750
rect 14648 25716 14724 25750
rect 14539 25678 14724 25716
rect 14539 25644 14614 25678
rect 14648 25644 14724 25678
rect 14539 25606 14724 25644
rect 14539 25572 14614 25606
rect 14648 25572 14724 25606
rect 14539 25534 14724 25572
rect 14539 25500 14614 25534
rect 14648 25500 14724 25534
rect 14539 25462 14724 25500
rect 14539 25428 14614 25462
rect 14648 25428 14724 25462
rect 14539 25390 14724 25428
rect 14539 25356 14614 25390
rect 14648 25356 14724 25390
rect 14539 25318 14724 25356
rect 14539 25284 14614 25318
rect 14648 25284 14724 25318
rect 14539 25246 14724 25284
rect 14539 25212 14614 25246
rect 14648 25212 14724 25246
rect 14539 25174 14724 25212
rect 14539 25140 14614 25174
rect 14648 25140 14724 25174
rect 14539 25102 14724 25140
rect 14539 25068 14614 25102
rect 14648 25068 14724 25102
rect 14539 25030 14724 25068
rect 14539 24996 14614 25030
rect 14648 24996 14724 25030
rect 14539 24958 14724 24996
rect 14539 24924 14614 24958
rect 14648 24924 14724 24958
rect 14539 24886 14724 24924
rect 14539 24852 14614 24886
rect 14648 24852 14724 24886
rect 14539 24814 14724 24852
rect 14539 24780 14614 24814
rect 14648 24780 14724 24814
rect 14539 24742 14724 24780
rect 14539 24708 14614 24742
rect 14648 24708 14724 24742
rect 14539 24670 14724 24708
rect 14539 24636 14614 24670
rect 14648 24636 14724 24670
rect 14539 24598 14724 24636
rect 14539 24564 14614 24598
rect 14648 24564 14724 24598
rect 14539 24526 14724 24564
rect 14539 24492 14614 24526
rect 14648 24492 14724 24526
rect 14539 24454 14724 24492
rect 14539 24420 14614 24454
rect 14648 24420 14724 24454
rect 14539 24382 14724 24420
rect 14539 24348 14614 24382
rect 14648 24348 14724 24382
rect 14539 24310 14724 24348
rect 14539 24276 14614 24310
rect 14648 24276 14724 24310
rect 14539 24238 14724 24276
rect 14539 24204 14614 24238
rect 14648 24204 14724 24238
rect 14539 24166 14724 24204
rect 14539 24132 14614 24166
rect 14648 24132 14724 24166
rect 14539 24094 14724 24132
rect 14539 24060 14614 24094
rect 14648 24060 14724 24094
rect 14539 24022 14724 24060
rect 14539 23988 14614 24022
rect 14648 23988 14724 24022
rect 14539 23950 14724 23988
rect 14539 23916 14614 23950
rect 14648 23916 14724 23950
rect 14539 23878 14724 23916
rect 14539 23844 14614 23878
rect 14648 23844 14724 23878
rect 14539 23806 14724 23844
rect 14539 23772 14614 23806
rect 14648 23772 14724 23806
rect 14539 23734 14724 23772
rect 14539 23700 14614 23734
rect 14648 23700 14724 23734
rect 14539 23662 14724 23700
rect 14539 23628 14614 23662
rect 14648 23628 14724 23662
rect 14539 23590 14724 23628
rect 14539 23556 14614 23590
rect 14648 23556 14724 23590
rect 14539 23518 14724 23556
rect 14539 23484 14614 23518
rect 14648 23484 14724 23518
rect 14539 23446 14724 23484
rect 14539 23412 14614 23446
rect 14648 23412 14724 23446
rect 14539 23374 14724 23412
rect 14539 23340 14614 23374
rect 14648 23340 14724 23374
rect 14539 23302 14724 23340
rect 14539 23268 14614 23302
rect 14648 23268 14724 23302
rect 14539 23230 14724 23268
rect 14539 23196 14614 23230
rect 14648 23196 14724 23230
rect 14539 23158 14724 23196
rect 14539 23124 14614 23158
rect 14648 23124 14724 23158
rect 14539 23086 14724 23124
rect 14539 23052 14614 23086
rect 14648 23052 14724 23086
rect 14539 23014 14724 23052
rect 14539 22980 14614 23014
rect 14648 22980 14724 23014
rect 14539 22942 14724 22980
rect 14539 22908 14614 22942
rect 14648 22908 14724 22942
rect 14539 22870 14724 22908
rect 14539 22836 14614 22870
rect 14648 22836 14724 22870
rect 14539 22798 14724 22836
rect 14539 22764 14614 22798
rect 14648 22764 14724 22798
rect 14539 22726 14724 22764
rect 14539 22692 14614 22726
rect 14648 22692 14724 22726
rect 14539 22654 14724 22692
rect 14539 22620 14614 22654
rect 14648 22620 14724 22654
rect 14539 22582 14724 22620
rect 14539 22548 14614 22582
rect 14648 22548 14724 22582
rect 14539 22510 14724 22548
rect 14539 22476 14614 22510
rect 14648 22476 14724 22510
rect 14539 22438 14724 22476
rect 14539 22404 14614 22438
rect 14648 22404 14724 22438
rect 14539 22366 14724 22404
rect 14539 22332 14614 22366
rect 14648 22332 14724 22366
rect 14539 22294 14724 22332
rect 14539 22260 14614 22294
rect 14648 22260 14724 22294
rect 14539 22222 14724 22260
rect 14539 22188 14614 22222
rect 14648 22188 14724 22222
rect 14539 22150 14724 22188
rect 14539 22116 14614 22150
rect 14648 22116 14724 22150
rect 14539 22078 14724 22116
rect 14539 22044 14614 22078
rect 14648 22044 14724 22078
rect 14539 22006 14724 22044
rect 14539 21972 14614 22006
rect 14648 21972 14724 22006
rect 14539 21934 14724 21972
rect 14539 21900 14614 21934
rect 14648 21900 14724 21934
rect 14539 21862 14724 21900
rect 14539 21828 14614 21862
rect 14648 21828 14724 21862
rect 14539 21790 14724 21828
rect 14539 21756 14614 21790
rect 14648 21756 14724 21790
rect 14539 21718 14724 21756
rect 14539 21684 14614 21718
rect 14648 21684 14724 21718
rect 14539 21646 14724 21684
rect 14539 21612 14614 21646
rect 14648 21612 14724 21646
rect 14539 21574 14724 21612
rect 14539 21540 14614 21574
rect 14648 21540 14724 21574
rect 14539 21502 14724 21540
rect 14539 21468 14614 21502
rect 14648 21468 14724 21502
rect 14539 21430 14724 21468
rect 14539 21396 14614 21430
rect 14648 21396 14724 21430
rect 14539 21358 14724 21396
rect 14539 21324 14614 21358
rect 14648 21324 14724 21358
rect 14539 21286 14724 21324
rect 14539 21252 14614 21286
rect 14648 21252 14724 21286
rect 14539 21214 14724 21252
rect 14539 21180 14614 21214
rect 14648 21180 14724 21214
rect 14539 21142 14724 21180
rect 14539 21108 14614 21142
rect 14648 21108 14724 21142
rect 14539 21070 14724 21108
rect 14539 21036 14614 21070
rect 14648 21036 14724 21070
rect 14539 20998 14724 21036
rect 14539 20964 14614 20998
rect 14648 20964 14724 20998
rect 14539 20926 14724 20964
rect 14539 20892 14614 20926
rect 14648 20892 14724 20926
rect 14539 20854 14724 20892
rect 14539 20820 14614 20854
rect 14648 20820 14724 20854
rect 14539 20782 14724 20820
rect 14539 20748 14614 20782
rect 14648 20748 14724 20782
rect 14539 20710 14724 20748
rect 14539 20676 14614 20710
rect 14648 20676 14724 20710
rect 14539 20638 14724 20676
rect 14539 20604 14614 20638
rect 14648 20604 14724 20638
rect 14539 20566 14724 20604
rect 14539 20532 14614 20566
rect 14648 20532 14724 20566
rect 14539 20494 14724 20532
rect 14539 20460 14614 20494
rect 14648 20460 14724 20494
rect 14539 20422 14724 20460
rect 14539 20388 14614 20422
rect 14648 20388 14724 20422
rect 14539 20350 14724 20388
rect 14539 20316 14614 20350
rect 14648 20316 14724 20350
rect 14539 20278 14724 20316
rect 14539 20244 14614 20278
rect 14648 20244 14724 20278
rect 14539 20206 14724 20244
rect 14539 20172 14614 20206
rect 14648 20172 14724 20206
rect 14539 20134 14724 20172
rect 14539 20100 14614 20134
rect 14648 20100 14724 20134
rect 14539 20062 14724 20100
rect 14539 20028 14614 20062
rect 14648 20028 14724 20062
rect 14539 19990 14724 20028
rect 14539 19956 14614 19990
rect 14648 19956 14724 19990
rect 14539 19918 14724 19956
rect 14539 19884 14614 19918
rect 14648 19884 14724 19918
rect 14539 19846 14724 19884
rect 14539 19812 14614 19846
rect 14648 19812 14724 19846
rect 14539 19774 14724 19812
rect 14539 19740 14614 19774
rect 14648 19740 14724 19774
rect 14539 19702 14724 19740
rect 14539 19668 14614 19702
rect 14648 19668 14724 19702
rect 14539 19630 14724 19668
rect 14539 19596 14614 19630
rect 14648 19596 14724 19630
rect 14539 19558 14724 19596
rect 14539 19524 14614 19558
rect 14648 19524 14724 19558
rect 14539 19486 14724 19524
rect 14539 19452 14614 19486
rect 14648 19452 14724 19486
rect 14539 19414 14724 19452
rect 14539 19380 14614 19414
rect 14648 19380 14724 19414
rect 14539 19342 14724 19380
rect 14539 19308 14614 19342
rect 14648 19308 14724 19342
rect 14539 19270 14724 19308
rect 14539 19236 14614 19270
rect 14648 19236 14724 19270
rect 14539 19198 14724 19236
rect 14539 19164 14614 19198
rect 14648 19164 14724 19198
rect 14539 19126 14724 19164
rect 14539 19092 14614 19126
rect 14648 19092 14724 19126
rect 14539 19054 14724 19092
rect 14539 19020 14614 19054
rect 14648 19020 14724 19054
rect 14539 18982 14724 19020
rect 14539 18948 14614 18982
rect 14648 18948 14724 18982
rect 14539 18910 14724 18948
rect 14539 18876 14614 18910
rect 14648 18876 14724 18910
rect 14539 18838 14724 18876
rect 14539 18804 14614 18838
rect 14648 18804 14724 18838
rect 14539 18766 14724 18804
rect 14539 18732 14614 18766
rect 14648 18732 14724 18766
rect 14539 18694 14724 18732
rect 14539 18660 14614 18694
rect 14648 18660 14724 18694
rect 14539 18622 14724 18660
rect 14539 18588 14614 18622
rect 14648 18588 14724 18622
rect 14539 18550 14724 18588
rect 14539 18516 14614 18550
rect 14648 18516 14724 18550
rect 14539 18478 14724 18516
rect 14539 18444 14614 18478
rect 14648 18444 14724 18478
rect 14539 18406 14724 18444
rect 14539 18372 14614 18406
rect 14648 18372 14724 18406
rect 14539 18334 14724 18372
rect 14539 18300 14614 18334
rect 14648 18300 14724 18334
rect 14539 18262 14724 18300
rect 14539 18228 14614 18262
rect 14648 18228 14724 18262
rect 14539 18190 14724 18228
rect 14539 18156 14614 18190
rect 14648 18156 14724 18190
rect 14539 18118 14724 18156
rect 14539 18084 14614 18118
rect 14648 18084 14724 18118
rect 14539 18046 14724 18084
rect 14539 18012 14614 18046
rect 14648 18012 14724 18046
rect 14539 17974 14724 18012
rect 14539 17940 14614 17974
rect 14648 17940 14724 17974
rect 14539 17902 14724 17940
rect 14539 17868 14614 17902
rect 14648 17868 14724 17902
rect 14539 17830 14724 17868
rect 14539 17796 14614 17830
rect 14648 17796 14724 17830
rect 14539 17758 14724 17796
rect 14539 17724 14614 17758
rect 14648 17724 14724 17758
rect 14539 17686 14724 17724
rect 14539 17652 14614 17686
rect 14648 17652 14724 17686
rect 14539 17614 14724 17652
rect 14539 17580 14614 17614
rect 14648 17580 14724 17614
rect 14539 17542 14724 17580
rect 14539 17508 14614 17542
rect 14648 17508 14724 17542
rect 14539 17470 14724 17508
rect 14539 17436 14614 17470
rect 14648 17436 14724 17470
rect 14539 17398 14724 17436
rect 14539 17364 14614 17398
rect 14648 17364 14724 17398
rect 14539 17326 14724 17364
rect 14539 17292 14614 17326
rect 14648 17292 14724 17326
rect 14539 17254 14724 17292
rect 14539 17220 14614 17254
rect 14648 17220 14724 17254
rect 14539 17182 14724 17220
rect 14539 17148 14614 17182
rect 14648 17148 14724 17182
rect 14539 17110 14724 17148
rect 14539 17076 14614 17110
rect 14648 17076 14724 17110
rect 14539 17038 14724 17076
rect 14539 17004 14614 17038
rect 14648 17004 14724 17038
rect 14539 16966 14724 17004
rect 14539 16932 14614 16966
rect 14648 16932 14724 16966
rect 14539 16894 14724 16932
rect 14539 16860 14614 16894
rect 14648 16860 14724 16894
rect 14539 16822 14724 16860
rect 14539 16788 14614 16822
rect 14648 16788 14724 16822
rect 14539 16750 14724 16788
rect 14539 16716 14614 16750
rect 14648 16716 14724 16750
rect 14539 16678 14724 16716
rect 14539 16644 14614 16678
rect 14648 16644 14724 16678
rect 14539 16606 14724 16644
rect 14539 16572 14614 16606
rect 14648 16572 14724 16606
rect 14539 16534 14724 16572
rect 14539 16500 14614 16534
rect 14648 16500 14724 16534
rect 14539 16462 14724 16500
rect 14539 16428 14614 16462
rect 14648 16428 14724 16462
rect 14539 16390 14724 16428
rect 14539 16356 14614 16390
rect 14648 16356 14724 16390
rect 14539 16318 14724 16356
rect 14539 16284 14614 16318
rect 14648 16284 14724 16318
rect 14539 16246 14724 16284
rect 14539 16212 14614 16246
rect 14648 16212 14724 16246
rect 14539 16174 14724 16212
rect 14539 16140 14614 16174
rect 14648 16140 14724 16174
rect 14539 16102 14724 16140
rect 14539 16068 14614 16102
rect 14648 16068 14724 16102
rect 14539 16030 14724 16068
rect 14539 15996 14614 16030
rect 14648 15996 14724 16030
rect 14539 15958 14724 15996
rect 14539 15924 14614 15958
rect 14648 15924 14724 15958
rect 14539 15886 14724 15924
rect 14539 15852 14614 15886
rect 14648 15852 14724 15886
rect 14539 15814 14724 15852
rect 14539 15780 14614 15814
rect 14648 15780 14724 15814
rect 14539 15742 14724 15780
rect 14539 15708 14614 15742
rect 14648 15708 14724 15742
rect 14539 15670 14724 15708
rect 14539 15636 14614 15670
rect 14648 15636 14724 15670
rect 14539 15598 14724 15636
rect 14539 15564 14614 15598
rect 14648 15564 14724 15598
rect 14539 15526 14724 15564
rect 14539 15492 14614 15526
rect 14648 15492 14724 15526
rect 14539 15454 14724 15492
rect 14539 15420 14614 15454
rect 14648 15420 14724 15454
rect 14539 15382 14724 15420
rect 14539 15348 14614 15382
rect 14648 15348 14724 15382
rect 14539 15310 14724 15348
rect 14539 15276 14614 15310
rect 14648 15276 14724 15310
rect 14539 15238 14724 15276
rect 14539 15204 14614 15238
rect 14648 15204 14724 15238
rect 14539 15166 14724 15204
rect 14539 15132 14614 15166
rect 14648 15132 14724 15166
rect 14539 15094 14724 15132
rect 14539 15060 14614 15094
rect 14648 15060 14724 15094
rect 14539 15022 14724 15060
rect 14539 14988 14614 15022
rect 14648 14988 14724 15022
rect 14539 14950 14724 14988
rect 14539 14916 14614 14950
rect 14648 14916 14724 14950
rect 14539 14878 14724 14916
rect 14539 14844 14614 14878
rect 14648 14844 14724 14878
rect 14539 14806 14724 14844
rect 14539 14772 14614 14806
rect 14648 14772 14724 14806
rect 14539 14734 14724 14772
rect 14539 14700 14614 14734
rect 14648 14700 14724 14734
rect 14539 14662 14724 14700
rect 14539 14628 14614 14662
rect 14648 14628 14724 14662
rect 14539 14590 14724 14628
rect 14539 14556 14614 14590
rect 14648 14556 14724 14590
rect 14539 14518 14724 14556
rect 14539 14484 14614 14518
rect 14648 14484 14724 14518
rect 14539 14446 14724 14484
rect 14539 14412 14614 14446
rect 14648 14412 14724 14446
rect 14539 14374 14724 14412
rect 14539 14340 14614 14374
rect 14648 14340 14724 14374
rect 14539 14302 14724 14340
rect 14539 14268 14614 14302
rect 14648 14268 14724 14302
rect 14539 14230 14724 14268
rect 14539 14196 14614 14230
rect 14648 14196 14724 14230
rect 14539 14158 14724 14196
rect 14539 14124 14614 14158
rect 14648 14124 14724 14158
rect 14539 14086 14724 14124
rect 14539 14052 14614 14086
rect 14648 14052 14724 14086
rect 14539 14014 14724 14052
rect 14539 13980 14614 14014
rect 14648 13980 14724 14014
rect 14539 13942 14724 13980
rect 14539 13908 14614 13942
rect 14648 13908 14724 13942
rect 14539 13870 14724 13908
rect 14539 13836 14614 13870
rect 14648 13836 14724 13870
rect 14539 13798 14724 13836
rect 14539 13764 14614 13798
rect 14648 13764 14724 13798
rect 14539 13726 14724 13764
rect 14539 13692 14614 13726
rect 14648 13692 14724 13726
rect 14539 13654 14724 13692
rect 14539 13620 14614 13654
rect 14648 13620 14724 13654
rect 14539 13582 14724 13620
rect 14539 13548 14614 13582
rect 14648 13548 14724 13582
rect 14539 13510 14724 13548
rect 14539 13476 14614 13510
rect 14648 13476 14724 13510
rect 14539 13438 14724 13476
rect 14539 13404 14614 13438
rect 14648 13404 14724 13438
rect 14539 13366 14724 13404
rect 14539 13332 14614 13366
rect 14648 13332 14724 13366
rect 14539 13294 14724 13332
rect 14539 13260 14614 13294
rect 14648 13260 14724 13294
rect 14539 13222 14724 13260
rect 14539 13188 14614 13222
rect 14648 13188 14724 13222
rect 14539 13150 14724 13188
rect 14539 13116 14614 13150
rect 14648 13116 14724 13150
rect 14539 13078 14724 13116
rect 14539 13044 14614 13078
rect 14648 13044 14724 13078
rect 14539 13006 14724 13044
rect 14539 12972 14614 13006
rect 14648 12972 14724 13006
rect 14539 12934 14724 12972
rect 14539 12900 14614 12934
rect 14648 12900 14724 12934
rect 14539 12862 14724 12900
rect 14539 12828 14614 12862
rect 14648 12828 14724 12862
rect 14539 12790 14724 12828
rect 14539 12756 14614 12790
rect 14648 12756 14724 12790
rect 14539 12718 14724 12756
rect 14539 12684 14614 12718
rect 14648 12684 14724 12718
rect 14539 12646 14724 12684
rect 14539 12612 14614 12646
rect 14648 12612 14724 12646
rect 14539 12574 14724 12612
rect 14539 12540 14614 12574
rect 14648 12540 14724 12574
rect 14539 12502 14724 12540
rect 14539 12468 14614 12502
rect 14648 12468 14724 12502
rect 14539 12430 14724 12468
rect 14539 12396 14614 12430
rect 14648 12396 14724 12430
rect 14539 12358 14724 12396
rect 14539 12324 14614 12358
rect 14648 12324 14724 12358
rect 14539 12286 14724 12324
rect 14539 12252 14614 12286
rect 14648 12252 14724 12286
rect 14539 12214 14724 12252
rect 14539 12180 14614 12214
rect 14648 12180 14724 12214
rect 14539 12142 14724 12180
rect 14539 12108 14614 12142
rect 14648 12108 14724 12142
rect 14539 12070 14724 12108
rect 14539 12036 14614 12070
rect 14648 12036 14724 12070
rect 14539 11998 14724 12036
rect 14539 11964 14614 11998
rect 14648 11964 14724 11998
rect 14539 11926 14724 11964
rect 14539 11892 14614 11926
rect 14648 11892 14724 11926
rect 14539 11854 14724 11892
rect 14539 11820 14614 11854
rect 14648 11820 14724 11854
rect 14539 11782 14724 11820
rect 14539 11748 14614 11782
rect 14648 11748 14724 11782
rect 14539 11710 14724 11748
rect 14539 11676 14614 11710
rect 14648 11676 14724 11710
rect 14539 11638 14724 11676
rect 14539 11604 14614 11638
rect 14648 11604 14724 11638
rect 14539 11566 14724 11604
rect 14539 11532 14614 11566
rect 14648 11532 14724 11566
rect 14539 11494 14724 11532
rect 14539 11460 14614 11494
rect 14648 11460 14724 11494
rect 14539 11422 14724 11460
rect 14539 11388 14614 11422
rect 14648 11388 14724 11422
rect 14539 11350 14724 11388
rect 14539 11316 14614 11350
rect 14648 11316 14724 11350
rect 14539 11278 14724 11316
rect 14539 11244 14614 11278
rect 14648 11244 14724 11278
rect 14539 11206 14724 11244
rect 14539 11172 14614 11206
rect 14648 11172 14724 11206
rect 14539 11134 14724 11172
rect 14539 11100 14614 11134
rect 14648 11100 14724 11134
rect 14539 11062 14724 11100
rect 14539 11028 14614 11062
rect 14648 11028 14724 11062
rect 14539 10990 14724 11028
rect 14539 10956 14614 10990
rect 14648 10956 14724 10990
rect 14539 10918 14724 10956
rect 14539 10884 14614 10918
rect 14648 10884 14724 10918
rect 14539 10846 14724 10884
rect 14539 10812 14614 10846
rect 14648 10812 14724 10846
rect 14539 10774 14724 10812
rect 14539 10740 14614 10774
rect 14648 10740 14724 10774
rect 14539 10702 14724 10740
rect 14539 10668 14614 10702
rect 14648 10668 14724 10702
rect 14539 10630 14724 10668
rect 14539 10596 14614 10630
rect 14648 10596 14724 10630
rect 14539 10558 14724 10596
rect 14539 10524 14614 10558
rect 14648 10524 14724 10558
rect 14539 10486 14724 10524
rect 14539 10452 14614 10486
rect 14648 10452 14724 10486
rect 14539 10414 14724 10452
rect 14539 10380 14614 10414
rect 14648 10380 14724 10414
rect 14539 10342 14724 10380
rect 14539 10308 14614 10342
rect 14648 10308 14724 10342
rect 14539 10270 14724 10308
rect 14539 10236 14614 10270
rect 14648 10236 14724 10270
rect 14539 10198 14724 10236
rect 14539 10164 14614 10198
rect 14648 10164 14724 10198
rect 14539 10126 14724 10164
rect 14539 10092 14614 10126
rect 14648 10092 14724 10126
rect 14539 10054 14724 10092
rect 14539 10020 14614 10054
rect 14648 10020 14724 10054
rect 14539 9982 14724 10020
rect 14539 9948 14614 9982
rect 14648 9948 14724 9982
rect 14539 9910 14724 9948
rect 14029 9908 14152 9910
tri 792 9907 793 9908 ne
rect 793 9907 14152 9908
rect 245 9841 430 9879
tri 793 9876 824 9907 ne
rect 824 9876 14152 9907
tri 14152 9876 14186 9910 nw
rect 14539 9876 14614 9910
rect 14648 9876 14724 9910
tri 824 9843 857 9876 ne
rect 857 9843 14119 9876
tri 14119 9843 14152 9876 nw
rect 245 9807 320 9841
rect 354 9807 430 9841
rect 245 9769 430 9807
rect 245 9735 320 9769
rect 354 9735 430 9769
rect 245 9697 430 9735
rect 245 9663 320 9697
rect 354 9663 430 9697
rect 245 9528 430 9663
rect 858 9775 2096 9843
rect 858 9741 883 9775
rect 917 9741 955 9775
rect 989 9741 1027 9775
rect 1061 9741 1099 9775
rect 1133 9741 1171 9775
rect 1205 9741 1243 9775
rect 1277 9741 1315 9775
rect 1349 9741 1387 9775
rect 1421 9741 1459 9775
rect 1493 9741 1531 9775
rect 1565 9741 1603 9775
rect 1637 9741 1675 9775
rect 1709 9741 1747 9775
rect 1781 9741 1819 9775
rect 1853 9741 1891 9775
rect 1925 9741 1963 9775
rect 1997 9741 2035 9775
rect 2069 9741 2096 9775
rect 858 9731 2096 9741
rect 245 9452 720 9528
rect 245 9418 320 9452
rect 354 9418 610 9452
rect 644 9418 720 9452
rect 245 9343 720 9418
rect 858 9295 908 9731
rect 2048 9295 2096 9731
rect 12858 9774 14096 9843
rect 12858 9740 12883 9774
rect 12917 9740 12955 9774
rect 12989 9740 13027 9774
rect 13061 9740 13099 9774
rect 13133 9740 13171 9774
rect 13205 9740 13243 9774
rect 13277 9740 13315 9774
rect 13349 9740 13387 9774
rect 13421 9740 13459 9774
rect 13493 9740 13531 9774
rect 13565 9740 13603 9774
rect 13637 9740 13675 9774
rect 13709 9740 13747 9774
rect 13781 9740 13819 9774
rect 13853 9740 13891 9774
rect 13925 9740 13963 9774
rect 13997 9740 14035 9774
rect 14069 9740 14096 9774
rect 12858 9731 14096 9740
rect 11273 9528 12512 9529
rect 2248 9484 12705 9528
rect 2248 9483 11322 9484
rect 2248 9452 2445 9483
rect 3585 9452 11322 9483
rect 12462 9452 12705 9484
rect 2248 9418 2311 9452
rect 2345 9418 2383 9452
rect 2417 9418 2445 9452
rect 3585 9418 3607 9452
rect 3641 9418 3679 9452
rect 3713 9418 3751 9452
rect 3785 9418 3823 9452
rect 3857 9418 3895 9452
rect 3929 9418 3967 9452
rect 4001 9418 4039 9452
rect 4073 9418 4111 9452
rect 4145 9418 4183 9452
rect 4217 9418 4255 9452
rect 4289 9418 4327 9452
rect 4361 9418 4399 9452
rect 4433 9418 4471 9452
rect 4505 9418 4543 9452
rect 4577 9418 4615 9452
rect 4649 9418 4687 9452
rect 4721 9418 4759 9452
rect 4793 9418 4831 9452
rect 4865 9418 4903 9452
rect 4937 9418 4975 9452
rect 5009 9418 5047 9452
rect 5081 9418 5119 9452
rect 5153 9418 5191 9452
rect 5225 9418 5263 9452
rect 5297 9418 5335 9452
rect 5369 9418 5407 9452
rect 5441 9418 5479 9452
rect 5513 9418 5551 9452
rect 5585 9418 5623 9452
rect 5657 9418 5695 9452
rect 5729 9418 5767 9452
rect 5801 9418 5839 9452
rect 5873 9418 5911 9452
rect 5945 9418 5983 9452
rect 6017 9418 6055 9452
rect 6089 9418 6127 9452
rect 6161 9418 6199 9452
rect 6233 9418 6271 9452
rect 6305 9418 6343 9452
rect 6377 9418 6415 9452
rect 6449 9418 6487 9452
rect 6521 9418 6559 9452
rect 6593 9418 6631 9452
rect 6665 9418 6703 9452
rect 6737 9418 6775 9452
rect 6809 9418 6847 9452
rect 6881 9418 6919 9452
rect 6953 9418 6991 9452
rect 7025 9418 7063 9452
rect 7097 9418 7135 9452
rect 7169 9418 7207 9452
rect 7241 9418 7279 9452
rect 7313 9418 7351 9452
rect 7385 9418 7423 9452
rect 7457 9418 7495 9452
rect 7529 9418 7567 9452
rect 7601 9418 7639 9452
rect 7673 9418 7711 9452
rect 7745 9418 7783 9452
rect 7817 9418 7855 9452
rect 7889 9418 7927 9452
rect 7961 9418 7999 9452
rect 8033 9418 8071 9452
rect 8105 9418 8143 9452
rect 8177 9418 8215 9452
rect 8249 9418 8287 9452
rect 8321 9418 8359 9452
rect 8393 9418 8431 9452
rect 8465 9418 8503 9452
rect 8537 9418 8575 9452
rect 8609 9418 8647 9452
rect 8681 9418 8719 9452
rect 8753 9418 8791 9452
rect 8825 9418 8863 9452
rect 8897 9418 8935 9452
rect 8969 9418 9007 9452
rect 9041 9418 9079 9452
rect 9113 9418 9151 9452
rect 9185 9418 9223 9452
rect 9257 9418 9295 9452
rect 9329 9418 9367 9452
rect 9401 9418 9439 9452
rect 9473 9418 9511 9452
rect 9545 9418 9583 9452
rect 9617 9418 9655 9452
rect 9689 9418 9727 9452
rect 9761 9418 9799 9452
rect 9833 9418 9871 9452
rect 9905 9418 9943 9452
rect 9977 9418 10015 9452
rect 10049 9418 10087 9452
rect 10121 9418 10159 9452
rect 10193 9418 10231 9452
rect 10265 9418 10303 9452
rect 10337 9418 10375 9452
rect 10409 9418 10447 9452
rect 10481 9418 10519 9452
rect 10553 9418 10591 9452
rect 10625 9418 10663 9452
rect 10697 9418 10735 9452
rect 10769 9418 10807 9452
rect 10841 9418 10879 9452
rect 10913 9418 10951 9452
rect 10985 9418 11023 9452
rect 11057 9418 11095 9452
rect 11129 9418 11167 9452
rect 11201 9418 11239 9452
rect 11273 9418 11311 9452
rect 12462 9418 12463 9452
rect 12497 9418 12535 9452
rect 12569 9418 12607 9452
rect 12641 9418 12705 9452
rect 2248 9343 2445 9418
rect 858 9252 2096 9295
rect 2396 8983 2445 9343
rect 3585 9343 11322 9418
rect 3585 8983 3635 9343
rect 2396 8939 3635 8983
rect 11273 8984 11322 9343
rect 12462 9343 12705 9418
rect 12462 8984 12512 9343
rect 12858 9295 12908 9731
rect 14048 9295 14096 9731
rect 14539 9838 14724 9876
rect 14539 9804 14614 9838
rect 14648 9804 14724 9838
rect 14539 9766 14724 9804
rect 14539 9732 14614 9766
rect 14648 9732 14724 9766
rect 14539 9694 14724 9732
rect 14539 9660 14614 9694
rect 14648 9660 14724 9694
rect 14539 9528 14724 9660
rect 14232 9452 14724 9528
rect 14232 9418 14314 9452
rect 14348 9418 14614 9452
rect 14648 9418 14724 9452
rect 14232 9343 14724 9418
rect 12858 9252 14096 9295
rect 11273 8940 12512 8984
<< via1 >>
rect 4944 31877 7236 32697
rect 7745 31877 10037 32697
rect 4939 30683 7231 30799
rect 7750 30683 10042 30799
rect 2509 30370 4481 30486
rect 10500 30370 12472 30486
rect 4939 30067 7231 30183
rect 7750 30067 10042 30183
rect 2509 29754 4481 29870
rect 10500 29754 12472 29870
rect 4939 29451 7231 29567
rect 7750 29451 10042 29567
rect 2509 29138 4481 29254
rect 10500 29138 12472 29254
rect 4939 28835 7231 28951
rect 7750 28835 10042 28951
rect 2509 28522 4481 28638
rect 10500 28522 12472 28638
rect 4939 28219 7231 28335
rect 7750 28219 10042 28335
rect 2509 27906 4481 28022
rect 10500 27906 12472 28022
rect 4939 27603 7231 27719
rect 7750 27603 10042 27719
rect 4933 26037 7225 26153
rect 7757 26037 10049 26153
rect 2546 25771 4454 25887
rect 10528 25771 12436 25887
rect 4933 25505 7225 25621
rect 7757 25505 10049 25621
rect 2546 25239 4454 25355
rect 10528 25239 12436 25355
rect 4933 24973 7225 25089
rect 7757 24973 10049 25089
rect 2546 24707 4454 24823
rect 10528 24707 12436 24823
rect 4933 24441 7225 24557
rect 7757 24441 10049 24557
rect 2546 24175 4454 24291
rect 10528 24175 12436 24291
rect 4933 23909 7225 24025
rect 7757 23909 10049 24025
rect 2546 23643 4454 23759
rect 10528 23643 12436 23759
rect 4933 23377 7225 23493
rect 7757 23377 10049 23493
rect 4945 21669 7237 22489
rect 7744 21669 10036 22489
rect 908 9295 2048 9731
rect 2445 9452 3585 9483
rect 11322 9452 12462 9484
rect 2445 9418 2455 9452
rect 2455 9418 2489 9452
rect 2489 9418 2527 9452
rect 2527 9418 2561 9452
rect 2561 9418 2599 9452
rect 2599 9418 2633 9452
rect 2633 9418 2671 9452
rect 2671 9418 2705 9452
rect 2705 9418 2743 9452
rect 2743 9418 2777 9452
rect 2777 9418 2815 9452
rect 2815 9418 2849 9452
rect 2849 9418 2887 9452
rect 2887 9418 2921 9452
rect 2921 9418 2959 9452
rect 2959 9418 2993 9452
rect 2993 9418 3031 9452
rect 3031 9418 3065 9452
rect 3065 9418 3103 9452
rect 3103 9418 3137 9452
rect 3137 9418 3175 9452
rect 3175 9418 3209 9452
rect 3209 9418 3247 9452
rect 3247 9418 3281 9452
rect 3281 9418 3319 9452
rect 3319 9418 3353 9452
rect 3353 9418 3391 9452
rect 3391 9418 3425 9452
rect 3425 9418 3463 9452
rect 3463 9418 3497 9452
rect 3497 9418 3535 9452
rect 3535 9418 3569 9452
rect 3569 9418 3585 9452
rect 11322 9418 11345 9452
rect 11345 9418 11383 9452
rect 11383 9418 11417 9452
rect 11417 9418 11455 9452
rect 11455 9418 11489 9452
rect 11489 9418 11527 9452
rect 11527 9418 11561 9452
rect 11561 9418 11599 9452
rect 11599 9418 11633 9452
rect 11633 9418 11671 9452
rect 11671 9418 11705 9452
rect 11705 9418 11743 9452
rect 11743 9418 11777 9452
rect 11777 9418 11815 9452
rect 11815 9418 11849 9452
rect 11849 9418 11887 9452
rect 11887 9418 11921 9452
rect 11921 9418 11959 9452
rect 11959 9418 11993 9452
rect 11993 9418 12031 9452
rect 12031 9418 12065 9452
rect 12065 9418 12103 9452
rect 12103 9418 12137 9452
rect 12137 9418 12175 9452
rect 12175 9418 12209 9452
rect 12209 9418 12247 9452
rect 12247 9418 12281 9452
rect 12281 9418 12319 9452
rect 12319 9418 12353 9452
rect 12353 9418 12391 9452
rect 12391 9418 12425 9452
rect 12425 9418 12462 9452
rect 2445 8983 3585 9418
rect 11322 8984 12462 9418
rect 12908 9295 14048 9731
<< metal2 >>
tri 4891 39322 4991 39422 se
rect 4991 39322 7191 39422
tri 7191 39322 7291 39422 sw
rect 4891 39213 7291 39322
rect 4891 35317 4979 39213
rect 7195 35317 7291 39213
rect 4891 32697 7291 35317
rect 4891 31877 4944 32697
rect 7236 31877 7291 32697
tri 301 31445 501 31645 se
rect 501 31445 4291 31645
tri 4291 31445 4491 31645 sw
rect 301 31344 4491 31445
rect 301 23288 466 31344
rect 2442 30486 4491 31344
rect 2442 30370 2509 30486
rect 4481 30370 4491 30486
rect 2442 29870 4491 30370
rect 2442 29754 2509 29870
rect 4481 29754 4491 29870
rect 2442 29254 4491 29754
rect 2442 29138 2509 29254
rect 4481 29138 4491 29254
rect 2442 28638 4491 29138
rect 2442 28522 2509 28638
rect 4481 28522 4491 28638
rect 2442 28022 4491 28522
rect 2442 27906 2509 28022
rect 4481 27906 4491 28022
rect 2442 25887 4491 27906
rect 4891 30799 7291 31877
rect 4891 30683 4939 30799
rect 7231 30683 7291 30799
rect 4891 30183 7291 30683
rect 4891 30067 4939 30183
rect 7231 30067 7291 30183
rect 4891 29567 7291 30067
rect 4891 29451 4939 29567
rect 7231 29451 7291 29567
rect 4891 28951 7291 29451
rect 4891 28835 4939 28951
rect 7231 28835 7291 28951
rect 4891 28335 7291 28835
rect 4891 28219 4939 28335
rect 7231 28219 7291 28335
rect 4891 27719 7291 28219
rect 4891 27603 4939 27719
rect 7231 27603 7291 27719
rect 4891 27317 7291 27603
tri 4891 27117 5091 27317 ne
rect 5091 27117 7091 27317
tri 7091 27117 7291 27317 nw
tri 7691 39322 7791 39422 se
rect 7791 39322 9991 39422
tri 9991 39322 10091 39422 sw
rect 7691 39213 10091 39322
rect 7691 35317 7779 39213
rect 9995 35317 10091 39213
rect 7691 32697 10091 35317
rect 7691 31877 7745 32697
rect 10037 31877 10091 32697
rect 7691 30799 10091 31877
rect 7691 30683 7750 30799
rect 10042 30683 10091 30799
rect 7691 30183 10091 30683
rect 7691 30067 7750 30183
rect 10042 30067 10091 30183
rect 7691 29567 10091 30067
rect 7691 29451 7750 29567
rect 10042 29451 10091 29567
rect 7691 28951 10091 29451
rect 7691 28835 7750 28951
rect 10042 28835 10091 28951
rect 7691 28335 10091 28835
rect 7691 28219 7750 28335
rect 10042 28219 10091 28335
rect 7691 27719 10091 28219
rect 7691 27603 7750 27719
rect 10042 27603 10091 27719
rect 7691 27317 10091 27603
tri 7691 27117 7891 27317 ne
rect 7891 27117 9891 27317
tri 9891 27117 10091 27317 nw
tri 10491 31445 10691 31645 se
rect 10691 31445 14431 31645
tri 14431 31445 14631 31645 sw
rect 10491 31392 14631 31445
rect 10491 30486 12455 31392
rect 10491 30370 10500 30486
rect 10491 29870 12455 30370
rect 10491 29754 10500 29870
rect 10491 29254 12455 29754
rect 10491 29138 10500 29254
rect 10491 28638 12455 29138
rect 10491 28522 10500 28638
rect 10491 28022 12455 28522
rect 10491 27906 10500 28022
rect 2442 25771 2546 25887
rect 4454 25771 4491 25887
rect 2442 25355 4491 25771
rect 2442 25239 2546 25355
rect 4454 25239 4491 25355
rect 2442 24823 4491 25239
rect 2442 24707 2546 24823
rect 4454 24707 4491 24823
rect 2442 24291 4491 24707
rect 2442 24175 2546 24291
rect 4454 24175 4491 24291
rect 2442 23759 4491 24175
rect 2442 23643 2546 23759
rect 4454 23643 4491 23759
rect 2442 23288 4491 23643
rect 301 23016 4491 23288
tri 301 22816 501 23016 ne
rect 501 22816 4291 23016
tri 4291 22816 4491 23016 nw
tri 4891 26278 5091 26478 se
rect 5091 26278 7091 26478
tri 7091 26278 7291 26478 sw
rect 4891 26153 7291 26278
rect 4891 26037 4933 26153
rect 7225 26037 7291 26153
rect 4891 25621 7291 26037
rect 4891 25505 4933 25621
rect 7225 25505 7291 25621
rect 4891 25089 7291 25505
rect 4891 24973 4933 25089
rect 7225 24973 7291 25089
rect 4891 24557 7291 24973
rect 4891 24441 4933 24557
rect 7225 24441 7291 24557
rect 4891 24025 7291 24441
rect 4891 23909 4933 24025
rect 7225 23909 7291 24025
rect 4891 23493 7291 23909
rect 4891 23377 4933 23493
rect 7225 23377 7291 23493
rect 4891 22489 7291 23377
rect 4891 21669 4945 22489
rect 7237 21669 7291 22489
rect 4891 18931 7291 21669
rect 4891 17275 4942 18931
rect 7238 17275 7291 18931
rect 4891 17214 7291 17275
rect 4891 17086 5103 17214
tri 4891 16986 4991 17086 ne
rect 4991 17078 5103 17086
rect 7239 17078 7291 17214
rect 4991 17056 7291 17078
rect 4991 16986 7221 17056
tri 7221 16986 7291 17056 nw
tri 7691 26278 7891 26478 se
rect 7891 26278 9891 26478
tri 9891 26278 10091 26478 sw
rect 7691 26153 10091 26278
rect 7691 26037 7757 26153
rect 10049 26037 10091 26153
rect 7691 25621 10091 26037
rect 7691 25505 7757 25621
rect 10049 25505 10091 25621
rect 7691 25089 10091 25505
rect 7691 24973 7757 25089
rect 10049 24973 10091 25089
rect 7691 24557 10091 24973
rect 7691 24441 7757 24557
rect 10049 24441 10091 24557
rect 7691 24025 10091 24441
rect 7691 23909 7757 24025
rect 10049 23909 10091 24025
rect 7691 23493 10091 23909
rect 7691 23377 7757 23493
rect 10049 23377 10091 23493
rect 7691 22489 10091 23377
rect 10491 25887 12455 27906
rect 10491 25771 10528 25887
rect 12436 25771 12455 25887
rect 10491 25355 12455 25771
rect 10491 25239 10528 25355
rect 12436 25239 12455 25355
rect 10491 24823 12455 25239
rect 10491 24707 10528 24823
rect 12436 24707 12455 24823
rect 10491 24291 12455 24707
rect 10491 24175 10528 24291
rect 12436 24175 12455 24291
rect 10491 23759 12455 24175
rect 10491 23643 10528 23759
rect 12436 23643 12455 23759
rect 10491 23336 12455 23643
rect 14431 23336 14631 31392
rect 10491 23016 14631 23336
tri 10491 22816 10691 23016 ne
rect 10691 22816 14431 23016
tri 14431 22816 14631 23016 nw
rect 7691 21669 7744 22489
rect 10036 21669 10091 22489
rect 7691 18931 10091 21669
rect 7691 17275 7742 18931
rect 10038 17275 10091 18931
rect 7691 17214 10091 17275
rect 7691 17078 7739 17214
rect 9875 17086 10091 17214
rect 9875 17078 9991 17086
rect 7691 17056 9991 17078
tri 7691 16986 7761 17056 ne
rect 7761 16986 9991 17056
tri 9991 16986 10091 17086 nw
rect 858 9741 2096 9772
rect 858 9285 890 9741
rect 2066 9285 2096 9741
rect 12858 9741 14096 9772
rect 858 9252 2096 9285
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 8939 3635 8965
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 12858 9285 12890 9741
rect 14066 9285 14096 9741
rect 12858 9252 14096 9285
rect 11273 8940 12512 8966
<< via2 >>
rect 4979 35317 7195 39213
rect 466 23288 2442 31344
rect 7779 35317 9995 39213
rect 12455 30486 14431 31392
rect 12455 30370 12472 30486
rect 12472 30370 14431 30486
rect 12455 29870 14431 30370
rect 12455 29754 12472 29870
rect 12472 29754 14431 29870
rect 12455 29254 14431 29754
rect 12455 29138 12472 29254
rect 12472 29138 14431 29254
rect 12455 28638 14431 29138
rect 12455 28522 12472 28638
rect 12472 28522 14431 28638
rect 12455 28022 14431 28522
rect 12455 27906 12472 28022
rect 12472 27906 14431 28022
rect 4942 17275 7238 18931
rect 5103 17078 7239 17214
rect 12455 23336 14431 27906
rect 7742 17275 10038 18931
rect 7739 17078 9875 17214
rect 890 9731 2066 9741
rect 890 9295 908 9731
rect 908 9295 2048 9731
rect 2048 9295 2066 9731
rect 890 9285 2066 9295
rect 2427 9483 3603 9501
rect 2427 8983 2445 9483
rect 2445 8983 3585 9483
rect 3585 8983 3603 9483
rect 2427 8965 3603 8983
rect 11304 9484 12480 9502
rect 11304 8984 11322 9484
rect 11322 8984 12462 9484
rect 12462 8984 12480 9484
rect 11304 8966 12480 8984
rect 12890 9731 14066 9741
rect 12890 9295 12908 9731
rect 12908 9295 14048 9731
rect 14048 9295 14066 9731
rect 12890 9285 14066 9295
<< metal3 >>
tri 4805 39522 5205 39922 se
rect 5205 39522 9786 39922
tri 9786 39522 10186 39922 sw
rect 4805 39217 10186 39522
rect 4805 35313 4975 39217
rect 7199 35313 7775 39217
rect 9999 35313 10186 39217
rect 4805 35266 10186 35313
tri 4805 35166 4905 35266 ne
rect 4905 35166 10086 35266
tri 10086 35166 10186 35266 nw
tri 99 33575 1155 34631 se
rect 1155 34618 13835 34631
rect 1155 34554 2276 34618
rect 2340 34554 2359 34618
rect 2423 34554 2443 34618
rect 2507 34554 2527 34618
rect 2591 34554 2611 34618
rect 2675 34554 12341 34618
rect 12405 34554 12425 34618
rect 12489 34554 12509 34618
rect 12573 34554 12593 34618
rect 12657 34554 12677 34618
rect 12741 34554 13835 34618
rect 1155 34524 13835 34554
rect 1155 34460 2276 34524
rect 2340 34460 2359 34524
rect 2423 34460 2443 34524
rect 2507 34460 2527 34524
rect 2591 34460 2611 34524
rect 2675 34460 12341 34524
rect 12405 34460 12425 34524
rect 12489 34460 12509 34524
rect 12573 34460 12593 34524
rect 12657 34460 12677 34524
rect 12741 34460 13835 34524
rect 1155 34441 13835 34460
rect 1155 34377 2148 34441
rect 2212 34430 12804 34441
rect 2212 34377 2276 34430
rect 1155 34366 2276 34377
rect 2340 34366 2359 34430
rect 2423 34366 2443 34430
rect 2507 34366 2527 34430
rect 2591 34366 2611 34430
rect 2675 34366 12341 34430
rect 12405 34366 12425 34430
rect 12489 34366 12509 34430
rect 12573 34366 12593 34430
rect 12657 34366 12677 34430
rect 12741 34377 12804 34430
rect 12868 34377 13835 34441
rect 12741 34366 13835 34377
rect 1155 34336 13835 34366
rect 1155 34316 2276 34336
rect 1155 34252 2004 34316
rect 2068 34252 2084 34316
rect 2148 34252 2164 34316
rect 2228 34272 2276 34316
rect 2340 34272 2359 34336
rect 2423 34272 2443 34336
rect 2507 34272 2527 34336
rect 2591 34272 2611 34336
rect 2675 34272 12341 34336
rect 12405 34272 12425 34336
rect 12489 34272 12509 34336
rect 12573 34272 12593 34336
rect 12657 34272 12677 34336
rect 12741 34316 13835 34336
rect 12741 34272 12788 34316
rect 2228 34252 12788 34272
rect 12852 34252 12868 34316
rect 12932 34252 12948 34316
rect 13012 34252 13835 34316
rect 1155 34242 13835 34252
rect 1155 34220 2276 34242
rect 1155 34183 2004 34220
rect 1155 34119 1890 34183
rect 1954 34156 2004 34183
rect 2068 34156 2084 34220
rect 2148 34156 2164 34220
rect 2228 34178 2276 34220
rect 2340 34178 2359 34242
rect 2423 34178 2443 34242
rect 2507 34178 2527 34242
rect 2591 34178 2611 34242
rect 2675 34178 12341 34242
rect 12405 34178 12425 34242
rect 12489 34178 12509 34242
rect 12573 34178 12593 34242
rect 12657 34178 12677 34242
rect 12741 34220 13835 34242
rect 12741 34178 12788 34220
rect 2228 34156 12788 34178
rect 12852 34156 12868 34220
rect 12932 34156 12948 34220
rect 13012 34183 13835 34220
rect 13012 34156 13062 34183
rect 1954 34148 13062 34156
rect 1954 34119 2276 34148
rect 1155 34084 2276 34119
rect 2340 34084 2359 34148
rect 2423 34084 2443 34148
rect 2507 34084 2527 34148
rect 2591 34084 2611 34148
rect 2675 34084 12341 34148
rect 12405 34084 12425 34148
rect 12489 34084 12509 34148
rect 12573 34084 12593 34148
rect 12657 34084 12677 34148
rect 12741 34119 13062 34148
rect 13126 34119 13835 34183
rect 12741 34084 13835 34119
rect 1155 34078 13835 34084
rect 1155 34014 1748 34078
rect 1812 34014 1837 34078
rect 1901 34014 1927 34078
rect 1991 34014 2017 34078
rect 2081 34014 2107 34078
rect 2171 34014 12845 34078
rect 12909 34014 12935 34078
rect 12999 34014 13025 34078
rect 13089 34014 13115 34078
rect 13179 34014 13204 34078
rect 13268 34014 13835 34078
rect 1155 34009 13835 34014
rect 1155 33962 2247 34009
rect 1155 33898 1748 33962
rect 1812 33898 1837 33962
rect 1901 33898 1927 33962
rect 1991 33898 2017 33962
rect 2081 33898 2107 33962
rect 2171 33945 2247 33962
rect 2311 33945 12705 34009
rect 12769 33962 13835 34009
rect 12769 33945 12845 33962
rect 2171 33898 12845 33945
rect 12909 33898 12935 33962
rect 12999 33898 13025 33962
rect 13089 33898 13115 33962
rect 13179 33898 13204 33962
rect 13268 33898 13835 33962
rect 1155 33886 13835 33898
rect 1155 33822 1644 33886
rect 1708 33848 13308 33886
rect 1708 33846 2700 33848
rect 1708 33822 1748 33846
rect 1155 33782 1748 33822
rect 1812 33782 1837 33846
rect 1901 33782 1927 33846
rect 1991 33782 2017 33846
rect 2081 33782 2107 33846
rect 2171 33782 2700 33846
rect 1155 33754 2700 33782
rect 1155 33690 1424 33754
rect 1488 33690 1513 33754
rect 1577 33690 1603 33754
rect 1667 33690 1693 33754
rect 1757 33690 1783 33754
rect 1847 33721 2700 33754
rect 1847 33690 1929 33721
rect 1155 33657 1929 33690
rect 1993 33657 2700 33721
rect 1155 33638 2700 33657
rect 1155 33575 1424 33638
rect 99 33574 1424 33575
rect 1488 33574 1513 33638
rect 1577 33574 1603 33638
rect 1667 33574 1693 33638
rect 1757 33574 1783 33638
rect 1847 33574 2700 33638
rect 99 33558 2700 33574
rect 99 33494 1316 33558
rect 1380 33522 2700 33558
rect 1380 33494 1424 33522
rect 99 33458 1424 33494
rect 1488 33458 1513 33522
rect 1577 33458 1603 33522
rect 1667 33458 1693 33522
rect 1757 33458 1783 33522
rect 1847 33458 2700 33522
rect 99 33434 2700 33458
tri 2700 33448 3100 33848 nw
tri 11900 33448 12300 33848 ne
rect 12300 33846 13308 33848
rect 12300 33782 12845 33846
rect 12909 33782 12935 33846
rect 12999 33782 13025 33846
rect 13089 33782 13115 33846
rect 13179 33782 13204 33846
rect 13268 33822 13308 33846
rect 13372 33822 13835 33886
rect 13268 33782 13835 33822
rect 12300 33754 13835 33782
rect 12300 33721 13169 33754
rect 12300 33657 13023 33721
rect 13087 33690 13169 33721
rect 13233 33690 13259 33754
rect 13323 33690 13349 33754
rect 13413 33690 13439 33754
rect 13503 33690 13528 33754
rect 13592 33690 13835 33754
rect 13087 33657 13835 33690
rect 12300 33638 13835 33657
rect 12300 33574 13169 33638
rect 13233 33574 13259 33638
rect 13323 33574 13349 33638
rect 13413 33574 13439 33638
rect 13503 33574 13528 33638
rect 13592 33608 13835 33638
tri 13835 33608 14858 34631 sw
rect 13592 33574 14858 33608
rect 12300 33558 14858 33574
rect 12300 33522 13636 33558
rect 12300 33458 13169 33522
rect 13233 33458 13259 33522
rect 13323 33458 13349 33522
rect 13413 33458 13439 33522
rect 13503 33458 13528 33522
rect 13592 33494 13636 33522
rect 13700 33494 14858 33558
rect 13592 33458 14858 33494
rect 99 33370 1104 33434
rect 1168 33370 1193 33434
rect 1257 33370 1283 33434
rect 1347 33370 1373 33434
rect 1437 33370 1463 33434
rect 1527 33396 2700 33434
rect 1527 33370 1604 33396
rect 99 33332 1604 33370
rect 1668 33332 2700 33396
rect 99 33318 2700 33332
rect 99 33254 1104 33318
rect 1168 33254 1193 33318
rect 1257 33254 1283 33318
rect 1347 33254 1373 33318
rect 1437 33254 1463 33318
rect 1527 33254 2700 33318
rect 99 33202 2700 33254
rect 99 33138 1104 33202
rect 1168 33138 1193 33202
rect 1257 33138 1283 33202
rect 1347 33138 1373 33202
rect 1437 33138 1463 33202
rect 1527 33138 2700 33202
rect 99 33109 2700 33138
rect 99 33045 982 33109
rect 1046 33045 1072 33109
rect 1136 33045 1162 33109
rect 1226 33045 1252 33109
rect 1316 33045 1342 33109
rect 1406 33045 1432 33109
rect 1496 33045 2700 33109
rect 99 33029 2700 33045
rect 99 32965 982 33029
rect 1046 32965 1072 33029
rect 1136 32965 1162 33029
rect 1226 32965 1252 33029
rect 1316 32965 1342 33029
rect 1406 32965 1432 33029
rect 1496 32965 2700 33029
rect 99 32949 2700 32965
rect 99 32885 982 32949
rect 1046 32885 1072 32949
rect 1136 32885 1162 32949
rect 1226 32885 1252 32949
rect 1316 32885 1342 32949
rect 1406 32885 1432 32949
rect 1496 32885 2700 32949
rect 99 32869 2700 32885
rect 99 32805 982 32869
rect 1046 32805 1072 32869
rect 1136 32805 1162 32869
rect 1226 32805 1252 32869
rect 1316 32805 1342 32869
rect 1406 32805 1432 32869
rect 1496 32805 2700 32869
rect 99 32789 2700 32805
rect 99 32725 982 32789
rect 1046 32725 1072 32789
rect 1136 32725 1162 32789
rect 1226 32725 1252 32789
rect 1316 32725 1342 32789
rect 1406 32725 1432 32789
rect 1496 32725 2700 32789
rect 99 32709 2700 32725
rect 99 32645 982 32709
rect 1046 32645 1072 32709
rect 1136 32645 1162 32709
rect 1226 32645 1252 32709
rect 1316 32645 1342 32709
rect 1406 32645 1432 32709
rect 1496 32645 2700 32709
rect 99 32629 2700 32645
rect 99 32565 982 32629
rect 1046 32565 1072 32629
rect 1136 32565 1162 32629
rect 1226 32565 1252 32629
rect 1316 32565 1342 32629
rect 1406 32565 1432 32629
rect 1496 32565 2700 32629
rect 99 32549 2700 32565
rect 99 32485 982 32549
rect 1046 32485 1072 32549
rect 1136 32485 1162 32549
rect 1226 32485 1252 32549
rect 1316 32485 1342 32549
rect 1406 32485 1432 32549
rect 1496 32485 2700 32549
rect 99 32469 2700 32485
rect 99 32405 982 32469
rect 1046 32405 1072 32469
rect 1136 32405 1162 32469
rect 1226 32405 1252 32469
rect 1316 32405 1342 32469
rect 1406 32405 1432 32469
rect 1496 32405 2700 32469
rect 99 32389 2700 32405
rect 99 32325 982 32389
rect 1046 32325 1072 32389
rect 1136 32325 1162 32389
rect 1226 32325 1252 32389
rect 1316 32325 1342 32389
rect 1406 32325 1432 32389
rect 1496 32325 2700 32389
rect 99 32309 2700 32325
rect 99 32245 982 32309
rect 1046 32245 1072 32309
rect 1136 32245 1162 32309
rect 1226 32245 1252 32309
rect 1316 32245 1342 32309
rect 1406 32245 1432 32309
rect 1496 32245 2700 32309
rect 99 32229 2700 32245
rect 99 32165 982 32229
rect 1046 32165 1072 32229
rect 1136 32165 1162 32229
rect 1226 32165 1252 32229
rect 1316 32165 1342 32229
rect 1406 32165 1432 32229
rect 1496 32165 2700 32229
rect 99 32149 2700 32165
rect 99 32085 982 32149
rect 1046 32085 1072 32149
rect 1136 32085 1162 32149
rect 1226 32085 1252 32149
rect 1316 32085 1342 32149
rect 1406 32085 1432 32149
rect 1496 32085 2700 32149
rect 99 32069 2700 32085
rect 99 32005 982 32069
rect 1046 32005 1072 32069
rect 1136 32005 1162 32069
rect 1226 32005 1252 32069
rect 1316 32005 1342 32069
rect 1406 32005 1432 32069
rect 1496 32005 2700 32069
rect 99 31989 2700 32005
rect 99 31925 982 31989
rect 1046 31925 1072 31989
rect 1136 31925 1162 31989
rect 1226 31925 1252 31989
rect 1316 31925 1342 31989
rect 1406 31925 1432 31989
rect 1496 31925 2700 31989
rect 99 31909 2700 31925
rect 99 31845 982 31909
rect 1046 31845 1072 31909
rect 1136 31845 1162 31909
rect 1226 31845 1252 31909
rect 1316 31845 1342 31909
rect 1406 31845 1432 31909
rect 1496 31845 2700 31909
rect 99 31829 2700 31845
rect 99 31765 982 31829
rect 1046 31765 1072 31829
rect 1136 31765 1162 31829
rect 1226 31765 1252 31829
rect 1316 31765 1342 31829
rect 1406 31765 1432 31829
rect 1496 31765 2700 31829
rect 99 31749 2700 31765
rect 99 31685 982 31749
rect 1046 31685 1072 31749
rect 1136 31685 1162 31749
rect 1226 31685 1252 31749
rect 1316 31685 1342 31749
rect 1406 31685 1432 31749
rect 1496 31685 2700 31749
rect 99 31669 2700 31685
rect 99 31605 982 31669
rect 1046 31605 1072 31669
rect 1136 31605 1162 31669
rect 1226 31605 1252 31669
rect 1316 31605 1342 31669
rect 1406 31605 1432 31669
rect 1496 31605 2700 31669
rect 99 31589 2700 31605
rect 99 31525 982 31589
rect 1046 31525 1072 31589
rect 1136 31525 1162 31589
rect 1226 31525 1252 31589
rect 1316 31525 1342 31589
rect 1406 31525 1432 31589
rect 1496 31525 2700 31589
rect 99 31509 2700 31525
rect 99 31445 982 31509
rect 1046 31445 1072 31509
rect 1136 31445 1162 31509
rect 1226 31445 1252 31509
rect 1316 31445 1342 31509
rect 1406 31445 1432 31509
rect 1496 31445 2700 31509
rect 99 31429 2700 31445
rect 99 31365 982 31429
rect 1046 31365 1072 31429
rect 1136 31365 1162 31429
rect 1226 31365 1252 31429
rect 1316 31365 1342 31429
rect 1406 31365 1432 31429
rect 1496 31365 2700 31429
rect 99 31349 2700 31365
rect 99 31344 982 31349
rect 1046 31344 1072 31349
rect 1136 31344 1162 31349
rect 1226 31344 1252 31349
rect 1316 31344 1342 31349
rect 1406 31344 1432 31349
rect 1496 31344 2700 31349
rect 99 23288 466 31344
rect 2442 23288 2700 31344
rect 99 23285 982 23288
rect 1046 23285 1072 23288
rect 1136 23285 1162 23288
rect 1226 23285 1252 23288
rect 1316 23285 1342 23288
rect 1406 23285 1432 23288
rect 1496 23285 2700 23288
rect 99 23268 2700 23285
rect 99 23204 982 23268
rect 1046 23204 1072 23268
rect 1136 23204 1162 23268
rect 1226 23204 1252 23268
rect 1316 23204 1342 23268
rect 1406 23204 1432 23268
rect 1496 23204 2700 23268
rect 99 23187 2700 23204
rect 99 23123 982 23187
rect 1046 23123 1072 23187
rect 1136 23123 1162 23187
rect 1226 23123 1252 23187
rect 1316 23123 1342 23187
rect 1406 23123 1432 23187
rect 1496 23123 2700 23187
rect 99 23106 2700 23123
rect 99 23042 982 23106
rect 1046 23042 1072 23106
rect 1136 23042 1162 23106
rect 1226 23042 1252 23106
rect 1316 23042 1342 23106
rect 1406 23042 1432 23106
rect 1496 23042 2700 23106
rect 99 23025 2700 23042
rect 99 22961 982 23025
rect 1046 22961 1072 23025
rect 1136 22961 1162 23025
rect 1226 22961 1252 23025
rect 1316 22961 1342 23025
rect 1406 22961 1432 23025
rect 1496 22961 2700 23025
rect 99 22944 2700 22961
rect 99 22880 982 22944
rect 1046 22880 1072 22944
rect 1136 22880 1162 22944
rect 1226 22880 1252 22944
rect 1316 22880 1342 22944
rect 1406 22880 1432 22944
rect 1496 22880 2700 22944
rect 99 22863 2700 22880
rect 99 22799 982 22863
rect 1046 22799 1072 22863
rect 1136 22799 1162 22863
rect 1226 22799 1252 22863
rect 1316 22799 1342 22863
rect 1406 22799 1432 22863
rect 1496 22799 2700 22863
rect 99 22782 2700 22799
rect 99 22718 982 22782
rect 1046 22718 1072 22782
rect 1136 22718 1162 22782
rect 1226 22718 1252 22782
rect 1316 22718 1342 22782
rect 1406 22718 1432 22782
rect 1496 22718 2700 22782
rect 99 22701 2700 22718
rect 99 22637 982 22701
rect 1046 22637 1072 22701
rect 1136 22637 1162 22701
rect 1226 22637 1252 22701
rect 1316 22637 1342 22701
rect 1406 22637 1432 22701
rect 1496 22637 2700 22701
rect 99 22620 2700 22637
rect 99 22556 982 22620
rect 1046 22556 1072 22620
rect 1136 22556 1162 22620
rect 1226 22556 1252 22620
rect 1316 22556 1342 22620
rect 1406 22556 1432 22620
rect 1496 22556 2700 22620
rect 99 22539 2700 22556
rect 99 22475 982 22539
rect 1046 22475 1072 22539
rect 1136 22475 1162 22539
rect 1226 22475 1252 22539
rect 1316 22475 1342 22539
rect 1406 22475 1432 22539
rect 1496 22475 2700 22539
rect 99 22458 2700 22475
rect 99 22394 982 22458
rect 1046 22394 1072 22458
rect 1136 22394 1162 22458
rect 1226 22394 1252 22458
rect 1316 22394 1342 22458
rect 1406 22394 1432 22458
rect 1496 22394 2700 22458
rect 99 22377 2700 22394
rect 99 22313 982 22377
rect 1046 22313 1072 22377
rect 1136 22313 1162 22377
rect 1226 22313 1252 22377
rect 1316 22313 1342 22377
rect 1406 22313 1432 22377
rect 1496 22313 2700 22377
rect 99 22296 2700 22313
rect 99 22232 982 22296
rect 1046 22232 1072 22296
rect 1136 22232 1162 22296
rect 1226 22232 1252 22296
rect 1316 22232 1342 22296
rect 1406 22232 1432 22296
rect 1496 22232 2700 22296
rect 99 22215 2700 22232
rect 99 22151 982 22215
rect 1046 22151 1072 22215
rect 1136 22151 1162 22215
rect 1226 22151 1252 22215
rect 1316 22151 1342 22215
rect 1406 22151 1432 22215
rect 1496 22151 2700 22215
rect 99 22134 2700 22151
rect 99 22070 982 22134
rect 1046 22070 1072 22134
rect 1136 22070 1162 22134
rect 1226 22070 1252 22134
rect 1316 22070 1342 22134
rect 1406 22070 1432 22134
rect 1496 22070 2700 22134
rect 99 22053 2700 22070
rect 99 21989 982 22053
rect 1046 21989 1072 22053
rect 1136 21989 1162 22053
rect 1226 21989 1252 22053
rect 1316 21989 1342 22053
rect 1406 21989 1432 22053
rect 1496 21989 2700 22053
rect 99 21972 2700 21989
rect 99 21908 982 21972
rect 1046 21908 1072 21972
rect 1136 21908 1162 21972
rect 1226 21908 1252 21972
rect 1316 21908 1342 21972
rect 1406 21908 1432 21972
rect 1496 21908 2700 21972
rect 99 21891 2700 21908
rect 99 21827 982 21891
rect 1046 21827 1072 21891
rect 1136 21827 1162 21891
rect 1226 21827 1252 21891
rect 1316 21827 1342 21891
rect 1406 21827 1432 21891
rect 1496 21827 2700 21891
rect 99 21810 2700 21827
rect 99 21746 982 21810
rect 1046 21746 1072 21810
rect 1136 21746 1162 21810
rect 1226 21746 1252 21810
rect 1316 21746 1342 21810
rect 1406 21746 1432 21810
rect 1496 21746 2700 21810
rect 99 21729 2700 21746
rect 99 21665 982 21729
rect 1046 21665 1072 21729
rect 1136 21665 1162 21729
rect 1226 21665 1252 21729
rect 1316 21665 1342 21729
rect 1406 21665 1432 21729
rect 1496 21665 2700 21729
rect 99 21648 2700 21665
rect 99 21584 982 21648
rect 1046 21584 1072 21648
rect 1136 21584 1162 21648
rect 1226 21584 1252 21648
rect 1316 21584 1342 21648
rect 1406 21584 1432 21648
rect 1496 21584 2700 21648
rect 99 21567 2700 21584
rect 99 21503 982 21567
rect 1046 21503 1072 21567
rect 1136 21503 1162 21567
rect 1226 21503 1252 21567
rect 1316 21503 1342 21567
rect 1406 21503 1432 21567
rect 1496 21503 2700 21567
rect 99 21486 2700 21503
rect 99 21422 982 21486
rect 1046 21422 1072 21486
rect 1136 21422 1162 21486
rect 1226 21422 1252 21486
rect 1316 21422 1342 21486
rect 1406 21422 1432 21486
rect 1496 21422 2700 21486
rect 99 21405 2700 21422
rect 99 21341 982 21405
rect 1046 21341 1072 21405
rect 1136 21341 1162 21405
rect 1226 21341 1252 21405
rect 1316 21341 1342 21405
rect 1406 21341 1432 21405
rect 1496 21341 2700 21405
rect 99 21324 2700 21341
rect 99 21260 982 21324
rect 1046 21260 1072 21324
rect 1136 21260 1162 21324
rect 1226 21260 1252 21324
rect 1316 21260 1342 21324
rect 1406 21260 1432 21324
rect 1496 21260 2700 21324
rect 99 21243 2700 21260
rect 99 21179 982 21243
rect 1046 21179 1072 21243
rect 1136 21179 1162 21243
rect 1226 21179 1252 21243
rect 1316 21179 1342 21243
rect 1406 21179 1432 21243
rect 1496 21179 2700 21243
rect 99 21162 2700 21179
rect 99 21098 982 21162
rect 1046 21098 1072 21162
rect 1136 21098 1162 21162
rect 1226 21098 1252 21162
rect 1316 21098 1342 21162
rect 1406 21098 1432 21162
rect 1496 21098 2700 21162
rect 99 21081 2700 21098
rect 99 21017 982 21081
rect 1046 21017 1072 21081
rect 1136 21017 1162 21081
rect 1226 21017 1252 21081
rect 1316 21017 1342 21081
rect 1406 21017 1432 21081
rect 1496 21017 2700 21081
rect 99 21000 2700 21017
rect 99 20936 982 21000
rect 1046 20936 1072 21000
rect 1136 20936 1162 21000
rect 1226 20936 1252 21000
rect 1316 20936 1342 21000
rect 1406 20936 1432 21000
rect 1496 20939 2700 21000
rect 1496 20936 1531 20939
rect 99 20919 1531 20936
rect 99 20855 982 20919
rect 1046 20855 1072 20919
rect 1136 20855 1162 20919
rect 1226 20855 1252 20919
rect 1316 20855 1342 20919
rect 1406 20855 1432 20919
rect 1496 20875 1531 20919
rect 1595 20875 2700 20939
rect 1496 20855 2700 20875
rect 99 20825 2700 20855
rect 99 20783 1312 20825
rect 99 20719 1141 20783
rect 1205 20761 1312 20783
rect 1376 20761 1401 20825
rect 1465 20761 1491 20825
rect 1555 20761 1581 20825
rect 1645 20761 1671 20825
rect 1735 20761 2700 20825
rect 1205 20719 2700 20761
rect 99 20709 2700 20719
rect 99 20645 1312 20709
rect 1376 20645 1401 20709
rect 1465 20645 1491 20709
rect 1555 20645 1581 20709
rect 1645 20645 1671 20709
rect 1735 20645 2700 20709
rect 99 20631 2700 20645
rect 99 20593 1812 20631
rect 99 20529 1312 20593
rect 1376 20529 1401 20593
rect 1465 20529 1491 20593
rect 1555 20529 1581 20593
rect 1645 20529 1671 20593
rect 1735 20567 1812 20593
rect 1876 20567 2700 20631
rect 1735 20529 2700 20567
rect 99 20505 2700 20529
rect 99 20469 1632 20505
rect 99 20405 1524 20469
rect 1588 20441 1632 20469
rect 1696 20441 1721 20505
rect 1785 20441 1811 20505
rect 1875 20441 1901 20505
rect 1965 20441 1991 20505
rect 2055 20441 2700 20505
rect 1588 20405 2700 20441
rect 99 20389 2700 20405
rect 99 20325 1632 20389
rect 1696 20325 1721 20389
rect 1785 20325 1811 20389
rect 1875 20325 1901 20389
rect 1965 20325 1991 20389
rect 2055 20325 2700 20389
rect 99 20306 2700 20325
rect 99 20273 2137 20306
rect 99 20209 1632 20273
rect 1696 20209 1721 20273
rect 1785 20209 1811 20273
rect 1875 20209 1901 20273
rect 1965 20209 1991 20273
rect 2055 20242 2137 20273
rect 2201 20242 2700 20306
rect 12300 33434 14858 33458
rect 12300 33396 13489 33434
rect 12300 33332 13348 33396
rect 13412 33370 13489 33396
rect 13553 33370 13579 33434
rect 13643 33370 13669 33434
rect 13733 33370 13759 33434
rect 13823 33370 13848 33434
rect 13912 33370 14858 33434
rect 13412 33332 14858 33370
rect 12300 33318 14858 33332
rect 12300 33254 13489 33318
rect 13553 33254 13579 33318
rect 13643 33254 13669 33318
rect 13733 33254 13759 33318
rect 13823 33254 13848 33318
rect 13912 33254 14858 33318
rect 12300 33202 14858 33254
rect 12300 33138 13489 33202
rect 13553 33138 13579 33202
rect 13643 33138 13669 33202
rect 13733 33138 13759 33202
rect 13823 33138 13848 33202
rect 13912 33138 14858 33202
rect 12300 33109 14858 33138
rect 12300 33045 13520 33109
rect 13584 33045 13610 33109
rect 13674 33045 13700 33109
rect 13764 33045 13790 33109
rect 13854 33045 13880 33109
rect 13944 33045 13970 33109
rect 14034 33045 14858 33109
rect 12300 33029 14858 33045
rect 12300 32965 13520 33029
rect 13584 32965 13610 33029
rect 13674 32965 13700 33029
rect 13764 32965 13790 33029
rect 13854 32965 13880 33029
rect 13944 32965 13970 33029
rect 14034 32965 14858 33029
rect 12300 32949 14858 32965
rect 12300 32885 13520 32949
rect 13584 32885 13610 32949
rect 13674 32885 13700 32949
rect 13764 32885 13790 32949
rect 13854 32885 13880 32949
rect 13944 32885 13970 32949
rect 14034 32885 14858 32949
rect 12300 32869 14858 32885
rect 12300 32805 13520 32869
rect 13584 32805 13610 32869
rect 13674 32805 13700 32869
rect 13764 32805 13790 32869
rect 13854 32805 13880 32869
rect 13944 32805 13970 32869
rect 14034 32805 14858 32869
rect 12300 32789 14858 32805
rect 12300 32725 13520 32789
rect 13584 32725 13610 32789
rect 13674 32725 13700 32789
rect 13764 32725 13790 32789
rect 13854 32725 13880 32789
rect 13944 32725 13970 32789
rect 14034 32725 14858 32789
rect 12300 32709 14858 32725
rect 12300 32645 13520 32709
rect 13584 32645 13610 32709
rect 13674 32645 13700 32709
rect 13764 32645 13790 32709
rect 13854 32645 13880 32709
rect 13944 32645 13970 32709
rect 14034 32645 14858 32709
rect 12300 32629 14858 32645
rect 12300 32565 13520 32629
rect 13584 32565 13610 32629
rect 13674 32565 13700 32629
rect 13764 32565 13790 32629
rect 13854 32565 13880 32629
rect 13944 32565 13970 32629
rect 14034 32565 14858 32629
rect 12300 32549 14858 32565
rect 12300 32485 13520 32549
rect 13584 32485 13610 32549
rect 13674 32485 13700 32549
rect 13764 32485 13790 32549
rect 13854 32485 13880 32549
rect 13944 32485 13970 32549
rect 14034 32485 14858 32549
rect 12300 32469 14858 32485
rect 12300 32405 13520 32469
rect 13584 32405 13610 32469
rect 13674 32405 13700 32469
rect 13764 32405 13790 32469
rect 13854 32405 13880 32469
rect 13944 32405 13970 32469
rect 14034 32405 14858 32469
rect 12300 32389 14858 32405
rect 12300 32325 13520 32389
rect 13584 32325 13610 32389
rect 13674 32325 13700 32389
rect 13764 32325 13790 32389
rect 13854 32325 13880 32389
rect 13944 32325 13970 32389
rect 14034 32325 14858 32389
rect 12300 32309 14858 32325
rect 12300 32245 13520 32309
rect 13584 32245 13610 32309
rect 13674 32245 13700 32309
rect 13764 32245 13790 32309
rect 13854 32245 13880 32309
rect 13944 32245 13970 32309
rect 14034 32245 14858 32309
rect 12300 32229 14858 32245
rect 12300 32165 13520 32229
rect 13584 32165 13610 32229
rect 13674 32165 13700 32229
rect 13764 32165 13790 32229
rect 13854 32165 13880 32229
rect 13944 32165 13970 32229
rect 14034 32165 14858 32229
rect 12300 32149 14858 32165
rect 12300 32085 13520 32149
rect 13584 32085 13610 32149
rect 13674 32085 13700 32149
rect 13764 32085 13790 32149
rect 13854 32085 13880 32149
rect 13944 32085 13970 32149
rect 14034 32085 14858 32149
rect 12300 32069 14858 32085
rect 12300 32005 13520 32069
rect 13584 32005 13610 32069
rect 13674 32005 13700 32069
rect 13764 32005 13790 32069
rect 13854 32005 13880 32069
rect 13944 32005 13970 32069
rect 14034 32005 14858 32069
rect 12300 31989 14858 32005
rect 12300 31925 13520 31989
rect 13584 31925 13610 31989
rect 13674 31925 13700 31989
rect 13764 31925 13790 31989
rect 13854 31925 13880 31989
rect 13944 31925 13970 31989
rect 14034 31925 14858 31989
rect 12300 31909 14858 31925
rect 12300 31845 13520 31909
rect 13584 31845 13610 31909
rect 13674 31845 13700 31909
rect 13764 31845 13790 31909
rect 13854 31845 13880 31909
rect 13944 31845 13970 31909
rect 14034 31845 14858 31909
rect 12300 31829 14858 31845
rect 12300 31765 13520 31829
rect 13584 31765 13610 31829
rect 13674 31765 13700 31829
rect 13764 31765 13790 31829
rect 13854 31765 13880 31829
rect 13944 31765 13970 31829
rect 14034 31765 14858 31829
rect 12300 31749 14858 31765
rect 12300 31685 13520 31749
rect 13584 31685 13610 31749
rect 13674 31685 13700 31749
rect 13764 31685 13790 31749
rect 13854 31685 13880 31749
rect 13944 31685 13970 31749
rect 14034 31685 14858 31749
rect 12300 31669 14858 31685
rect 12300 31605 13520 31669
rect 13584 31605 13610 31669
rect 13674 31605 13700 31669
rect 13764 31605 13790 31669
rect 13854 31605 13880 31669
rect 13944 31605 13970 31669
rect 14034 31605 14858 31669
rect 12300 31589 14858 31605
rect 12300 31525 13520 31589
rect 13584 31525 13610 31589
rect 13674 31525 13700 31589
rect 13764 31525 13790 31589
rect 13854 31525 13880 31589
rect 13944 31525 13970 31589
rect 14034 31525 14858 31589
rect 12300 31509 14858 31525
rect 12300 31445 13520 31509
rect 13584 31445 13610 31509
rect 13674 31445 13700 31509
rect 13764 31445 13790 31509
rect 13854 31445 13880 31509
rect 13944 31445 13970 31509
rect 14034 31445 14858 31509
rect 12300 31429 14858 31445
rect 12300 31392 13520 31429
rect 13584 31392 13610 31429
rect 13674 31392 13700 31429
rect 13764 31392 13790 31429
rect 13854 31392 13880 31429
rect 13944 31392 13970 31429
rect 14034 31392 14858 31429
rect 12300 23336 12455 31392
rect 14431 23336 14858 31392
rect 12300 23285 13520 23336
rect 13584 23285 13610 23336
rect 13674 23285 13700 23336
rect 13764 23285 13790 23336
rect 13854 23285 13880 23336
rect 13944 23285 13970 23336
rect 14034 23285 14858 23336
rect 12300 23268 14858 23285
rect 12300 23204 13520 23268
rect 13584 23204 13610 23268
rect 13674 23204 13700 23268
rect 13764 23204 13790 23268
rect 13854 23204 13880 23268
rect 13944 23204 13970 23268
rect 14034 23204 14858 23268
rect 12300 23187 14858 23204
rect 12300 23123 13520 23187
rect 13584 23123 13610 23187
rect 13674 23123 13700 23187
rect 13764 23123 13790 23187
rect 13854 23123 13880 23187
rect 13944 23123 13970 23187
rect 14034 23123 14858 23187
rect 12300 23106 14858 23123
rect 12300 23042 13520 23106
rect 13584 23042 13610 23106
rect 13674 23042 13700 23106
rect 13764 23042 13790 23106
rect 13854 23042 13880 23106
rect 13944 23042 13970 23106
rect 14034 23042 14858 23106
rect 12300 23025 14858 23042
rect 12300 22961 13520 23025
rect 13584 22961 13610 23025
rect 13674 22961 13700 23025
rect 13764 22961 13790 23025
rect 13854 22961 13880 23025
rect 13944 22961 13970 23025
rect 14034 22961 14858 23025
rect 12300 22944 14858 22961
rect 12300 22880 13520 22944
rect 13584 22880 13610 22944
rect 13674 22880 13700 22944
rect 13764 22880 13790 22944
rect 13854 22880 13880 22944
rect 13944 22880 13970 22944
rect 14034 22880 14858 22944
rect 12300 22863 14858 22880
rect 12300 22799 13520 22863
rect 13584 22799 13610 22863
rect 13674 22799 13700 22863
rect 13764 22799 13790 22863
rect 13854 22799 13880 22863
rect 13944 22799 13970 22863
rect 14034 22799 14858 22863
rect 12300 22782 14858 22799
rect 12300 22718 13520 22782
rect 13584 22718 13610 22782
rect 13674 22718 13700 22782
rect 13764 22718 13790 22782
rect 13854 22718 13880 22782
rect 13944 22718 13970 22782
rect 14034 22718 14858 22782
rect 12300 22701 14858 22718
rect 12300 22637 13520 22701
rect 13584 22637 13610 22701
rect 13674 22637 13700 22701
rect 13764 22637 13790 22701
rect 13854 22637 13880 22701
rect 13944 22637 13970 22701
rect 14034 22637 14858 22701
rect 12300 22620 14858 22637
rect 12300 22556 13520 22620
rect 13584 22556 13610 22620
rect 13674 22556 13700 22620
rect 13764 22556 13790 22620
rect 13854 22556 13880 22620
rect 13944 22556 13970 22620
rect 14034 22556 14858 22620
rect 12300 22539 14858 22556
rect 12300 22475 13520 22539
rect 13584 22475 13610 22539
rect 13674 22475 13700 22539
rect 13764 22475 13790 22539
rect 13854 22475 13880 22539
rect 13944 22475 13970 22539
rect 14034 22475 14858 22539
rect 12300 22458 14858 22475
rect 12300 22394 13520 22458
rect 13584 22394 13610 22458
rect 13674 22394 13700 22458
rect 13764 22394 13790 22458
rect 13854 22394 13880 22458
rect 13944 22394 13970 22458
rect 14034 22394 14858 22458
rect 12300 22377 14858 22394
rect 12300 22313 13520 22377
rect 13584 22313 13610 22377
rect 13674 22313 13700 22377
rect 13764 22313 13790 22377
rect 13854 22313 13880 22377
rect 13944 22313 13970 22377
rect 14034 22313 14858 22377
rect 12300 22296 14858 22313
rect 12300 22232 13520 22296
rect 13584 22232 13610 22296
rect 13674 22232 13700 22296
rect 13764 22232 13790 22296
rect 13854 22232 13880 22296
rect 13944 22232 13970 22296
rect 14034 22232 14858 22296
rect 12300 22215 14858 22232
rect 12300 22151 13520 22215
rect 13584 22151 13610 22215
rect 13674 22151 13700 22215
rect 13764 22151 13790 22215
rect 13854 22151 13880 22215
rect 13944 22151 13970 22215
rect 14034 22151 14858 22215
rect 12300 22134 14858 22151
rect 12300 22070 13520 22134
rect 13584 22070 13610 22134
rect 13674 22070 13700 22134
rect 13764 22070 13790 22134
rect 13854 22070 13880 22134
rect 13944 22070 13970 22134
rect 14034 22070 14858 22134
rect 12300 22053 14858 22070
rect 12300 21989 13520 22053
rect 13584 21989 13610 22053
rect 13674 21989 13700 22053
rect 13764 21989 13790 22053
rect 13854 21989 13880 22053
rect 13944 21989 13970 22053
rect 14034 21989 14858 22053
rect 12300 21972 14858 21989
rect 12300 21908 13520 21972
rect 13584 21908 13610 21972
rect 13674 21908 13700 21972
rect 13764 21908 13790 21972
rect 13854 21908 13880 21972
rect 13944 21908 13970 21972
rect 14034 21908 14858 21972
rect 12300 21891 14858 21908
rect 12300 21827 13520 21891
rect 13584 21827 13610 21891
rect 13674 21827 13700 21891
rect 13764 21827 13790 21891
rect 13854 21827 13880 21891
rect 13944 21827 13970 21891
rect 14034 21827 14858 21891
rect 12300 21810 14858 21827
rect 12300 21746 13520 21810
rect 13584 21746 13610 21810
rect 13674 21746 13700 21810
rect 13764 21746 13790 21810
rect 13854 21746 13880 21810
rect 13944 21746 13970 21810
rect 14034 21746 14858 21810
rect 12300 21729 14858 21746
rect 12300 21665 13520 21729
rect 13584 21665 13610 21729
rect 13674 21665 13700 21729
rect 13764 21665 13790 21729
rect 13854 21665 13880 21729
rect 13944 21665 13970 21729
rect 14034 21665 14858 21729
rect 12300 21648 14858 21665
rect 12300 21584 13520 21648
rect 13584 21584 13610 21648
rect 13674 21584 13700 21648
rect 13764 21584 13790 21648
rect 13854 21584 13880 21648
rect 13944 21584 13970 21648
rect 14034 21584 14858 21648
rect 12300 21567 14858 21584
rect 12300 21503 13520 21567
rect 13584 21503 13610 21567
rect 13674 21503 13700 21567
rect 13764 21503 13790 21567
rect 13854 21503 13880 21567
rect 13944 21503 13970 21567
rect 14034 21503 14858 21567
rect 12300 21486 14858 21503
rect 12300 21422 13520 21486
rect 13584 21422 13610 21486
rect 13674 21422 13700 21486
rect 13764 21422 13790 21486
rect 13854 21422 13880 21486
rect 13944 21422 13970 21486
rect 14034 21422 14858 21486
rect 12300 21405 14858 21422
rect 12300 21341 13520 21405
rect 13584 21341 13610 21405
rect 13674 21341 13700 21405
rect 13764 21341 13790 21405
rect 13854 21341 13880 21405
rect 13944 21341 13970 21405
rect 14034 21341 14858 21405
rect 12300 21324 14858 21341
rect 12300 21260 13520 21324
rect 13584 21260 13610 21324
rect 13674 21260 13700 21324
rect 13764 21260 13790 21324
rect 13854 21260 13880 21324
rect 13944 21260 13970 21324
rect 14034 21260 14858 21324
rect 12300 21243 14858 21260
rect 12300 21179 13520 21243
rect 13584 21179 13610 21243
rect 13674 21179 13700 21243
rect 13764 21179 13790 21243
rect 13854 21179 13880 21243
rect 13944 21179 13970 21243
rect 14034 21179 14858 21243
rect 12300 21162 14858 21179
rect 12300 21098 13520 21162
rect 13584 21098 13610 21162
rect 13674 21098 13700 21162
rect 13764 21098 13790 21162
rect 13854 21098 13880 21162
rect 13944 21098 13970 21162
rect 14034 21098 14858 21162
rect 12300 21081 14858 21098
rect 12300 21017 13520 21081
rect 13584 21017 13610 21081
rect 13674 21017 13700 21081
rect 13764 21017 13790 21081
rect 13854 21017 13880 21081
rect 13944 21017 13970 21081
rect 14034 21017 14858 21081
rect 12300 21000 14858 21017
rect 12300 20939 13520 21000
rect 12300 20875 13421 20939
rect 13485 20936 13520 20939
rect 13584 20936 13610 21000
rect 13674 20936 13700 21000
rect 13764 20936 13790 21000
rect 13854 20936 13880 21000
rect 13944 20936 13970 21000
rect 14034 20936 14858 21000
rect 13485 20919 14858 20936
rect 13485 20875 13520 20919
rect 12300 20855 13520 20875
rect 13584 20855 13610 20919
rect 13674 20855 13700 20919
rect 13764 20855 13790 20919
rect 13854 20855 13880 20919
rect 13944 20855 13970 20919
rect 14034 20855 14858 20919
rect 12300 20825 14858 20855
rect 12300 20761 13281 20825
rect 13345 20761 13371 20825
rect 13435 20761 13461 20825
rect 13525 20761 13551 20825
rect 13615 20761 13640 20825
rect 13704 20823 14858 20825
rect 13704 20761 13749 20823
rect 12300 20759 13749 20761
rect 13813 20816 14858 20823
rect 13813 20759 13851 20816
rect 12300 20752 13851 20759
rect 13915 20752 14858 20816
rect 12300 20712 14858 20752
rect 12300 20709 13749 20712
rect 12300 20645 13281 20709
rect 13345 20645 13371 20709
rect 13435 20645 13461 20709
rect 13525 20645 13551 20709
rect 13615 20645 13640 20709
rect 13704 20648 13749 20709
rect 13813 20648 14858 20712
rect 13704 20645 14858 20648
rect 12300 20631 14858 20645
rect 12300 20567 13140 20631
rect 13204 20593 14858 20631
rect 13204 20567 13281 20593
rect 12300 20529 13281 20567
rect 13345 20529 13371 20593
rect 13435 20529 13461 20593
rect 13525 20529 13551 20593
rect 13615 20529 13640 20593
rect 13704 20529 14858 20593
rect 12300 20505 14858 20529
rect 12300 20441 12961 20505
rect 13025 20441 13051 20505
rect 13115 20441 13141 20505
rect 13205 20441 13231 20505
rect 13295 20441 13320 20505
rect 13384 20469 14858 20505
rect 13384 20441 13428 20469
rect 12300 20405 13428 20441
rect 13492 20405 14858 20469
rect 12300 20389 14858 20405
rect 12300 20325 12961 20389
rect 13025 20325 13051 20389
rect 13115 20325 13141 20389
rect 13205 20325 13231 20389
rect 13295 20325 13320 20389
rect 13384 20325 14858 20389
rect 12300 20306 14858 20325
rect 2055 20209 2700 20242
rect 99 20181 2700 20209
rect 99 20141 1956 20181
rect 99 20077 1852 20141
rect 1916 20117 1956 20141
rect 2020 20117 2045 20181
rect 2109 20117 2135 20181
rect 2199 20117 2225 20181
rect 2289 20117 2315 20181
rect 2379 20117 2700 20181
rect 1916 20077 2700 20117
rect 99 20070 2700 20077
tri 2700 20070 2909 20279 sw
tri 12111 20070 12300 20259 se
rect 12300 20242 12815 20306
rect 12879 20273 14858 20306
rect 12879 20242 12961 20273
rect 12300 20209 12961 20242
rect 13025 20209 13051 20273
rect 13115 20209 13141 20273
rect 13205 20209 13231 20273
rect 13295 20209 13320 20273
rect 13384 20209 14858 20273
rect 12300 20181 14858 20209
rect 12300 20117 12637 20181
rect 12701 20117 12727 20181
rect 12791 20117 12817 20181
rect 12881 20117 12907 20181
rect 12971 20117 12996 20181
rect 13060 20141 14858 20181
rect 13060 20117 13100 20141
rect 12300 20077 13100 20117
rect 13164 20077 14858 20141
rect 12300 20070 14858 20077
rect 99 20065 2456 20070
rect 99 20001 1956 20065
rect 2020 20001 2045 20065
rect 2109 20001 2135 20065
rect 2199 20001 2225 20065
rect 2289 20001 2315 20065
rect 2379 20006 2456 20065
rect 2520 20006 2571 20070
rect 2635 20006 2686 20070
rect 2750 20006 2802 20070
rect 2866 20006 2909 20070
rect 2379 20005 2909 20006
tri 2909 20005 2974 20070 sw
tri 12110 20069 12111 20070 se
rect 12111 20069 12150 20070
tri 12046 20005 12110 20069 se
rect 12110 20006 12150 20069
rect 12214 20006 12266 20070
rect 12330 20006 12381 20070
rect 12445 20006 12496 20070
rect 12560 20065 14858 20070
rect 12560 20006 12637 20065
rect 12110 20005 12637 20006
rect 2379 20001 2974 20005
rect 99 19955 2974 20001
rect 99 19950 2906 19955
rect 99 19949 2456 19950
rect 99 19885 1956 19949
rect 2020 19885 2045 19949
rect 2109 19885 2135 19949
rect 2199 19885 2225 19949
rect 2289 19885 2315 19949
rect 2379 19886 2456 19949
rect 2520 19886 2571 19950
rect 2635 19886 2686 19950
rect 2750 19886 2802 19950
rect 2866 19891 2906 19950
rect 2970 19891 2974 19955
rect 2866 19886 2974 19891
rect 2379 19885 2974 19886
rect 99 19844 2974 19885
tri 2974 19844 3135 20005 sw
tri 12027 19986 12046 20005 se
rect 12046 20001 12637 20005
rect 12701 20001 12727 20065
rect 12791 20001 12817 20065
rect 12881 20001 12907 20065
rect 12971 20001 12996 20065
rect 13060 20001 14858 20065
rect 12046 19986 14858 20001
tri 11885 19844 12027 19986 se
rect 12027 19955 14858 19986
rect 12027 19891 12046 19955
rect 12110 19950 14858 19955
rect 12110 19891 12150 19950
rect 12027 19886 12150 19891
rect 12214 19886 12266 19950
rect 12330 19886 12381 19950
rect 12445 19886 12496 19950
rect 12560 19949 14858 19950
rect 12560 19886 12637 19949
rect 12027 19885 12637 19886
rect 12701 19885 12727 19949
rect 12791 19885 12817 19949
rect 12881 19885 12907 19949
rect 12971 19885 12996 19949
rect 13060 19885 14858 19949
rect 12027 19844 14858 19885
rect 99 19800 2293 19844
rect 99 19736 2193 19800
rect 2257 19780 2293 19800
rect 2357 19780 2377 19844
rect 2441 19780 2461 19844
rect 2525 19780 2545 19844
rect 2609 19780 2629 19844
rect 2693 19780 2713 19844
rect 2777 19780 2797 19844
rect 2861 19780 2881 19844
rect 2945 19780 2965 19844
rect 3029 19780 3049 19844
rect 3113 19780 3135 19844
rect 2257 19736 3135 19780
rect 99 19728 3135 19736
rect 99 19664 2293 19728
rect 2357 19664 2377 19728
rect 2441 19664 2461 19728
rect 2525 19664 2545 19728
rect 2609 19664 2629 19728
rect 2693 19664 2713 19728
rect 2777 19664 2797 19728
rect 2861 19664 2881 19728
rect 2945 19664 2965 19728
rect 3029 19664 3049 19728
rect 3113 19707 3135 19728
tri 3135 19707 3272 19844 sw
tri 11753 19712 11885 19844 se
rect 11885 19780 11903 19844
rect 11967 19780 11987 19844
rect 12051 19780 12071 19844
rect 12135 19780 12155 19844
rect 12219 19780 12239 19844
rect 12303 19780 12323 19844
rect 12387 19780 12407 19844
rect 12471 19780 12491 19844
rect 12555 19780 12575 19844
rect 12639 19780 12659 19844
rect 12723 19800 14858 19844
rect 12723 19780 12759 19800
rect 11885 19736 12759 19780
rect 12823 19736 14858 19800
rect 11885 19728 14858 19736
rect 11885 19712 11903 19728
tri 11748 19707 11753 19712 se
rect 11753 19707 11903 19712
rect 3113 19664 3153 19707
rect 99 19643 3153 19664
rect 3217 19643 3272 19707
rect 99 19614 3272 19643
rect 99 19612 3153 19614
rect 99 19548 2293 19612
rect 2357 19548 2377 19612
rect 2441 19548 2461 19612
rect 2525 19548 2545 19612
rect 2609 19548 2629 19612
rect 2693 19548 2713 19612
rect 2777 19548 2797 19612
rect 2861 19548 2881 19612
rect 2945 19548 2965 19612
rect 3029 19548 3049 19612
rect 3113 19550 3153 19612
rect 3217 19550 3272 19614
rect 3113 19548 3272 19550
rect 99 18934 3272 19548
tri 3272 18934 4045 19707 sw
tri 11237 19196 11748 19707 se
rect 11748 19643 11799 19707
rect 11863 19664 11903 19707
rect 11967 19664 11987 19728
rect 12051 19664 12071 19728
rect 12135 19664 12155 19728
rect 12219 19664 12239 19728
rect 12303 19664 12323 19728
rect 12387 19664 12407 19728
rect 12471 19664 12491 19728
rect 12555 19664 12575 19728
rect 12639 19664 12659 19728
rect 12723 19664 14858 19728
rect 11863 19643 14858 19664
rect 11748 19614 14858 19643
rect 11748 19550 11799 19614
rect 11863 19612 14858 19614
rect 11863 19550 11903 19612
rect 11748 19548 11903 19550
rect 11967 19548 11987 19612
rect 12051 19548 12071 19612
rect 12135 19548 12155 19612
rect 12219 19548 12239 19612
rect 12303 19548 12323 19612
rect 12387 19548 12407 19612
rect 12471 19548 12491 19612
rect 12555 19548 12575 19612
rect 12639 19548 12659 19612
rect 12723 19548 14858 19612
rect 11748 19196 14858 19548
tri 4842 18996 5042 19196 se
rect 5042 18996 9935 19196
tri 9935 18996 10135 19196 sw
rect 99 18931 4045 18934
tri 4045 18931 4048 18934 sw
rect 4842 18931 10135 18996
rect 99 18871 4048 18931
tri 4048 18871 4108 18931 sw
rect 99 17061 4108 18871
rect 4842 18895 4942 18931
rect 7238 18895 7742 18931
rect 10038 18895 10135 18931
rect 4842 17311 4938 18895
rect 7242 17311 7738 18895
rect 10042 17311 10135 18895
rect 4842 17275 4942 17311
rect 7238 17275 7742 17311
rect 10038 17275 10135 17311
rect 4842 17230 10135 17275
tri 4842 17214 4858 17230 ne
rect 4858 17218 9935 17230
rect 4858 17214 5099 17218
tri 4858 17078 4994 17214 ne
rect 4994 17078 5099 17214
tri 4994 17071 5001 17078 ne
rect 5001 17074 5099 17078
rect 7243 17074 7735 17218
rect 9879 17074 9935 17218
rect 5001 17071 9935 17074
tri 4108 17061 4118 17071 sw
tri 5001 17061 5011 17071 ne
rect 5011 17061 9935 17071
rect 99 16575 4118 17061
tri 99 14722 1952 16575 ne
rect 1952 16471 4118 16575
tri 4118 16471 4708 17061 sw
tri 5011 17030 5042 17061 ne
rect 5042 17030 9935 17061
tri 9935 17030 10135 17230 nw
tri 10912 18871 11237 19196 se
rect 11237 18871 14858 19196
tri 10872 17030 10912 17070 se
rect 10912 17030 14858 18871
tri 10313 16471 10872 17030 se
rect 10872 16628 14858 17030
rect 10872 16471 12952 16628
rect 1952 14722 12952 16471
tri 12952 14722 14858 16628 nw
tri 1952 11722 4952 14722 ne
rect 858 9741 2098 9774
rect 858 9285 890 9741
rect 2066 9285 2098 9741
rect 858 4811 2098 9285
rect 2396 9501 3635 9528
rect 2396 8965 2427 9501
rect 3603 8965 3635 9501
rect 2396 6025 3635 8965
rect 2396 5241 2423 6025
rect 3607 5241 3635 6025
rect 2396 5122 3635 5241
rect 858 4027 887 4811
rect 2071 4027 2098 4811
rect 858 3955 2098 4027
rect 4952 1 9952 14722
tri 9952 11722 12952 14722 nw
rect 12858 9741 14098 9774
rect 11273 9502 12512 9529
rect 11273 8966 11304 9502
rect 12480 8966 12512 9502
rect 11273 6024 12512 8966
rect 11273 5240 11297 6024
rect 12481 5240 12512 6024
rect 11273 5122 12512 5240
rect 12858 9285 12890 9741
rect 14066 9285 14098 9741
rect 12858 4811 14098 9285
rect 12858 4027 12887 4811
rect 14071 4027 14098 4811
rect 12858 3955 14098 4027
<< via3 >>
rect 4975 39213 7199 39217
rect 4975 35317 4979 39213
rect 4979 35317 7195 39213
rect 7195 35317 7199 39213
rect 4975 35313 7199 35317
rect 7775 39213 9999 39217
rect 7775 35317 7779 39213
rect 7779 35317 9995 39213
rect 9995 35317 9999 39213
rect 7775 35313 9999 35317
rect 2276 34554 2340 34618
rect 2359 34554 2423 34618
rect 2443 34554 2507 34618
rect 2527 34554 2591 34618
rect 2611 34554 2675 34618
rect 12341 34554 12405 34618
rect 12425 34554 12489 34618
rect 12509 34554 12573 34618
rect 12593 34554 12657 34618
rect 12677 34554 12741 34618
rect 2276 34460 2340 34524
rect 2359 34460 2423 34524
rect 2443 34460 2507 34524
rect 2527 34460 2591 34524
rect 2611 34460 2675 34524
rect 12341 34460 12405 34524
rect 12425 34460 12489 34524
rect 12509 34460 12573 34524
rect 12593 34460 12657 34524
rect 12677 34460 12741 34524
rect 2148 34377 2212 34441
rect 2276 34366 2340 34430
rect 2359 34366 2423 34430
rect 2443 34366 2507 34430
rect 2527 34366 2591 34430
rect 2611 34366 2675 34430
rect 12341 34366 12405 34430
rect 12425 34366 12489 34430
rect 12509 34366 12573 34430
rect 12593 34366 12657 34430
rect 12677 34366 12741 34430
rect 12804 34377 12868 34441
rect 2004 34252 2068 34316
rect 2084 34252 2148 34316
rect 2164 34252 2228 34316
rect 2276 34272 2340 34336
rect 2359 34272 2423 34336
rect 2443 34272 2507 34336
rect 2527 34272 2591 34336
rect 2611 34272 2675 34336
rect 12341 34272 12405 34336
rect 12425 34272 12489 34336
rect 12509 34272 12573 34336
rect 12593 34272 12657 34336
rect 12677 34272 12741 34336
rect 12788 34252 12852 34316
rect 12868 34252 12932 34316
rect 12948 34252 13012 34316
rect 1890 34119 1954 34183
rect 2004 34156 2068 34220
rect 2084 34156 2148 34220
rect 2164 34156 2228 34220
rect 2276 34178 2340 34242
rect 2359 34178 2423 34242
rect 2443 34178 2507 34242
rect 2527 34178 2591 34242
rect 2611 34178 2675 34242
rect 12341 34178 12405 34242
rect 12425 34178 12489 34242
rect 12509 34178 12573 34242
rect 12593 34178 12657 34242
rect 12677 34178 12741 34242
rect 12788 34156 12852 34220
rect 12868 34156 12932 34220
rect 12948 34156 13012 34220
rect 2276 34084 2340 34148
rect 2359 34084 2423 34148
rect 2443 34084 2507 34148
rect 2527 34084 2591 34148
rect 2611 34084 2675 34148
rect 12341 34084 12405 34148
rect 12425 34084 12489 34148
rect 12509 34084 12573 34148
rect 12593 34084 12657 34148
rect 12677 34084 12741 34148
rect 13062 34119 13126 34183
rect 1748 34014 1812 34078
rect 1837 34014 1901 34078
rect 1927 34014 1991 34078
rect 2017 34014 2081 34078
rect 2107 34014 2171 34078
rect 12845 34014 12909 34078
rect 12935 34014 12999 34078
rect 13025 34014 13089 34078
rect 13115 34014 13179 34078
rect 13204 34014 13268 34078
rect 1748 33898 1812 33962
rect 1837 33898 1901 33962
rect 1927 33898 1991 33962
rect 2017 33898 2081 33962
rect 2107 33898 2171 33962
rect 2247 33945 2311 34009
rect 12705 33945 12769 34009
rect 12845 33898 12909 33962
rect 12935 33898 12999 33962
rect 13025 33898 13089 33962
rect 13115 33898 13179 33962
rect 13204 33898 13268 33962
rect 1644 33822 1708 33886
rect 1748 33782 1812 33846
rect 1837 33782 1901 33846
rect 1927 33782 1991 33846
rect 2017 33782 2081 33846
rect 2107 33782 2171 33846
rect 1424 33690 1488 33754
rect 1513 33690 1577 33754
rect 1603 33690 1667 33754
rect 1693 33690 1757 33754
rect 1783 33690 1847 33754
rect 1929 33657 1993 33721
rect 1424 33574 1488 33638
rect 1513 33574 1577 33638
rect 1603 33574 1667 33638
rect 1693 33574 1757 33638
rect 1783 33574 1847 33638
rect 1316 33494 1380 33558
rect 1424 33458 1488 33522
rect 1513 33458 1577 33522
rect 1603 33458 1667 33522
rect 1693 33458 1757 33522
rect 1783 33458 1847 33522
rect 12845 33782 12909 33846
rect 12935 33782 12999 33846
rect 13025 33782 13089 33846
rect 13115 33782 13179 33846
rect 13204 33782 13268 33846
rect 13308 33822 13372 33886
rect 13023 33657 13087 33721
rect 13169 33690 13233 33754
rect 13259 33690 13323 33754
rect 13349 33690 13413 33754
rect 13439 33690 13503 33754
rect 13528 33690 13592 33754
rect 13169 33574 13233 33638
rect 13259 33574 13323 33638
rect 13349 33574 13413 33638
rect 13439 33574 13503 33638
rect 13528 33574 13592 33638
rect 13169 33458 13233 33522
rect 13259 33458 13323 33522
rect 13349 33458 13413 33522
rect 13439 33458 13503 33522
rect 13528 33458 13592 33522
rect 13636 33494 13700 33558
rect 1104 33370 1168 33434
rect 1193 33370 1257 33434
rect 1283 33370 1347 33434
rect 1373 33370 1437 33434
rect 1463 33370 1527 33434
rect 1604 33332 1668 33396
rect 1104 33254 1168 33318
rect 1193 33254 1257 33318
rect 1283 33254 1347 33318
rect 1373 33254 1437 33318
rect 1463 33254 1527 33318
rect 1104 33138 1168 33202
rect 1193 33138 1257 33202
rect 1283 33138 1347 33202
rect 1373 33138 1437 33202
rect 1463 33138 1527 33202
rect 982 33045 1046 33109
rect 1072 33045 1136 33109
rect 1162 33045 1226 33109
rect 1252 33045 1316 33109
rect 1342 33045 1406 33109
rect 1432 33045 1496 33109
rect 982 32965 1046 33029
rect 1072 32965 1136 33029
rect 1162 32965 1226 33029
rect 1252 32965 1316 33029
rect 1342 32965 1406 33029
rect 1432 32965 1496 33029
rect 982 32885 1046 32949
rect 1072 32885 1136 32949
rect 1162 32885 1226 32949
rect 1252 32885 1316 32949
rect 1342 32885 1406 32949
rect 1432 32885 1496 32949
rect 982 32805 1046 32869
rect 1072 32805 1136 32869
rect 1162 32805 1226 32869
rect 1252 32805 1316 32869
rect 1342 32805 1406 32869
rect 1432 32805 1496 32869
rect 982 32725 1046 32789
rect 1072 32725 1136 32789
rect 1162 32725 1226 32789
rect 1252 32725 1316 32789
rect 1342 32725 1406 32789
rect 1432 32725 1496 32789
rect 982 32645 1046 32709
rect 1072 32645 1136 32709
rect 1162 32645 1226 32709
rect 1252 32645 1316 32709
rect 1342 32645 1406 32709
rect 1432 32645 1496 32709
rect 982 32565 1046 32629
rect 1072 32565 1136 32629
rect 1162 32565 1226 32629
rect 1252 32565 1316 32629
rect 1342 32565 1406 32629
rect 1432 32565 1496 32629
rect 982 32485 1046 32549
rect 1072 32485 1136 32549
rect 1162 32485 1226 32549
rect 1252 32485 1316 32549
rect 1342 32485 1406 32549
rect 1432 32485 1496 32549
rect 982 32405 1046 32469
rect 1072 32405 1136 32469
rect 1162 32405 1226 32469
rect 1252 32405 1316 32469
rect 1342 32405 1406 32469
rect 1432 32405 1496 32469
rect 982 32325 1046 32389
rect 1072 32325 1136 32389
rect 1162 32325 1226 32389
rect 1252 32325 1316 32389
rect 1342 32325 1406 32389
rect 1432 32325 1496 32389
rect 982 32245 1046 32309
rect 1072 32245 1136 32309
rect 1162 32245 1226 32309
rect 1252 32245 1316 32309
rect 1342 32245 1406 32309
rect 1432 32245 1496 32309
rect 982 32165 1046 32229
rect 1072 32165 1136 32229
rect 1162 32165 1226 32229
rect 1252 32165 1316 32229
rect 1342 32165 1406 32229
rect 1432 32165 1496 32229
rect 982 32085 1046 32149
rect 1072 32085 1136 32149
rect 1162 32085 1226 32149
rect 1252 32085 1316 32149
rect 1342 32085 1406 32149
rect 1432 32085 1496 32149
rect 982 32005 1046 32069
rect 1072 32005 1136 32069
rect 1162 32005 1226 32069
rect 1252 32005 1316 32069
rect 1342 32005 1406 32069
rect 1432 32005 1496 32069
rect 982 31925 1046 31989
rect 1072 31925 1136 31989
rect 1162 31925 1226 31989
rect 1252 31925 1316 31989
rect 1342 31925 1406 31989
rect 1432 31925 1496 31989
rect 982 31845 1046 31909
rect 1072 31845 1136 31909
rect 1162 31845 1226 31909
rect 1252 31845 1316 31909
rect 1342 31845 1406 31909
rect 1432 31845 1496 31909
rect 982 31765 1046 31829
rect 1072 31765 1136 31829
rect 1162 31765 1226 31829
rect 1252 31765 1316 31829
rect 1342 31765 1406 31829
rect 1432 31765 1496 31829
rect 982 31685 1046 31749
rect 1072 31685 1136 31749
rect 1162 31685 1226 31749
rect 1252 31685 1316 31749
rect 1342 31685 1406 31749
rect 1432 31685 1496 31749
rect 982 31605 1046 31669
rect 1072 31605 1136 31669
rect 1162 31605 1226 31669
rect 1252 31605 1316 31669
rect 1342 31605 1406 31669
rect 1432 31605 1496 31669
rect 982 31525 1046 31589
rect 1072 31525 1136 31589
rect 1162 31525 1226 31589
rect 1252 31525 1316 31589
rect 1342 31525 1406 31589
rect 1432 31525 1496 31589
rect 982 31445 1046 31509
rect 1072 31445 1136 31509
rect 1162 31445 1226 31509
rect 1252 31445 1316 31509
rect 1342 31445 1406 31509
rect 1432 31445 1496 31509
rect 982 31365 1046 31429
rect 1072 31365 1136 31429
rect 1162 31365 1226 31429
rect 1252 31365 1316 31429
rect 1342 31365 1406 31429
rect 1432 31365 1496 31429
rect 982 31344 1046 31349
rect 1072 31344 1136 31349
rect 1162 31344 1226 31349
rect 1252 31344 1316 31349
rect 1342 31344 1406 31349
rect 1432 31344 1496 31349
rect 982 31285 1046 31344
rect 1072 31285 1136 31344
rect 1162 31285 1226 31344
rect 1252 31285 1316 31344
rect 1342 31285 1406 31344
rect 1432 31285 1496 31344
rect 982 31205 1046 31269
rect 1072 31205 1136 31269
rect 1162 31205 1226 31269
rect 1252 31205 1316 31269
rect 1342 31205 1406 31269
rect 1432 31205 1496 31269
rect 982 31125 1046 31189
rect 1072 31125 1136 31189
rect 1162 31125 1226 31189
rect 1252 31125 1316 31189
rect 1342 31125 1406 31189
rect 1432 31125 1496 31189
rect 982 31045 1046 31109
rect 1072 31045 1136 31109
rect 1162 31045 1226 31109
rect 1252 31045 1316 31109
rect 1342 31045 1406 31109
rect 1432 31045 1496 31109
rect 982 30965 1046 31029
rect 1072 30965 1136 31029
rect 1162 30965 1226 31029
rect 1252 30965 1316 31029
rect 1342 30965 1406 31029
rect 1432 30965 1496 31029
rect 982 30885 1046 30949
rect 1072 30885 1136 30949
rect 1162 30885 1226 30949
rect 1252 30885 1316 30949
rect 1342 30885 1406 30949
rect 1432 30885 1496 30949
rect 982 30805 1046 30869
rect 1072 30805 1136 30869
rect 1162 30805 1226 30869
rect 1252 30805 1316 30869
rect 1342 30805 1406 30869
rect 1432 30805 1496 30869
rect 982 30725 1046 30789
rect 1072 30725 1136 30789
rect 1162 30725 1226 30789
rect 1252 30725 1316 30789
rect 1342 30725 1406 30789
rect 1432 30725 1496 30789
rect 982 30645 1046 30709
rect 1072 30645 1136 30709
rect 1162 30645 1226 30709
rect 1252 30645 1316 30709
rect 1342 30645 1406 30709
rect 1432 30645 1496 30709
rect 982 30565 1046 30629
rect 1072 30565 1136 30629
rect 1162 30565 1226 30629
rect 1252 30565 1316 30629
rect 1342 30565 1406 30629
rect 1432 30565 1496 30629
rect 982 30485 1046 30549
rect 1072 30485 1136 30549
rect 1162 30485 1226 30549
rect 1252 30485 1316 30549
rect 1342 30485 1406 30549
rect 1432 30485 1496 30549
rect 982 30405 1046 30469
rect 1072 30405 1136 30469
rect 1162 30405 1226 30469
rect 1252 30405 1316 30469
rect 1342 30405 1406 30469
rect 1432 30405 1496 30469
rect 982 30325 1046 30389
rect 1072 30325 1136 30389
rect 1162 30325 1226 30389
rect 1252 30325 1316 30389
rect 1342 30325 1406 30389
rect 1432 30325 1496 30389
rect 982 30245 1046 30309
rect 1072 30245 1136 30309
rect 1162 30245 1226 30309
rect 1252 30245 1316 30309
rect 1342 30245 1406 30309
rect 1432 30245 1496 30309
rect 982 30165 1046 30229
rect 1072 30165 1136 30229
rect 1162 30165 1226 30229
rect 1252 30165 1316 30229
rect 1342 30165 1406 30229
rect 1432 30165 1496 30229
rect 982 30085 1046 30149
rect 1072 30085 1136 30149
rect 1162 30085 1226 30149
rect 1252 30085 1316 30149
rect 1342 30085 1406 30149
rect 1432 30085 1496 30149
rect 982 30005 1046 30069
rect 1072 30005 1136 30069
rect 1162 30005 1226 30069
rect 1252 30005 1316 30069
rect 1342 30005 1406 30069
rect 1432 30005 1496 30069
rect 982 29925 1046 29989
rect 1072 29925 1136 29989
rect 1162 29925 1226 29989
rect 1252 29925 1316 29989
rect 1342 29925 1406 29989
rect 1432 29925 1496 29989
rect 982 29845 1046 29909
rect 1072 29845 1136 29909
rect 1162 29845 1226 29909
rect 1252 29845 1316 29909
rect 1342 29845 1406 29909
rect 1432 29845 1496 29909
rect 982 29765 1046 29829
rect 1072 29765 1136 29829
rect 1162 29765 1226 29829
rect 1252 29765 1316 29829
rect 1342 29765 1406 29829
rect 1432 29765 1496 29829
rect 982 29685 1046 29749
rect 1072 29685 1136 29749
rect 1162 29685 1226 29749
rect 1252 29685 1316 29749
rect 1342 29685 1406 29749
rect 1432 29685 1496 29749
rect 982 29605 1046 29669
rect 1072 29605 1136 29669
rect 1162 29605 1226 29669
rect 1252 29605 1316 29669
rect 1342 29605 1406 29669
rect 1432 29605 1496 29669
rect 982 29525 1046 29589
rect 1072 29525 1136 29589
rect 1162 29525 1226 29589
rect 1252 29525 1316 29589
rect 1342 29525 1406 29589
rect 1432 29525 1496 29589
rect 982 29445 1046 29509
rect 1072 29445 1136 29509
rect 1162 29445 1226 29509
rect 1252 29445 1316 29509
rect 1342 29445 1406 29509
rect 1432 29445 1496 29509
rect 982 29365 1046 29429
rect 1072 29365 1136 29429
rect 1162 29365 1226 29429
rect 1252 29365 1316 29429
rect 1342 29365 1406 29429
rect 1432 29365 1496 29429
rect 982 29285 1046 29349
rect 1072 29285 1136 29349
rect 1162 29285 1226 29349
rect 1252 29285 1316 29349
rect 1342 29285 1406 29349
rect 1432 29285 1496 29349
rect 982 29205 1046 29269
rect 1072 29205 1136 29269
rect 1162 29205 1226 29269
rect 1252 29205 1316 29269
rect 1342 29205 1406 29269
rect 1432 29205 1496 29269
rect 982 29125 1046 29189
rect 1072 29125 1136 29189
rect 1162 29125 1226 29189
rect 1252 29125 1316 29189
rect 1342 29125 1406 29189
rect 1432 29125 1496 29189
rect 982 29045 1046 29109
rect 1072 29045 1136 29109
rect 1162 29045 1226 29109
rect 1252 29045 1316 29109
rect 1342 29045 1406 29109
rect 1432 29045 1496 29109
rect 982 28965 1046 29029
rect 1072 28965 1136 29029
rect 1162 28965 1226 29029
rect 1252 28965 1316 29029
rect 1342 28965 1406 29029
rect 1432 28965 1496 29029
rect 982 28885 1046 28949
rect 1072 28885 1136 28949
rect 1162 28885 1226 28949
rect 1252 28885 1316 28949
rect 1342 28885 1406 28949
rect 1432 28885 1496 28949
rect 982 28805 1046 28869
rect 1072 28805 1136 28869
rect 1162 28805 1226 28869
rect 1252 28805 1316 28869
rect 1342 28805 1406 28869
rect 1432 28805 1496 28869
rect 982 28725 1046 28789
rect 1072 28725 1136 28789
rect 1162 28725 1226 28789
rect 1252 28725 1316 28789
rect 1342 28725 1406 28789
rect 1432 28725 1496 28789
rect 982 28645 1046 28709
rect 1072 28645 1136 28709
rect 1162 28645 1226 28709
rect 1252 28645 1316 28709
rect 1342 28645 1406 28709
rect 1432 28645 1496 28709
rect 982 28565 1046 28629
rect 1072 28565 1136 28629
rect 1162 28565 1226 28629
rect 1252 28565 1316 28629
rect 1342 28565 1406 28629
rect 1432 28565 1496 28629
rect 982 28485 1046 28549
rect 1072 28485 1136 28549
rect 1162 28485 1226 28549
rect 1252 28485 1316 28549
rect 1342 28485 1406 28549
rect 1432 28485 1496 28549
rect 982 28405 1046 28469
rect 1072 28405 1136 28469
rect 1162 28405 1226 28469
rect 1252 28405 1316 28469
rect 1342 28405 1406 28469
rect 1432 28405 1496 28469
rect 982 28325 1046 28389
rect 1072 28325 1136 28389
rect 1162 28325 1226 28389
rect 1252 28325 1316 28389
rect 1342 28325 1406 28389
rect 1432 28325 1496 28389
rect 982 28245 1046 28309
rect 1072 28245 1136 28309
rect 1162 28245 1226 28309
rect 1252 28245 1316 28309
rect 1342 28245 1406 28309
rect 1432 28245 1496 28309
rect 982 28165 1046 28229
rect 1072 28165 1136 28229
rect 1162 28165 1226 28229
rect 1252 28165 1316 28229
rect 1342 28165 1406 28229
rect 1432 28165 1496 28229
rect 982 28085 1046 28149
rect 1072 28085 1136 28149
rect 1162 28085 1226 28149
rect 1252 28085 1316 28149
rect 1342 28085 1406 28149
rect 1432 28085 1496 28149
rect 982 28005 1046 28069
rect 1072 28005 1136 28069
rect 1162 28005 1226 28069
rect 1252 28005 1316 28069
rect 1342 28005 1406 28069
rect 1432 28005 1496 28069
rect 982 27925 1046 27989
rect 1072 27925 1136 27989
rect 1162 27925 1226 27989
rect 1252 27925 1316 27989
rect 1342 27925 1406 27989
rect 1432 27925 1496 27989
rect 982 27845 1046 27909
rect 1072 27845 1136 27909
rect 1162 27845 1226 27909
rect 1252 27845 1316 27909
rect 1342 27845 1406 27909
rect 1432 27845 1496 27909
rect 982 27765 1046 27829
rect 1072 27765 1136 27829
rect 1162 27765 1226 27829
rect 1252 27765 1316 27829
rect 1342 27765 1406 27829
rect 1432 27765 1496 27829
rect 982 27685 1046 27749
rect 1072 27685 1136 27749
rect 1162 27685 1226 27749
rect 1252 27685 1316 27749
rect 1342 27685 1406 27749
rect 1432 27685 1496 27749
rect 982 27605 1046 27669
rect 1072 27605 1136 27669
rect 1162 27605 1226 27669
rect 1252 27605 1316 27669
rect 1342 27605 1406 27669
rect 1432 27605 1496 27669
rect 982 27525 1046 27589
rect 1072 27525 1136 27589
rect 1162 27525 1226 27589
rect 1252 27525 1316 27589
rect 1342 27525 1406 27589
rect 1432 27525 1496 27589
rect 982 27445 1046 27509
rect 1072 27445 1136 27509
rect 1162 27445 1226 27509
rect 1252 27445 1316 27509
rect 1342 27445 1406 27509
rect 1432 27445 1496 27509
rect 982 27365 1046 27429
rect 1072 27365 1136 27429
rect 1162 27365 1226 27429
rect 1252 27365 1316 27429
rect 1342 27365 1406 27429
rect 1432 27365 1496 27429
rect 982 27285 1046 27349
rect 1072 27285 1136 27349
rect 1162 27285 1226 27349
rect 1252 27285 1316 27349
rect 1342 27285 1406 27349
rect 1432 27285 1496 27349
rect 982 27205 1046 27269
rect 1072 27205 1136 27269
rect 1162 27205 1226 27269
rect 1252 27205 1316 27269
rect 1342 27205 1406 27269
rect 1432 27205 1496 27269
rect 982 27125 1046 27189
rect 1072 27125 1136 27189
rect 1162 27125 1226 27189
rect 1252 27125 1316 27189
rect 1342 27125 1406 27189
rect 1432 27125 1496 27189
rect 982 27045 1046 27109
rect 1072 27045 1136 27109
rect 1162 27045 1226 27109
rect 1252 27045 1316 27109
rect 1342 27045 1406 27109
rect 1432 27045 1496 27109
rect 982 26965 1046 27029
rect 1072 26965 1136 27029
rect 1162 26965 1226 27029
rect 1252 26965 1316 27029
rect 1342 26965 1406 27029
rect 1432 26965 1496 27029
rect 982 26885 1046 26949
rect 1072 26885 1136 26949
rect 1162 26885 1226 26949
rect 1252 26885 1316 26949
rect 1342 26885 1406 26949
rect 1432 26885 1496 26949
rect 982 26805 1046 26869
rect 1072 26805 1136 26869
rect 1162 26805 1226 26869
rect 1252 26805 1316 26869
rect 1342 26805 1406 26869
rect 1432 26805 1496 26869
rect 982 26725 1046 26789
rect 1072 26725 1136 26789
rect 1162 26725 1226 26789
rect 1252 26725 1316 26789
rect 1342 26725 1406 26789
rect 1432 26725 1496 26789
rect 982 26645 1046 26709
rect 1072 26645 1136 26709
rect 1162 26645 1226 26709
rect 1252 26645 1316 26709
rect 1342 26645 1406 26709
rect 1432 26645 1496 26709
rect 982 26565 1046 26629
rect 1072 26565 1136 26629
rect 1162 26565 1226 26629
rect 1252 26565 1316 26629
rect 1342 26565 1406 26629
rect 1432 26565 1496 26629
rect 982 26485 1046 26549
rect 1072 26485 1136 26549
rect 1162 26485 1226 26549
rect 1252 26485 1316 26549
rect 1342 26485 1406 26549
rect 1432 26485 1496 26549
rect 982 26405 1046 26469
rect 1072 26405 1136 26469
rect 1162 26405 1226 26469
rect 1252 26405 1316 26469
rect 1342 26405 1406 26469
rect 1432 26405 1496 26469
rect 982 26325 1046 26389
rect 1072 26325 1136 26389
rect 1162 26325 1226 26389
rect 1252 26325 1316 26389
rect 1342 26325 1406 26389
rect 1432 26325 1496 26389
rect 982 26245 1046 26309
rect 1072 26245 1136 26309
rect 1162 26245 1226 26309
rect 1252 26245 1316 26309
rect 1342 26245 1406 26309
rect 1432 26245 1496 26309
rect 982 26165 1046 26229
rect 1072 26165 1136 26229
rect 1162 26165 1226 26229
rect 1252 26165 1316 26229
rect 1342 26165 1406 26229
rect 1432 26165 1496 26229
rect 982 26085 1046 26149
rect 1072 26085 1136 26149
rect 1162 26085 1226 26149
rect 1252 26085 1316 26149
rect 1342 26085 1406 26149
rect 1432 26085 1496 26149
rect 982 26005 1046 26069
rect 1072 26005 1136 26069
rect 1162 26005 1226 26069
rect 1252 26005 1316 26069
rect 1342 26005 1406 26069
rect 1432 26005 1496 26069
rect 982 25925 1046 25989
rect 1072 25925 1136 25989
rect 1162 25925 1226 25989
rect 1252 25925 1316 25989
rect 1342 25925 1406 25989
rect 1432 25925 1496 25989
rect 982 25845 1046 25909
rect 1072 25845 1136 25909
rect 1162 25845 1226 25909
rect 1252 25845 1316 25909
rect 1342 25845 1406 25909
rect 1432 25845 1496 25909
rect 982 25765 1046 25829
rect 1072 25765 1136 25829
rect 1162 25765 1226 25829
rect 1252 25765 1316 25829
rect 1342 25765 1406 25829
rect 1432 25765 1496 25829
rect 982 25685 1046 25749
rect 1072 25685 1136 25749
rect 1162 25685 1226 25749
rect 1252 25685 1316 25749
rect 1342 25685 1406 25749
rect 1432 25685 1496 25749
rect 982 25605 1046 25669
rect 1072 25605 1136 25669
rect 1162 25605 1226 25669
rect 1252 25605 1316 25669
rect 1342 25605 1406 25669
rect 1432 25605 1496 25669
rect 982 25525 1046 25589
rect 1072 25525 1136 25589
rect 1162 25525 1226 25589
rect 1252 25525 1316 25589
rect 1342 25525 1406 25589
rect 1432 25525 1496 25589
rect 982 25445 1046 25509
rect 1072 25445 1136 25509
rect 1162 25445 1226 25509
rect 1252 25445 1316 25509
rect 1342 25445 1406 25509
rect 1432 25445 1496 25509
rect 982 25365 1046 25429
rect 1072 25365 1136 25429
rect 1162 25365 1226 25429
rect 1252 25365 1316 25429
rect 1342 25365 1406 25429
rect 1432 25365 1496 25429
rect 982 25285 1046 25349
rect 1072 25285 1136 25349
rect 1162 25285 1226 25349
rect 1252 25285 1316 25349
rect 1342 25285 1406 25349
rect 1432 25285 1496 25349
rect 982 25205 1046 25269
rect 1072 25205 1136 25269
rect 1162 25205 1226 25269
rect 1252 25205 1316 25269
rect 1342 25205 1406 25269
rect 1432 25205 1496 25269
rect 982 25125 1046 25189
rect 1072 25125 1136 25189
rect 1162 25125 1226 25189
rect 1252 25125 1316 25189
rect 1342 25125 1406 25189
rect 1432 25125 1496 25189
rect 982 25045 1046 25109
rect 1072 25045 1136 25109
rect 1162 25045 1226 25109
rect 1252 25045 1316 25109
rect 1342 25045 1406 25109
rect 1432 25045 1496 25109
rect 982 24965 1046 25029
rect 1072 24965 1136 25029
rect 1162 24965 1226 25029
rect 1252 24965 1316 25029
rect 1342 24965 1406 25029
rect 1432 24965 1496 25029
rect 982 24885 1046 24949
rect 1072 24885 1136 24949
rect 1162 24885 1226 24949
rect 1252 24885 1316 24949
rect 1342 24885 1406 24949
rect 1432 24885 1496 24949
rect 982 24805 1046 24869
rect 1072 24805 1136 24869
rect 1162 24805 1226 24869
rect 1252 24805 1316 24869
rect 1342 24805 1406 24869
rect 1432 24805 1496 24869
rect 982 24725 1046 24789
rect 1072 24725 1136 24789
rect 1162 24725 1226 24789
rect 1252 24725 1316 24789
rect 1342 24725 1406 24789
rect 1432 24725 1496 24789
rect 982 24645 1046 24709
rect 1072 24645 1136 24709
rect 1162 24645 1226 24709
rect 1252 24645 1316 24709
rect 1342 24645 1406 24709
rect 1432 24645 1496 24709
rect 982 24565 1046 24629
rect 1072 24565 1136 24629
rect 1162 24565 1226 24629
rect 1252 24565 1316 24629
rect 1342 24565 1406 24629
rect 1432 24565 1496 24629
rect 982 24485 1046 24549
rect 1072 24485 1136 24549
rect 1162 24485 1226 24549
rect 1252 24485 1316 24549
rect 1342 24485 1406 24549
rect 1432 24485 1496 24549
rect 982 24405 1046 24469
rect 1072 24405 1136 24469
rect 1162 24405 1226 24469
rect 1252 24405 1316 24469
rect 1342 24405 1406 24469
rect 1432 24405 1496 24469
rect 982 24325 1046 24389
rect 1072 24325 1136 24389
rect 1162 24325 1226 24389
rect 1252 24325 1316 24389
rect 1342 24325 1406 24389
rect 1432 24325 1496 24389
rect 982 24245 1046 24309
rect 1072 24245 1136 24309
rect 1162 24245 1226 24309
rect 1252 24245 1316 24309
rect 1342 24245 1406 24309
rect 1432 24245 1496 24309
rect 982 24165 1046 24229
rect 1072 24165 1136 24229
rect 1162 24165 1226 24229
rect 1252 24165 1316 24229
rect 1342 24165 1406 24229
rect 1432 24165 1496 24229
rect 982 24085 1046 24149
rect 1072 24085 1136 24149
rect 1162 24085 1226 24149
rect 1252 24085 1316 24149
rect 1342 24085 1406 24149
rect 1432 24085 1496 24149
rect 982 24005 1046 24069
rect 1072 24005 1136 24069
rect 1162 24005 1226 24069
rect 1252 24005 1316 24069
rect 1342 24005 1406 24069
rect 1432 24005 1496 24069
rect 982 23925 1046 23989
rect 1072 23925 1136 23989
rect 1162 23925 1226 23989
rect 1252 23925 1316 23989
rect 1342 23925 1406 23989
rect 1432 23925 1496 23989
rect 982 23845 1046 23909
rect 1072 23845 1136 23909
rect 1162 23845 1226 23909
rect 1252 23845 1316 23909
rect 1342 23845 1406 23909
rect 1432 23845 1496 23909
rect 982 23765 1046 23829
rect 1072 23765 1136 23829
rect 1162 23765 1226 23829
rect 1252 23765 1316 23829
rect 1342 23765 1406 23829
rect 1432 23765 1496 23829
rect 982 23685 1046 23749
rect 1072 23685 1136 23749
rect 1162 23685 1226 23749
rect 1252 23685 1316 23749
rect 1342 23685 1406 23749
rect 1432 23685 1496 23749
rect 982 23605 1046 23669
rect 1072 23605 1136 23669
rect 1162 23605 1226 23669
rect 1252 23605 1316 23669
rect 1342 23605 1406 23669
rect 1432 23605 1496 23669
rect 982 23525 1046 23589
rect 1072 23525 1136 23589
rect 1162 23525 1226 23589
rect 1252 23525 1316 23589
rect 1342 23525 1406 23589
rect 1432 23525 1496 23589
rect 982 23445 1046 23509
rect 1072 23445 1136 23509
rect 1162 23445 1226 23509
rect 1252 23445 1316 23509
rect 1342 23445 1406 23509
rect 1432 23445 1496 23509
rect 982 23365 1046 23429
rect 1072 23365 1136 23429
rect 1162 23365 1226 23429
rect 1252 23365 1316 23429
rect 1342 23365 1406 23429
rect 1432 23365 1496 23429
rect 982 23288 1046 23349
rect 1072 23288 1136 23349
rect 1162 23288 1226 23349
rect 1252 23288 1316 23349
rect 1342 23288 1406 23349
rect 1432 23288 1496 23349
rect 982 23285 1046 23288
rect 1072 23285 1136 23288
rect 1162 23285 1226 23288
rect 1252 23285 1316 23288
rect 1342 23285 1406 23288
rect 1432 23285 1496 23288
rect 982 23204 1046 23268
rect 1072 23204 1136 23268
rect 1162 23204 1226 23268
rect 1252 23204 1316 23268
rect 1342 23204 1406 23268
rect 1432 23204 1496 23268
rect 982 23123 1046 23187
rect 1072 23123 1136 23187
rect 1162 23123 1226 23187
rect 1252 23123 1316 23187
rect 1342 23123 1406 23187
rect 1432 23123 1496 23187
rect 982 23042 1046 23106
rect 1072 23042 1136 23106
rect 1162 23042 1226 23106
rect 1252 23042 1316 23106
rect 1342 23042 1406 23106
rect 1432 23042 1496 23106
rect 982 22961 1046 23025
rect 1072 22961 1136 23025
rect 1162 22961 1226 23025
rect 1252 22961 1316 23025
rect 1342 22961 1406 23025
rect 1432 22961 1496 23025
rect 982 22880 1046 22944
rect 1072 22880 1136 22944
rect 1162 22880 1226 22944
rect 1252 22880 1316 22944
rect 1342 22880 1406 22944
rect 1432 22880 1496 22944
rect 982 22799 1046 22863
rect 1072 22799 1136 22863
rect 1162 22799 1226 22863
rect 1252 22799 1316 22863
rect 1342 22799 1406 22863
rect 1432 22799 1496 22863
rect 982 22718 1046 22782
rect 1072 22718 1136 22782
rect 1162 22718 1226 22782
rect 1252 22718 1316 22782
rect 1342 22718 1406 22782
rect 1432 22718 1496 22782
rect 982 22637 1046 22701
rect 1072 22637 1136 22701
rect 1162 22637 1226 22701
rect 1252 22637 1316 22701
rect 1342 22637 1406 22701
rect 1432 22637 1496 22701
rect 982 22556 1046 22620
rect 1072 22556 1136 22620
rect 1162 22556 1226 22620
rect 1252 22556 1316 22620
rect 1342 22556 1406 22620
rect 1432 22556 1496 22620
rect 982 22475 1046 22539
rect 1072 22475 1136 22539
rect 1162 22475 1226 22539
rect 1252 22475 1316 22539
rect 1342 22475 1406 22539
rect 1432 22475 1496 22539
rect 982 22394 1046 22458
rect 1072 22394 1136 22458
rect 1162 22394 1226 22458
rect 1252 22394 1316 22458
rect 1342 22394 1406 22458
rect 1432 22394 1496 22458
rect 982 22313 1046 22377
rect 1072 22313 1136 22377
rect 1162 22313 1226 22377
rect 1252 22313 1316 22377
rect 1342 22313 1406 22377
rect 1432 22313 1496 22377
rect 982 22232 1046 22296
rect 1072 22232 1136 22296
rect 1162 22232 1226 22296
rect 1252 22232 1316 22296
rect 1342 22232 1406 22296
rect 1432 22232 1496 22296
rect 982 22151 1046 22215
rect 1072 22151 1136 22215
rect 1162 22151 1226 22215
rect 1252 22151 1316 22215
rect 1342 22151 1406 22215
rect 1432 22151 1496 22215
rect 982 22070 1046 22134
rect 1072 22070 1136 22134
rect 1162 22070 1226 22134
rect 1252 22070 1316 22134
rect 1342 22070 1406 22134
rect 1432 22070 1496 22134
rect 982 21989 1046 22053
rect 1072 21989 1136 22053
rect 1162 21989 1226 22053
rect 1252 21989 1316 22053
rect 1342 21989 1406 22053
rect 1432 21989 1496 22053
rect 982 21908 1046 21972
rect 1072 21908 1136 21972
rect 1162 21908 1226 21972
rect 1252 21908 1316 21972
rect 1342 21908 1406 21972
rect 1432 21908 1496 21972
rect 982 21827 1046 21891
rect 1072 21827 1136 21891
rect 1162 21827 1226 21891
rect 1252 21827 1316 21891
rect 1342 21827 1406 21891
rect 1432 21827 1496 21891
rect 982 21746 1046 21810
rect 1072 21746 1136 21810
rect 1162 21746 1226 21810
rect 1252 21746 1316 21810
rect 1342 21746 1406 21810
rect 1432 21746 1496 21810
rect 982 21665 1046 21729
rect 1072 21665 1136 21729
rect 1162 21665 1226 21729
rect 1252 21665 1316 21729
rect 1342 21665 1406 21729
rect 1432 21665 1496 21729
rect 982 21584 1046 21648
rect 1072 21584 1136 21648
rect 1162 21584 1226 21648
rect 1252 21584 1316 21648
rect 1342 21584 1406 21648
rect 1432 21584 1496 21648
rect 982 21503 1046 21567
rect 1072 21503 1136 21567
rect 1162 21503 1226 21567
rect 1252 21503 1316 21567
rect 1342 21503 1406 21567
rect 1432 21503 1496 21567
rect 982 21422 1046 21486
rect 1072 21422 1136 21486
rect 1162 21422 1226 21486
rect 1252 21422 1316 21486
rect 1342 21422 1406 21486
rect 1432 21422 1496 21486
rect 982 21341 1046 21405
rect 1072 21341 1136 21405
rect 1162 21341 1226 21405
rect 1252 21341 1316 21405
rect 1342 21341 1406 21405
rect 1432 21341 1496 21405
rect 982 21260 1046 21324
rect 1072 21260 1136 21324
rect 1162 21260 1226 21324
rect 1252 21260 1316 21324
rect 1342 21260 1406 21324
rect 1432 21260 1496 21324
rect 982 21179 1046 21243
rect 1072 21179 1136 21243
rect 1162 21179 1226 21243
rect 1252 21179 1316 21243
rect 1342 21179 1406 21243
rect 1432 21179 1496 21243
rect 982 21098 1046 21162
rect 1072 21098 1136 21162
rect 1162 21098 1226 21162
rect 1252 21098 1316 21162
rect 1342 21098 1406 21162
rect 1432 21098 1496 21162
rect 982 21017 1046 21081
rect 1072 21017 1136 21081
rect 1162 21017 1226 21081
rect 1252 21017 1316 21081
rect 1342 21017 1406 21081
rect 1432 21017 1496 21081
rect 982 20936 1046 21000
rect 1072 20936 1136 21000
rect 1162 20936 1226 21000
rect 1252 20936 1316 21000
rect 1342 20936 1406 21000
rect 1432 20936 1496 21000
rect 982 20855 1046 20919
rect 1072 20855 1136 20919
rect 1162 20855 1226 20919
rect 1252 20855 1316 20919
rect 1342 20855 1406 20919
rect 1432 20855 1496 20919
rect 1531 20875 1595 20939
rect 1141 20719 1205 20783
rect 1312 20761 1376 20825
rect 1401 20761 1465 20825
rect 1491 20761 1555 20825
rect 1581 20761 1645 20825
rect 1671 20761 1735 20825
rect 1312 20645 1376 20709
rect 1401 20645 1465 20709
rect 1491 20645 1555 20709
rect 1581 20645 1645 20709
rect 1671 20645 1735 20709
rect 1312 20529 1376 20593
rect 1401 20529 1465 20593
rect 1491 20529 1555 20593
rect 1581 20529 1645 20593
rect 1671 20529 1735 20593
rect 1812 20567 1876 20631
rect 1524 20405 1588 20469
rect 1632 20441 1696 20505
rect 1721 20441 1785 20505
rect 1811 20441 1875 20505
rect 1901 20441 1965 20505
rect 1991 20441 2055 20505
rect 1632 20325 1696 20389
rect 1721 20325 1785 20389
rect 1811 20325 1875 20389
rect 1901 20325 1965 20389
rect 1991 20325 2055 20389
rect 1632 20209 1696 20273
rect 1721 20209 1785 20273
rect 1811 20209 1875 20273
rect 1901 20209 1965 20273
rect 1991 20209 2055 20273
rect 2137 20242 2201 20306
rect 13348 33332 13412 33396
rect 13489 33370 13553 33434
rect 13579 33370 13643 33434
rect 13669 33370 13733 33434
rect 13759 33370 13823 33434
rect 13848 33370 13912 33434
rect 13489 33254 13553 33318
rect 13579 33254 13643 33318
rect 13669 33254 13733 33318
rect 13759 33254 13823 33318
rect 13848 33254 13912 33318
rect 13489 33138 13553 33202
rect 13579 33138 13643 33202
rect 13669 33138 13733 33202
rect 13759 33138 13823 33202
rect 13848 33138 13912 33202
rect 13520 33045 13584 33109
rect 13610 33045 13674 33109
rect 13700 33045 13764 33109
rect 13790 33045 13854 33109
rect 13880 33045 13944 33109
rect 13970 33045 14034 33109
rect 13520 32965 13584 33029
rect 13610 32965 13674 33029
rect 13700 32965 13764 33029
rect 13790 32965 13854 33029
rect 13880 32965 13944 33029
rect 13970 32965 14034 33029
rect 13520 32885 13584 32949
rect 13610 32885 13674 32949
rect 13700 32885 13764 32949
rect 13790 32885 13854 32949
rect 13880 32885 13944 32949
rect 13970 32885 14034 32949
rect 13520 32805 13584 32869
rect 13610 32805 13674 32869
rect 13700 32805 13764 32869
rect 13790 32805 13854 32869
rect 13880 32805 13944 32869
rect 13970 32805 14034 32869
rect 13520 32725 13584 32789
rect 13610 32725 13674 32789
rect 13700 32725 13764 32789
rect 13790 32725 13854 32789
rect 13880 32725 13944 32789
rect 13970 32725 14034 32789
rect 13520 32645 13584 32709
rect 13610 32645 13674 32709
rect 13700 32645 13764 32709
rect 13790 32645 13854 32709
rect 13880 32645 13944 32709
rect 13970 32645 14034 32709
rect 13520 32565 13584 32629
rect 13610 32565 13674 32629
rect 13700 32565 13764 32629
rect 13790 32565 13854 32629
rect 13880 32565 13944 32629
rect 13970 32565 14034 32629
rect 13520 32485 13584 32549
rect 13610 32485 13674 32549
rect 13700 32485 13764 32549
rect 13790 32485 13854 32549
rect 13880 32485 13944 32549
rect 13970 32485 14034 32549
rect 13520 32405 13584 32469
rect 13610 32405 13674 32469
rect 13700 32405 13764 32469
rect 13790 32405 13854 32469
rect 13880 32405 13944 32469
rect 13970 32405 14034 32469
rect 13520 32325 13584 32389
rect 13610 32325 13674 32389
rect 13700 32325 13764 32389
rect 13790 32325 13854 32389
rect 13880 32325 13944 32389
rect 13970 32325 14034 32389
rect 13520 32245 13584 32309
rect 13610 32245 13674 32309
rect 13700 32245 13764 32309
rect 13790 32245 13854 32309
rect 13880 32245 13944 32309
rect 13970 32245 14034 32309
rect 13520 32165 13584 32229
rect 13610 32165 13674 32229
rect 13700 32165 13764 32229
rect 13790 32165 13854 32229
rect 13880 32165 13944 32229
rect 13970 32165 14034 32229
rect 13520 32085 13584 32149
rect 13610 32085 13674 32149
rect 13700 32085 13764 32149
rect 13790 32085 13854 32149
rect 13880 32085 13944 32149
rect 13970 32085 14034 32149
rect 13520 32005 13584 32069
rect 13610 32005 13674 32069
rect 13700 32005 13764 32069
rect 13790 32005 13854 32069
rect 13880 32005 13944 32069
rect 13970 32005 14034 32069
rect 13520 31925 13584 31989
rect 13610 31925 13674 31989
rect 13700 31925 13764 31989
rect 13790 31925 13854 31989
rect 13880 31925 13944 31989
rect 13970 31925 14034 31989
rect 13520 31845 13584 31909
rect 13610 31845 13674 31909
rect 13700 31845 13764 31909
rect 13790 31845 13854 31909
rect 13880 31845 13944 31909
rect 13970 31845 14034 31909
rect 13520 31765 13584 31829
rect 13610 31765 13674 31829
rect 13700 31765 13764 31829
rect 13790 31765 13854 31829
rect 13880 31765 13944 31829
rect 13970 31765 14034 31829
rect 13520 31685 13584 31749
rect 13610 31685 13674 31749
rect 13700 31685 13764 31749
rect 13790 31685 13854 31749
rect 13880 31685 13944 31749
rect 13970 31685 14034 31749
rect 13520 31605 13584 31669
rect 13610 31605 13674 31669
rect 13700 31605 13764 31669
rect 13790 31605 13854 31669
rect 13880 31605 13944 31669
rect 13970 31605 14034 31669
rect 13520 31525 13584 31589
rect 13610 31525 13674 31589
rect 13700 31525 13764 31589
rect 13790 31525 13854 31589
rect 13880 31525 13944 31589
rect 13970 31525 14034 31589
rect 13520 31445 13584 31509
rect 13610 31445 13674 31509
rect 13700 31445 13764 31509
rect 13790 31445 13854 31509
rect 13880 31445 13944 31509
rect 13970 31445 14034 31509
rect 13520 31392 13584 31429
rect 13610 31392 13674 31429
rect 13700 31392 13764 31429
rect 13790 31392 13854 31429
rect 13880 31392 13944 31429
rect 13970 31392 14034 31429
rect 13520 31365 13584 31392
rect 13610 31365 13674 31392
rect 13700 31365 13764 31392
rect 13790 31365 13854 31392
rect 13880 31365 13944 31392
rect 13970 31365 14034 31392
rect 13520 31285 13584 31349
rect 13610 31285 13674 31349
rect 13700 31285 13764 31349
rect 13790 31285 13854 31349
rect 13880 31285 13944 31349
rect 13970 31285 14034 31349
rect 13520 31205 13584 31269
rect 13610 31205 13674 31269
rect 13700 31205 13764 31269
rect 13790 31205 13854 31269
rect 13880 31205 13944 31269
rect 13970 31205 14034 31269
rect 13520 31125 13584 31189
rect 13610 31125 13674 31189
rect 13700 31125 13764 31189
rect 13790 31125 13854 31189
rect 13880 31125 13944 31189
rect 13970 31125 14034 31189
rect 13520 31045 13584 31109
rect 13610 31045 13674 31109
rect 13700 31045 13764 31109
rect 13790 31045 13854 31109
rect 13880 31045 13944 31109
rect 13970 31045 14034 31109
rect 13520 30965 13584 31029
rect 13610 30965 13674 31029
rect 13700 30965 13764 31029
rect 13790 30965 13854 31029
rect 13880 30965 13944 31029
rect 13970 30965 14034 31029
rect 13520 30885 13584 30949
rect 13610 30885 13674 30949
rect 13700 30885 13764 30949
rect 13790 30885 13854 30949
rect 13880 30885 13944 30949
rect 13970 30885 14034 30949
rect 13520 30805 13584 30869
rect 13610 30805 13674 30869
rect 13700 30805 13764 30869
rect 13790 30805 13854 30869
rect 13880 30805 13944 30869
rect 13970 30805 14034 30869
rect 13520 30725 13584 30789
rect 13610 30725 13674 30789
rect 13700 30725 13764 30789
rect 13790 30725 13854 30789
rect 13880 30725 13944 30789
rect 13970 30725 14034 30789
rect 13520 30645 13584 30709
rect 13610 30645 13674 30709
rect 13700 30645 13764 30709
rect 13790 30645 13854 30709
rect 13880 30645 13944 30709
rect 13970 30645 14034 30709
rect 13520 30565 13584 30629
rect 13610 30565 13674 30629
rect 13700 30565 13764 30629
rect 13790 30565 13854 30629
rect 13880 30565 13944 30629
rect 13970 30565 14034 30629
rect 13520 30485 13584 30549
rect 13610 30485 13674 30549
rect 13700 30485 13764 30549
rect 13790 30485 13854 30549
rect 13880 30485 13944 30549
rect 13970 30485 14034 30549
rect 13520 30405 13584 30469
rect 13610 30405 13674 30469
rect 13700 30405 13764 30469
rect 13790 30405 13854 30469
rect 13880 30405 13944 30469
rect 13970 30405 14034 30469
rect 13520 30325 13584 30389
rect 13610 30325 13674 30389
rect 13700 30325 13764 30389
rect 13790 30325 13854 30389
rect 13880 30325 13944 30389
rect 13970 30325 14034 30389
rect 13520 30245 13584 30309
rect 13610 30245 13674 30309
rect 13700 30245 13764 30309
rect 13790 30245 13854 30309
rect 13880 30245 13944 30309
rect 13970 30245 14034 30309
rect 13520 30165 13584 30229
rect 13610 30165 13674 30229
rect 13700 30165 13764 30229
rect 13790 30165 13854 30229
rect 13880 30165 13944 30229
rect 13970 30165 14034 30229
rect 13520 30085 13584 30149
rect 13610 30085 13674 30149
rect 13700 30085 13764 30149
rect 13790 30085 13854 30149
rect 13880 30085 13944 30149
rect 13970 30085 14034 30149
rect 13520 30005 13584 30069
rect 13610 30005 13674 30069
rect 13700 30005 13764 30069
rect 13790 30005 13854 30069
rect 13880 30005 13944 30069
rect 13970 30005 14034 30069
rect 13520 29925 13584 29989
rect 13610 29925 13674 29989
rect 13700 29925 13764 29989
rect 13790 29925 13854 29989
rect 13880 29925 13944 29989
rect 13970 29925 14034 29989
rect 13520 29845 13584 29909
rect 13610 29845 13674 29909
rect 13700 29845 13764 29909
rect 13790 29845 13854 29909
rect 13880 29845 13944 29909
rect 13970 29845 14034 29909
rect 13520 29765 13584 29829
rect 13610 29765 13674 29829
rect 13700 29765 13764 29829
rect 13790 29765 13854 29829
rect 13880 29765 13944 29829
rect 13970 29765 14034 29829
rect 13520 29685 13584 29749
rect 13610 29685 13674 29749
rect 13700 29685 13764 29749
rect 13790 29685 13854 29749
rect 13880 29685 13944 29749
rect 13970 29685 14034 29749
rect 13520 29605 13584 29669
rect 13610 29605 13674 29669
rect 13700 29605 13764 29669
rect 13790 29605 13854 29669
rect 13880 29605 13944 29669
rect 13970 29605 14034 29669
rect 13520 29525 13584 29589
rect 13610 29525 13674 29589
rect 13700 29525 13764 29589
rect 13790 29525 13854 29589
rect 13880 29525 13944 29589
rect 13970 29525 14034 29589
rect 13520 29445 13584 29509
rect 13610 29445 13674 29509
rect 13700 29445 13764 29509
rect 13790 29445 13854 29509
rect 13880 29445 13944 29509
rect 13970 29445 14034 29509
rect 13520 29365 13584 29429
rect 13610 29365 13674 29429
rect 13700 29365 13764 29429
rect 13790 29365 13854 29429
rect 13880 29365 13944 29429
rect 13970 29365 14034 29429
rect 13520 29285 13584 29349
rect 13610 29285 13674 29349
rect 13700 29285 13764 29349
rect 13790 29285 13854 29349
rect 13880 29285 13944 29349
rect 13970 29285 14034 29349
rect 13520 29205 13584 29269
rect 13610 29205 13674 29269
rect 13700 29205 13764 29269
rect 13790 29205 13854 29269
rect 13880 29205 13944 29269
rect 13970 29205 14034 29269
rect 13520 29125 13584 29189
rect 13610 29125 13674 29189
rect 13700 29125 13764 29189
rect 13790 29125 13854 29189
rect 13880 29125 13944 29189
rect 13970 29125 14034 29189
rect 13520 29045 13584 29109
rect 13610 29045 13674 29109
rect 13700 29045 13764 29109
rect 13790 29045 13854 29109
rect 13880 29045 13944 29109
rect 13970 29045 14034 29109
rect 13520 28965 13584 29029
rect 13610 28965 13674 29029
rect 13700 28965 13764 29029
rect 13790 28965 13854 29029
rect 13880 28965 13944 29029
rect 13970 28965 14034 29029
rect 13520 28885 13584 28949
rect 13610 28885 13674 28949
rect 13700 28885 13764 28949
rect 13790 28885 13854 28949
rect 13880 28885 13944 28949
rect 13970 28885 14034 28949
rect 13520 28805 13584 28869
rect 13610 28805 13674 28869
rect 13700 28805 13764 28869
rect 13790 28805 13854 28869
rect 13880 28805 13944 28869
rect 13970 28805 14034 28869
rect 13520 28725 13584 28789
rect 13610 28725 13674 28789
rect 13700 28725 13764 28789
rect 13790 28725 13854 28789
rect 13880 28725 13944 28789
rect 13970 28725 14034 28789
rect 13520 28645 13584 28709
rect 13610 28645 13674 28709
rect 13700 28645 13764 28709
rect 13790 28645 13854 28709
rect 13880 28645 13944 28709
rect 13970 28645 14034 28709
rect 13520 28565 13584 28629
rect 13610 28565 13674 28629
rect 13700 28565 13764 28629
rect 13790 28565 13854 28629
rect 13880 28565 13944 28629
rect 13970 28565 14034 28629
rect 13520 28485 13584 28549
rect 13610 28485 13674 28549
rect 13700 28485 13764 28549
rect 13790 28485 13854 28549
rect 13880 28485 13944 28549
rect 13970 28485 14034 28549
rect 13520 28405 13584 28469
rect 13610 28405 13674 28469
rect 13700 28405 13764 28469
rect 13790 28405 13854 28469
rect 13880 28405 13944 28469
rect 13970 28405 14034 28469
rect 13520 28325 13584 28389
rect 13610 28325 13674 28389
rect 13700 28325 13764 28389
rect 13790 28325 13854 28389
rect 13880 28325 13944 28389
rect 13970 28325 14034 28389
rect 13520 28245 13584 28309
rect 13610 28245 13674 28309
rect 13700 28245 13764 28309
rect 13790 28245 13854 28309
rect 13880 28245 13944 28309
rect 13970 28245 14034 28309
rect 13520 28165 13584 28229
rect 13610 28165 13674 28229
rect 13700 28165 13764 28229
rect 13790 28165 13854 28229
rect 13880 28165 13944 28229
rect 13970 28165 14034 28229
rect 13520 28085 13584 28149
rect 13610 28085 13674 28149
rect 13700 28085 13764 28149
rect 13790 28085 13854 28149
rect 13880 28085 13944 28149
rect 13970 28085 14034 28149
rect 13520 28005 13584 28069
rect 13610 28005 13674 28069
rect 13700 28005 13764 28069
rect 13790 28005 13854 28069
rect 13880 28005 13944 28069
rect 13970 28005 14034 28069
rect 13520 27925 13584 27989
rect 13610 27925 13674 27989
rect 13700 27925 13764 27989
rect 13790 27925 13854 27989
rect 13880 27925 13944 27989
rect 13970 27925 14034 27989
rect 13520 27845 13584 27909
rect 13610 27845 13674 27909
rect 13700 27845 13764 27909
rect 13790 27845 13854 27909
rect 13880 27845 13944 27909
rect 13970 27845 14034 27909
rect 13520 27765 13584 27829
rect 13610 27765 13674 27829
rect 13700 27765 13764 27829
rect 13790 27765 13854 27829
rect 13880 27765 13944 27829
rect 13970 27765 14034 27829
rect 13520 27685 13584 27749
rect 13610 27685 13674 27749
rect 13700 27685 13764 27749
rect 13790 27685 13854 27749
rect 13880 27685 13944 27749
rect 13970 27685 14034 27749
rect 13520 27605 13584 27669
rect 13610 27605 13674 27669
rect 13700 27605 13764 27669
rect 13790 27605 13854 27669
rect 13880 27605 13944 27669
rect 13970 27605 14034 27669
rect 13520 27525 13584 27589
rect 13610 27525 13674 27589
rect 13700 27525 13764 27589
rect 13790 27525 13854 27589
rect 13880 27525 13944 27589
rect 13970 27525 14034 27589
rect 13520 27445 13584 27509
rect 13610 27445 13674 27509
rect 13700 27445 13764 27509
rect 13790 27445 13854 27509
rect 13880 27445 13944 27509
rect 13970 27445 14034 27509
rect 13520 27365 13584 27429
rect 13610 27365 13674 27429
rect 13700 27365 13764 27429
rect 13790 27365 13854 27429
rect 13880 27365 13944 27429
rect 13970 27365 14034 27429
rect 13520 27285 13584 27349
rect 13610 27285 13674 27349
rect 13700 27285 13764 27349
rect 13790 27285 13854 27349
rect 13880 27285 13944 27349
rect 13970 27285 14034 27349
rect 13520 27205 13584 27269
rect 13610 27205 13674 27269
rect 13700 27205 13764 27269
rect 13790 27205 13854 27269
rect 13880 27205 13944 27269
rect 13970 27205 14034 27269
rect 13520 27125 13584 27189
rect 13610 27125 13674 27189
rect 13700 27125 13764 27189
rect 13790 27125 13854 27189
rect 13880 27125 13944 27189
rect 13970 27125 14034 27189
rect 13520 27045 13584 27109
rect 13610 27045 13674 27109
rect 13700 27045 13764 27109
rect 13790 27045 13854 27109
rect 13880 27045 13944 27109
rect 13970 27045 14034 27109
rect 13520 26965 13584 27029
rect 13610 26965 13674 27029
rect 13700 26965 13764 27029
rect 13790 26965 13854 27029
rect 13880 26965 13944 27029
rect 13970 26965 14034 27029
rect 13520 26885 13584 26949
rect 13610 26885 13674 26949
rect 13700 26885 13764 26949
rect 13790 26885 13854 26949
rect 13880 26885 13944 26949
rect 13970 26885 14034 26949
rect 13520 26805 13584 26869
rect 13610 26805 13674 26869
rect 13700 26805 13764 26869
rect 13790 26805 13854 26869
rect 13880 26805 13944 26869
rect 13970 26805 14034 26869
rect 13520 26725 13584 26789
rect 13610 26725 13674 26789
rect 13700 26725 13764 26789
rect 13790 26725 13854 26789
rect 13880 26725 13944 26789
rect 13970 26725 14034 26789
rect 13520 26645 13584 26709
rect 13610 26645 13674 26709
rect 13700 26645 13764 26709
rect 13790 26645 13854 26709
rect 13880 26645 13944 26709
rect 13970 26645 14034 26709
rect 13520 26565 13584 26629
rect 13610 26565 13674 26629
rect 13700 26565 13764 26629
rect 13790 26565 13854 26629
rect 13880 26565 13944 26629
rect 13970 26565 14034 26629
rect 13520 26485 13584 26549
rect 13610 26485 13674 26549
rect 13700 26485 13764 26549
rect 13790 26485 13854 26549
rect 13880 26485 13944 26549
rect 13970 26485 14034 26549
rect 13520 26405 13584 26469
rect 13610 26405 13674 26469
rect 13700 26405 13764 26469
rect 13790 26405 13854 26469
rect 13880 26405 13944 26469
rect 13970 26405 14034 26469
rect 13520 26325 13584 26389
rect 13610 26325 13674 26389
rect 13700 26325 13764 26389
rect 13790 26325 13854 26389
rect 13880 26325 13944 26389
rect 13970 26325 14034 26389
rect 13520 26245 13584 26309
rect 13610 26245 13674 26309
rect 13700 26245 13764 26309
rect 13790 26245 13854 26309
rect 13880 26245 13944 26309
rect 13970 26245 14034 26309
rect 13520 26165 13584 26229
rect 13610 26165 13674 26229
rect 13700 26165 13764 26229
rect 13790 26165 13854 26229
rect 13880 26165 13944 26229
rect 13970 26165 14034 26229
rect 13520 26085 13584 26149
rect 13610 26085 13674 26149
rect 13700 26085 13764 26149
rect 13790 26085 13854 26149
rect 13880 26085 13944 26149
rect 13970 26085 14034 26149
rect 13520 26005 13584 26069
rect 13610 26005 13674 26069
rect 13700 26005 13764 26069
rect 13790 26005 13854 26069
rect 13880 26005 13944 26069
rect 13970 26005 14034 26069
rect 13520 25925 13584 25989
rect 13610 25925 13674 25989
rect 13700 25925 13764 25989
rect 13790 25925 13854 25989
rect 13880 25925 13944 25989
rect 13970 25925 14034 25989
rect 13520 25845 13584 25909
rect 13610 25845 13674 25909
rect 13700 25845 13764 25909
rect 13790 25845 13854 25909
rect 13880 25845 13944 25909
rect 13970 25845 14034 25909
rect 13520 25765 13584 25829
rect 13610 25765 13674 25829
rect 13700 25765 13764 25829
rect 13790 25765 13854 25829
rect 13880 25765 13944 25829
rect 13970 25765 14034 25829
rect 13520 25685 13584 25749
rect 13610 25685 13674 25749
rect 13700 25685 13764 25749
rect 13790 25685 13854 25749
rect 13880 25685 13944 25749
rect 13970 25685 14034 25749
rect 13520 25605 13584 25669
rect 13610 25605 13674 25669
rect 13700 25605 13764 25669
rect 13790 25605 13854 25669
rect 13880 25605 13944 25669
rect 13970 25605 14034 25669
rect 13520 25525 13584 25589
rect 13610 25525 13674 25589
rect 13700 25525 13764 25589
rect 13790 25525 13854 25589
rect 13880 25525 13944 25589
rect 13970 25525 14034 25589
rect 13520 25445 13584 25509
rect 13610 25445 13674 25509
rect 13700 25445 13764 25509
rect 13790 25445 13854 25509
rect 13880 25445 13944 25509
rect 13970 25445 14034 25509
rect 13520 25365 13584 25429
rect 13610 25365 13674 25429
rect 13700 25365 13764 25429
rect 13790 25365 13854 25429
rect 13880 25365 13944 25429
rect 13970 25365 14034 25429
rect 13520 25285 13584 25349
rect 13610 25285 13674 25349
rect 13700 25285 13764 25349
rect 13790 25285 13854 25349
rect 13880 25285 13944 25349
rect 13970 25285 14034 25349
rect 13520 25205 13584 25269
rect 13610 25205 13674 25269
rect 13700 25205 13764 25269
rect 13790 25205 13854 25269
rect 13880 25205 13944 25269
rect 13970 25205 14034 25269
rect 13520 25125 13584 25189
rect 13610 25125 13674 25189
rect 13700 25125 13764 25189
rect 13790 25125 13854 25189
rect 13880 25125 13944 25189
rect 13970 25125 14034 25189
rect 13520 25045 13584 25109
rect 13610 25045 13674 25109
rect 13700 25045 13764 25109
rect 13790 25045 13854 25109
rect 13880 25045 13944 25109
rect 13970 25045 14034 25109
rect 13520 24965 13584 25029
rect 13610 24965 13674 25029
rect 13700 24965 13764 25029
rect 13790 24965 13854 25029
rect 13880 24965 13944 25029
rect 13970 24965 14034 25029
rect 13520 24885 13584 24949
rect 13610 24885 13674 24949
rect 13700 24885 13764 24949
rect 13790 24885 13854 24949
rect 13880 24885 13944 24949
rect 13970 24885 14034 24949
rect 13520 24805 13584 24869
rect 13610 24805 13674 24869
rect 13700 24805 13764 24869
rect 13790 24805 13854 24869
rect 13880 24805 13944 24869
rect 13970 24805 14034 24869
rect 13520 24725 13584 24789
rect 13610 24725 13674 24789
rect 13700 24725 13764 24789
rect 13790 24725 13854 24789
rect 13880 24725 13944 24789
rect 13970 24725 14034 24789
rect 13520 24645 13584 24709
rect 13610 24645 13674 24709
rect 13700 24645 13764 24709
rect 13790 24645 13854 24709
rect 13880 24645 13944 24709
rect 13970 24645 14034 24709
rect 13520 24565 13584 24629
rect 13610 24565 13674 24629
rect 13700 24565 13764 24629
rect 13790 24565 13854 24629
rect 13880 24565 13944 24629
rect 13970 24565 14034 24629
rect 13520 24485 13584 24549
rect 13610 24485 13674 24549
rect 13700 24485 13764 24549
rect 13790 24485 13854 24549
rect 13880 24485 13944 24549
rect 13970 24485 14034 24549
rect 13520 24405 13584 24469
rect 13610 24405 13674 24469
rect 13700 24405 13764 24469
rect 13790 24405 13854 24469
rect 13880 24405 13944 24469
rect 13970 24405 14034 24469
rect 13520 24325 13584 24389
rect 13610 24325 13674 24389
rect 13700 24325 13764 24389
rect 13790 24325 13854 24389
rect 13880 24325 13944 24389
rect 13970 24325 14034 24389
rect 13520 24245 13584 24309
rect 13610 24245 13674 24309
rect 13700 24245 13764 24309
rect 13790 24245 13854 24309
rect 13880 24245 13944 24309
rect 13970 24245 14034 24309
rect 13520 24165 13584 24229
rect 13610 24165 13674 24229
rect 13700 24165 13764 24229
rect 13790 24165 13854 24229
rect 13880 24165 13944 24229
rect 13970 24165 14034 24229
rect 13520 24085 13584 24149
rect 13610 24085 13674 24149
rect 13700 24085 13764 24149
rect 13790 24085 13854 24149
rect 13880 24085 13944 24149
rect 13970 24085 14034 24149
rect 13520 24005 13584 24069
rect 13610 24005 13674 24069
rect 13700 24005 13764 24069
rect 13790 24005 13854 24069
rect 13880 24005 13944 24069
rect 13970 24005 14034 24069
rect 13520 23925 13584 23989
rect 13610 23925 13674 23989
rect 13700 23925 13764 23989
rect 13790 23925 13854 23989
rect 13880 23925 13944 23989
rect 13970 23925 14034 23989
rect 13520 23845 13584 23909
rect 13610 23845 13674 23909
rect 13700 23845 13764 23909
rect 13790 23845 13854 23909
rect 13880 23845 13944 23909
rect 13970 23845 14034 23909
rect 13520 23765 13584 23829
rect 13610 23765 13674 23829
rect 13700 23765 13764 23829
rect 13790 23765 13854 23829
rect 13880 23765 13944 23829
rect 13970 23765 14034 23829
rect 13520 23685 13584 23749
rect 13610 23685 13674 23749
rect 13700 23685 13764 23749
rect 13790 23685 13854 23749
rect 13880 23685 13944 23749
rect 13970 23685 14034 23749
rect 13520 23605 13584 23669
rect 13610 23605 13674 23669
rect 13700 23605 13764 23669
rect 13790 23605 13854 23669
rect 13880 23605 13944 23669
rect 13970 23605 14034 23669
rect 13520 23525 13584 23589
rect 13610 23525 13674 23589
rect 13700 23525 13764 23589
rect 13790 23525 13854 23589
rect 13880 23525 13944 23589
rect 13970 23525 14034 23589
rect 13520 23445 13584 23509
rect 13610 23445 13674 23509
rect 13700 23445 13764 23509
rect 13790 23445 13854 23509
rect 13880 23445 13944 23509
rect 13970 23445 14034 23509
rect 13520 23365 13584 23429
rect 13610 23365 13674 23429
rect 13700 23365 13764 23429
rect 13790 23365 13854 23429
rect 13880 23365 13944 23429
rect 13970 23365 14034 23429
rect 13520 23336 13584 23349
rect 13610 23336 13674 23349
rect 13700 23336 13764 23349
rect 13790 23336 13854 23349
rect 13880 23336 13944 23349
rect 13970 23336 14034 23349
rect 13520 23285 13584 23336
rect 13610 23285 13674 23336
rect 13700 23285 13764 23336
rect 13790 23285 13854 23336
rect 13880 23285 13944 23336
rect 13970 23285 14034 23336
rect 13520 23204 13584 23268
rect 13610 23204 13674 23268
rect 13700 23204 13764 23268
rect 13790 23204 13854 23268
rect 13880 23204 13944 23268
rect 13970 23204 14034 23268
rect 13520 23123 13584 23187
rect 13610 23123 13674 23187
rect 13700 23123 13764 23187
rect 13790 23123 13854 23187
rect 13880 23123 13944 23187
rect 13970 23123 14034 23187
rect 13520 23042 13584 23106
rect 13610 23042 13674 23106
rect 13700 23042 13764 23106
rect 13790 23042 13854 23106
rect 13880 23042 13944 23106
rect 13970 23042 14034 23106
rect 13520 22961 13584 23025
rect 13610 22961 13674 23025
rect 13700 22961 13764 23025
rect 13790 22961 13854 23025
rect 13880 22961 13944 23025
rect 13970 22961 14034 23025
rect 13520 22880 13584 22944
rect 13610 22880 13674 22944
rect 13700 22880 13764 22944
rect 13790 22880 13854 22944
rect 13880 22880 13944 22944
rect 13970 22880 14034 22944
rect 13520 22799 13584 22863
rect 13610 22799 13674 22863
rect 13700 22799 13764 22863
rect 13790 22799 13854 22863
rect 13880 22799 13944 22863
rect 13970 22799 14034 22863
rect 13520 22718 13584 22782
rect 13610 22718 13674 22782
rect 13700 22718 13764 22782
rect 13790 22718 13854 22782
rect 13880 22718 13944 22782
rect 13970 22718 14034 22782
rect 13520 22637 13584 22701
rect 13610 22637 13674 22701
rect 13700 22637 13764 22701
rect 13790 22637 13854 22701
rect 13880 22637 13944 22701
rect 13970 22637 14034 22701
rect 13520 22556 13584 22620
rect 13610 22556 13674 22620
rect 13700 22556 13764 22620
rect 13790 22556 13854 22620
rect 13880 22556 13944 22620
rect 13970 22556 14034 22620
rect 13520 22475 13584 22539
rect 13610 22475 13674 22539
rect 13700 22475 13764 22539
rect 13790 22475 13854 22539
rect 13880 22475 13944 22539
rect 13970 22475 14034 22539
rect 13520 22394 13584 22458
rect 13610 22394 13674 22458
rect 13700 22394 13764 22458
rect 13790 22394 13854 22458
rect 13880 22394 13944 22458
rect 13970 22394 14034 22458
rect 13520 22313 13584 22377
rect 13610 22313 13674 22377
rect 13700 22313 13764 22377
rect 13790 22313 13854 22377
rect 13880 22313 13944 22377
rect 13970 22313 14034 22377
rect 13520 22232 13584 22296
rect 13610 22232 13674 22296
rect 13700 22232 13764 22296
rect 13790 22232 13854 22296
rect 13880 22232 13944 22296
rect 13970 22232 14034 22296
rect 13520 22151 13584 22215
rect 13610 22151 13674 22215
rect 13700 22151 13764 22215
rect 13790 22151 13854 22215
rect 13880 22151 13944 22215
rect 13970 22151 14034 22215
rect 13520 22070 13584 22134
rect 13610 22070 13674 22134
rect 13700 22070 13764 22134
rect 13790 22070 13854 22134
rect 13880 22070 13944 22134
rect 13970 22070 14034 22134
rect 13520 21989 13584 22053
rect 13610 21989 13674 22053
rect 13700 21989 13764 22053
rect 13790 21989 13854 22053
rect 13880 21989 13944 22053
rect 13970 21989 14034 22053
rect 13520 21908 13584 21972
rect 13610 21908 13674 21972
rect 13700 21908 13764 21972
rect 13790 21908 13854 21972
rect 13880 21908 13944 21972
rect 13970 21908 14034 21972
rect 13520 21827 13584 21891
rect 13610 21827 13674 21891
rect 13700 21827 13764 21891
rect 13790 21827 13854 21891
rect 13880 21827 13944 21891
rect 13970 21827 14034 21891
rect 13520 21746 13584 21810
rect 13610 21746 13674 21810
rect 13700 21746 13764 21810
rect 13790 21746 13854 21810
rect 13880 21746 13944 21810
rect 13970 21746 14034 21810
rect 13520 21665 13584 21729
rect 13610 21665 13674 21729
rect 13700 21665 13764 21729
rect 13790 21665 13854 21729
rect 13880 21665 13944 21729
rect 13970 21665 14034 21729
rect 13520 21584 13584 21648
rect 13610 21584 13674 21648
rect 13700 21584 13764 21648
rect 13790 21584 13854 21648
rect 13880 21584 13944 21648
rect 13970 21584 14034 21648
rect 13520 21503 13584 21567
rect 13610 21503 13674 21567
rect 13700 21503 13764 21567
rect 13790 21503 13854 21567
rect 13880 21503 13944 21567
rect 13970 21503 14034 21567
rect 13520 21422 13584 21486
rect 13610 21422 13674 21486
rect 13700 21422 13764 21486
rect 13790 21422 13854 21486
rect 13880 21422 13944 21486
rect 13970 21422 14034 21486
rect 13520 21341 13584 21405
rect 13610 21341 13674 21405
rect 13700 21341 13764 21405
rect 13790 21341 13854 21405
rect 13880 21341 13944 21405
rect 13970 21341 14034 21405
rect 13520 21260 13584 21324
rect 13610 21260 13674 21324
rect 13700 21260 13764 21324
rect 13790 21260 13854 21324
rect 13880 21260 13944 21324
rect 13970 21260 14034 21324
rect 13520 21179 13584 21243
rect 13610 21179 13674 21243
rect 13700 21179 13764 21243
rect 13790 21179 13854 21243
rect 13880 21179 13944 21243
rect 13970 21179 14034 21243
rect 13520 21098 13584 21162
rect 13610 21098 13674 21162
rect 13700 21098 13764 21162
rect 13790 21098 13854 21162
rect 13880 21098 13944 21162
rect 13970 21098 14034 21162
rect 13520 21017 13584 21081
rect 13610 21017 13674 21081
rect 13700 21017 13764 21081
rect 13790 21017 13854 21081
rect 13880 21017 13944 21081
rect 13970 21017 14034 21081
rect 13421 20875 13485 20939
rect 13520 20936 13584 21000
rect 13610 20936 13674 21000
rect 13700 20936 13764 21000
rect 13790 20936 13854 21000
rect 13880 20936 13944 21000
rect 13970 20936 14034 21000
rect 13520 20855 13584 20919
rect 13610 20855 13674 20919
rect 13700 20855 13764 20919
rect 13790 20855 13854 20919
rect 13880 20855 13944 20919
rect 13970 20855 14034 20919
rect 13281 20761 13345 20825
rect 13371 20761 13435 20825
rect 13461 20761 13525 20825
rect 13551 20761 13615 20825
rect 13640 20761 13704 20825
rect 13749 20759 13813 20823
rect 13851 20752 13915 20816
rect 13281 20645 13345 20709
rect 13371 20645 13435 20709
rect 13461 20645 13525 20709
rect 13551 20645 13615 20709
rect 13640 20645 13704 20709
rect 13749 20648 13813 20712
rect 13140 20567 13204 20631
rect 13281 20529 13345 20593
rect 13371 20529 13435 20593
rect 13461 20529 13525 20593
rect 13551 20529 13615 20593
rect 13640 20529 13704 20593
rect 12961 20441 13025 20505
rect 13051 20441 13115 20505
rect 13141 20441 13205 20505
rect 13231 20441 13295 20505
rect 13320 20441 13384 20505
rect 13428 20405 13492 20469
rect 12961 20325 13025 20389
rect 13051 20325 13115 20389
rect 13141 20325 13205 20389
rect 13231 20325 13295 20389
rect 13320 20325 13384 20389
rect 1852 20077 1916 20141
rect 1956 20117 2020 20181
rect 2045 20117 2109 20181
rect 2135 20117 2199 20181
rect 2225 20117 2289 20181
rect 2315 20117 2379 20181
rect 12815 20242 12879 20306
rect 12961 20209 13025 20273
rect 13051 20209 13115 20273
rect 13141 20209 13205 20273
rect 13231 20209 13295 20273
rect 13320 20209 13384 20273
rect 12637 20117 12701 20181
rect 12727 20117 12791 20181
rect 12817 20117 12881 20181
rect 12907 20117 12971 20181
rect 12996 20117 13060 20181
rect 13100 20077 13164 20141
rect 1956 20001 2020 20065
rect 2045 20001 2109 20065
rect 2135 20001 2199 20065
rect 2225 20001 2289 20065
rect 2315 20001 2379 20065
rect 2456 20006 2520 20070
rect 2571 20006 2635 20070
rect 2686 20006 2750 20070
rect 2802 20006 2866 20070
rect 12150 20006 12214 20070
rect 12266 20006 12330 20070
rect 12381 20006 12445 20070
rect 12496 20006 12560 20070
rect 1956 19885 2020 19949
rect 2045 19885 2109 19949
rect 2135 19885 2199 19949
rect 2225 19885 2289 19949
rect 2315 19885 2379 19949
rect 2456 19886 2520 19950
rect 2571 19886 2635 19950
rect 2686 19886 2750 19950
rect 2802 19886 2866 19950
rect 2906 19891 2970 19955
rect 12637 20001 12701 20065
rect 12727 20001 12791 20065
rect 12817 20001 12881 20065
rect 12907 20001 12971 20065
rect 12996 20001 13060 20065
rect 12046 19891 12110 19955
rect 12150 19886 12214 19950
rect 12266 19886 12330 19950
rect 12381 19886 12445 19950
rect 12496 19886 12560 19950
rect 12637 19885 12701 19949
rect 12727 19885 12791 19949
rect 12817 19885 12881 19949
rect 12907 19885 12971 19949
rect 12996 19885 13060 19949
rect 2193 19736 2257 19800
rect 2293 19780 2357 19844
rect 2377 19780 2441 19844
rect 2461 19780 2525 19844
rect 2545 19780 2609 19844
rect 2629 19780 2693 19844
rect 2713 19780 2777 19844
rect 2797 19780 2861 19844
rect 2881 19780 2945 19844
rect 2965 19780 3029 19844
rect 3049 19780 3113 19844
rect 2293 19664 2357 19728
rect 2377 19664 2441 19728
rect 2461 19664 2525 19728
rect 2545 19664 2609 19728
rect 2629 19664 2693 19728
rect 2713 19664 2777 19728
rect 2797 19664 2861 19728
rect 2881 19664 2945 19728
rect 2965 19664 3029 19728
rect 3049 19664 3113 19728
rect 11903 19780 11967 19844
rect 11987 19780 12051 19844
rect 12071 19780 12135 19844
rect 12155 19780 12219 19844
rect 12239 19780 12303 19844
rect 12323 19780 12387 19844
rect 12407 19780 12471 19844
rect 12491 19780 12555 19844
rect 12575 19780 12639 19844
rect 12659 19780 12723 19844
rect 12759 19736 12823 19800
rect 3153 19643 3217 19707
rect 2293 19548 2357 19612
rect 2377 19548 2441 19612
rect 2461 19548 2525 19612
rect 2545 19548 2609 19612
rect 2629 19548 2693 19612
rect 2713 19548 2777 19612
rect 2797 19548 2861 19612
rect 2881 19548 2945 19612
rect 2965 19548 3029 19612
rect 3049 19548 3113 19612
rect 3153 19550 3217 19614
rect 11799 19643 11863 19707
rect 11903 19664 11967 19728
rect 11987 19664 12051 19728
rect 12071 19664 12135 19728
rect 12155 19664 12219 19728
rect 12239 19664 12303 19728
rect 12323 19664 12387 19728
rect 12407 19664 12471 19728
rect 12491 19664 12555 19728
rect 12575 19664 12639 19728
rect 12659 19664 12723 19728
rect 11799 19550 11863 19614
rect 11903 19548 11967 19612
rect 11987 19548 12051 19612
rect 12071 19548 12135 19612
rect 12155 19548 12219 19612
rect 12239 19548 12303 19612
rect 12323 19548 12387 19612
rect 12407 19548 12471 19612
rect 12491 19548 12555 19612
rect 12575 19548 12639 19612
rect 12659 19548 12723 19612
rect 4938 17311 4942 18895
rect 4942 17311 7238 18895
rect 7238 17311 7242 18895
rect 7738 17311 7742 18895
rect 7742 17311 10038 18895
rect 10038 17311 10042 18895
rect 5099 17214 7243 17218
rect 5099 17078 5103 17214
rect 5103 17078 7239 17214
rect 7239 17078 7243 17214
rect 5099 17074 7243 17078
rect 7735 17214 9879 17218
rect 7735 17078 7739 17214
rect 7739 17078 9875 17214
rect 9875 17078 9879 17214
rect 7735 17074 9879 17078
rect 2423 5241 3607 6025
rect 887 4027 2071 4811
rect 11297 5240 12481 6024
rect 12887 4027 14071 4811
<< metal4 >>
rect 4949 39217 7225 39241
rect 767 36409 1727 37008
rect 4949 35313 4975 39217
rect 7199 35313 7225 39217
rect 4949 35290 7225 35313
rect 7749 39217 10025 39241
rect 7749 35313 7775 39217
rect 9999 35313 10025 39217
rect 13204 36409 14164 37008
rect 7749 35290 10025 35313
rect 2275 34618 2676 34621
rect 2275 34554 2276 34618
rect 2340 34554 2359 34618
rect 2423 34554 2443 34618
rect 2507 34554 2527 34618
rect 2591 34554 2611 34618
rect 2675 34554 2676 34618
rect 2275 34524 2676 34554
rect 2131 34441 2213 34474
rect 2131 34377 2148 34441
rect 2212 34377 2213 34441
rect 2131 34344 2213 34377
rect 2275 34460 2276 34524
rect 2340 34460 2359 34524
rect 2423 34460 2443 34524
rect 2507 34460 2527 34524
rect 2591 34460 2611 34524
rect 2675 34460 2676 34524
rect 2275 34430 2676 34460
rect 2275 34366 2276 34430
rect 2340 34366 2359 34430
rect 2423 34366 2443 34430
rect 2507 34366 2527 34430
rect 2591 34366 2611 34430
rect 2675 34366 2676 34430
rect 2275 34336 2676 34366
rect 2002 34316 2230 34317
rect 2002 34252 2004 34316
rect 2068 34252 2084 34316
rect 2148 34252 2164 34316
rect 2228 34252 2230 34316
rect 2002 34220 2230 34252
rect 1873 34183 1955 34216
rect 1873 34119 1890 34183
rect 1954 34119 1955 34183
rect 2002 34156 2004 34220
rect 2068 34156 2084 34220
rect 2148 34156 2164 34220
rect 2228 34156 2230 34220
rect 2002 34155 2230 34156
rect 2275 34272 2276 34336
rect 2340 34272 2359 34336
rect 2423 34272 2443 34336
rect 2507 34272 2527 34336
rect 2591 34272 2611 34336
rect 2675 34272 2676 34336
rect 2275 34242 2676 34272
rect 2275 34178 2276 34242
rect 2340 34178 2359 34242
rect 2423 34178 2443 34242
rect 2507 34178 2527 34242
rect 2591 34178 2611 34242
rect 2675 34178 2676 34242
rect 1873 34086 1955 34119
rect 2275 34148 2676 34178
rect 2275 34084 2276 34148
rect 2340 34084 2359 34148
rect 2423 34084 2443 34148
rect 2507 34084 2527 34148
rect 2591 34084 2611 34148
rect 2675 34084 2676 34148
rect 2275 34081 2676 34084
rect 12340 34618 12742 34621
rect 12340 34554 12341 34618
rect 12405 34554 12425 34618
rect 12489 34554 12509 34618
rect 12573 34554 12593 34618
rect 12657 34554 12677 34618
rect 12741 34554 12742 34618
rect 12340 34524 12742 34554
rect 12340 34460 12341 34524
rect 12405 34460 12425 34524
rect 12489 34460 12509 34524
rect 12573 34460 12593 34524
rect 12657 34460 12677 34524
rect 12741 34460 12742 34524
rect 12340 34430 12742 34460
rect 12340 34366 12341 34430
rect 12405 34366 12425 34430
rect 12489 34366 12509 34430
rect 12573 34366 12593 34430
rect 12657 34366 12677 34430
rect 12741 34366 12742 34430
rect 12340 34336 12742 34366
rect 12803 34441 12885 34474
rect 12803 34377 12804 34441
rect 12868 34377 12885 34441
rect 12803 34344 12885 34377
rect 12340 34272 12341 34336
rect 12405 34272 12425 34336
rect 12489 34272 12509 34336
rect 12573 34272 12593 34336
rect 12657 34272 12677 34336
rect 12741 34272 12742 34336
rect 12340 34242 12742 34272
rect 12340 34178 12341 34242
rect 12405 34178 12425 34242
rect 12489 34178 12509 34242
rect 12573 34178 12593 34242
rect 12657 34178 12677 34242
rect 12741 34178 12742 34242
rect 12340 34148 12742 34178
rect 12786 34316 13014 34317
rect 12786 34252 12788 34316
rect 12852 34252 12868 34316
rect 12932 34252 12948 34316
rect 13012 34252 13014 34316
rect 12786 34220 13014 34252
rect 12786 34156 12788 34220
rect 12852 34156 12868 34220
rect 12932 34156 12948 34220
rect 13012 34156 13014 34220
rect 12786 34155 13014 34156
rect 13061 34183 13143 34216
rect 12340 34084 12341 34148
rect 12405 34084 12425 34148
rect 12489 34084 12509 34148
rect 12573 34084 12593 34148
rect 12657 34084 12677 34148
rect 12741 34084 12742 34148
rect 13061 34119 13062 34183
rect 13126 34119 13143 34183
rect 13061 34086 13143 34119
rect 12340 34081 12742 34084
rect 1747 34078 2172 34080
rect 1747 34014 1748 34078
rect 1812 34014 1837 34078
rect 1901 34014 1927 34078
rect 1991 34014 2017 34078
rect 2081 34014 2107 34078
rect 2171 34014 2172 34078
rect 12844 34078 13269 34080
rect 1747 33962 2172 34014
rect 1584 33886 1709 33919
rect 1584 33822 1644 33886
rect 1708 33822 1709 33886
rect 1584 33789 1709 33822
rect 1747 33898 1748 33962
rect 1812 33898 1837 33962
rect 1901 33898 1927 33962
rect 1991 33898 2017 33962
rect 2081 33898 2107 33962
rect 2171 33898 2172 33962
rect 2187 34009 2312 34042
rect 2187 33945 2247 34009
rect 2311 33945 2312 34009
rect 2187 33912 2312 33945
rect 12704 34009 12829 34042
rect 12704 33945 12705 34009
rect 12769 33945 12829 34009
rect 12704 33912 12829 33945
rect 12844 34014 12845 34078
rect 12909 34014 12935 34078
rect 12999 34014 13025 34078
rect 13089 34014 13115 34078
rect 13179 34014 13204 34078
rect 13268 34014 13269 34078
rect 12844 33962 13269 34014
rect 1747 33846 2172 33898
rect 1747 33782 1748 33846
rect 1812 33782 1837 33846
rect 1901 33782 1927 33846
rect 1991 33782 2017 33846
rect 2081 33782 2107 33846
rect 2171 33782 2172 33846
rect 1747 33780 2172 33782
rect 12844 33898 12845 33962
rect 12909 33898 12935 33962
rect 12999 33898 13025 33962
rect 13089 33898 13115 33962
rect 13179 33898 13204 33962
rect 13268 33898 13269 33962
rect 12844 33846 13269 33898
rect 12844 33782 12845 33846
rect 12909 33782 12935 33846
rect 12999 33782 13025 33846
rect 13089 33782 13115 33846
rect 13179 33782 13204 33846
rect 13268 33782 13269 33846
rect 13307 33886 13432 33919
rect 13307 33822 13308 33886
rect 13372 33822 13432 33886
rect 13307 33789 13432 33822
rect 12844 33780 13269 33782
rect 1423 33754 1848 33756
rect 13168 33754 13593 33756
rect 1423 33690 1424 33754
rect 1488 33690 1513 33754
rect 1577 33690 1603 33754
rect 1667 33690 1693 33754
rect 1757 33690 1783 33754
rect 1847 33690 1848 33754
rect 1423 33638 1848 33690
rect 1256 33558 1381 33591
rect 1256 33494 1316 33558
rect 1380 33494 1381 33558
rect 1256 33461 1381 33494
rect 1423 33574 1424 33638
rect 1488 33574 1513 33638
rect 1577 33574 1603 33638
rect 1667 33574 1693 33638
rect 1757 33574 1783 33638
rect 1847 33574 1848 33638
rect 1869 33721 1994 33754
rect 1869 33657 1929 33721
rect 1993 33657 1994 33721
rect 1869 33624 1994 33657
rect 13022 33721 13147 33754
rect 13022 33657 13023 33721
rect 13087 33657 13147 33721
rect 13022 33624 13147 33657
rect 13168 33690 13169 33754
rect 13233 33690 13259 33754
rect 13323 33690 13349 33754
rect 13413 33690 13439 33754
rect 13503 33690 13528 33754
rect 13592 33690 13593 33754
rect 13168 33638 13593 33690
rect 1423 33522 1848 33574
rect 1423 33458 1424 33522
rect 1488 33458 1513 33522
rect 1577 33458 1603 33522
rect 1667 33458 1693 33522
rect 1757 33458 1783 33522
rect 1847 33458 1848 33522
rect 1423 33456 1848 33458
rect 13168 33574 13169 33638
rect 13233 33574 13259 33638
rect 13323 33574 13349 33638
rect 13413 33574 13439 33638
rect 13503 33574 13528 33638
rect 13592 33574 13593 33638
rect 13168 33522 13593 33574
rect 13168 33458 13169 33522
rect 13233 33458 13259 33522
rect 13323 33458 13349 33522
rect 13413 33458 13439 33522
rect 13503 33458 13528 33522
rect 13592 33458 13593 33522
rect 13635 33558 13760 33591
rect 13635 33494 13636 33558
rect 13700 33494 13760 33558
rect 13635 33461 13760 33494
rect 13168 33456 13593 33458
rect 1103 33434 1528 33436
rect 1103 33370 1104 33434
rect 1168 33370 1193 33434
rect 1257 33370 1283 33434
rect 1347 33370 1373 33434
rect 1437 33370 1463 33434
rect 1527 33370 1528 33434
rect 13488 33434 13913 33436
rect 1103 33318 1528 33370
rect 1103 33254 1104 33318
rect 1168 33254 1193 33318
rect 1257 33254 1283 33318
rect 1347 33254 1373 33318
rect 1437 33254 1463 33318
rect 1527 33254 1528 33318
rect 1544 33396 1669 33429
rect 1544 33332 1604 33396
rect 1668 33332 1669 33396
rect 1544 33299 1669 33332
rect 13347 33396 13472 33429
rect 13347 33332 13348 33396
rect 13412 33332 13472 33396
rect 13347 33299 13472 33332
rect 13488 33370 13489 33434
rect 13553 33370 13579 33434
rect 13643 33370 13669 33434
rect 13733 33370 13759 33434
rect 13823 33370 13848 33434
rect 13912 33370 13913 33434
rect 13488 33318 13913 33370
rect 1103 33202 1528 33254
rect 1103 33138 1104 33202
rect 1168 33138 1193 33202
rect 1257 33138 1283 33202
rect 1347 33138 1373 33202
rect 1437 33138 1463 33202
rect 1527 33138 1528 33202
rect 1103 33136 1528 33138
rect 13488 33254 13489 33318
rect 13553 33254 13579 33318
rect 13643 33254 13669 33318
rect 13733 33254 13759 33318
rect 13823 33254 13848 33318
rect 13912 33254 13913 33318
rect 13488 33202 13913 33254
rect 13488 33138 13489 33202
rect 13553 33138 13579 33202
rect 13643 33138 13669 33202
rect 13733 33138 13759 33202
rect 13823 33138 13848 33202
rect 13912 33138 13913 33202
rect 13488 33136 13913 33138
rect 977 33109 1501 33110
rect 977 33045 982 33109
rect 1046 33045 1072 33109
rect 1136 33045 1162 33109
rect 1226 33045 1252 33109
rect 1316 33045 1342 33109
rect 1406 33045 1432 33109
rect 1496 33045 1501 33109
rect 977 33029 1501 33045
rect 977 32965 982 33029
rect 1046 32965 1072 33029
rect 1136 32965 1162 33029
rect 1226 32965 1252 33029
rect 1316 32965 1342 33029
rect 1406 32965 1432 33029
rect 1496 32965 1501 33029
rect 977 32949 1501 32965
rect 977 32885 982 32949
rect 1046 32885 1072 32949
rect 1136 32885 1162 32949
rect 1226 32885 1252 32949
rect 1316 32885 1342 32949
rect 1406 32885 1432 32949
rect 1496 32885 1501 32949
rect 977 32869 1501 32885
rect 977 32805 982 32869
rect 1046 32805 1072 32869
rect 1136 32805 1162 32869
rect 1226 32805 1252 32869
rect 1316 32805 1342 32869
rect 1406 32805 1432 32869
rect 1496 32805 1501 32869
rect 977 32789 1501 32805
rect 977 32725 982 32789
rect 1046 32725 1072 32789
rect 1136 32725 1162 32789
rect 1226 32725 1252 32789
rect 1316 32725 1342 32789
rect 1406 32725 1432 32789
rect 1496 32725 1501 32789
rect 977 32709 1501 32725
rect 977 32645 982 32709
rect 1046 32645 1072 32709
rect 1136 32645 1162 32709
rect 1226 32645 1252 32709
rect 1316 32645 1342 32709
rect 1406 32645 1432 32709
rect 1496 32645 1501 32709
rect 977 32629 1501 32645
rect 977 32565 982 32629
rect 1046 32565 1072 32629
rect 1136 32565 1162 32629
rect 1226 32565 1252 32629
rect 1316 32565 1342 32629
rect 1406 32565 1432 32629
rect 1496 32565 1501 32629
rect 977 32549 1501 32565
rect 977 32485 982 32549
rect 1046 32485 1072 32549
rect 1136 32485 1162 32549
rect 1226 32485 1252 32549
rect 1316 32485 1342 32549
rect 1406 32485 1432 32549
rect 1496 32485 1501 32549
rect 977 32469 1501 32485
rect 977 32405 982 32469
rect 1046 32405 1072 32469
rect 1136 32405 1162 32469
rect 1226 32405 1252 32469
rect 1316 32405 1342 32469
rect 1406 32405 1432 32469
rect 1496 32405 1501 32469
rect 977 32389 1501 32405
rect 977 32325 982 32389
rect 1046 32325 1072 32389
rect 1136 32325 1162 32389
rect 1226 32325 1252 32389
rect 1316 32325 1342 32389
rect 1406 32325 1432 32389
rect 1496 32325 1501 32389
rect 977 32309 1501 32325
rect 977 32245 982 32309
rect 1046 32245 1072 32309
rect 1136 32245 1162 32309
rect 1226 32245 1252 32309
rect 1316 32245 1342 32309
rect 1406 32245 1432 32309
rect 1496 32245 1501 32309
rect 977 32229 1501 32245
rect 977 32165 982 32229
rect 1046 32165 1072 32229
rect 1136 32165 1162 32229
rect 1226 32165 1252 32229
rect 1316 32165 1342 32229
rect 1406 32165 1432 32229
rect 1496 32165 1501 32229
rect 977 32149 1501 32165
rect 977 32085 982 32149
rect 1046 32085 1072 32149
rect 1136 32085 1162 32149
rect 1226 32085 1252 32149
rect 1316 32085 1342 32149
rect 1406 32085 1432 32149
rect 1496 32085 1501 32149
rect 977 32069 1501 32085
rect 977 32005 982 32069
rect 1046 32005 1072 32069
rect 1136 32005 1162 32069
rect 1226 32005 1252 32069
rect 1316 32005 1342 32069
rect 1406 32005 1432 32069
rect 1496 32005 1501 32069
rect 977 31989 1501 32005
rect 977 31925 982 31989
rect 1046 31925 1072 31989
rect 1136 31925 1162 31989
rect 1226 31925 1252 31989
rect 1316 31925 1342 31989
rect 1406 31925 1432 31989
rect 1496 31925 1501 31989
rect 977 31909 1501 31925
rect 977 31845 982 31909
rect 1046 31845 1072 31909
rect 1136 31845 1162 31909
rect 1226 31845 1252 31909
rect 1316 31845 1342 31909
rect 1406 31845 1432 31909
rect 1496 31845 1501 31909
rect 977 31829 1501 31845
rect 977 31765 982 31829
rect 1046 31765 1072 31829
rect 1136 31765 1162 31829
rect 1226 31765 1252 31829
rect 1316 31765 1342 31829
rect 1406 31765 1432 31829
rect 1496 31765 1501 31829
rect 977 31749 1501 31765
rect 977 31685 982 31749
rect 1046 31685 1072 31749
rect 1136 31685 1162 31749
rect 1226 31685 1252 31749
rect 1316 31685 1342 31749
rect 1406 31685 1432 31749
rect 1496 31685 1501 31749
rect 977 31669 1501 31685
rect 977 31605 982 31669
rect 1046 31605 1072 31669
rect 1136 31605 1162 31669
rect 1226 31605 1252 31669
rect 1316 31605 1342 31669
rect 1406 31605 1432 31669
rect 1496 31605 1501 31669
rect 977 31589 1501 31605
rect 977 31525 982 31589
rect 1046 31525 1072 31589
rect 1136 31525 1162 31589
rect 1226 31525 1252 31589
rect 1316 31525 1342 31589
rect 1406 31525 1432 31589
rect 1496 31525 1501 31589
rect 977 31509 1501 31525
rect 977 31445 982 31509
rect 1046 31445 1072 31509
rect 1136 31445 1162 31509
rect 1226 31445 1252 31509
rect 1316 31445 1342 31509
rect 1406 31445 1432 31509
rect 1496 31445 1501 31509
rect 977 31429 1501 31445
rect 977 31365 982 31429
rect 1046 31365 1072 31429
rect 1136 31365 1162 31429
rect 1226 31365 1252 31429
rect 1316 31365 1342 31429
rect 1406 31365 1432 31429
rect 1496 31365 1501 31429
rect 977 31349 1501 31365
rect 977 31285 982 31349
rect 1046 31285 1072 31349
rect 1136 31285 1162 31349
rect 1226 31285 1252 31349
rect 1316 31285 1342 31349
rect 1406 31285 1432 31349
rect 1496 31285 1501 31349
rect 977 31269 1501 31285
rect 977 31205 982 31269
rect 1046 31205 1072 31269
rect 1136 31205 1162 31269
rect 1226 31205 1252 31269
rect 1316 31205 1342 31269
rect 1406 31205 1432 31269
rect 1496 31205 1501 31269
rect 977 31189 1501 31205
rect 977 31125 982 31189
rect 1046 31125 1072 31189
rect 1136 31125 1162 31189
rect 1226 31125 1252 31189
rect 1316 31125 1342 31189
rect 1406 31125 1432 31189
rect 1496 31125 1501 31189
rect 977 31109 1501 31125
rect 977 31045 982 31109
rect 1046 31045 1072 31109
rect 1136 31045 1162 31109
rect 1226 31045 1252 31109
rect 1316 31045 1342 31109
rect 1406 31045 1432 31109
rect 1496 31045 1501 31109
rect 977 31029 1501 31045
rect 977 30965 982 31029
rect 1046 30965 1072 31029
rect 1136 30965 1162 31029
rect 1226 30965 1252 31029
rect 1316 30965 1342 31029
rect 1406 30965 1432 31029
rect 1496 30965 1501 31029
rect 977 30949 1501 30965
rect 977 30885 982 30949
rect 1046 30885 1072 30949
rect 1136 30885 1162 30949
rect 1226 30885 1252 30949
rect 1316 30885 1342 30949
rect 1406 30885 1432 30949
rect 1496 30885 1501 30949
rect 977 30869 1501 30885
rect 977 30805 982 30869
rect 1046 30805 1072 30869
rect 1136 30805 1162 30869
rect 1226 30805 1252 30869
rect 1316 30805 1342 30869
rect 1406 30805 1432 30869
rect 1496 30805 1501 30869
rect 977 30789 1501 30805
rect 977 30725 982 30789
rect 1046 30725 1072 30789
rect 1136 30725 1162 30789
rect 1226 30725 1252 30789
rect 1316 30725 1342 30789
rect 1406 30725 1432 30789
rect 1496 30725 1501 30789
rect 977 30709 1501 30725
rect 977 30645 982 30709
rect 1046 30645 1072 30709
rect 1136 30645 1162 30709
rect 1226 30645 1252 30709
rect 1316 30645 1342 30709
rect 1406 30645 1432 30709
rect 1496 30645 1501 30709
rect 977 30629 1501 30645
rect 977 30565 982 30629
rect 1046 30565 1072 30629
rect 1136 30565 1162 30629
rect 1226 30565 1252 30629
rect 1316 30565 1342 30629
rect 1406 30565 1432 30629
rect 1496 30565 1501 30629
rect 977 30549 1501 30565
rect 977 30485 982 30549
rect 1046 30485 1072 30549
rect 1136 30485 1162 30549
rect 1226 30485 1252 30549
rect 1316 30485 1342 30549
rect 1406 30485 1432 30549
rect 1496 30485 1501 30549
rect 977 30469 1501 30485
rect 977 30405 982 30469
rect 1046 30405 1072 30469
rect 1136 30405 1162 30469
rect 1226 30405 1252 30469
rect 1316 30405 1342 30469
rect 1406 30405 1432 30469
rect 1496 30405 1501 30469
rect 977 30389 1501 30405
rect 977 30325 982 30389
rect 1046 30325 1072 30389
rect 1136 30325 1162 30389
rect 1226 30325 1252 30389
rect 1316 30325 1342 30389
rect 1406 30325 1432 30389
rect 1496 30325 1501 30389
rect 977 30309 1501 30325
rect 977 30245 982 30309
rect 1046 30245 1072 30309
rect 1136 30245 1162 30309
rect 1226 30245 1252 30309
rect 1316 30245 1342 30309
rect 1406 30245 1432 30309
rect 1496 30245 1501 30309
rect 977 30229 1501 30245
rect 977 30165 982 30229
rect 1046 30165 1072 30229
rect 1136 30165 1162 30229
rect 1226 30165 1252 30229
rect 1316 30165 1342 30229
rect 1406 30165 1432 30229
rect 1496 30165 1501 30229
rect 977 30149 1501 30165
rect 977 30085 982 30149
rect 1046 30085 1072 30149
rect 1136 30085 1162 30149
rect 1226 30085 1252 30149
rect 1316 30085 1342 30149
rect 1406 30085 1432 30149
rect 1496 30085 1501 30149
rect 977 30069 1501 30085
rect 977 30005 982 30069
rect 1046 30005 1072 30069
rect 1136 30005 1162 30069
rect 1226 30005 1252 30069
rect 1316 30005 1342 30069
rect 1406 30005 1432 30069
rect 1496 30005 1501 30069
rect 977 29989 1501 30005
rect 977 29925 982 29989
rect 1046 29925 1072 29989
rect 1136 29925 1162 29989
rect 1226 29925 1252 29989
rect 1316 29925 1342 29989
rect 1406 29925 1432 29989
rect 1496 29925 1501 29989
rect 977 29909 1501 29925
rect 977 29845 982 29909
rect 1046 29845 1072 29909
rect 1136 29845 1162 29909
rect 1226 29845 1252 29909
rect 1316 29845 1342 29909
rect 1406 29845 1432 29909
rect 1496 29845 1501 29909
rect 977 29829 1501 29845
rect 977 29765 982 29829
rect 1046 29765 1072 29829
rect 1136 29765 1162 29829
rect 1226 29765 1252 29829
rect 1316 29765 1342 29829
rect 1406 29765 1432 29829
rect 1496 29765 1501 29829
rect 977 29749 1501 29765
rect 977 29685 982 29749
rect 1046 29685 1072 29749
rect 1136 29685 1162 29749
rect 1226 29685 1252 29749
rect 1316 29685 1342 29749
rect 1406 29685 1432 29749
rect 1496 29685 1501 29749
rect 977 29669 1501 29685
rect 977 29605 982 29669
rect 1046 29605 1072 29669
rect 1136 29605 1162 29669
rect 1226 29605 1252 29669
rect 1316 29605 1342 29669
rect 1406 29605 1432 29669
rect 1496 29605 1501 29669
rect 977 29589 1501 29605
rect 977 29525 982 29589
rect 1046 29525 1072 29589
rect 1136 29525 1162 29589
rect 1226 29525 1252 29589
rect 1316 29525 1342 29589
rect 1406 29525 1432 29589
rect 1496 29525 1501 29589
rect 977 29509 1501 29525
rect 977 29445 982 29509
rect 1046 29445 1072 29509
rect 1136 29445 1162 29509
rect 1226 29445 1252 29509
rect 1316 29445 1342 29509
rect 1406 29445 1432 29509
rect 1496 29445 1501 29509
rect 977 29429 1501 29445
rect 977 29365 982 29429
rect 1046 29365 1072 29429
rect 1136 29365 1162 29429
rect 1226 29365 1252 29429
rect 1316 29365 1342 29429
rect 1406 29365 1432 29429
rect 1496 29365 1501 29429
rect 977 29349 1501 29365
rect 977 29285 982 29349
rect 1046 29285 1072 29349
rect 1136 29285 1162 29349
rect 1226 29285 1252 29349
rect 1316 29285 1342 29349
rect 1406 29285 1432 29349
rect 1496 29285 1501 29349
rect 977 29269 1501 29285
rect 977 29205 982 29269
rect 1046 29205 1072 29269
rect 1136 29205 1162 29269
rect 1226 29205 1252 29269
rect 1316 29205 1342 29269
rect 1406 29205 1432 29269
rect 1496 29205 1501 29269
rect 977 29189 1501 29205
rect 977 29125 982 29189
rect 1046 29125 1072 29189
rect 1136 29125 1162 29189
rect 1226 29125 1252 29189
rect 1316 29125 1342 29189
rect 1406 29125 1432 29189
rect 1496 29125 1501 29189
rect 977 29109 1501 29125
rect 977 29045 982 29109
rect 1046 29045 1072 29109
rect 1136 29045 1162 29109
rect 1226 29045 1252 29109
rect 1316 29045 1342 29109
rect 1406 29045 1432 29109
rect 1496 29045 1501 29109
rect 977 29029 1501 29045
rect 977 28965 982 29029
rect 1046 28965 1072 29029
rect 1136 28965 1162 29029
rect 1226 28965 1252 29029
rect 1316 28965 1342 29029
rect 1406 28965 1432 29029
rect 1496 28965 1501 29029
rect 977 28949 1501 28965
rect 977 28885 982 28949
rect 1046 28885 1072 28949
rect 1136 28885 1162 28949
rect 1226 28885 1252 28949
rect 1316 28885 1342 28949
rect 1406 28885 1432 28949
rect 1496 28885 1501 28949
rect 977 28869 1501 28885
rect 977 28805 982 28869
rect 1046 28805 1072 28869
rect 1136 28805 1162 28869
rect 1226 28805 1252 28869
rect 1316 28805 1342 28869
rect 1406 28805 1432 28869
rect 1496 28805 1501 28869
rect 977 28789 1501 28805
rect 977 28725 982 28789
rect 1046 28725 1072 28789
rect 1136 28725 1162 28789
rect 1226 28725 1252 28789
rect 1316 28725 1342 28789
rect 1406 28725 1432 28789
rect 1496 28725 1501 28789
rect 977 28709 1501 28725
rect 977 28645 982 28709
rect 1046 28645 1072 28709
rect 1136 28645 1162 28709
rect 1226 28645 1252 28709
rect 1316 28645 1342 28709
rect 1406 28645 1432 28709
rect 1496 28645 1501 28709
rect 977 28629 1501 28645
rect 977 28565 982 28629
rect 1046 28565 1072 28629
rect 1136 28565 1162 28629
rect 1226 28565 1252 28629
rect 1316 28565 1342 28629
rect 1406 28565 1432 28629
rect 1496 28565 1501 28629
rect 977 28549 1501 28565
rect 977 28485 982 28549
rect 1046 28485 1072 28549
rect 1136 28485 1162 28549
rect 1226 28485 1252 28549
rect 1316 28485 1342 28549
rect 1406 28485 1432 28549
rect 1496 28485 1501 28549
rect 977 28469 1501 28485
rect 977 28405 982 28469
rect 1046 28405 1072 28469
rect 1136 28405 1162 28469
rect 1226 28405 1252 28469
rect 1316 28405 1342 28469
rect 1406 28405 1432 28469
rect 1496 28405 1501 28469
rect 977 28389 1501 28405
rect 977 28325 982 28389
rect 1046 28325 1072 28389
rect 1136 28325 1162 28389
rect 1226 28325 1252 28389
rect 1316 28325 1342 28389
rect 1406 28325 1432 28389
rect 1496 28325 1501 28389
rect 977 28309 1501 28325
rect 977 28245 982 28309
rect 1046 28245 1072 28309
rect 1136 28245 1162 28309
rect 1226 28245 1252 28309
rect 1316 28245 1342 28309
rect 1406 28245 1432 28309
rect 1496 28245 1501 28309
rect 977 28229 1501 28245
rect 977 28165 982 28229
rect 1046 28165 1072 28229
rect 1136 28165 1162 28229
rect 1226 28165 1252 28229
rect 1316 28165 1342 28229
rect 1406 28165 1432 28229
rect 1496 28165 1501 28229
rect 977 28149 1501 28165
rect 977 28085 982 28149
rect 1046 28085 1072 28149
rect 1136 28085 1162 28149
rect 1226 28085 1252 28149
rect 1316 28085 1342 28149
rect 1406 28085 1432 28149
rect 1496 28085 1501 28149
rect 977 28069 1501 28085
rect 977 28005 982 28069
rect 1046 28005 1072 28069
rect 1136 28005 1162 28069
rect 1226 28005 1252 28069
rect 1316 28005 1342 28069
rect 1406 28005 1432 28069
rect 1496 28005 1501 28069
rect 977 27989 1501 28005
rect 977 27925 982 27989
rect 1046 27925 1072 27989
rect 1136 27925 1162 27989
rect 1226 27925 1252 27989
rect 1316 27925 1342 27989
rect 1406 27925 1432 27989
rect 1496 27925 1501 27989
rect 977 27909 1501 27925
rect 977 27845 982 27909
rect 1046 27845 1072 27909
rect 1136 27845 1162 27909
rect 1226 27845 1252 27909
rect 1316 27845 1342 27909
rect 1406 27845 1432 27909
rect 1496 27845 1501 27909
rect 977 27829 1501 27845
rect 977 27765 982 27829
rect 1046 27765 1072 27829
rect 1136 27765 1162 27829
rect 1226 27765 1252 27829
rect 1316 27765 1342 27829
rect 1406 27765 1432 27829
rect 1496 27765 1501 27829
rect 977 27749 1501 27765
rect 977 27685 982 27749
rect 1046 27685 1072 27749
rect 1136 27685 1162 27749
rect 1226 27685 1252 27749
rect 1316 27685 1342 27749
rect 1406 27685 1432 27749
rect 1496 27685 1501 27749
rect 977 27669 1501 27685
rect 977 27605 982 27669
rect 1046 27605 1072 27669
rect 1136 27605 1162 27669
rect 1226 27605 1252 27669
rect 1316 27605 1342 27669
rect 1406 27605 1432 27669
rect 1496 27605 1501 27669
rect 977 27589 1501 27605
rect 977 27525 982 27589
rect 1046 27525 1072 27589
rect 1136 27525 1162 27589
rect 1226 27525 1252 27589
rect 1316 27525 1342 27589
rect 1406 27525 1432 27589
rect 1496 27525 1501 27589
rect 977 27509 1501 27525
rect 977 27445 982 27509
rect 1046 27445 1072 27509
rect 1136 27445 1162 27509
rect 1226 27445 1252 27509
rect 1316 27445 1342 27509
rect 977 27429 1384 27445
rect 977 27365 982 27429
rect 1046 27365 1072 27429
rect 1136 27365 1162 27429
rect 1226 27365 1252 27429
rect 1316 27365 1342 27429
rect 977 27349 1384 27365
rect 977 27285 982 27349
rect 1046 27285 1072 27349
rect 1136 27285 1162 27349
rect 1226 27285 1252 27349
rect 1316 27285 1342 27349
rect 977 27269 1384 27285
rect 977 27205 982 27269
rect 1046 27205 1072 27269
rect 1136 27205 1162 27269
rect 1226 27205 1252 27269
rect 1316 27205 1342 27269
rect 977 27189 1384 27205
rect 977 27125 982 27189
rect 1046 27125 1072 27189
rect 1136 27125 1162 27189
rect 1226 27125 1252 27189
rect 1316 27125 1342 27189
rect 977 27109 1384 27125
rect 977 27045 982 27109
rect 1046 27045 1072 27109
rect 1136 27045 1162 27109
rect 1226 27045 1252 27109
rect 1316 27045 1342 27109
rect 977 27029 1384 27045
rect 977 26965 982 27029
rect 1046 26965 1072 27029
rect 1136 26965 1162 27029
rect 1226 26965 1252 27029
rect 1316 26965 1342 27029
rect 977 26949 1384 26965
rect 977 26885 982 26949
rect 1046 26885 1072 26949
rect 1136 26885 1162 26949
rect 1226 26885 1252 26949
rect 1316 26885 1342 26949
rect 977 26869 1384 26885
rect 977 26805 982 26869
rect 1046 26805 1072 26869
rect 1136 26805 1162 26869
rect 1226 26805 1252 26869
rect 1316 26805 1342 26869
rect 977 26789 1384 26805
rect 977 26725 982 26789
rect 1046 26725 1072 26789
rect 1136 26725 1162 26789
rect 1226 26725 1252 26789
rect 1316 26725 1342 26789
rect 977 26709 1384 26725
rect 977 26645 982 26709
rect 1046 26645 1072 26709
rect 1136 26645 1162 26709
rect 1226 26645 1252 26709
rect 1316 26645 1342 26709
rect 1406 26645 1432 27509
rect 1496 26645 1501 27509
rect 977 26629 1501 26645
rect 977 26565 982 26629
rect 1046 26565 1072 26629
rect 1136 26565 1162 26629
rect 1226 26565 1252 26629
rect 1316 26565 1342 26629
rect 1406 26565 1432 26629
rect 1496 26565 1501 26629
rect 977 26549 1501 26565
rect 977 26485 982 26549
rect 1046 26485 1072 26549
rect 1136 26485 1162 26549
rect 1226 26485 1252 26549
rect 1316 26485 1342 26549
rect 1406 26485 1432 26549
rect 1496 26485 1501 26549
rect 977 26469 1501 26485
rect 977 26405 982 26469
rect 1046 26405 1072 26469
rect 1136 26405 1162 26469
rect 1226 26405 1252 26469
rect 1316 26405 1342 26469
rect 1406 26405 1432 26469
rect 1496 26405 1501 26469
rect 977 26389 1501 26405
rect 977 26325 982 26389
rect 1046 26325 1072 26389
rect 1136 26325 1162 26389
rect 1226 26325 1252 26389
rect 1316 26325 1342 26389
rect 1406 26325 1432 26389
rect 1496 26325 1501 26389
rect 977 26309 1501 26325
rect 977 26245 982 26309
rect 1046 26245 1072 26309
rect 1136 26245 1162 26309
rect 1226 26245 1252 26309
rect 1316 26245 1342 26309
rect 1406 26245 1432 26309
rect 1496 26245 1501 26309
rect 977 26229 1501 26245
rect 977 26165 982 26229
rect 1046 26165 1072 26229
rect 1136 26165 1162 26229
rect 1226 26165 1252 26229
rect 1316 26165 1342 26229
rect 1406 26165 1432 26229
rect 1496 26165 1501 26229
rect 977 26149 1501 26165
rect 977 26085 982 26149
rect 1046 26085 1072 26149
rect 1136 26085 1162 26149
rect 1226 26085 1252 26149
rect 1316 26085 1342 26149
rect 1406 26085 1432 26149
rect 1496 26085 1501 26149
rect 977 26069 1501 26085
rect 977 26005 982 26069
rect 1046 26005 1072 26069
rect 1136 26005 1162 26069
rect 1226 26005 1252 26069
rect 1316 26005 1342 26069
rect 1406 26005 1432 26069
rect 1496 26005 1501 26069
rect 977 25989 1501 26005
rect 977 25925 982 25989
rect 1046 25925 1072 25989
rect 1136 25925 1162 25989
rect 1226 25925 1252 25989
rect 1316 25925 1342 25989
rect 1406 25925 1432 25989
rect 1496 25925 1501 25989
rect 977 25909 1501 25925
rect 977 25845 982 25909
rect 1046 25845 1072 25909
rect 1136 25845 1162 25909
rect 1226 25845 1252 25909
rect 1316 25845 1342 25909
rect 1406 25845 1432 25909
rect 1496 25845 1501 25909
rect 977 25829 1501 25845
rect 977 25765 982 25829
rect 1046 25765 1072 25829
rect 1136 25765 1162 25829
rect 1226 25765 1252 25829
rect 1316 25765 1342 25829
rect 1406 25765 1432 25829
rect 1496 25765 1501 25829
rect 977 25749 1501 25765
rect 977 25685 982 25749
rect 1046 25685 1072 25749
rect 1136 25685 1162 25749
rect 1226 25685 1252 25749
rect 1316 25685 1342 25749
rect 1406 25685 1432 25749
rect 1496 25685 1501 25749
rect 977 25669 1501 25685
rect 977 25605 982 25669
rect 1046 25605 1072 25669
rect 1136 25605 1162 25669
rect 1226 25605 1252 25669
rect 1316 25605 1342 25669
rect 1406 25605 1432 25669
rect 1496 25605 1501 25669
rect 977 25589 1501 25605
rect 977 25525 982 25589
rect 1046 25525 1072 25589
rect 1136 25525 1162 25589
rect 1226 25525 1252 25589
rect 1316 25525 1342 25589
rect 1406 25525 1432 25589
rect 1496 25525 1501 25589
rect 977 25509 1501 25525
rect 977 25445 982 25509
rect 1046 25445 1072 25509
rect 1136 25445 1162 25509
rect 1226 25445 1252 25509
rect 1316 25445 1342 25509
rect 1406 25445 1432 25509
rect 1496 25445 1501 25509
rect 977 25429 1501 25445
rect 977 25365 982 25429
rect 1046 25365 1072 25429
rect 1136 25365 1162 25429
rect 1226 25365 1252 25429
rect 1316 25365 1342 25429
rect 1406 25365 1432 25429
rect 1496 25365 1501 25429
rect 977 25349 1501 25365
rect 977 25285 982 25349
rect 1046 25285 1072 25349
rect 1136 25285 1162 25349
rect 1226 25285 1252 25349
rect 1316 25285 1342 25349
rect 1406 25285 1432 25349
rect 1496 25285 1501 25349
rect 977 25269 1501 25285
rect 977 25205 982 25269
rect 1046 25205 1072 25269
rect 1136 25205 1162 25269
rect 1226 25205 1252 25269
rect 1316 25205 1342 25269
rect 1406 25205 1432 25269
rect 1496 25205 1501 25269
rect 977 25189 1501 25205
rect 977 25125 982 25189
rect 1046 25125 1072 25189
rect 1136 25125 1162 25189
rect 1226 25125 1252 25189
rect 1316 25125 1342 25189
rect 1406 25125 1432 25189
rect 1496 25125 1501 25189
rect 977 25109 1501 25125
rect 977 25045 982 25109
rect 1046 25045 1072 25109
rect 1136 25045 1162 25109
rect 1226 25045 1252 25109
rect 1316 25045 1342 25109
rect 1406 25045 1432 25109
rect 1496 25045 1501 25109
rect 977 25029 1501 25045
rect 977 24965 982 25029
rect 1046 24965 1072 25029
rect 1136 24965 1162 25029
rect 1226 24965 1252 25029
rect 1316 24965 1342 25029
rect 1406 24965 1432 25029
rect 1496 24965 1501 25029
rect 977 24949 1501 24965
rect 977 24885 982 24949
rect 1046 24885 1072 24949
rect 1136 24885 1162 24949
rect 1226 24885 1252 24949
rect 1316 24885 1342 24949
rect 1406 24885 1432 24949
rect 1496 24885 1501 24949
rect 977 24869 1501 24885
rect 977 24805 982 24869
rect 1046 24805 1072 24869
rect 1136 24805 1162 24869
rect 1226 24805 1252 24869
rect 1316 24805 1342 24869
rect 1406 24805 1432 24869
rect 1496 24805 1501 24869
rect 977 24789 1501 24805
rect 977 24725 982 24789
rect 1046 24725 1072 24789
rect 1136 24725 1162 24789
rect 1226 24725 1252 24789
rect 1316 24725 1342 24789
rect 1406 24725 1432 24789
rect 1496 24725 1501 24789
rect 977 24709 1501 24725
rect 977 24645 982 24709
rect 1046 24645 1072 24709
rect 1136 24645 1162 24709
rect 1226 24645 1252 24709
rect 1316 24645 1342 24709
rect 1406 24645 1432 24709
rect 1496 24645 1501 24709
rect 977 24629 1501 24645
rect 977 24565 982 24629
rect 1046 24565 1072 24629
rect 1136 24565 1162 24629
rect 1226 24565 1252 24629
rect 1316 24565 1342 24629
rect 1406 24565 1432 24629
rect 1496 24565 1501 24629
rect 977 24549 1501 24565
rect 977 24485 982 24549
rect 1046 24485 1072 24549
rect 1136 24485 1162 24549
rect 1226 24485 1252 24549
rect 1316 24485 1342 24549
rect 1406 24485 1432 24549
rect 1496 24485 1501 24549
rect 977 24469 1501 24485
rect 977 24405 982 24469
rect 1046 24405 1072 24469
rect 1136 24405 1162 24469
rect 1226 24405 1252 24469
rect 1316 24405 1342 24469
rect 1406 24405 1432 24469
rect 1496 24405 1501 24469
rect 977 24389 1501 24405
rect 977 24325 982 24389
rect 1046 24325 1072 24389
rect 1136 24325 1162 24389
rect 1226 24325 1252 24389
rect 1316 24325 1342 24389
rect 1406 24325 1432 24389
rect 1496 24325 1501 24389
rect 977 24309 1501 24325
rect 977 24245 982 24309
rect 1046 24245 1072 24309
rect 1136 24245 1162 24309
rect 1226 24245 1252 24309
rect 1316 24245 1342 24309
rect 1406 24245 1432 24309
rect 1496 24245 1501 24309
rect 977 24229 1501 24245
rect 977 24165 982 24229
rect 1046 24165 1072 24229
rect 1136 24165 1162 24229
rect 1226 24165 1252 24229
rect 1316 24165 1342 24229
rect 1406 24165 1432 24229
rect 1496 24165 1501 24229
rect 977 24149 1501 24165
rect 977 24085 982 24149
rect 1046 24085 1072 24149
rect 1136 24085 1162 24149
rect 1226 24085 1252 24149
rect 1316 24085 1342 24149
rect 1406 24085 1432 24149
rect 1496 24085 1501 24149
rect 977 24069 1501 24085
rect 977 24005 982 24069
rect 1046 24005 1072 24069
rect 1136 24005 1162 24069
rect 1226 24005 1252 24069
rect 1316 24005 1342 24069
rect 1406 24005 1432 24069
rect 1496 24005 1501 24069
rect 977 23989 1501 24005
rect 977 23925 982 23989
rect 1046 23925 1072 23989
rect 1136 23925 1162 23989
rect 1226 23925 1252 23989
rect 1316 23925 1342 23989
rect 1406 23925 1432 23989
rect 1496 23925 1501 23989
rect 977 23909 1501 23925
rect 977 23845 982 23909
rect 1046 23845 1072 23909
rect 1136 23845 1162 23909
rect 1226 23845 1252 23909
rect 1316 23845 1342 23909
rect 1406 23845 1432 23909
rect 1496 23845 1501 23909
rect 977 23829 1501 23845
rect 977 23765 982 23829
rect 1046 23765 1072 23829
rect 1136 23765 1162 23829
rect 1226 23765 1252 23829
rect 1316 23765 1342 23829
rect 1406 23765 1432 23829
rect 1496 23765 1501 23829
rect 977 23749 1501 23765
rect 977 23685 982 23749
rect 1046 23685 1072 23749
rect 1136 23685 1162 23749
rect 1226 23685 1252 23749
rect 1316 23685 1342 23749
rect 1406 23685 1432 23749
rect 1496 23685 1501 23749
rect 977 23669 1501 23685
rect 977 23605 982 23669
rect 1046 23605 1072 23669
rect 1136 23605 1162 23669
rect 1226 23605 1252 23669
rect 1316 23605 1342 23669
rect 1406 23605 1432 23669
rect 1496 23605 1501 23669
rect 977 23589 1501 23605
rect 977 23525 982 23589
rect 1046 23525 1072 23589
rect 1136 23525 1162 23589
rect 1226 23525 1252 23589
rect 1316 23525 1342 23589
rect 1406 23525 1432 23589
rect 1496 23525 1501 23589
rect 977 23509 1501 23525
rect 977 23445 982 23509
rect 1046 23445 1072 23509
rect 1136 23445 1162 23509
rect 1226 23445 1252 23509
rect 1316 23445 1342 23509
rect 1406 23445 1432 23509
rect 1496 23445 1501 23509
rect 977 23429 1501 23445
rect 977 23365 982 23429
rect 1046 23365 1072 23429
rect 1136 23365 1162 23429
rect 1226 23365 1252 23429
rect 1316 23365 1342 23429
rect 1406 23365 1432 23429
rect 1496 23365 1501 23429
rect 977 23349 1501 23365
rect 977 23285 982 23349
rect 1046 23285 1072 23349
rect 1136 23285 1162 23349
rect 1226 23285 1252 23349
rect 1316 23285 1342 23349
rect 1406 23285 1432 23349
rect 1496 23285 1501 23349
rect 977 23268 1501 23285
rect 977 23204 982 23268
rect 1046 23204 1072 23268
rect 1136 23204 1162 23268
rect 1226 23204 1252 23268
rect 1316 23204 1342 23268
rect 1406 23204 1432 23268
rect 1496 23204 1501 23268
rect 977 23187 1501 23204
rect 977 23123 982 23187
rect 1046 23123 1072 23187
rect 1136 23123 1162 23187
rect 1226 23123 1252 23187
rect 1316 23123 1342 23187
rect 1406 23123 1432 23187
rect 1496 23123 1501 23187
rect 977 23106 1501 23123
rect 977 23042 982 23106
rect 1046 23042 1072 23106
rect 1136 23042 1162 23106
rect 1226 23042 1252 23106
rect 1316 23042 1342 23106
rect 1406 23042 1432 23106
rect 1496 23042 1501 23106
rect 977 23025 1501 23042
rect 977 22961 982 23025
rect 1046 22961 1072 23025
rect 1136 22961 1162 23025
rect 1226 22961 1252 23025
rect 1316 22961 1342 23025
rect 1406 22961 1432 23025
rect 1496 22961 1501 23025
rect 977 22944 1501 22961
rect 977 22880 982 22944
rect 1046 22880 1072 22944
rect 1136 22880 1162 22944
rect 1226 22880 1252 22944
rect 1316 22880 1342 22944
rect 1406 22880 1432 22944
rect 1496 22880 1501 22944
rect 977 22863 1501 22880
rect 977 22799 982 22863
rect 1046 22799 1072 22863
rect 1136 22799 1162 22863
rect 1226 22799 1252 22863
rect 1316 22799 1342 22863
rect 1406 22799 1432 22863
rect 1496 22799 1501 22863
rect 977 22782 1501 22799
rect 977 22718 982 22782
rect 1046 22718 1072 22782
rect 1136 22718 1162 22782
rect 1226 22718 1252 22782
rect 1316 22718 1342 22782
rect 1406 22718 1432 22782
rect 1496 22718 1501 22782
rect 977 22701 1501 22718
rect 977 22637 982 22701
rect 1046 22637 1072 22701
rect 1136 22637 1162 22701
rect 1226 22637 1252 22701
rect 1316 22637 1342 22701
rect 1406 22637 1432 22701
rect 1496 22637 1501 22701
rect 977 22620 1501 22637
rect 977 22556 982 22620
rect 1046 22556 1072 22620
rect 1136 22556 1162 22620
rect 1226 22556 1252 22620
rect 1316 22556 1342 22620
rect 1406 22556 1432 22620
rect 1496 22556 1501 22620
rect 977 22539 1501 22556
rect 977 22475 982 22539
rect 1046 22475 1072 22539
rect 1136 22475 1162 22539
rect 1226 22475 1252 22539
rect 1316 22475 1342 22539
rect 1406 22475 1432 22539
rect 1496 22475 1501 22539
rect 977 22458 1501 22475
rect 977 22394 982 22458
rect 1046 22394 1072 22458
rect 1136 22394 1162 22458
rect 1226 22394 1252 22458
rect 1316 22394 1342 22458
rect 1406 22394 1432 22458
rect 1496 22394 1501 22458
rect 977 22377 1501 22394
rect 977 22313 982 22377
rect 1046 22313 1072 22377
rect 1136 22313 1162 22377
rect 1226 22313 1252 22377
rect 1316 22313 1342 22377
rect 1406 22313 1432 22377
rect 1496 22313 1501 22377
rect 977 22296 1501 22313
rect 977 22232 982 22296
rect 1046 22232 1072 22296
rect 1136 22232 1162 22296
rect 1226 22232 1252 22296
rect 1316 22232 1342 22296
rect 1406 22232 1432 22296
rect 1496 22232 1501 22296
rect 977 22215 1501 22232
rect 977 22151 982 22215
rect 1046 22151 1072 22215
rect 1136 22151 1162 22215
rect 1226 22151 1252 22215
rect 1316 22151 1342 22215
rect 1406 22151 1432 22215
rect 1496 22151 1501 22215
rect 977 22134 1501 22151
rect 977 22070 982 22134
rect 1046 22070 1072 22134
rect 1136 22070 1162 22134
rect 1226 22070 1252 22134
rect 1316 22070 1342 22134
rect 1406 22070 1432 22134
rect 1496 22070 1501 22134
rect 977 22053 1501 22070
rect 977 21989 982 22053
rect 1046 21989 1072 22053
rect 1136 21989 1162 22053
rect 1226 21989 1252 22053
rect 1316 21989 1342 22053
rect 1406 21989 1432 22053
rect 1496 21989 1501 22053
rect 977 21972 1501 21989
rect 977 21908 982 21972
rect 1046 21908 1072 21972
rect 1136 21908 1162 21972
rect 1226 21908 1252 21972
rect 1316 21908 1342 21972
rect 1406 21908 1432 21972
rect 1496 21908 1501 21972
rect 977 21891 1501 21908
rect 977 21827 982 21891
rect 1046 21827 1072 21891
rect 1136 21827 1162 21891
rect 1226 21827 1252 21891
rect 1316 21827 1342 21891
rect 1406 21827 1432 21891
rect 1496 21827 1501 21891
rect 977 21810 1501 21827
rect 977 21746 982 21810
rect 1046 21746 1072 21810
rect 1136 21746 1162 21810
rect 1226 21746 1252 21810
rect 1316 21746 1342 21810
rect 1406 21746 1432 21810
rect 1496 21746 1501 21810
rect 977 21729 1501 21746
rect 977 21665 982 21729
rect 1046 21665 1072 21729
rect 1136 21665 1162 21729
rect 1226 21665 1252 21729
rect 1316 21665 1342 21729
rect 1406 21665 1432 21729
rect 1496 21665 1501 21729
rect 977 21648 1501 21665
rect 977 21584 982 21648
rect 1046 21584 1072 21648
rect 1136 21584 1162 21648
rect 1226 21584 1252 21648
rect 1316 21584 1342 21648
rect 1406 21584 1432 21648
rect 1496 21584 1501 21648
rect 977 21567 1501 21584
rect 977 21503 982 21567
rect 1046 21503 1072 21567
rect 1136 21503 1162 21567
rect 1226 21503 1252 21567
rect 1316 21503 1342 21567
rect 1406 21503 1432 21567
rect 1496 21503 1501 21567
rect 977 21486 1501 21503
rect 977 21422 982 21486
rect 1046 21422 1072 21486
rect 1136 21422 1162 21486
rect 1226 21422 1252 21486
rect 1316 21422 1342 21486
rect 1406 21422 1432 21486
rect 1496 21422 1501 21486
rect 977 21405 1501 21422
rect 977 21341 982 21405
rect 1046 21341 1072 21405
rect 1136 21341 1162 21405
rect 1226 21341 1252 21405
rect 1316 21341 1342 21405
rect 1406 21341 1432 21405
rect 1496 21341 1501 21405
rect 977 21324 1501 21341
rect 977 21260 982 21324
rect 1046 21260 1072 21324
rect 1136 21260 1162 21324
rect 1226 21260 1252 21324
rect 1316 21260 1342 21324
rect 1406 21260 1432 21324
rect 1496 21260 1501 21324
rect 977 21243 1501 21260
rect 977 21179 982 21243
rect 1046 21179 1072 21243
rect 1136 21179 1162 21243
rect 1226 21179 1252 21243
rect 1316 21179 1342 21243
rect 1406 21179 1432 21243
rect 1496 21179 1501 21243
rect 977 21162 1501 21179
rect 977 21098 982 21162
rect 1046 21098 1072 21162
rect 1136 21098 1162 21162
rect 1226 21098 1252 21162
rect 1316 21098 1342 21162
rect 1406 21098 1432 21162
rect 1496 21098 1501 21162
rect 977 21081 1501 21098
rect 977 21017 982 21081
rect 1046 21017 1072 21081
rect 1136 21017 1162 21081
rect 1226 21017 1252 21081
rect 1316 21017 1342 21081
rect 1406 21017 1432 21081
rect 1496 21017 1501 21081
rect 977 21000 1501 21017
rect 977 20936 982 21000
rect 1046 20936 1072 21000
rect 1136 20936 1162 21000
rect 1226 20936 1252 21000
rect 1316 20936 1342 21000
rect 1406 20936 1432 21000
rect 1496 20972 1501 21000
rect 13515 33109 14039 33110
rect 13515 33045 13520 33109
rect 13584 33045 13610 33109
rect 13674 33045 13700 33109
rect 13764 33045 13790 33109
rect 13854 33045 13880 33109
rect 13944 33045 13970 33109
rect 14034 33045 14039 33109
rect 13515 33029 14039 33045
rect 13515 32965 13520 33029
rect 13584 32965 13610 33029
rect 13674 32965 13700 33029
rect 13764 32965 13790 33029
rect 13854 32965 13880 33029
rect 13944 32965 13970 33029
rect 14034 32965 14039 33029
rect 13515 32949 14039 32965
rect 13515 32885 13520 32949
rect 13584 32885 13610 32949
rect 13674 32885 13700 32949
rect 13764 32885 13790 32949
rect 13854 32885 13880 32949
rect 13944 32885 13970 32949
rect 14034 32885 14039 32949
rect 13515 32869 14039 32885
rect 13515 32805 13520 32869
rect 13584 32805 13610 32869
rect 13674 32805 13700 32869
rect 13764 32805 13790 32869
rect 13854 32805 13880 32869
rect 13944 32805 13970 32869
rect 14034 32805 14039 32869
rect 13515 32789 14039 32805
rect 13515 32725 13520 32789
rect 13584 32725 13610 32789
rect 13674 32725 13700 32789
rect 13764 32725 13790 32789
rect 13854 32725 13880 32789
rect 13944 32725 13970 32789
rect 14034 32725 14039 32789
rect 13515 32709 14039 32725
rect 13515 32645 13520 32709
rect 13584 32645 13610 32709
rect 13674 32645 13700 32709
rect 13764 32645 13790 32709
rect 13854 32645 13880 32709
rect 13944 32645 13970 32709
rect 14034 32645 14039 32709
rect 13515 32629 14039 32645
rect 13515 32565 13520 32629
rect 13584 32565 13610 32629
rect 13674 32565 13700 32629
rect 13764 32565 13790 32629
rect 13854 32565 13880 32629
rect 13944 32565 13970 32629
rect 14034 32565 14039 32629
rect 13515 32549 14039 32565
rect 13515 32485 13520 32549
rect 13584 32485 13610 32549
rect 13674 32485 13700 32549
rect 13764 32485 13790 32549
rect 13854 32485 13880 32549
rect 13944 32485 13970 32549
rect 14034 32485 14039 32549
rect 13515 32469 14039 32485
rect 13515 32405 13520 32469
rect 13584 32405 13610 32469
rect 13674 32405 13700 32469
rect 13764 32405 13790 32469
rect 13854 32405 13880 32469
rect 13944 32405 13970 32469
rect 14034 32405 14039 32469
rect 13515 32389 14039 32405
rect 13515 32325 13520 32389
rect 13584 32325 13610 32389
rect 13674 32325 13700 32389
rect 13764 32325 13790 32389
rect 13854 32325 13880 32389
rect 13944 32325 13970 32389
rect 14034 32325 14039 32389
rect 13515 32309 14039 32325
rect 13515 32245 13520 32309
rect 13584 32245 13610 32309
rect 13674 32245 13700 32309
rect 13764 32245 13790 32309
rect 13854 32245 13880 32309
rect 13944 32245 13970 32309
rect 14034 32245 14039 32309
rect 13515 32229 14039 32245
rect 13515 32165 13520 32229
rect 13584 32165 13610 32229
rect 13674 32165 13700 32229
rect 13764 32165 13790 32229
rect 13854 32165 13880 32229
rect 13944 32165 13970 32229
rect 14034 32165 14039 32229
rect 13515 32149 14039 32165
rect 13515 32085 13520 32149
rect 13584 32085 13610 32149
rect 13674 32085 13700 32149
rect 13764 32085 13790 32149
rect 13854 32085 13880 32149
rect 13944 32085 13970 32149
rect 14034 32085 14039 32149
rect 13515 32069 14039 32085
rect 13515 32005 13520 32069
rect 13584 32005 13610 32069
rect 13674 32005 13700 32069
rect 13764 32005 13790 32069
rect 13854 32005 13880 32069
rect 13944 32005 13970 32069
rect 14034 32005 14039 32069
rect 13515 31989 14039 32005
rect 13515 31925 13520 31989
rect 13584 31925 13610 31989
rect 13674 31925 13700 31989
rect 13764 31925 13790 31989
rect 13854 31925 13880 31989
rect 13944 31925 13970 31989
rect 14034 31925 14039 31989
rect 13515 31909 14039 31925
rect 13515 31845 13520 31909
rect 13584 31845 13610 31909
rect 13674 31845 13700 31909
rect 13764 31845 13790 31909
rect 13854 31845 13880 31909
rect 13944 31845 13970 31909
rect 14034 31845 14039 31909
rect 13515 31829 14039 31845
rect 13515 31765 13520 31829
rect 13584 31765 13610 31829
rect 13674 31765 13700 31829
rect 13764 31765 13790 31829
rect 13854 31765 13880 31829
rect 13944 31765 13970 31829
rect 14034 31765 14039 31829
rect 13515 31749 14039 31765
rect 13515 31685 13520 31749
rect 13584 31685 13610 31749
rect 13674 31685 13700 31749
rect 13764 31685 13790 31749
rect 13854 31685 13880 31749
rect 13944 31685 13970 31749
rect 14034 31685 14039 31749
rect 13515 31669 14039 31685
rect 13515 31605 13520 31669
rect 13584 31605 13610 31669
rect 13674 31605 13700 31669
rect 13764 31605 13790 31669
rect 13854 31605 13880 31669
rect 13944 31605 13970 31669
rect 14034 31605 14039 31669
rect 13515 31589 14039 31605
rect 13515 31525 13520 31589
rect 13584 31525 13610 31589
rect 13674 31525 13700 31589
rect 13764 31525 13790 31589
rect 13854 31525 13880 31589
rect 13944 31525 13970 31589
rect 14034 31525 14039 31589
rect 13515 31509 14039 31525
rect 13515 31445 13520 31509
rect 13584 31445 13610 31509
rect 13674 31445 13700 31509
rect 13764 31445 13790 31509
rect 13854 31445 13880 31509
rect 13944 31445 13970 31509
rect 14034 31445 14039 31509
rect 13515 31429 14039 31445
rect 13515 31365 13520 31429
rect 13584 31365 13610 31429
rect 13674 31365 13700 31429
rect 13764 31365 13790 31429
rect 13854 31365 13880 31429
rect 13944 31365 13970 31429
rect 14034 31365 14039 31429
rect 13515 31349 14039 31365
rect 13515 31285 13520 31349
rect 13584 31285 13610 31349
rect 13674 31285 13700 31349
rect 13764 31285 13790 31349
rect 13854 31285 13880 31349
rect 13944 31285 13970 31349
rect 14034 31285 14039 31349
rect 13515 31269 14039 31285
rect 13515 31205 13520 31269
rect 13584 31205 13610 31269
rect 13674 31205 13700 31269
rect 13764 31205 13790 31269
rect 13854 31205 13880 31269
rect 13944 31205 13970 31269
rect 14034 31205 14039 31269
rect 13515 31189 14039 31205
rect 13515 31125 13520 31189
rect 13584 31125 13610 31189
rect 13674 31125 13700 31189
rect 13764 31125 13790 31189
rect 13854 31125 13880 31189
rect 13944 31125 13970 31189
rect 14034 31125 14039 31189
rect 13515 31109 14039 31125
rect 13515 31045 13520 31109
rect 13584 31045 13610 31109
rect 13674 31045 13700 31109
rect 13764 31045 13790 31109
rect 13854 31045 13880 31109
rect 13944 31045 13970 31109
rect 14034 31045 14039 31109
rect 13515 31029 14039 31045
rect 13515 30965 13520 31029
rect 13584 30965 13610 31029
rect 13674 30965 13700 31029
rect 13764 30965 13790 31029
rect 13854 30965 13880 31029
rect 13944 30965 13970 31029
rect 14034 30965 14039 31029
rect 13515 30949 14039 30965
rect 13515 30885 13520 30949
rect 13584 30885 13610 30949
rect 13674 30885 13700 30949
rect 13764 30885 13790 30949
rect 13854 30885 13880 30949
rect 13944 30885 13970 30949
rect 14034 30885 14039 30949
rect 13515 30869 14039 30885
rect 13515 30805 13520 30869
rect 13584 30805 13610 30869
rect 13674 30805 13700 30869
rect 13764 30805 13790 30869
rect 13854 30805 13880 30869
rect 13944 30805 13970 30869
rect 14034 30805 14039 30869
rect 13515 30789 14039 30805
rect 13515 30725 13520 30789
rect 13584 30725 13610 30789
rect 13674 30725 13700 30789
rect 13764 30725 13790 30789
rect 13854 30725 13880 30789
rect 13944 30725 13970 30789
rect 14034 30725 14039 30789
rect 13515 30709 14039 30725
rect 13515 30645 13520 30709
rect 13584 30645 13610 30709
rect 13674 30645 13700 30709
rect 13764 30645 13790 30709
rect 13854 30645 13880 30709
rect 13944 30645 13970 30709
rect 14034 30645 14039 30709
rect 13515 30629 14039 30645
rect 13515 30565 13520 30629
rect 13584 30565 13610 30629
rect 13674 30565 13700 30629
rect 13764 30565 13790 30629
rect 13854 30565 13880 30629
rect 13944 30565 13970 30629
rect 14034 30565 14039 30629
rect 13515 30549 14039 30565
rect 13515 30485 13520 30549
rect 13584 30485 13610 30549
rect 13674 30485 13700 30549
rect 13764 30485 13790 30549
rect 13854 30485 13880 30549
rect 13944 30485 13970 30549
rect 14034 30485 14039 30549
rect 13515 30469 14039 30485
rect 13515 30405 13520 30469
rect 13584 30405 13610 30469
rect 13674 30405 13700 30469
rect 13764 30405 13790 30469
rect 13854 30405 13880 30469
rect 13944 30405 13970 30469
rect 14034 30405 14039 30469
rect 13515 30389 14039 30405
rect 13515 30325 13520 30389
rect 13584 30325 13610 30389
rect 13674 30325 13700 30389
rect 13764 30325 13790 30389
rect 13854 30325 13880 30389
rect 13944 30325 13970 30389
rect 14034 30325 14039 30389
rect 13515 30309 14039 30325
rect 13515 30245 13520 30309
rect 13584 30245 13610 30309
rect 13674 30245 13700 30309
rect 13764 30245 13790 30309
rect 13854 30245 13880 30309
rect 13944 30245 13970 30309
rect 14034 30245 14039 30309
rect 13515 30229 14039 30245
rect 13515 30165 13520 30229
rect 13584 30165 13610 30229
rect 13674 30165 13700 30229
rect 13764 30165 13790 30229
rect 13854 30165 13880 30229
rect 13944 30165 13970 30229
rect 14034 30165 14039 30229
rect 13515 30149 14039 30165
rect 13515 30085 13520 30149
rect 13584 30085 13610 30149
rect 13674 30085 13700 30149
rect 13764 30085 13790 30149
rect 13854 30085 13880 30149
rect 13944 30085 13970 30149
rect 14034 30085 14039 30149
rect 13515 30069 14039 30085
rect 13515 30005 13520 30069
rect 13584 30005 13610 30069
rect 13674 30005 13700 30069
rect 13764 30005 13790 30069
rect 13854 30005 13880 30069
rect 13944 30005 13970 30069
rect 14034 30005 14039 30069
rect 13515 29989 14039 30005
rect 13515 29925 13520 29989
rect 13584 29925 13610 29989
rect 13674 29925 13700 29989
rect 13764 29925 13790 29989
rect 13854 29925 13880 29989
rect 13944 29925 13970 29989
rect 14034 29925 14039 29989
rect 13515 29909 14039 29925
rect 13515 29845 13520 29909
rect 13584 29845 13610 29909
rect 13674 29845 13700 29909
rect 13764 29845 13790 29909
rect 13854 29845 13880 29909
rect 13944 29845 13970 29909
rect 14034 29845 14039 29909
rect 13515 29829 14039 29845
rect 13515 29765 13520 29829
rect 13584 29765 13610 29829
rect 13674 29765 13700 29829
rect 13764 29765 13790 29829
rect 13854 29765 13880 29829
rect 13944 29765 13970 29829
rect 14034 29765 14039 29829
rect 13515 29749 14039 29765
rect 13515 29685 13520 29749
rect 13584 29685 13610 29749
rect 13674 29685 13700 29749
rect 13764 29685 13790 29749
rect 13854 29685 13880 29749
rect 13944 29685 13970 29749
rect 14034 29685 14039 29749
rect 13515 29669 14039 29685
rect 13515 29605 13520 29669
rect 13584 29605 13610 29669
rect 13674 29605 13700 29669
rect 13764 29605 13790 29669
rect 13854 29605 13880 29669
rect 13944 29605 13970 29669
rect 14034 29605 14039 29669
rect 13515 29589 14039 29605
rect 13515 29525 13520 29589
rect 13584 29525 13610 29589
rect 13674 29525 13700 29589
rect 13764 29525 13790 29589
rect 13854 29525 13880 29589
rect 13944 29525 13970 29589
rect 14034 29525 14039 29589
rect 13515 29509 14039 29525
rect 13515 29445 13520 29509
rect 13584 29445 13610 29509
rect 13674 29445 13700 29509
rect 13764 29445 13790 29509
rect 13854 29445 13880 29509
rect 13944 29445 13970 29509
rect 14034 29445 14039 29509
rect 13515 29429 14039 29445
rect 13515 29365 13520 29429
rect 13584 29365 13610 29429
rect 13674 29365 13700 29429
rect 13764 29365 13790 29429
rect 13854 29365 13880 29429
rect 13944 29365 13970 29429
rect 14034 29365 14039 29429
rect 13515 29349 14039 29365
rect 13515 29285 13520 29349
rect 13584 29285 13610 29349
rect 13674 29285 13700 29349
rect 13764 29285 13790 29349
rect 13854 29285 13880 29349
rect 13944 29285 13970 29349
rect 14034 29285 14039 29349
rect 13515 29269 14039 29285
rect 13515 29205 13520 29269
rect 13584 29205 13610 29269
rect 13674 29205 13700 29269
rect 13764 29205 13790 29269
rect 13854 29205 13880 29269
rect 13944 29205 13970 29269
rect 14034 29205 14039 29269
rect 13515 29189 14039 29205
rect 13515 29125 13520 29189
rect 13584 29125 13610 29189
rect 13674 29125 13700 29189
rect 13764 29125 13790 29189
rect 13854 29125 13880 29189
rect 13944 29125 13970 29189
rect 14034 29125 14039 29189
rect 13515 29109 14039 29125
rect 13515 29045 13520 29109
rect 13584 29045 13610 29109
rect 13674 29045 13700 29109
rect 13764 29045 13790 29109
rect 13854 29045 13880 29109
rect 13944 29045 13970 29109
rect 14034 29045 14039 29109
rect 13515 29029 14039 29045
rect 13515 28965 13520 29029
rect 13584 28965 13610 29029
rect 13674 28965 13700 29029
rect 13764 28965 13790 29029
rect 13854 28965 13880 29029
rect 13944 28965 13970 29029
rect 14034 28965 14039 29029
rect 13515 28949 14039 28965
rect 13515 28885 13520 28949
rect 13584 28885 13610 28949
rect 13674 28885 13700 28949
rect 13764 28885 13790 28949
rect 13854 28885 13880 28949
rect 13944 28885 13970 28949
rect 14034 28885 14039 28949
rect 13515 28869 14039 28885
rect 13515 28805 13520 28869
rect 13584 28805 13610 28869
rect 13674 28805 13700 28869
rect 13764 28805 13790 28869
rect 13854 28805 13880 28869
rect 13944 28805 13970 28869
rect 14034 28805 14039 28869
rect 13515 28789 14039 28805
rect 13515 28725 13520 28789
rect 13584 28725 13610 28789
rect 13674 28725 13700 28789
rect 13764 28725 13790 28789
rect 13854 28725 13880 28789
rect 13944 28725 13970 28789
rect 14034 28725 14039 28789
rect 13515 28709 14039 28725
rect 13515 28645 13520 28709
rect 13584 28645 13610 28709
rect 13674 28645 13700 28709
rect 13764 28645 13790 28709
rect 13854 28645 13880 28709
rect 13944 28645 13970 28709
rect 14034 28645 14039 28709
rect 13515 28629 14039 28645
rect 13515 28565 13520 28629
rect 13584 28565 13610 28629
rect 13674 28565 13700 28629
rect 13764 28565 13790 28629
rect 13854 28565 13880 28629
rect 13944 28565 13970 28629
rect 14034 28565 14039 28629
rect 13515 28549 14039 28565
rect 13515 28485 13520 28549
rect 13584 28485 13610 28549
rect 13674 28485 13700 28549
rect 13764 28485 13790 28549
rect 13854 28485 13880 28549
rect 13944 28485 13970 28549
rect 14034 28485 14039 28549
rect 13515 28469 14039 28485
rect 13515 28405 13520 28469
rect 13584 28405 13610 28469
rect 13674 28405 13700 28469
rect 13764 28405 13790 28469
rect 13854 28405 13880 28469
rect 13944 28405 13970 28469
rect 14034 28405 14039 28469
rect 13515 28389 14039 28405
rect 13515 28325 13520 28389
rect 13584 28325 13610 28389
rect 13674 28325 13700 28389
rect 13764 28325 13790 28389
rect 13854 28325 13880 28389
rect 13944 28325 13970 28389
rect 14034 28325 14039 28389
rect 13515 28309 14039 28325
rect 13515 28245 13520 28309
rect 13584 28245 13610 28309
rect 13674 28245 13700 28309
rect 13764 28245 13790 28309
rect 13854 28245 13880 28309
rect 13944 28245 13970 28309
rect 14034 28245 14039 28309
rect 13515 28229 14039 28245
rect 13515 28165 13520 28229
rect 13584 28165 13610 28229
rect 13674 28165 13700 28229
rect 13764 28165 13790 28229
rect 13854 28165 13880 28229
rect 13944 28165 13970 28229
rect 14034 28165 14039 28229
rect 13515 28149 14039 28165
rect 13515 28085 13520 28149
rect 13584 28085 13610 28149
rect 13674 28085 13700 28149
rect 13764 28085 13790 28149
rect 13854 28085 13880 28149
rect 13944 28085 13970 28149
rect 14034 28085 14039 28149
rect 13515 28069 14039 28085
rect 13515 28005 13520 28069
rect 13584 28005 13610 28069
rect 13674 28005 13700 28069
rect 13764 28005 13790 28069
rect 13854 28005 13880 28069
rect 13944 28005 13970 28069
rect 14034 28005 14039 28069
rect 13515 27989 14039 28005
rect 13515 27925 13520 27989
rect 13584 27925 13610 27989
rect 13674 27925 13700 27989
rect 13764 27925 13790 27989
rect 13854 27925 13880 27989
rect 13944 27925 13970 27989
rect 14034 27925 14039 27989
rect 13515 27909 14039 27925
rect 13515 27845 13520 27909
rect 13584 27845 13610 27909
rect 13674 27845 13700 27909
rect 13764 27845 13790 27909
rect 13854 27845 13880 27909
rect 13944 27845 13970 27909
rect 14034 27845 14039 27909
rect 13515 27829 14039 27845
rect 13515 27765 13520 27829
rect 13584 27765 13610 27829
rect 13674 27765 13700 27829
rect 13764 27765 13790 27829
rect 13854 27765 13880 27829
rect 13944 27765 13970 27829
rect 14034 27765 14039 27829
rect 13515 27749 14039 27765
rect 13515 27685 13520 27749
rect 13584 27685 13610 27749
rect 13674 27685 13700 27749
rect 13764 27685 13790 27749
rect 13854 27685 13880 27749
rect 13944 27685 13970 27749
rect 14034 27685 14039 27749
rect 13515 27669 14039 27685
rect 13515 27605 13520 27669
rect 13584 27605 13610 27669
rect 13674 27605 13700 27669
rect 13764 27605 13790 27669
rect 13854 27605 13880 27669
rect 13944 27605 13970 27669
rect 14034 27605 14039 27669
rect 13515 27589 14039 27605
rect 13515 27525 13520 27589
rect 13584 27525 13610 27589
rect 13674 27525 13700 27589
rect 13764 27525 13790 27589
rect 13854 27525 13880 27589
rect 13944 27525 13970 27589
rect 14034 27525 14039 27589
rect 13515 27509 14039 27525
rect 13515 27445 13520 27509
rect 13584 27445 13610 27509
rect 13674 27445 13700 27509
rect 13764 27445 13790 27509
rect 13854 27445 13880 27509
rect 13944 27445 13970 27509
rect 14034 27445 14039 27509
rect 13515 27429 14039 27445
rect 13515 27365 13520 27429
rect 13584 27365 13610 27429
rect 13674 27365 13700 27429
rect 13764 27365 13790 27429
rect 13854 27365 13880 27429
rect 13944 27365 13970 27429
rect 14034 27365 14039 27429
rect 13515 27349 14039 27365
rect 13515 27285 13520 27349
rect 13584 27285 13610 27349
rect 13674 27285 13700 27349
rect 13764 27285 13790 27349
rect 13854 27285 13880 27349
rect 13944 27285 13970 27349
rect 14034 27285 14039 27349
rect 13515 27269 14039 27285
rect 13515 27205 13520 27269
rect 13584 27205 13610 27269
rect 13674 27205 13700 27269
rect 13764 27205 13790 27269
rect 13854 27205 13880 27269
rect 13944 27205 13970 27269
rect 14034 27205 14039 27269
rect 13515 27189 14039 27205
rect 13515 27125 13520 27189
rect 13584 27125 13610 27189
rect 13674 27125 13700 27189
rect 13764 27125 13790 27189
rect 13854 27125 13880 27189
rect 13944 27125 13970 27189
rect 14034 27125 14039 27189
rect 13515 27109 14039 27125
rect 13515 27045 13520 27109
rect 13584 27045 13610 27109
rect 13674 27045 13700 27109
rect 13764 27045 13790 27109
rect 13854 27045 13880 27109
rect 13944 27045 13970 27109
rect 14034 27045 14039 27109
rect 13515 27029 14039 27045
rect 13515 26965 13520 27029
rect 13584 26965 13610 27029
rect 13674 26965 13700 27029
rect 13764 26965 13790 27029
rect 13854 26965 13880 27029
rect 13944 26965 13970 27029
rect 14034 26965 14039 27029
rect 13515 26949 14039 26965
rect 13515 26885 13520 26949
rect 13584 26885 13610 26949
rect 13674 26885 13700 26949
rect 13764 26885 13790 26949
rect 13854 26885 13880 26949
rect 13944 26885 13970 26949
rect 14034 26885 14039 26949
rect 13515 26869 14039 26885
rect 13515 26805 13520 26869
rect 13584 26805 13610 26869
rect 13674 26805 13700 26869
rect 13764 26805 13790 26869
rect 13854 26805 13880 26869
rect 13944 26805 13970 26869
rect 14034 26805 14039 26869
rect 13515 26789 14039 26805
rect 13515 26725 13520 26789
rect 13584 26725 13610 26789
rect 13674 26725 13700 26789
rect 13764 26725 13790 26789
rect 13854 26725 13880 26789
rect 13944 26725 13970 26789
rect 14034 26725 14039 26789
rect 13515 26709 14039 26725
rect 13515 26645 13520 26709
rect 13584 26645 13610 26709
rect 13674 26645 13700 26709
rect 13764 26645 13790 26709
rect 13854 26645 13880 26709
rect 13944 26645 13970 26709
rect 14034 26645 14039 26709
rect 13515 26629 14039 26645
rect 13515 26565 13520 26629
rect 13584 26565 13610 26629
rect 13674 26565 13700 26629
rect 13764 26565 13790 26629
rect 13854 26565 13880 26629
rect 13944 26565 13970 26629
rect 14034 26565 14039 26629
rect 13515 26549 14039 26565
rect 13515 26485 13520 26549
rect 13584 26485 13610 26549
rect 13674 26485 13700 26549
rect 13764 26485 13790 26549
rect 13854 26485 13880 26549
rect 13944 26485 13970 26549
rect 14034 26485 14039 26549
rect 13515 26469 14039 26485
rect 13515 26405 13520 26469
rect 13584 26405 13610 26469
rect 13674 26405 13700 26469
rect 13764 26405 13790 26469
rect 13854 26405 13880 26469
rect 13944 26405 13970 26469
rect 14034 26405 14039 26469
rect 13515 26389 14039 26405
rect 13515 26325 13520 26389
rect 13584 26325 13610 26389
rect 13674 26325 13700 26389
rect 13764 26325 13790 26389
rect 13854 26325 13880 26389
rect 13944 26325 13970 26389
rect 14034 26325 14039 26389
rect 13515 26309 14039 26325
rect 13515 26245 13520 26309
rect 13584 26245 13610 26309
rect 13674 26245 13700 26309
rect 13764 26245 13790 26309
rect 13854 26245 13880 26309
rect 13944 26245 13970 26309
rect 14034 26245 14039 26309
rect 13515 26229 14039 26245
rect 13515 26165 13520 26229
rect 13584 26165 13610 26229
rect 13674 26165 13700 26229
rect 13764 26165 13790 26229
rect 13854 26165 13880 26229
rect 13944 26165 13970 26229
rect 14034 26165 14039 26229
rect 13515 26149 14039 26165
rect 13515 26085 13520 26149
rect 13584 26085 13610 26149
rect 13674 26085 13700 26149
rect 13764 26085 13790 26149
rect 13854 26085 13880 26149
rect 13944 26085 13970 26149
rect 14034 26085 14039 26149
rect 13515 26069 14039 26085
rect 13515 26005 13520 26069
rect 13584 26005 13610 26069
rect 13674 26005 13700 26069
rect 13764 26005 13790 26069
rect 13854 26005 13880 26069
rect 13944 26005 13970 26069
rect 14034 26005 14039 26069
rect 13515 25989 14039 26005
rect 13515 25925 13520 25989
rect 13584 25925 13610 25989
rect 13674 25925 13700 25989
rect 13764 25925 13790 25989
rect 13854 25925 13880 25989
rect 13944 25925 13970 25989
rect 14034 25925 14039 25989
rect 13515 25909 14039 25925
rect 13515 25845 13520 25909
rect 13584 25845 13610 25909
rect 13674 25845 13700 25909
rect 13764 25845 13790 25909
rect 13854 25845 13880 25909
rect 13944 25845 13970 25909
rect 14034 25845 14039 25909
rect 13515 25829 14039 25845
rect 13515 25765 13520 25829
rect 13584 25765 13610 25829
rect 13674 25765 13700 25829
rect 13764 25765 13790 25829
rect 13854 25765 13880 25829
rect 13944 25765 13970 25829
rect 14034 25765 14039 25829
rect 13515 25749 14039 25765
rect 13515 25685 13520 25749
rect 13584 25685 13610 25749
rect 13674 25685 13700 25749
rect 13764 25685 13790 25749
rect 13854 25685 13880 25749
rect 13944 25685 13970 25749
rect 14034 25685 14039 25749
rect 13515 25669 14039 25685
rect 13515 25605 13520 25669
rect 13584 25605 13610 25669
rect 13674 25605 13700 25669
rect 13764 25605 13790 25669
rect 13854 25605 13880 25669
rect 13944 25605 13970 25669
rect 14034 25605 14039 25669
rect 13515 25589 14039 25605
rect 13515 25525 13520 25589
rect 13584 25525 13610 25589
rect 13674 25525 13700 25589
rect 13764 25525 13790 25589
rect 13854 25525 13880 25589
rect 13944 25525 13970 25589
rect 14034 25525 14039 25589
rect 13515 25509 14039 25525
rect 13515 25445 13520 25509
rect 13584 25445 13610 25509
rect 13674 25445 13700 25509
rect 13764 25445 13790 25509
rect 13854 25445 13880 25509
rect 13944 25445 13970 25509
rect 14034 25445 14039 25509
rect 13515 25429 14039 25445
rect 13515 25365 13520 25429
rect 13584 25365 13610 25429
rect 13674 25365 13700 25429
rect 13764 25365 13790 25429
rect 13854 25365 13880 25429
rect 13944 25365 13970 25429
rect 14034 25365 14039 25429
rect 13515 25349 14039 25365
rect 13515 25285 13520 25349
rect 13584 25285 13610 25349
rect 13674 25285 13700 25349
rect 13764 25285 13790 25349
rect 13854 25285 13880 25349
rect 13944 25285 13970 25349
rect 14034 25285 14039 25349
rect 13515 25269 14039 25285
rect 13515 25205 13520 25269
rect 13584 25205 13610 25269
rect 13674 25205 13700 25269
rect 13764 25205 13790 25269
rect 13854 25205 13880 25269
rect 13944 25205 13970 25269
rect 14034 25205 14039 25269
rect 13515 25189 14039 25205
rect 13515 25125 13520 25189
rect 13584 25125 13610 25189
rect 13674 25125 13700 25189
rect 13764 25125 13790 25189
rect 13854 25125 13880 25189
rect 13944 25125 13970 25189
rect 14034 25125 14039 25189
rect 13515 25109 14039 25125
rect 13515 25045 13520 25109
rect 13584 25045 13610 25109
rect 13674 25045 13700 25109
rect 13764 25045 13790 25109
rect 13854 25045 13880 25109
rect 13944 25045 13970 25109
rect 14034 25045 14039 25109
rect 13515 25029 14039 25045
rect 13515 24965 13520 25029
rect 13584 24965 13610 25029
rect 13674 24965 13700 25029
rect 13764 24965 13790 25029
rect 13854 24965 13880 25029
rect 13944 24965 13970 25029
rect 14034 24965 14039 25029
rect 13515 24949 14039 24965
rect 13515 24885 13520 24949
rect 13584 24885 13610 24949
rect 13674 24885 13700 24949
rect 13764 24885 13790 24949
rect 13854 24885 13880 24949
rect 13944 24885 13970 24949
rect 14034 24885 14039 24949
rect 13515 24869 14039 24885
rect 13515 24805 13520 24869
rect 13584 24805 13610 24869
rect 13674 24805 13700 24869
rect 13764 24805 13790 24869
rect 13854 24805 13880 24869
rect 13944 24805 13970 24869
rect 14034 24805 14039 24869
rect 13515 24789 14039 24805
rect 13515 24725 13520 24789
rect 13584 24725 13610 24789
rect 13674 24725 13700 24789
rect 13764 24725 13790 24789
rect 13854 24725 13880 24789
rect 13944 24725 13970 24789
rect 14034 24725 14039 24789
rect 13515 24709 14039 24725
rect 13515 24645 13520 24709
rect 13584 24645 13610 24709
rect 13674 24645 13700 24709
rect 13764 24645 13790 24709
rect 13854 24645 13880 24709
rect 13944 24645 13970 24709
rect 14034 24645 14039 24709
rect 13515 24629 14039 24645
rect 13515 24565 13520 24629
rect 13584 24565 13610 24629
rect 13674 24565 13700 24629
rect 13764 24565 13790 24629
rect 13854 24565 13880 24629
rect 13944 24565 13970 24629
rect 14034 24565 14039 24629
rect 13515 24549 14039 24565
rect 13515 24485 13520 24549
rect 13584 24485 13610 24549
rect 13674 24485 13700 24549
rect 13764 24485 13790 24549
rect 13854 24485 13880 24549
rect 13944 24485 13970 24549
rect 14034 24485 14039 24549
rect 13515 24469 14039 24485
rect 13515 24405 13520 24469
rect 13584 24405 13610 24469
rect 13674 24405 13700 24469
rect 13764 24405 13790 24469
rect 13854 24405 13880 24469
rect 13944 24405 13970 24469
rect 14034 24405 14039 24469
rect 13515 24389 14039 24405
rect 13515 24325 13520 24389
rect 13584 24325 13610 24389
rect 13674 24325 13700 24389
rect 13764 24325 13790 24389
rect 13854 24325 13880 24389
rect 13944 24325 13970 24389
rect 14034 24325 14039 24389
rect 13515 24309 14039 24325
rect 13515 24245 13520 24309
rect 13584 24245 13610 24309
rect 13674 24245 13700 24309
rect 13764 24245 13790 24309
rect 13854 24245 13880 24309
rect 13944 24245 13970 24309
rect 14034 24245 14039 24309
rect 13515 24229 14039 24245
rect 13515 24165 13520 24229
rect 13584 24165 13610 24229
rect 13674 24165 13700 24229
rect 13764 24165 13790 24229
rect 13854 24165 13880 24229
rect 13944 24165 13970 24229
rect 14034 24165 14039 24229
rect 13515 24149 14039 24165
rect 13515 24085 13520 24149
rect 13584 24085 13610 24149
rect 13674 24085 13700 24149
rect 13764 24085 13790 24149
rect 13854 24085 13880 24149
rect 13944 24085 13970 24149
rect 14034 24085 14039 24149
rect 13515 24069 14039 24085
rect 13515 24005 13520 24069
rect 13584 24005 13610 24069
rect 13674 24005 13700 24069
rect 13764 24005 13790 24069
rect 13854 24005 13880 24069
rect 13944 24005 13970 24069
rect 14034 24005 14039 24069
rect 13515 23989 14039 24005
rect 13515 23925 13520 23989
rect 13584 23925 13610 23989
rect 13674 23925 13700 23989
rect 13764 23925 13790 23989
rect 13854 23925 13880 23989
rect 13944 23925 13970 23989
rect 14034 23925 14039 23989
rect 13515 23909 14039 23925
rect 13515 23845 13520 23909
rect 13584 23845 13610 23909
rect 13674 23845 13700 23909
rect 13764 23845 13790 23909
rect 13854 23845 13880 23909
rect 13944 23845 13970 23909
rect 14034 23845 14039 23909
rect 13515 23829 14039 23845
rect 13515 23765 13520 23829
rect 13584 23765 13610 23829
rect 13674 23765 13700 23829
rect 13764 23765 13790 23829
rect 13854 23765 13880 23829
rect 13944 23765 13970 23829
rect 14034 23765 14039 23829
rect 13515 23749 14039 23765
rect 13515 23685 13520 23749
rect 13584 23685 13610 23749
rect 13674 23685 13700 23749
rect 13764 23685 13790 23749
rect 13854 23685 13880 23749
rect 13944 23685 13970 23749
rect 14034 23685 14039 23749
rect 13515 23669 14039 23685
rect 13515 23605 13520 23669
rect 13584 23605 13610 23669
rect 13674 23605 13700 23669
rect 13764 23605 13790 23669
rect 13854 23605 13880 23669
rect 13944 23605 13970 23669
rect 14034 23605 14039 23669
rect 13515 23589 14039 23605
rect 13515 23525 13520 23589
rect 13584 23525 13610 23589
rect 13674 23525 13700 23589
rect 13764 23525 13790 23589
rect 13854 23525 13880 23589
rect 13944 23525 13970 23589
rect 14034 23525 14039 23589
rect 13515 23509 14039 23525
rect 13515 23445 13520 23509
rect 13584 23445 13610 23509
rect 13674 23445 13700 23509
rect 13764 23445 13790 23509
rect 13854 23445 13880 23509
rect 13944 23445 13970 23509
rect 14034 23445 14039 23509
rect 13515 23429 14039 23445
rect 13515 23365 13520 23429
rect 13584 23365 13610 23429
rect 13674 23365 13700 23429
rect 13764 23365 13790 23429
rect 13854 23365 13880 23429
rect 13944 23365 13970 23429
rect 14034 23365 14039 23429
rect 13515 23349 14039 23365
rect 13515 23285 13520 23349
rect 13584 23285 13610 23349
rect 13674 23285 13700 23349
rect 13764 23285 13790 23349
rect 13854 23285 13880 23349
rect 13944 23285 13970 23349
rect 14034 23285 14039 23349
rect 13515 23268 14039 23285
rect 13515 23204 13520 23268
rect 13584 23204 13610 23268
rect 13674 23204 13700 23268
rect 13764 23204 13790 23268
rect 13854 23204 13880 23268
rect 13944 23204 13970 23268
rect 14034 23204 14039 23268
rect 13515 23187 14039 23204
rect 13515 23123 13520 23187
rect 13584 23123 13610 23187
rect 13674 23123 13700 23187
rect 13764 23123 13790 23187
rect 13854 23123 13880 23187
rect 13944 23123 13970 23187
rect 14034 23123 14039 23187
rect 13515 23106 14039 23123
rect 13515 23042 13520 23106
rect 13584 23042 13610 23106
rect 13674 23042 13700 23106
rect 13764 23042 13790 23106
rect 13854 23042 13880 23106
rect 13944 23042 13970 23106
rect 14034 23042 14039 23106
rect 13515 23025 14039 23042
rect 13515 22961 13520 23025
rect 13584 22961 13610 23025
rect 13674 22961 13700 23025
rect 13764 22961 13790 23025
rect 13854 22961 13880 23025
rect 13944 22961 13970 23025
rect 14034 22961 14039 23025
rect 13515 22944 14039 22961
rect 13515 22880 13520 22944
rect 13584 22880 13610 22944
rect 13674 22880 13700 22944
rect 13764 22880 13790 22944
rect 13854 22880 13880 22944
rect 13944 22880 13970 22944
rect 14034 22880 14039 22944
rect 13515 22863 14039 22880
rect 13515 22799 13520 22863
rect 13584 22799 13610 22863
rect 13674 22799 13700 22863
rect 13764 22799 13790 22863
rect 13854 22799 13880 22863
rect 13944 22799 13970 22863
rect 14034 22799 14039 22863
rect 13515 22782 14039 22799
rect 13515 22718 13520 22782
rect 13584 22718 13610 22782
rect 13674 22718 13700 22782
rect 13764 22718 13790 22782
rect 13854 22718 13880 22782
rect 13944 22718 13970 22782
rect 14034 22718 14039 22782
rect 13515 22701 14039 22718
rect 13515 22637 13520 22701
rect 13584 22637 13610 22701
rect 13674 22637 13700 22701
rect 13764 22637 13790 22701
rect 13854 22637 13880 22701
rect 13944 22637 13970 22701
rect 14034 22637 14039 22701
rect 13515 22620 14039 22637
rect 13515 22556 13520 22620
rect 13584 22556 13610 22620
rect 13674 22556 13700 22620
rect 13764 22556 13790 22620
rect 13854 22556 13880 22620
rect 13944 22556 13970 22620
rect 14034 22556 14039 22620
rect 13515 22539 14039 22556
rect 13515 22475 13520 22539
rect 13584 22475 13610 22539
rect 13674 22475 13700 22539
rect 13764 22475 13790 22539
rect 13854 22475 13880 22539
rect 13944 22475 13970 22539
rect 14034 22475 14039 22539
rect 13515 22458 14039 22475
rect 13515 22394 13520 22458
rect 13584 22394 13610 22458
rect 13674 22394 13700 22458
rect 13764 22394 13790 22458
rect 13854 22394 13880 22458
rect 13944 22394 13970 22458
rect 14034 22394 14039 22458
rect 13515 22377 14039 22394
rect 13515 22313 13520 22377
rect 13584 22313 13610 22377
rect 13674 22313 13700 22377
rect 13764 22313 13790 22377
rect 13854 22313 13880 22377
rect 13944 22313 13970 22377
rect 14034 22313 14039 22377
rect 13515 22296 14039 22313
rect 13515 22232 13520 22296
rect 13584 22232 13610 22296
rect 13674 22232 13700 22296
rect 13764 22232 13790 22296
rect 13854 22232 13880 22296
rect 13944 22232 13970 22296
rect 14034 22232 14039 22296
rect 13515 22215 14039 22232
rect 13515 22151 13520 22215
rect 13584 22151 13610 22215
rect 13674 22151 13700 22215
rect 13764 22151 13790 22215
rect 13854 22151 13880 22215
rect 13944 22151 13970 22215
rect 14034 22151 14039 22215
rect 13515 22134 14039 22151
rect 13515 22070 13520 22134
rect 13584 22070 13610 22134
rect 13674 22070 13700 22134
rect 13764 22070 13790 22134
rect 13854 22070 13880 22134
rect 13944 22070 13970 22134
rect 14034 22070 14039 22134
rect 13515 22053 14039 22070
rect 13515 21989 13520 22053
rect 13584 21989 13610 22053
rect 13674 21989 13700 22053
rect 13764 21989 13790 22053
rect 13854 21989 13880 22053
rect 13944 21989 13970 22053
rect 14034 21989 14039 22053
rect 13515 21972 14039 21989
rect 13515 21908 13520 21972
rect 13584 21908 13610 21972
rect 13674 21908 13700 21972
rect 13764 21908 13790 21972
rect 13854 21908 13880 21972
rect 13944 21908 13970 21972
rect 14034 21908 14039 21972
rect 13515 21891 14039 21908
rect 13515 21827 13520 21891
rect 13584 21827 13610 21891
rect 13674 21827 13700 21891
rect 13764 21827 13790 21891
rect 13854 21827 13880 21891
rect 13944 21827 13970 21891
rect 14034 21827 14039 21891
rect 13515 21810 14039 21827
rect 13515 21746 13520 21810
rect 13584 21746 13610 21810
rect 13674 21746 13700 21810
rect 13764 21746 13790 21810
rect 13854 21746 13880 21810
rect 13944 21746 13970 21810
rect 14034 21746 14039 21810
rect 13515 21729 14039 21746
rect 13515 21665 13520 21729
rect 13584 21665 13610 21729
rect 13674 21665 13700 21729
rect 13764 21665 13790 21729
rect 13854 21665 13880 21729
rect 13944 21665 13970 21729
rect 14034 21665 14039 21729
rect 13515 21648 14039 21665
rect 13515 21584 13520 21648
rect 13584 21584 13610 21648
rect 13674 21584 13700 21648
rect 13764 21584 13790 21648
rect 13854 21584 13880 21648
rect 13944 21584 13970 21648
rect 14034 21584 14039 21648
rect 13515 21567 14039 21584
rect 13515 21503 13520 21567
rect 13584 21503 13610 21567
rect 13674 21503 13700 21567
rect 13764 21503 13790 21567
rect 13854 21503 13880 21567
rect 13944 21503 13970 21567
rect 14034 21503 14039 21567
rect 13515 21486 14039 21503
rect 13515 21422 13520 21486
rect 13584 21422 13610 21486
rect 13674 21422 13700 21486
rect 13764 21422 13790 21486
rect 13854 21422 13880 21486
rect 13944 21422 13970 21486
rect 14034 21422 14039 21486
rect 13515 21405 14039 21422
rect 13515 21341 13520 21405
rect 13584 21341 13610 21405
rect 13674 21341 13700 21405
rect 13764 21341 13790 21405
rect 13854 21341 13880 21405
rect 13944 21341 13970 21405
rect 14034 21341 14039 21405
rect 13515 21324 14039 21341
rect 13515 21260 13520 21324
rect 13584 21260 13610 21324
rect 13674 21260 13700 21324
rect 13764 21260 13790 21324
rect 13854 21260 13880 21324
rect 13944 21260 13970 21324
rect 14034 21260 14039 21324
rect 13515 21243 14039 21260
rect 13515 21179 13520 21243
rect 13584 21179 13610 21243
rect 13674 21179 13700 21243
rect 13764 21179 13790 21243
rect 13854 21179 13880 21243
rect 13944 21179 13970 21243
rect 14034 21179 14039 21243
rect 13515 21162 14039 21179
rect 13515 21098 13520 21162
rect 13584 21098 13610 21162
rect 13674 21098 13700 21162
rect 13764 21098 13790 21162
rect 13854 21098 13880 21162
rect 13944 21098 13970 21162
rect 14034 21098 14039 21162
rect 13515 21081 14039 21098
rect 13515 21017 13520 21081
rect 13584 21017 13610 21081
rect 13674 21017 13700 21081
rect 13764 21017 13790 21081
rect 13854 21017 13880 21081
rect 13944 21017 13970 21081
rect 14034 21017 14039 21081
rect 13515 21000 14039 21017
rect 13515 20972 13520 21000
rect 1496 20939 1596 20972
rect 1496 20936 1531 20939
rect 977 20919 1531 20936
rect 977 20855 982 20919
rect 1046 20855 1072 20919
rect 1136 20855 1162 20919
rect 1226 20855 1252 20919
rect 1316 20855 1342 20919
rect 1406 20855 1432 20919
rect 1496 20875 1531 20919
rect 1595 20875 1596 20939
rect 1496 20855 1596 20875
rect 977 20854 1596 20855
rect 1471 20842 1596 20854
rect 13420 20939 13520 20972
rect 13420 20875 13421 20939
rect 13485 20936 13520 20939
rect 13584 20936 13610 21000
rect 13674 20936 13700 21000
rect 13764 20936 13790 21000
rect 13854 20936 13880 21000
rect 13944 20936 13970 21000
rect 14034 20936 14039 21000
rect 13485 20919 14039 20936
rect 13485 20875 13520 20919
rect 13420 20855 13520 20875
rect 13584 20855 13610 20919
rect 13674 20855 13700 20919
rect 13764 20855 13790 20919
rect 13854 20855 13880 20919
rect 13944 20855 13970 20919
rect 14034 20855 14039 20919
rect 13420 20854 14039 20855
rect 13420 20842 13545 20854
rect 1311 20825 1736 20827
rect 1140 20783 1265 20816
rect 1140 20719 1141 20783
rect 1205 20719 1265 20783
rect 1140 20686 1265 20719
rect 1311 20761 1312 20825
rect 1376 20761 1401 20825
rect 1465 20761 1491 20825
rect 1555 20761 1581 20825
rect 1645 20761 1671 20825
rect 1735 20761 1736 20825
rect 1311 20709 1736 20761
rect 1311 20645 1312 20709
rect 1376 20645 1401 20709
rect 1465 20645 1491 20709
rect 1555 20645 1581 20709
rect 1645 20645 1671 20709
rect 1735 20645 1736 20709
rect 13280 20825 13705 20827
rect 13280 20761 13281 20825
rect 13345 20761 13371 20825
rect 13435 20761 13461 20825
rect 13525 20761 13551 20825
rect 13615 20761 13640 20825
rect 13704 20761 13705 20825
rect 13280 20709 13705 20761
rect 1311 20593 1736 20645
rect 1311 20529 1312 20593
rect 1376 20529 1401 20593
rect 1465 20529 1491 20593
rect 1555 20529 1581 20593
rect 1645 20529 1671 20593
rect 1735 20529 1736 20593
rect 1752 20631 1877 20664
rect 1752 20567 1812 20631
rect 1876 20567 1877 20631
rect 1752 20534 1877 20567
rect 13139 20631 13264 20664
rect 13139 20567 13140 20631
rect 13204 20567 13264 20631
rect 13139 20534 13264 20567
rect 13280 20645 13281 20709
rect 13345 20645 13371 20709
rect 13435 20645 13461 20709
rect 13525 20645 13551 20709
rect 13615 20645 13640 20709
rect 13704 20645 13705 20709
rect 13719 20823 13843 20824
rect 13719 20759 13749 20823
rect 13813 20759 13843 20823
rect 13719 20712 13843 20759
rect 13849 20816 13916 20849
rect 13849 20752 13851 20816
rect 13915 20752 13916 20816
rect 13849 20719 13916 20752
rect 13719 20648 13749 20712
rect 13813 20648 13843 20712
rect 13719 20647 13843 20648
rect 13280 20593 13705 20645
rect 1311 20527 1736 20529
rect 13280 20529 13281 20593
rect 13345 20529 13371 20593
rect 13435 20529 13461 20593
rect 13525 20529 13551 20593
rect 13615 20529 13640 20593
rect 13704 20529 13705 20593
rect 13280 20527 13705 20529
rect 1631 20505 2056 20507
rect 1464 20469 1589 20502
rect 1464 20405 1524 20469
rect 1588 20405 1589 20469
rect 1464 20372 1589 20405
rect 1631 20441 1632 20505
rect 1696 20441 1721 20505
rect 1785 20441 1811 20505
rect 1875 20441 1901 20505
rect 1965 20441 1991 20505
rect 2055 20441 2056 20505
rect 1631 20389 2056 20441
rect 1631 20325 1632 20389
rect 1696 20325 1721 20389
rect 1785 20325 1811 20389
rect 1875 20325 1901 20389
rect 1965 20325 1991 20389
rect 2055 20325 2056 20389
rect 12960 20505 13385 20507
rect 12960 20441 12961 20505
rect 13025 20441 13051 20505
rect 13115 20441 13141 20505
rect 13205 20441 13231 20505
rect 13295 20441 13320 20505
rect 13384 20441 13385 20505
rect 12960 20389 13385 20441
rect 1631 20273 2056 20325
rect 1631 20209 1632 20273
rect 1696 20209 1721 20273
rect 1785 20209 1811 20273
rect 1875 20209 1901 20273
rect 1965 20209 1991 20273
rect 2055 20209 2056 20273
rect 2077 20306 2202 20339
rect 2077 20242 2137 20306
rect 2201 20242 2202 20306
rect 2077 20209 2202 20242
rect 12814 20306 12939 20339
rect 12814 20242 12815 20306
rect 12879 20242 12939 20306
rect 12814 20209 12939 20242
rect 12960 20325 12961 20389
rect 13025 20325 13051 20389
rect 13115 20325 13141 20389
rect 13205 20325 13231 20389
rect 13295 20325 13320 20389
rect 13384 20325 13385 20389
rect 13427 20469 13552 20502
rect 13427 20405 13428 20469
rect 13492 20405 13552 20469
rect 13427 20372 13552 20405
rect 12960 20273 13385 20325
rect 12960 20209 12961 20273
rect 13025 20209 13051 20273
rect 13115 20209 13141 20273
rect 13205 20209 13231 20273
rect 13295 20209 13320 20273
rect 13384 20209 13385 20273
rect 1631 20207 2056 20209
rect 12960 20207 13385 20209
rect 1955 20181 2380 20183
rect 1792 20141 1917 20174
rect 1792 20077 1852 20141
rect 1916 20077 1917 20141
rect 1792 20044 1917 20077
rect 1955 20117 1956 20181
rect 2020 20117 2045 20181
rect 2109 20117 2135 20181
rect 2199 20117 2225 20181
rect 2289 20117 2315 20181
rect 2379 20117 2380 20181
rect 1955 20065 2380 20117
rect 12636 20181 13061 20183
rect 12636 20117 12637 20181
rect 12701 20117 12727 20181
rect 12791 20117 12817 20181
rect 12881 20117 12907 20181
rect 12971 20117 12996 20181
rect 13060 20117 13061 20181
rect 1955 20001 1956 20065
rect 2020 20001 2045 20065
rect 2109 20001 2135 20065
rect 2199 20001 2225 20065
rect 2289 20001 2315 20065
rect 2379 20001 2380 20065
rect 1955 19949 2380 20001
rect 1955 19885 1956 19949
rect 2020 19885 2045 19949
rect 2109 19885 2135 19949
rect 2199 19885 2225 19949
rect 2289 19885 2315 19949
rect 2379 19885 2380 19949
rect 2455 20070 2867 20071
rect 2455 20006 2456 20070
rect 2520 20006 2571 20070
rect 2635 20006 2686 20070
rect 2750 20006 2802 20070
rect 2866 20006 2867 20070
rect 2455 19950 2867 20006
rect 12149 20070 12561 20071
rect 12149 20006 12150 20070
rect 12214 20006 12266 20070
rect 12330 20006 12381 20070
rect 12445 20006 12496 20070
rect 12560 20006 12561 20070
rect 2455 19886 2456 19950
rect 2520 19886 2571 19950
rect 2635 19886 2686 19950
rect 2750 19886 2802 19950
rect 2866 19886 2867 19950
rect 2455 19885 2867 19886
rect 2881 19955 2971 19988
rect 2881 19891 2906 19955
rect 2970 19891 2971 19955
rect 1955 19883 2380 19885
rect 2881 19858 2971 19891
rect 12045 19955 12135 19988
rect 12045 19891 12046 19955
rect 12110 19891 12135 19955
rect 12045 19858 12135 19891
rect 12149 19950 12561 20006
rect 12149 19886 12150 19950
rect 12214 19886 12266 19950
rect 12330 19886 12381 19950
rect 12445 19886 12496 19950
rect 12560 19886 12561 19950
rect 12149 19885 12561 19886
rect 12636 20065 13061 20117
rect 12636 20001 12637 20065
rect 12701 20001 12727 20065
rect 12791 20001 12817 20065
rect 12881 20001 12907 20065
rect 12971 20001 12996 20065
rect 13060 20001 13061 20065
rect 13099 20141 13224 20174
rect 13099 20077 13100 20141
rect 13164 20077 13224 20141
rect 13099 20044 13224 20077
rect 12636 19949 13061 20001
rect 12636 19885 12637 19949
rect 12701 19885 12727 19949
rect 12791 19885 12817 19949
rect 12881 19885 12907 19949
rect 12971 19885 12996 19949
rect 13060 19885 13061 19949
rect 12636 19883 13061 19885
rect 2292 19844 3114 19846
rect 2133 19800 2258 19833
rect 2133 19736 2193 19800
rect 2257 19736 2258 19800
rect 2133 19703 2258 19736
rect 2292 19780 2293 19844
rect 2357 19780 2377 19844
rect 2441 19780 2461 19844
rect 2525 19780 2545 19844
rect 2609 19780 2629 19844
rect 2693 19780 2713 19844
rect 2777 19780 2797 19844
rect 2861 19780 2881 19844
rect 2945 19780 2965 19844
rect 3029 19780 3049 19844
rect 3113 19780 3114 19844
rect 2292 19728 3114 19780
rect 2292 19664 2293 19728
rect 2357 19664 2377 19728
rect 2441 19664 2461 19728
rect 2525 19664 2545 19728
rect 2609 19664 2629 19728
rect 2693 19664 2713 19728
rect 2777 19664 2797 19728
rect 2861 19664 2881 19728
rect 2945 19664 2965 19728
rect 3029 19664 3049 19728
rect 3113 19664 3114 19728
rect 11902 19844 12724 19846
rect 11902 19780 11903 19844
rect 11967 19780 11987 19844
rect 12051 19780 12071 19844
rect 12135 19780 12155 19844
rect 12219 19780 12239 19844
rect 12303 19780 12323 19844
rect 12387 19780 12407 19844
rect 12471 19780 12491 19844
rect 12555 19780 12575 19844
rect 12639 19780 12659 19844
rect 12723 19780 12724 19844
rect 11902 19728 12724 19780
rect 2292 19612 3114 19664
rect 2292 19548 2293 19612
rect 2357 19548 2377 19612
rect 2441 19548 2461 19612
rect 2525 19548 2545 19612
rect 2609 19548 2629 19612
rect 2693 19548 2713 19612
rect 2777 19548 2797 19612
rect 2861 19548 2881 19612
rect 2945 19548 2965 19612
rect 3029 19548 3049 19612
rect 3113 19548 3114 19612
rect 3123 19707 3247 19708
rect 3123 19643 3153 19707
rect 3217 19643 3247 19707
rect 3123 19614 3247 19643
rect 3123 19550 3153 19614
rect 3217 19550 3247 19614
rect 3123 19549 3247 19550
rect 11769 19707 11893 19708
rect 11769 19643 11799 19707
rect 11863 19643 11893 19707
rect 11769 19614 11893 19643
rect 11769 19550 11799 19614
rect 11863 19550 11893 19614
rect 11769 19549 11893 19550
rect 11902 19664 11903 19728
rect 11967 19664 11987 19728
rect 12051 19664 12071 19728
rect 12135 19664 12155 19728
rect 12219 19664 12239 19728
rect 12303 19664 12323 19728
rect 12387 19664 12407 19728
rect 12471 19664 12491 19728
rect 12555 19664 12575 19728
rect 12639 19664 12659 19728
rect 12723 19664 12724 19728
rect 12758 19800 12883 19833
rect 12758 19736 12759 19800
rect 12823 19736 12883 19800
rect 12758 19703 12883 19736
rect 11902 19612 12724 19664
rect 2292 19546 3114 19548
rect 11902 19548 11903 19612
rect 11967 19548 11987 19612
rect 12051 19548 12071 19612
rect 12135 19548 12155 19612
rect 12219 19548 12239 19612
rect 12303 19548 12323 19612
rect 12387 19548 12407 19612
rect 12471 19548 12491 19612
rect 12555 19548 12575 19612
rect 12639 19548 12659 19612
rect 12723 19548 12724 19612
rect 11902 19546 12724 19548
rect 4912 18895 7268 18934
rect 4912 17311 4938 18895
rect 7242 17311 7268 18895
rect 4912 17273 7268 17311
rect 7712 18895 10068 18934
rect 7712 17311 7738 18895
rect 10042 17311 10068 18895
rect 7712 17273 10068 17311
rect 5077 17218 7265 17231
rect 5077 17074 5099 17218
rect 7243 17074 7265 17218
rect 5077 17061 7265 17074
rect 7713 17218 9901 17231
rect 7713 17074 7735 17218
rect 9879 17074 9901 17218
rect 7713 17061 9901 17074
rect 2423 6025 3607 6053
rect 2423 5213 3607 5241
rect 11297 6024 12481 6052
rect 11297 5212 12481 5240
rect 886 4811 2072 4856
rect 886 4027 887 4811
rect 2071 4027 2072 4811
rect 886 3983 2072 4027
rect 12886 4811 14072 4856
rect 12886 4027 12887 4811
rect 14071 4027 14072 4811
rect 12886 3983 14072 4027
use sky130_ef_io__esd_ndiode_11v0_array  sky130_ef_io__esd_vddio
timestamp 1694700623
transform 0 1 7494 1 0 24764
box -1962 -5766 1962 5766
use sky130_ef_io__esd_pdiode_11v0_array  sky130_ef_io__esd_vssio
timestamp 1694700623
transform 0 1 7508 1 0 29198
box -1566 -5188 1566 5188
use sky130_fd_io__com_busses_esd  sky130_fd_io__com_busses_esd_0
timestamp 1694700623
transform 1 0 8 0 1 550
box 0 -142 15000 39451
<< properties >>
string GDS_END 4173624
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 2065562
<< end >>
