magic
tech sky130B
timestamp 1694700623
<< properties >>
string GDS_END 39966826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39966122
<< end >>
