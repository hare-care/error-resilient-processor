magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 315 157 1193 203
rect 1 21 1193 157
rect 29 -17 63 21
<< locali >>
rect 17 214 66 323
rect 122 268 178 323
rect 112 234 178 268
rect 122 214 178 234
rect 417 333 467 493
rect 585 333 651 493
rect 857 333 923 493
rect 1025 333 1091 493
rect 417 289 1091 333
rect 417 131 483 289
rect 649 215 710 289
rect 744 215 923 255
rect 989 215 1175 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 396 74 488
rect 108 439 153 527
rect 187 430 315 493
rect 17 357 246 396
rect 212 180 246 357
rect 17 146 246 180
rect 280 282 315 430
rect 349 299 383 527
rect 501 367 551 527
rect 685 367 823 527
rect 957 367 991 527
rect 1125 289 1179 527
rect 17 51 69 146
rect 280 143 316 282
rect 280 112 315 143
rect 549 215 615 255
rect 585 131 923 181
rect 957 147 1179 181
rect 103 17 153 109
rect 187 51 315 112
rect 349 97 383 117
rect 957 97 1007 147
rect 349 51 735 97
rect 773 51 1007 97
rect 1041 17 1075 113
rect 1109 51 1179 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 200 215 627 261
<< labels >>
rlabel locali s 122 214 178 234 6 A_N
port 1 nsew signal input
rlabel locali s 112 234 178 268 6 A_N
port 1 nsew signal input
rlabel locali s 122 268 178 323 6 A_N
port 1 nsew signal input
rlabel locali s 17 214 66 323 6 B_N
port 2 nsew signal input
rlabel locali s 744 215 923 255 6 C
port 3 nsew signal input
rlabel locali s 989 215 1175 255 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1193 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 315 157 1193 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 649 215 710 289 6 Y
port 9 nsew signal output
rlabel locali s 417 131 483 289 6 Y
port 9 nsew signal output
rlabel locali s 417 289 1091 333 6 Y
port 9 nsew signal output
rlabel locali s 1025 333 1091 493 6 Y
port 9 nsew signal output
rlabel locali s 857 333 923 493 6 Y
port 9 nsew signal output
rlabel locali s 585 333 651 493 6 Y
port 9 nsew signal output
rlabel locali s 417 333 467 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1943734
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1933346
<< end >>
