magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 930 897
<< pwell >>
rect 4 283 266 289
rect 4 43 859 283
rect -26 -43 890 43
<< mvnmos >>
rect 83 113 183 263
rect 360 107 460 257
rect 516 107 616 257
rect 676 107 776 257
<< mvpmos >>
rect 130 443 230 743
rect 330 443 430 743
rect 502 443 602 743
rect 658 443 758 743
<< mvndiff >>
rect 30 251 83 263
rect 30 217 38 251
rect 72 217 83 251
rect 30 159 83 217
rect 30 125 38 159
rect 72 125 83 159
rect 30 113 83 125
rect 183 255 240 263
rect 183 221 194 255
rect 228 221 240 255
rect 183 155 240 221
rect 183 121 194 155
rect 228 121 240 155
rect 183 113 240 121
rect 303 249 360 257
rect 303 215 315 249
rect 349 215 360 249
rect 303 149 360 215
rect 303 115 315 149
rect 349 115 360 149
rect 303 107 360 115
rect 460 249 516 257
rect 460 215 471 249
rect 505 215 516 249
rect 460 149 516 215
rect 460 115 471 149
rect 505 115 516 149
rect 460 107 516 115
rect 616 167 676 257
rect 616 133 627 167
rect 661 133 676 167
rect 616 107 676 133
rect 776 249 833 257
rect 776 215 787 249
rect 821 215 833 249
rect 776 149 833 215
rect 776 115 787 149
rect 821 115 833 149
rect 776 107 833 115
<< mvpdiff >>
rect 73 735 130 743
rect 73 701 85 735
rect 119 701 130 735
rect 73 652 130 701
rect 73 618 85 652
rect 119 618 130 652
rect 73 568 130 618
rect 73 534 85 568
rect 119 534 130 568
rect 73 485 130 534
rect 73 451 85 485
rect 119 451 130 485
rect 73 443 130 451
rect 230 735 330 743
rect 230 701 241 735
rect 275 701 330 735
rect 230 655 330 701
rect 230 621 241 655
rect 275 621 330 655
rect 230 574 330 621
rect 230 540 241 574
rect 275 540 330 574
rect 230 494 330 540
rect 230 460 241 494
rect 275 460 330 494
rect 230 443 330 460
rect 430 735 502 743
rect 430 701 441 735
rect 475 701 502 735
rect 430 652 502 701
rect 430 618 441 652
rect 475 618 502 652
rect 430 568 502 618
rect 430 534 441 568
rect 475 534 502 568
rect 430 485 502 534
rect 430 451 441 485
rect 475 451 502 485
rect 430 443 502 451
rect 602 443 658 743
rect 758 735 815 743
rect 758 701 769 735
rect 803 701 815 735
rect 758 652 815 701
rect 758 618 769 652
rect 803 618 815 652
rect 758 568 815 618
rect 758 534 769 568
rect 803 534 815 568
rect 758 485 815 534
rect 758 451 769 485
rect 803 451 815 485
rect 758 443 815 451
<< mvndiffc >>
rect 38 217 72 251
rect 38 125 72 159
rect 194 221 228 255
rect 194 121 228 155
rect 315 215 349 249
rect 315 115 349 149
rect 471 215 505 249
rect 471 115 505 149
rect 627 133 661 167
rect 787 215 821 249
rect 787 115 821 149
<< mvpdiffc >>
rect 85 701 119 735
rect 85 618 119 652
rect 85 534 119 568
rect 85 451 119 485
rect 241 701 275 735
rect 241 621 275 655
rect 241 540 275 574
rect 241 460 275 494
rect 441 701 475 735
rect 441 618 475 652
rect 441 534 475 568
rect 441 451 475 485
rect 769 701 803 735
rect 769 618 803 652
rect 769 534 803 568
rect 769 451 803 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
<< poly >>
rect 130 743 230 769
rect 330 743 430 769
rect 502 743 602 769
rect 658 743 758 769
rect 130 417 230 443
rect 83 343 230 417
rect 83 309 117 343
rect 151 317 230 343
rect 330 417 430 443
rect 330 395 460 417
rect 330 361 350 395
rect 384 361 460 395
rect 151 309 183 317
rect 83 263 183 309
rect 330 283 460 361
rect 502 383 602 443
rect 658 417 758 443
rect 502 360 616 383
rect 502 326 522 360
rect 556 326 616 360
rect 502 283 616 326
rect 658 351 776 417
rect 658 317 678 351
rect 712 317 776 351
rect 658 283 776 317
rect 360 257 460 283
rect 516 257 616 283
rect 676 257 776 283
rect 83 87 183 113
rect 360 81 460 107
rect 516 81 616 107
rect 676 81 776 107
<< polycont >>
rect 117 309 151 343
rect 350 361 384 395
rect 522 326 556 360
rect 678 317 712 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
rect 25 735 119 751
rect 25 701 85 735
rect 25 652 119 701
rect 25 618 85 652
rect 25 568 119 618
rect 25 534 85 568
rect 25 485 119 534
rect 25 451 85 485
rect 155 735 405 751
rect 189 701 227 735
rect 275 701 299 735
rect 333 701 371 735
rect 155 655 405 701
rect 155 621 241 655
rect 275 621 405 655
rect 155 574 405 621
rect 155 540 241 574
rect 275 540 405 574
rect 155 494 405 540
rect 155 460 241 494
rect 275 460 405 494
rect 441 735 475 751
rect 441 652 475 701
rect 593 735 846 751
rect 593 701 594 735
rect 628 701 666 735
rect 700 701 738 735
rect 803 701 810 735
rect 844 701 846 735
rect 593 652 846 701
rect 441 568 475 618
rect 441 485 475 534
rect 25 395 119 451
rect 217 395 400 424
rect 25 251 76 395
rect 217 361 350 395
rect 384 361 400 395
rect 110 343 167 359
rect 110 309 117 343
rect 151 325 167 343
rect 441 325 475 451
rect 151 309 475 325
rect 511 360 557 652
rect 593 618 769 652
rect 803 618 846 652
rect 593 568 846 618
rect 593 534 769 568
rect 803 534 846 568
rect 593 485 846 534
rect 593 451 769 485
rect 803 451 846 485
rect 593 435 846 451
rect 511 326 522 360
rect 556 326 557 360
rect 511 310 557 326
rect 601 351 839 367
rect 601 317 678 351
rect 712 317 839 351
rect 110 291 475 309
rect 601 301 839 317
rect 25 217 38 251
rect 72 217 76 251
rect 25 159 76 217
rect 25 125 38 159
rect 72 125 76 159
rect 25 105 76 125
rect 110 221 194 255
rect 228 221 263 255
rect 110 155 263 221
rect 110 121 194 155
rect 228 121 263 155
rect 110 113 263 121
rect 110 79 120 113
rect 154 79 221 113
rect 255 79 263 113
rect 299 249 365 291
rect 771 255 837 265
rect 299 215 315 249
rect 349 215 365 249
rect 299 149 365 215
rect 299 115 315 149
rect 349 115 365 149
rect 299 99 365 115
rect 455 249 837 255
rect 455 215 471 249
rect 505 221 787 249
rect 505 215 521 221
rect 455 149 521 215
rect 771 215 787 221
rect 821 215 837 249
rect 455 115 471 149
rect 505 115 521 149
rect 455 99 521 115
rect 557 167 735 185
rect 557 133 627 167
rect 661 133 735 167
rect 557 113 735 133
rect 110 73 263 79
rect 591 79 629 113
rect 663 79 701 113
rect 771 149 837 215
rect 771 115 787 149
rect 821 115 837 149
rect 771 99 837 115
rect 557 73 735 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 155 701 189 735
rect 227 701 241 735
rect 241 701 261 735
rect 299 701 333 735
rect 371 701 405 735
rect 594 701 628 735
rect 666 701 700 735
rect 738 701 769 735
rect 769 701 772 735
rect 810 701 844 735
rect 120 79 154 113
rect 221 79 255 113
rect 557 79 591 113
rect 629 79 663 113
rect 701 79 735 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 831 864 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 864 831
rect 0 791 864 797
rect 0 735 864 763
rect 0 701 155 735
rect 189 701 227 735
rect 261 701 299 735
rect 333 701 371 735
rect 405 701 594 735
rect 628 701 666 735
rect 700 701 738 735
rect 772 701 810 735
rect 844 701 864 735
rect 0 689 864 701
rect 0 113 864 125
rect 0 79 120 113
rect 154 79 221 113
rect 255 79 557 113
rect 591 79 629 113
rect 663 79 701 113
rect 735 79 864 113
rect 0 51 864 79
rect 0 17 864 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -23 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21a_1
flabel metal1 s 0 51 864 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 864 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 864 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 864 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 612 545 646 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 612 65 646 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 864 814
string GDS_END 179726
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 167972
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
