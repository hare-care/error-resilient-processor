magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< obsli1 >>
rect 34 2492 1958 2558
rect 34 100 100 2492
rect 260 2266 1732 2332
rect 260 326 326 2266
rect 662 1864 1330 1930
rect 662 728 728 1864
rect 895 895 1097 1697
rect 1264 728 1330 1864
rect 662 662 1330 728
rect 1666 326 1732 2266
rect 260 260 1732 326
rect 1892 100 1958 2492
rect 34 34 1958 100
<< obsm1 >>
rect 38 2496 1954 2554
rect 38 96 96 2496
rect 264 2270 1728 2328
rect 264 322 322 2270
rect 666 1868 1326 1926
rect 666 724 724 1868
rect 895 907 1097 1685
rect 1268 724 1326 1868
rect 666 666 1326 724
rect 1670 322 1728 2270
rect 264 264 1728 322
rect 1896 96 1954 2496
rect 38 38 1954 96
<< properties >>
string FIXED_BBOX 26 26 1966 2566
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8779906
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8732342
<< end >>
