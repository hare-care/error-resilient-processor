magic
tech sky130B
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_0
timestamp 1694700623
transform 1 0 581 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_1
timestamp 1694700623
transform 1 0 1501 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_2
timestamp 1694700623
transform 1 0 2421 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_3
timestamp 1694700623
transform 1 0 3341 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_4
timestamp 1694700623
transform 1 0 4261 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_5
timestamp 1694700623
transform 1 0 5181 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_6
timestamp 1694700623
transform 1 0 6101 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_7
timestamp 1694700623
transform 1 0 7021 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_8
timestamp 1694700623
transform 1 0 7941 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_9
timestamp 1694700623
transform 1 0 8861 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808675  sky130_fd_pr__hvdftpl1s__example_55959141808675_0
timestamp 1694700623
transform -1 0 -79 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808675  sky130_fd_pr__hvdftpl1s__example_55959141808675_1
timestamp 1694700623
transform 1 0 9781 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 11221224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11209504
<< end >>
