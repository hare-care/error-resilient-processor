magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< dnwell >>
rect -915 14603 5413 15797
rect -915 9930 85 14603
<< nwell >>
rect 1 15589 15172 16593
rect 1 15507 5496 15589
rect 1 14893 588 15507
rect 5328 14893 5496 15507
rect 1 14711 5496 14893
rect 12570 14777 15172 15589
rect 14350 14723 15172 14777
rect 218 14523 5496 14711
rect 8293 8874 15173 8875
rect -32 6931 15173 8874
rect 3462 109 6890 1131
<< pwell >>
rect 648 14953 5268 15447
rect -973 8935 15143 9711
rect 18 6661 7134 6869
rect 12467 6661 15143 6869
rect 18 6025 15143 6661
rect 14891 5962 15143 6025
rect 14951 1314 15143 5962
rect 7018 1308 15143 1314
rect 42 1225 15143 1308
rect 3511 1191 15143 1225
rect 6962 962 15143 1191
rect 6962 395 7780 962
rect 9661 702 15143 962
rect 9661 395 11682 702
rect 14439 395 15143 702
rect 6962 49 15143 395
rect 3519 -7 15143 49
rect 3519 -37 7048 -7
<< mvnmos >>
rect 782 15140 1782 15260
rect 1892 15140 2892 15260
rect 3013 15140 4013 15260
rect 4134 15140 5134 15260
<< mvpmos >>
rect 3726 804 5126 904
rect 5256 804 6656 904
rect 3726 648 5126 748
rect 5256 648 6656 748
rect 3726 492 5126 592
rect 5256 492 6656 592
rect 3726 336 5126 436
rect 5256 336 6656 436
<< mvndiff >>
rect 782 15305 1782 15313
rect 782 15271 794 15305
rect 828 15271 862 15305
rect 896 15271 930 15305
rect 964 15271 998 15305
rect 1032 15271 1066 15305
rect 1100 15271 1134 15305
rect 1168 15271 1202 15305
rect 1236 15271 1270 15305
rect 1304 15271 1338 15305
rect 1372 15271 1406 15305
rect 1440 15271 1474 15305
rect 1508 15271 1542 15305
rect 1576 15271 1610 15305
rect 1644 15271 1678 15305
rect 1712 15271 1782 15305
rect 782 15260 1782 15271
rect 1892 15305 2892 15313
rect 1892 15271 1962 15305
rect 1996 15271 2030 15305
rect 2064 15271 2098 15305
rect 2132 15271 2166 15305
rect 2200 15271 2234 15305
rect 2268 15271 2302 15305
rect 2336 15271 2370 15305
rect 2404 15271 2438 15305
rect 2472 15271 2506 15305
rect 2540 15271 2574 15305
rect 2608 15271 2642 15305
rect 2676 15271 2710 15305
rect 2744 15271 2778 15305
rect 2812 15271 2846 15305
rect 2880 15271 2892 15305
rect 1892 15260 2892 15271
rect 3013 15305 4013 15313
rect 3013 15271 3083 15305
rect 3117 15271 3151 15305
rect 3185 15271 3219 15305
rect 3253 15271 3287 15305
rect 3321 15271 3355 15305
rect 3389 15271 3423 15305
rect 3457 15271 3491 15305
rect 3525 15271 3559 15305
rect 3593 15271 3627 15305
rect 3661 15271 3695 15305
rect 3729 15271 3763 15305
rect 3797 15271 3831 15305
rect 3865 15271 3899 15305
rect 3933 15271 3967 15305
rect 4001 15271 4013 15305
rect 3013 15260 4013 15271
rect 4134 15305 5134 15313
rect 4134 15271 4204 15305
rect 4238 15271 4272 15305
rect 4306 15271 4340 15305
rect 4374 15271 4408 15305
rect 4442 15271 4476 15305
rect 4510 15271 4544 15305
rect 4578 15271 4612 15305
rect 4646 15271 4680 15305
rect 4714 15271 4748 15305
rect 4782 15271 4816 15305
rect 4850 15271 4884 15305
rect 4918 15271 4952 15305
rect 4986 15271 5020 15305
rect 5054 15271 5088 15305
rect 5122 15271 5134 15305
rect 4134 15260 5134 15271
rect 782 15129 1782 15140
rect 782 15095 794 15129
rect 828 15095 862 15129
rect 896 15095 930 15129
rect 964 15095 998 15129
rect 1032 15095 1066 15129
rect 1100 15095 1134 15129
rect 1168 15095 1202 15129
rect 1236 15095 1270 15129
rect 1304 15095 1338 15129
rect 1372 15095 1406 15129
rect 1440 15095 1474 15129
rect 1508 15095 1542 15129
rect 1576 15095 1610 15129
rect 1644 15095 1678 15129
rect 1712 15095 1782 15129
rect 782 15087 1782 15095
rect 1892 15129 2892 15140
rect 1892 15095 1962 15129
rect 1996 15095 2030 15129
rect 2064 15095 2098 15129
rect 2132 15095 2166 15129
rect 2200 15095 2234 15129
rect 2268 15095 2302 15129
rect 2336 15095 2370 15129
rect 2404 15095 2438 15129
rect 2472 15095 2506 15129
rect 2540 15095 2574 15129
rect 2608 15095 2642 15129
rect 2676 15095 2710 15129
rect 2744 15095 2778 15129
rect 2812 15095 2846 15129
rect 2880 15095 2892 15129
rect 1892 15087 2892 15095
rect 3013 15129 4013 15140
rect 3013 15095 3083 15129
rect 3117 15095 3151 15129
rect 3185 15095 3219 15129
rect 3253 15095 3287 15129
rect 3321 15095 3355 15129
rect 3389 15095 3423 15129
rect 3457 15095 3491 15129
rect 3525 15095 3559 15129
rect 3593 15095 3627 15129
rect 3661 15095 3695 15129
rect 3729 15095 3763 15129
rect 3797 15095 3831 15129
rect 3865 15095 3899 15129
rect 3933 15095 3967 15129
rect 4001 15095 4013 15129
rect 3013 15087 4013 15095
rect 4134 15129 5134 15140
rect 4134 15095 4204 15129
rect 4238 15095 4272 15129
rect 4306 15095 4340 15129
rect 4374 15095 4408 15129
rect 4442 15095 4476 15129
rect 4510 15095 4544 15129
rect 4578 15095 4612 15129
rect 4646 15095 4680 15129
rect 4714 15095 4748 15129
rect 4782 15095 4816 15129
rect 4850 15095 4884 15129
rect 4918 15095 4952 15129
rect 4986 15095 5020 15129
rect 5054 15095 5088 15129
rect 5122 15095 5134 15129
rect 4134 15087 5134 15095
<< mvpdiff >>
rect 3726 949 5126 957
rect 3726 915 3738 949
rect 3772 915 3806 949
rect 3840 915 3874 949
rect 3908 915 3942 949
rect 3976 915 4010 949
rect 4044 915 4078 949
rect 4112 915 4146 949
rect 4180 915 4214 949
rect 4248 915 4282 949
rect 4316 915 4350 949
rect 4384 915 4418 949
rect 4452 915 4486 949
rect 4520 915 4554 949
rect 4588 915 4622 949
rect 4656 915 4690 949
rect 4724 915 4758 949
rect 4792 915 4826 949
rect 4860 915 4894 949
rect 4928 915 4962 949
rect 4996 915 5030 949
rect 5064 915 5126 949
rect 3726 904 5126 915
rect 5256 949 6656 957
rect 5256 915 5268 949
rect 5302 915 5336 949
rect 5370 915 5404 949
rect 5438 915 5472 949
rect 5506 915 5540 949
rect 5574 915 5608 949
rect 5642 915 5676 949
rect 5710 915 5744 949
rect 5778 915 5812 949
rect 5846 915 5880 949
rect 5914 915 5948 949
rect 5982 915 6016 949
rect 6050 915 6084 949
rect 6118 915 6152 949
rect 6186 915 6220 949
rect 6254 915 6288 949
rect 6322 915 6356 949
rect 6390 915 6424 949
rect 6458 915 6492 949
rect 6526 915 6560 949
rect 6594 915 6656 949
rect 5256 904 6656 915
rect 3726 793 5126 804
rect 3726 759 3738 793
rect 3772 759 3806 793
rect 3840 759 3874 793
rect 3908 759 3942 793
rect 3976 759 4010 793
rect 4044 759 4078 793
rect 4112 759 4146 793
rect 4180 759 4214 793
rect 4248 759 4282 793
rect 4316 759 4350 793
rect 4384 759 4418 793
rect 4452 759 4486 793
rect 4520 759 4554 793
rect 4588 759 4622 793
rect 4656 759 4690 793
rect 4724 759 4758 793
rect 4792 759 4826 793
rect 4860 759 4894 793
rect 4928 759 4962 793
rect 4996 759 5030 793
rect 5064 759 5126 793
rect 3726 748 5126 759
rect 5256 793 6656 804
rect 5256 759 5268 793
rect 5302 759 5336 793
rect 5370 759 5404 793
rect 5438 759 5472 793
rect 5506 759 5540 793
rect 5574 759 5608 793
rect 5642 759 5676 793
rect 5710 759 5744 793
rect 5778 759 5812 793
rect 5846 759 5880 793
rect 5914 759 5948 793
rect 5982 759 6016 793
rect 6050 759 6084 793
rect 6118 759 6152 793
rect 6186 759 6220 793
rect 6254 759 6288 793
rect 6322 759 6356 793
rect 6390 759 6424 793
rect 6458 759 6492 793
rect 6526 759 6560 793
rect 6594 759 6656 793
rect 5256 748 6656 759
rect 3726 637 5126 648
rect 3726 603 3738 637
rect 3772 603 3806 637
rect 3840 603 3874 637
rect 3908 603 3942 637
rect 3976 603 4010 637
rect 4044 603 4078 637
rect 4112 603 4146 637
rect 4180 603 4214 637
rect 4248 603 4282 637
rect 4316 603 4350 637
rect 4384 603 4418 637
rect 4452 603 4486 637
rect 4520 603 4554 637
rect 4588 603 4622 637
rect 4656 603 4690 637
rect 4724 603 4758 637
rect 4792 603 4826 637
rect 4860 603 4894 637
rect 4928 603 4962 637
rect 4996 603 5030 637
rect 5064 603 5126 637
rect 3726 592 5126 603
rect 5256 637 6656 648
rect 5256 603 5268 637
rect 5302 603 5336 637
rect 5370 603 5404 637
rect 5438 603 5472 637
rect 5506 603 5540 637
rect 5574 603 5608 637
rect 5642 603 5676 637
rect 5710 603 5744 637
rect 5778 603 5812 637
rect 5846 603 5880 637
rect 5914 603 5948 637
rect 5982 603 6016 637
rect 6050 603 6084 637
rect 6118 603 6152 637
rect 6186 603 6220 637
rect 6254 603 6288 637
rect 6322 603 6356 637
rect 6390 603 6424 637
rect 6458 603 6492 637
rect 6526 603 6560 637
rect 6594 603 6656 637
rect 5256 592 6656 603
rect 3726 481 5126 492
rect 3726 447 3738 481
rect 3772 447 3806 481
rect 3840 447 3874 481
rect 3908 447 3942 481
rect 3976 447 4010 481
rect 4044 447 4078 481
rect 4112 447 4146 481
rect 4180 447 4214 481
rect 4248 447 4282 481
rect 4316 447 4350 481
rect 4384 447 4418 481
rect 4452 447 4486 481
rect 4520 447 4554 481
rect 4588 447 4622 481
rect 4656 447 4690 481
rect 4724 447 4758 481
rect 4792 447 4826 481
rect 4860 447 4894 481
rect 4928 447 4962 481
rect 4996 447 5030 481
rect 5064 447 5126 481
rect 3726 436 5126 447
rect 5256 481 6656 492
rect 5256 447 5268 481
rect 5302 447 5336 481
rect 5370 447 5404 481
rect 5438 447 5472 481
rect 5506 447 5540 481
rect 5574 447 5608 481
rect 5642 447 5676 481
rect 5710 447 5744 481
rect 5778 447 5812 481
rect 5846 447 5880 481
rect 5914 447 5948 481
rect 5982 447 6016 481
rect 6050 447 6084 481
rect 6118 447 6152 481
rect 6186 447 6220 481
rect 6254 447 6288 481
rect 6322 447 6356 481
rect 6390 447 6424 481
rect 6458 447 6492 481
rect 6526 447 6560 481
rect 6594 447 6656 481
rect 5256 436 6656 447
rect 3726 325 5126 336
rect 3726 291 3738 325
rect 3772 291 3806 325
rect 3840 291 3874 325
rect 3908 291 3942 325
rect 3976 291 4010 325
rect 4044 291 4078 325
rect 4112 291 4146 325
rect 4180 291 4214 325
rect 4248 291 4282 325
rect 4316 291 4350 325
rect 4384 291 4418 325
rect 4452 291 4486 325
rect 4520 291 4554 325
rect 4588 291 4622 325
rect 4656 291 4690 325
rect 4724 291 4758 325
rect 4792 291 4826 325
rect 4860 291 4894 325
rect 4928 291 4962 325
rect 4996 291 5030 325
rect 5064 291 5126 325
rect 3726 283 5126 291
rect 5256 325 6656 336
rect 5256 291 5268 325
rect 5302 291 5336 325
rect 5370 291 5404 325
rect 5438 291 5472 325
rect 5506 291 5540 325
rect 5574 291 5608 325
rect 5642 291 5676 325
rect 5710 291 5744 325
rect 5778 291 5812 325
rect 5846 291 5880 325
rect 5914 291 5948 325
rect 5982 291 6016 325
rect 6050 291 6084 325
rect 6118 291 6152 325
rect 6186 291 6220 325
rect 6254 291 6288 325
rect 6322 291 6356 325
rect 6390 291 6424 325
rect 6458 291 6492 325
rect 6526 291 6560 325
rect 6594 291 6656 325
rect 5256 283 6656 291
<< mvndiffc >>
rect 794 15271 828 15305
rect 862 15271 896 15305
rect 930 15271 964 15305
rect 998 15271 1032 15305
rect 1066 15271 1100 15305
rect 1134 15271 1168 15305
rect 1202 15271 1236 15305
rect 1270 15271 1304 15305
rect 1338 15271 1372 15305
rect 1406 15271 1440 15305
rect 1474 15271 1508 15305
rect 1542 15271 1576 15305
rect 1610 15271 1644 15305
rect 1678 15271 1712 15305
rect 1962 15271 1996 15305
rect 2030 15271 2064 15305
rect 2098 15271 2132 15305
rect 2166 15271 2200 15305
rect 2234 15271 2268 15305
rect 2302 15271 2336 15305
rect 2370 15271 2404 15305
rect 2438 15271 2472 15305
rect 2506 15271 2540 15305
rect 2574 15271 2608 15305
rect 2642 15271 2676 15305
rect 2710 15271 2744 15305
rect 2778 15271 2812 15305
rect 2846 15271 2880 15305
rect 3083 15271 3117 15305
rect 3151 15271 3185 15305
rect 3219 15271 3253 15305
rect 3287 15271 3321 15305
rect 3355 15271 3389 15305
rect 3423 15271 3457 15305
rect 3491 15271 3525 15305
rect 3559 15271 3593 15305
rect 3627 15271 3661 15305
rect 3695 15271 3729 15305
rect 3763 15271 3797 15305
rect 3831 15271 3865 15305
rect 3899 15271 3933 15305
rect 3967 15271 4001 15305
rect 4204 15271 4238 15305
rect 4272 15271 4306 15305
rect 4340 15271 4374 15305
rect 4408 15271 4442 15305
rect 4476 15271 4510 15305
rect 4544 15271 4578 15305
rect 4612 15271 4646 15305
rect 4680 15271 4714 15305
rect 4748 15271 4782 15305
rect 4816 15271 4850 15305
rect 4884 15271 4918 15305
rect 4952 15271 4986 15305
rect 5020 15271 5054 15305
rect 5088 15271 5122 15305
rect 794 15095 828 15129
rect 862 15095 896 15129
rect 930 15095 964 15129
rect 998 15095 1032 15129
rect 1066 15095 1100 15129
rect 1134 15095 1168 15129
rect 1202 15095 1236 15129
rect 1270 15095 1304 15129
rect 1338 15095 1372 15129
rect 1406 15095 1440 15129
rect 1474 15095 1508 15129
rect 1542 15095 1576 15129
rect 1610 15095 1644 15129
rect 1678 15095 1712 15129
rect 1962 15095 1996 15129
rect 2030 15095 2064 15129
rect 2098 15095 2132 15129
rect 2166 15095 2200 15129
rect 2234 15095 2268 15129
rect 2302 15095 2336 15129
rect 2370 15095 2404 15129
rect 2438 15095 2472 15129
rect 2506 15095 2540 15129
rect 2574 15095 2608 15129
rect 2642 15095 2676 15129
rect 2710 15095 2744 15129
rect 2778 15095 2812 15129
rect 2846 15095 2880 15129
rect 3083 15095 3117 15129
rect 3151 15095 3185 15129
rect 3219 15095 3253 15129
rect 3287 15095 3321 15129
rect 3355 15095 3389 15129
rect 3423 15095 3457 15129
rect 3491 15095 3525 15129
rect 3559 15095 3593 15129
rect 3627 15095 3661 15129
rect 3695 15095 3729 15129
rect 3763 15095 3797 15129
rect 3831 15095 3865 15129
rect 3899 15095 3933 15129
rect 3967 15095 4001 15129
rect 4204 15095 4238 15129
rect 4272 15095 4306 15129
rect 4340 15095 4374 15129
rect 4408 15095 4442 15129
rect 4476 15095 4510 15129
rect 4544 15095 4578 15129
rect 4612 15095 4646 15129
rect 4680 15095 4714 15129
rect 4748 15095 4782 15129
rect 4816 15095 4850 15129
rect 4884 15095 4918 15129
rect 4952 15095 4986 15129
rect 5020 15095 5054 15129
rect 5088 15095 5122 15129
<< mvpdiffc >>
rect 3738 915 3772 949
rect 3806 915 3840 949
rect 3874 915 3908 949
rect 3942 915 3976 949
rect 4010 915 4044 949
rect 4078 915 4112 949
rect 4146 915 4180 949
rect 4214 915 4248 949
rect 4282 915 4316 949
rect 4350 915 4384 949
rect 4418 915 4452 949
rect 4486 915 4520 949
rect 4554 915 4588 949
rect 4622 915 4656 949
rect 4690 915 4724 949
rect 4758 915 4792 949
rect 4826 915 4860 949
rect 4894 915 4928 949
rect 4962 915 4996 949
rect 5030 915 5064 949
rect 5268 915 5302 949
rect 5336 915 5370 949
rect 5404 915 5438 949
rect 5472 915 5506 949
rect 5540 915 5574 949
rect 5608 915 5642 949
rect 5676 915 5710 949
rect 5744 915 5778 949
rect 5812 915 5846 949
rect 5880 915 5914 949
rect 5948 915 5982 949
rect 6016 915 6050 949
rect 6084 915 6118 949
rect 6152 915 6186 949
rect 6220 915 6254 949
rect 6288 915 6322 949
rect 6356 915 6390 949
rect 6424 915 6458 949
rect 6492 915 6526 949
rect 6560 915 6594 949
rect 3738 759 3772 793
rect 3806 759 3840 793
rect 3874 759 3908 793
rect 3942 759 3976 793
rect 4010 759 4044 793
rect 4078 759 4112 793
rect 4146 759 4180 793
rect 4214 759 4248 793
rect 4282 759 4316 793
rect 4350 759 4384 793
rect 4418 759 4452 793
rect 4486 759 4520 793
rect 4554 759 4588 793
rect 4622 759 4656 793
rect 4690 759 4724 793
rect 4758 759 4792 793
rect 4826 759 4860 793
rect 4894 759 4928 793
rect 4962 759 4996 793
rect 5030 759 5064 793
rect 5268 759 5302 793
rect 5336 759 5370 793
rect 5404 759 5438 793
rect 5472 759 5506 793
rect 5540 759 5574 793
rect 5608 759 5642 793
rect 5676 759 5710 793
rect 5744 759 5778 793
rect 5812 759 5846 793
rect 5880 759 5914 793
rect 5948 759 5982 793
rect 6016 759 6050 793
rect 6084 759 6118 793
rect 6152 759 6186 793
rect 6220 759 6254 793
rect 6288 759 6322 793
rect 6356 759 6390 793
rect 6424 759 6458 793
rect 6492 759 6526 793
rect 6560 759 6594 793
rect 3738 603 3772 637
rect 3806 603 3840 637
rect 3874 603 3908 637
rect 3942 603 3976 637
rect 4010 603 4044 637
rect 4078 603 4112 637
rect 4146 603 4180 637
rect 4214 603 4248 637
rect 4282 603 4316 637
rect 4350 603 4384 637
rect 4418 603 4452 637
rect 4486 603 4520 637
rect 4554 603 4588 637
rect 4622 603 4656 637
rect 4690 603 4724 637
rect 4758 603 4792 637
rect 4826 603 4860 637
rect 4894 603 4928 637
rect 4962 603 4996 637
rect 5030 603 5064 637
rect 5268 603 5302 637
rect 5336 603 5370 637
rect 5404 603 5438 637
rect 5472 603 5506 637
rect 5540 603 5574 637
rect 5608 603 5642 637
rect 5676 603 5710 637
rect 5744 603 5778 637
rect 5812 603 5846 637
rect 5880 603 5914 637
rect 5948 603 5982 637
rect 6016 603 6050 637
rect 6084 603 6118 637
rect 6152 603 6186 637
rect 6220 603 6254 637
rect 6288 603 6322 637
rect 6356 603 6390 637
rect 6424 603 6458 637
rect 6492 603 6526 637
rect 6560 603 6594 637
rect 3738 447 3772 481
rect 3806 447 3840 481
rect 3874 447 3908 481
rect 3942 447 3976 481
rect 4010 447 4044 481
rect 4078 447 4112 481
rect 4146 447 4180 481
rect 4214 447 4248 481
rect 4282 447 4316 481
rect 4350 447 4384 481
rect 4418 447 4452 481
rect 4486 447 4520 481
rect 4554 447 4588 481
rect 4622 447 4656 481
rect 4690 447 4724 481
rect 4758 447 4792 481
rect 4826 447 4860 481
rect 4894 447 4928 481
rect 4962 447 4996 481
rect 5030 447 5064 481
rect 5268 447 5302 481
rect 5336 447 5370 481
rect 5404 447 5438 481
rect 5472 447 5506 481
rect 5540 447 5574 481
rect 5608 447 5642 481
rect 5676 447 5710 481
rect 5744 447 5778 481
rect 5812 447 5846 481
rect 5880 447 5914 481
rect 5948 447 5982 481
rect 6016 447 6050 481
rect 6084 447 6118 481
rect 6152 447 6186 481
rect 6220 447 6254 481
rect 6288 447 6322 481
rect 6356 447 6390 481
rect 6424 447 6458 481
rect 6492 447 6526 481
rect 6560 447 6594 481
rect 3738 291 3772 325
rect 3806 291 3840 325
rect 3874 291 3908 325
rect 3942 291 3976 325
rect 4010 291 4044 325
rect 4078 291 4112 325
rect 4146 291 4180 325
rect 4214 291 4248 325
rect 4282 291 4316 325
rect 4350 291 4384 325
rect 4418 291 4452 325
rect 4486 291 4520 325
rect 4554 291 4588 325
rect 4622 291 4656 325
rect 4690 291 4724 325
rect 4758 291 4792 325
rect 4826 291 4860 325
rect 4894 291 4928 325
rect 4962 291 4996 325
rect 5030 291 5064 325
rect 5268 291 5302 325
rect 5336 291 5370 325
rect 5404 291 5438 325
rect 5472 291 5506 325
rect 5540 291 5574 325
rect 5608 291 5642 325
rect 5676 291 5710 325
rect 5744 291 5778 325
rect 5812 291 5846 325
rect 5880 291 5914 325
rect 5948 291 5982 325
rect 6016 291 6050 325
rect 6084 291 6118 325
rect 6152 291 6186 325
rect 6220 291 6254 325
rect 6288 291 6322 325
rect 6356 291 6390 325
rect 6424 291 6458 325
rect 6492 291 6526 325
rect 6560 291 6594 325
<< mvpsubdiff >>
rect 674 15387 698 15421
rect 732 15387 767 15421
rect 801 15387 836 15421
rect 870 15387 905 15421
rect 939 15387 974 15421
rect 1008 15387 1043 15421
rect 1077 15387 1112 15421
rect 1146 15387 1181 15421
rect 1215 15387 1250 15421
rect 1284 15387 1319 15421
rect 1353 15387 1388 15421
rect 1422 15387 1457 15421
rect 1491 15387 1526 15421
rect 1560 15387 1595 15421
rect 1629 15387 1664 15421
rect 1698 15387 1733 15421
rect 1767 15387 1802 15421
rect 1836 15387 1871 15421
rect 1905 15387 1940 15421
rect 1974 15387 2009 15421
rect 2043 15387 2078 15421
rect 2112 15387 2147 15421
rect 2181 15387 2216 15421
rect 2250 15387 2285 15421
rect 2319 15387 2354 15421
rect 2388 15387 2423 15421
rect 2457 15387 2492 15421
rect 2526 15387 2561 15421
rect 2595 15387 2630 15421
rect 2664 15387 2699 15421
rect 2733 15387 2768 15421
rect 2802 15387 2837 15421
rect 2871 15387 2906 15421
rect 2940 15387 2975 15421
rect 3009 15387 3044 15421
rect 3078 15387 3113 15421
rect 3147 15387 3182 15421
rect 3216 15387 3251 15421
rect 3285 15387 3320 15421
rect 3354 15387 3389 15421
rect 3423 15387 3458 15421
rect 3492 15387 3527 15421
rect 3561 15387 3596 15421
rect 3630 15387 3665 15421
rect 3699 15387 3734 15421
rect 3768 15387 3803 15421
rect 3837 15387 3872 15421
rect 3906 15387 3941 15421
rect 3975 15387 4010 15421
rect 4044 15387 4079 15421
rect 4113 15387 4148 15421
rect 4182 15387 4217 15421
rect 4251 15387 4286 15421
rect 4320 15387 4355 15421
rect 4389 15387 4424 15421
rect 4458 15387 4493 15421
rect 4527 15387 4562 15421
rect 4596 15387 4631 15421
rect 4665 15387 4700 15421
rect 4734 15387 4769 15421
rect 4803 15387 4838 15421
rect 4872 15387 4907 15421
rect 4941 15387 4976 15421
rect 5010 15387 5045 15421
rect 5079 15387 5114 15421
rect 5148 15397 5242 15421
rect 5148 15387 5208 15397
rect 674 15323 708 15387
rect 674 15252 708 15289
rect 5208 15284 5242 15363
rect 674 15181 708 15218
rect 674 15109 708 15147
rect 5208 15150 5242 15250
rect 674 15037 708 15075
rect 5208 15013 5242 15116
rect 708 15003 768 15013
rect 674 14979 768 15003
rect 802 14979 837 15013
rect 871 14979 906 15013
rect 940 14979 975 15013
rect 1009 14979 1044 15013
rect 1078 14979 1113 15013
rect 1147 14979 1182 15013
rect 1216 14979 1251 15013
rect 1285 14979 1320 15013
rect 1354 14979 1389 15013
rect 1423 14979 1458 15013
rect 1492 14979 1527 15013
rect 1561 14979 1596 15013
rect 1630 14979 1665 15013
rect 1699 14979 1734 15013
rect 1768 14979 1803 15013
rect 1837 14979 1872 15013
rect 1906 14979 1941 15013
rect 1975 14979 2010 15013
rect 2044 14979 2079 15013
rect 2113 14979 2148 15013
rect 2182 14979 2217 15013
rect 2251 14979 2286 15013
rect 2320 14979 2355 15013
rect 2389 14979 2424 15013
rect 2458 14979 2493 15013
rect 2527 14979 2562 15013
rect 2596 14979 2631 15013
rect 2665 14979 2700 15013
rect 2734 14979 2769 15013
rect 2803 14979 2838 15013
rect 2872 14979 2907 15013
rect 2941 14979 2976 15013
rect 3010 14979 3045 15013
rect 3079 14979 3114 15013
rect 3148 14979 3183 15013
rect 3217 14979 3252 15013
rect 3286 14979 3321 15013
rect 3355 14979 3390 15013
rect 3424 14979 3459 15013
rect 3493 14979 3528 15013
rect 3562 14979 3597 15013
rect 3631 14979 3666 15013
rect 3700 14979 3735 15013
rect 3769 14979 3804 15013
rect 3838 14979 3873 15013
rect 3907 14979 3942 15013
rect 3976 14979 4011 15013
rect 4045 14979 4080 15013
rect 4114 14979 4149 15013
rect 4183 14979 4218 15013
rect 4252 14979 4287 15013
rect 4321 14979 4356 15013
rect 4390 14979 4425 15013
rect 4459 14979 4494 15013
rect 4528 14979 4563 15013
rect 4597 14979 4632 15013
rect 4666 14979 4701 15013
rect 4735 14979 4770 15013
rect 4804 14979 4839 15013
rect 4873 14979 4908 15013
rect 4942 14979 4977 15013
rect 5011 14979 5046 15013
rect 5080 14979 5115 15013
rect 5149 14979 5184 15013
rect 5218 14979 5242 15013
rect -947 9680 15117 9685
rect -947 9647 -723 9680
rect -947 9613 -932 9647
rect -898 9613 -864 9647
rect -830 9613 -796 9647
rect -762 9646 -723 9647
rect -689 9646 -654 9680
rect -620 9646 -585 9680
rect -551 9646 -516 9680
rect -482 9646 -447 9680
rect -413 9646 -378 9680
rect -344 9646 -309 9680
rect -275 9646 -240 9680
rect -206 9646 -171 9680
rect -137 9646 -102 9680
rect -68 9646 -33 9680
rect -762 9613 -33 9646
rect -947 9612 -33 9613
rect -947 9578 -723 9612
rect -689 9578 -654 9612
rect -620 9578 -585 9612
rect -551 9578 -516 9612
rect -482 9578 -447 9612
rect -413 9578 -378 9612
rect -344 9578 -309 9612
rect -275 9578 -240 9612
rect -206 9578 -171 9612
rect -137 9578 -102 9612
rect -68 9578 -33 9612
rect -947 9571 -33 9578
rect -947 9537 -932 9571
rect -898 9537 -864 9571
rect -830 9537 -796 9571
rect -762 9544 -33 9571
rect -762 9537 -723 9544
rect -947 9510 -723 9537
rect -689 9510 -654 9544
rect -620 9510 -585 9544
rect -551 9510 -516 9544
rect -482 9510 -447 9544
rect -413 9510 -378 9544
rect -344 9510 -309 9544
rect -275 9510 -240 9544
rect -206 9510 -171 9544
rect -137 9510 -102 9544
rect -68 9510 -33 9544
rect -947 9495 -33 9510
rect -947 9461 -932 9495
rect -898 9461 -864 9495
rect -830 9461 -796 9495
rect -762 9476 -33 9495
rect -762 9461 -723 9476
rect -947 9442 -723 9461
rect -689 9442 -654 9476
rect -620 9442 -585 9476
rect -551 9442 -516 9476
rect -482 9442 -447 9476
rect -413 9442 -378 9476
rect -344 9442 -309 9476
rect -275 9442 -240 9476
rect -206 9442 -171 9476
rect -137 9442 -102 9476
rect -68 9442 -33 9476
rect -947 9418 -33 9442
rect -947 9384 -932 9418
rect -898 9384 -864 9418
rect -830 9384 -796 9418
rect -762 9408 -33 9418
rect -762 9384 -723 9408
rect -947 9374 -723 9384
rect -689 9374 -654 9408
rect -620 9374 -585 9408
rect -551 9374 -516 9408
rect -482 9374 -447 9408
rect -413 9374 -378 9408
rect -344 9374 -309 9408
rect -275 9374 -240 9408
rect -206 9374 -171 9408
rect -137 9374 -102 9408
rect -68 9374 -33 9408
rect -947 9341 -33 9374
rect -947 9307 -932 9341
rect -898 9307 -864 9341
rect -830 9307 -796 9341
rect -762 9340 -33 9341
rect -762 9307 -723 9340
rect -947 9306 -723 9307
rect -689 9306 -654 9340
rect -620 9306 -585 9340
rect -551 9306 -516 9340
rect -482 9306 -447 9340
rect -413 9306 -378 9340
rect -344 9306 -309 9340
rect -275 9306 -240 9340
rect -206 9306 -171 9340
rect -137 9306 -102 9340
rect -68 9306 -33 9340
rect -947 9272 -33 9306
rect -947 9264 -723 9272
rect -947 9230 -932 9264
rect -898 9230 -864 9264
rect -830 9230 -796 9264
rect -762 9238 -723 9264
rect -689 9238 -654 9272
rect -620 9238 -585 9272
rect -551 9238 -516 9272
rect -482 9238 -447 9272
rect -413 9238 -378 9272
rect -344 9238 -309 9272
rect -275 9238 -240 9272
rect -206 9238 -171 9272
rect -137 9238 -102 9272
rect -68 9238 -33 9272
rect -762 9230 -33 9238
rect -947 9204 -33 9230
rect -947 9187 -723 9204
rect -947 9153 -932 9187
rect -898 9153 -864 9187
rect -830 9153 -796 9187
rect -762 9170 -723 9187
rect -689 9170 -654 9204
rect -620 9170 -585 9204
rect -551 9170 -516 9204
rect -482 9170 -447 9204
rect -413 9170 -378 9204
rect -344 9170 -309 9204
rect -275 9170 -240 9204
rect -206 9170 -171 9204
rect -137 9170 -102 9204
rect -68 9170 -33 9204
rect -762 9153 -33 9170
rect -947 9136 -33 9153
rect -947 9110 -723 9136
rect -947 9076 -932 9110
rect -898 9076 -864 9110
rect -830 9076 -796 9110
rect -762 9102 -723 9110
rect -689 9102 -654 9136
rect -620 9102 -585 9136
rect -551 9102 -516 9136
rect -482 9102 -447 9136
rect -413 9102 -378 9136
rect -344 9102 -309 9136
rect -275 9102 -240 9136
rect -206 9102 -171 9136
rect -137 9102 -102 9136
rect -68 9102 -33 9136
rect -762 9076 -33 9102
rect -947 9068 -33 9076
rect -947 9034 -723 9068
rect -689 9034 -654 9068
rect -620 9034 -585 9068
rect -551 9034 -516 9068
rect -482 9034 -447 9068
rect -413 9034 -378 9068
rect -344 9034 -309 9068
rect -275 9034 -240 9068
rect -206 9034 -171 9068
rect -137 9034 -102 9068
rect -68 9034 -33 9068
rect -947 9033 -33 9034
rect -947 8999 -932 9033
rect -898 8999 -864 9033
rect -830 8999 -796 9033
rect -762 9000 -33 9033
rect -762 8999 -723 9000
rect -947 8966 -723 8999
rect -689 8966 -654 9000
rect -620 8966 -585 9000
rect -551 8966 -516 9000
rect -482 8966 -447 9000
rect -413 8966 -378 9000
rect -344 8966 -309 9000
rect -275 8966 -240 9000
rect -206 8966 -171 9000
rect -137 8966 -102 9000
rect -68 8966 -33 9000
rect 14893 9647 15117 9680
rect 14893 9613 14932 9647
rect 14966 9613 15000 9647
rect 15034 9613 15068 9647
rect 15102 9613 15117 9647
rect 14893 9571 15117 9613
rect 14893 9537 14932 9571
rect 14966 9537 15000 9571
rect 15034 9537 15068 9571
rect 15102 9537 15117 9571
rect 14893 9495 15117 9537
rect 14893 9461 14932 9495
rect 14966 9461 15000 9495
rect 15034 9461 15068 9495
rect 15102 9461 15117 9495
rect 14893 9418 15117 9461
rect 14893 9384 14932 9418
rect 14966 9384 15000 9418
rect 15034 9384 15068 9418
rect 15102 9384 15117 9418
rect 14893 9341 15117 9384
rect 14893 9307 14932 9341
rect 14966 9307 15000 9341
rect 15034 9307 15068 9341
rect 15102 9307 15117 9341
rect 14893 9264 15117 9307
rect 14893 9230 14932 9264
rect 14966 9230 15000 9264
rect 15034 9230 15068 9264
rect 15102 9230 15117 9264
rect 14893 9187 15117 9230
rect 14893 9153 14932 9187
rect 14966 9153 15000 9187
rect 15034 9153 15068 9187
rect 15102 9153 15117 9187
rect 14893 9110 15117 9153
rect 14893 9076 14932 9110
rect 14966 9076 15000 9110
rect 15034 9076 15068 9110
rect 15102 9076 15117 9110
rect 14893 9033 15117 9076
rect 14893 8999 14932 9033
rect 14966 8999 15000 9033
rect 15034 8999 15068 9033
rect 15102 8999 15117 9033
rect 14893 8966 15117 8999
rect -947 8961 15117 8966
rect 44 6809 68 6843
rect 102 6809 137 6843
rect 171 6809 206 6843
rect 240 6809 275 6843
rect 309 6809 344 6843
rect 378 6809 413 6843
rect 447 6809 482 6843
rect 516 6809 551 6843
rect 585 6809 620 6843
rect 654 6809 689 6843
rect 723 6809 758 6843
rect 792 6809 827 6843
rect 861 6809 896 6843
rect 930 6809 965 6843
rect 999 6809 1034 6843
rect 1068 6809 1103 6843
rect 1137 6809 1172 6843
rect 1206 6809 1241 6843
rect 1275 6809 1310 6843
rect 1344 6809 1379 6843
rect 1413 6809 1448 6843
rect 1482 6809 1517 6843
rect 1551 6809 1586 6843
rect 1620 6809 1655 6843
rect 1689 6809 1724 6843
rect 1758 6809 1793 6843
rect 1827 6809 1862 6843
rect 1896 6809 1931 6843
rect 1965 6809 2000 6843
rect 2034 6809 2069 6843
rect 2103 6809 2138 6843
rect 2172 6809 2207 6843
rect 2241 6809 2276 6843
rect 2310 6809 2345 6843
rect 2379 6809 2414 6843
rect 2448 6809 2483 6843
rect 2517 6809 2552 6843
rect 2586 6809 2621 6843
rect 2655 6809 2690 6843
rect 2724 6809 2759 6843
rect 2793 6809 2828 6843
rect 2862 6809 2897 6843
rect 2931 6809 2966 6843
rect 3000 6809 3035 6843
rect 3069 6809 3104 6843
rect 3138 6809 3173 6843
rect 3207 6809 3242 6843
rect 3276 6809 3310 6843
rect 3344 6809 3378 6843
rect 3412 6809 3446 6843
rect 3480 6809 3514 6843
rect 3548 6809 3582 6843
rect 3616 6809 3650 6843
rect 3684 6809 3718 6843
rect 3752 6809 3786 6843
rect 3820 6809 3854 6843
rect 3888 6809 3922 6843
rect 3956 6809 3990 6843
rect 4024 6809 4058 6843
rect 4092 6809 4126 6843
rect 4160 6809 4194 6843
rect 4228 6809 4262 6843
rect 4296 6809 4330 6843
rect 4364 6809 4398 6843
rect 4432 6809 4466 6843
rect 4500 6809 4534 6843
rect 4568 6809 4602 6843
rect 4636 6809 4670 6843
rect 4704 6809 4738 6843
rect 4772 6809 4806 6843
rect 4840 6809 4874 6843
rect 4908 6809 4942 6843
rect 4976 6809 5010 6843
rect 5044 6809 5078 6843
rect 5112 6809 5146 6843
rect 5180 6809 5214 6843
rect 5248 6809 5282 6843
rect 5316 6809 5350 6843
rect 5384 6809 5418 6843
rect 5452 6809 5486 6843
rect 5520 6809 5554 6843
rect 5588 6809 5622 6843
rect 5656 6809 5690 6843
rect 5724 6809 5758 6843
rect 5792 6809 5826 6843
rect 5860 6809 5894 6843
rect 5928 6809 5962 6843
rect 5996 6809 6030 6843
rect 6064 6809 6098 6843
rect 6132 6809 6166 6843
rect 6200 6809 6234 6843
rect 6268 6809 6302 6843
rect 6336 6809 6370 6843
rect 6404 6809 6438 6843
rect 6472 6809 6506 6843
rect 6540 6809 6574 6843
rect 6608 6809 6642 6843
rect 6676 6809 6710 6843
rect 6744 6809 6778 6843
rect 6812 6809 6846 6843
rect 6880 6809 6914 6843
rect 6948 6809 6982 6843
rect 7016 6809 7050 6843
rect 7084 6809 7108 6843
rect 44 6756 7108 6809
rect 44 6722 68 6756
rect 102 6722 137 6756
rect 171 6722 206 6756
rect 240 6722 275 6756
rect 309 6722 344 6756
rect 378 6722 413 6756
rect 447 6722 482 6756
rect 516 6722 551 6756
rect 585 6722 620 6756
rect 654 6722 689 6756
rect 723 6722 758 6756
rect 792 6722 827 6756
rect 861 6722 896 6756
rect 930 6722 965 6756
rect 999 6722 1034 6756
rect 1068 6722 1103 6756
rect 1137 6722 1172 6756
rect 1206 6722 1241 6756
rect 1275 6722 1310 6756
rect 1344 6722 1379 6756
rect 1413 6722 1448 6756
rect 1482 6722 1517 6756
rect 1551 6722 1586 6756
rect 1620 6722 1655 6756
rect 1689 6722 1724 6756
rect 1758 6722 1793 6756
rect 1827 6722 1862 6756
rect 1896 6722 1931 6756
rect 1965 6722 2000 6756
rect 2034 6722 2069 6756
rect 2103 6722 2138 6756
rect 2172 6722 2207 6756
rect 2241 6722 2276 6756
rect 2310 6722 2345 6756
rect 2379 6722 2414 6756
rect 2448 6722 2483 6756
rect 2517 6722 2552 6756
rect 2586 6722 2621 6756
rect 2655 6722 2690 6756
rect 2724 6722 2759 6756
rect 2793 6722 2828 6756
rect 2862 6722 2897 6756
rect 2931 6722 2966 6756
rect 3000 6722 3035 6756
rect 3069 6722 3104 6756
rect 3138 6722 3173 6756
rect 3207 6722 3242 6756
rect 3276 6722 3310 6756
rect 3344 6722 3378 6756
rect 3412 6722 3446 6756
rect 3480 6722 3514 6756
rect 3548 6722 3582 6756
rect 3616 6722 3650 6756
rect 3684 6722 3718 6756
rect 3752 6722 3786 6756
rect 3820 6722 3854 6756
rect 3888 6722 3922 6756
rect 3956 6722 3990 6756
rect 4024 6722 4058 6756
rect 4092 6722 4126 6756
rect 4160 6722 4194 6756
rect 4228 6722 4262 6756
rect 4296 6722 4330 6756
rect 4364 6722 4398 6756
rect 4432 6722 4466 6756
rect 4500 6722 4534 6756
rect 4568 6722 4602 6756
rect 4636 6722 4670 6756
rect 4704 6722 4738 6756
rect 4772 6722 4806 6756
rect 4840 6722 4874 6756
rect 4908 6722 4942 6756
rect 4976 6722 5010 6756
rect 5044 6722 5078 6756
rect 5112 6722 5146 6756
rect 5180 6722 5214 6756
rect 5248 6722 5282 6756
rect 5316 6722 5350 6756
rect 5384 6722 5418 6756
rect 5452 6722 5486 6756
rect 5520 6722 5554 6756
rect 5588 6722 5622 6756
rect 5656 6722 5690 6756
rect 5724 6722 5758 6756
rect 5792 6722 5826 6756
rect 5860 6722 5894 6756
rect 5928 6722 5962 6756
rect 5996 6722 6030 6756
rect 6064 6722 6098 6756
rect 6132 6722 6166 6756
rect 6200 6722 6234 6756
rect 6268 6722 6302 6756
rect 6336 6722 6370 6756
rect 6404 6722 6438 6756
rect 6472 6722 6506 6756
rect 6540 6722 6574 6756
rect 6608 6722 6642 6756
rect 6676 6722 6710 6756
rect 6744 6722 6778 6756
rect 6812 6722 6846 6756
rect 6880 6722 6914 6756
rect 6948 6722 6982 6756
rect 7016 6722 7050 6756
rect 7084 6722 7108 6756
rect 44 6669 7108 6722
rect 44 6635 68 6669
rect 102 6635 137 6669
rect 171 6635 206 6669
rect 240 6635 275 6669
rect 309 6635 344 6669
rect 378 6635 413 6669
rect 447 6635 482 6669
rect 516 6635 551 6669
rect 585 6635 620 6669
rect 654 6635 689 6669
rect 723 6635 758 6669
rect 792 6635 827 6669
rect 861 6635 896 6669
rect 930 6635 965 6669
rect 999 6635 1034 6669
rect 1068 6635 1103 6669
rect 1137 6635 1172 6669
rect 1206 6635 1241 6669
rect 1275 6635 1310 6669
rect 1344 6635 1379 6669
rect 1413 6635 1448 6669
rect 1482 6635 1517 6669
rect 1551 6635 1586 6669
rect 1620 6635 1655 6669
rect 1689 6635 1724 6669
rect 1758 6635 1793 6669
rect 1827 6635 1862 6669
rect 1896 6635 1931 6669
rect 1965 6635 2000 6669
rect 2034 6635 2069 6669
rect 2103 6635 2138 6669
rect 2172 6635 2207 6669
rect 2241 6635 2276 6669
rect 2310 6635 2345 6669
rect 2379 6635 2414 6669
rect 2448 6635 2483 6669
rect 2517 6635 2552 6669
rect 2586 6635 2621 6669
rect 2655 6635 2690 6669
rect 2724 6635 2759 6669
rect 2793 6635 2828 6669
rect 2862 6635 2897 6669
rect 2931 6635 2966 6669
rect 3000 6635 3035 6669
rect 3069 6635 3104 6669
rect 3138 6635 3173 6669
rect 3207 6635 3242 6669
rect 3276 6635 3310 6669
rect 3344 6635 3378 6669
rect 3412 6635 3446 6669
rect 3480 6635 3514 6669
rect 3548 6635 3582 6669
rect 3616 6635 3650 6669
rect 3684 6635 3718 6669
rect 3752 6635 3786 6669
rect 3820 6635 3854 6669
rect 3888 6635 3922 6669
rect 3956 6635 3990 6669
rect 4024 6635 4058 6669
rect 4092 6635 4126 6669
rect 4160 6635 4194 6669
rect 4228 6635 4262 6669
rect 4296 6635 4330 6669
rect 4364 6635 4398 6669
rect 4432 6635 4466 6669
rect 4500 6635 4534 6669
rect 4568 6635 4602 6669
rect 4636 6635 4670 6669
rect 4704 6635 4738 6669
rect 4772 6635 4806 6669
rect 4840 6635 4874 6669
rect 4908 6635 4942 6669
rect 4976 6635 5010 6669
rect 5044 6635 5078 6669
rect 5112 6635 5146 6669
rect 5180 6635 5214 6669
rect 5248 6635 5282 6669
rect 5316 6635 5350 6669
rect 5384 6635 5418 6669
rect 5452 6635 5486 6669
rect 5520 6635 5554 6669
rect 5588 6635 5622 6669
rect 5656 6635 5690 6669
rect 5724 6635 5758 6669
rect 5792 6635 5826 6669
rect 5860 6635 5894 6669
rect 5928 6635 5962 6669
rect 5996 6635 6030 6669
rect 6064 6635 6098 6669
rect 6132 6635 6166 6669
rect 6200 6635 6234 6669
rect 6268 6635 6302 6669
rect 6336 6635 6370 6669
rect 6404 6635 6438 6669
rect 6472 6635 6506 6669
rect 6540 6635 6574 6669
rect 6608 6635 6642 6669
rect 6676 6635 6710 6669
rect 6744 6635 6778 6669
rect 6812 6635 6846 6669
rect 6880 6635 6914 6669
rect 6948 6635 6982 6669
rect 7016 6635 7050 6669
rect 7084 6635 7108 6669
rect 12493 6809 12517 6843
rect 12551 6809 12586 6843
rect 12620 6809 12655 6843
rect 12689 6809 12724 6843
rect 12758 6809 12793 6843
rect 12827 6809 12862 6843
rect 12896 6809 12931 6843
rect 12965 6809 13000 6843
rect 13034 6809 13069 6843
rect 13103 6809 13138 6843
rect 13172 6809 13207 6843
rect 13241 6809 13276 6843
rect 13310 6809 13345 6843
rect 13379 6809 13414 6843
rect 13448 6809 13483 6843
rect 13517 6809 13552 6843
rect 13586 6809 13621 6843
rect 13655 6809 13690 6843
rect 13724 6809 13759 6843
rect 13793 6809 13828 6843
rect 13862 6809 13897 6843
rect 13931 6809 13966 6843
rect 14000 6809 14035 6843
rect 14069 6809 14104 6843
rect 14138 6809 14173 6843
rect 14207 6809 14242 6843
rect 14276 6809 14311 6843
rect 14345 6809 14380 6843
rect 14414 6809 14449 6843
rect 14483 6809 14518 6843
rect 14552 6809 14587 6843
rect 14621 6809 14655 6843
rect 14689 6809 14723 6843
rect 14757 6809 14791 6843
rect 14825 6809 14859 6843
rect 14893 6809 15117 6843
rect 12493 6805 15117 6809
rect 12493 6771 14932 6805
rect 14966 6771 15000 6805
rect 15034 6771 15068 6805
rect 15102 6771 15117 6805
rect 12493 6756 15117 6771
rect 12493 6722 12517 6756
rect 12551 6722 12586 6756
rect 12620 6722 12655 6756
rect 12689 6722 12724 6756
rect 12758 6722 12793 6756
rect 12827 6722 12862 6756
rect 12896 6722 12931 6756
rect 12965 6722 13000 6756
rect 13034 6722 13069 6756
rect 13103 6722 13138 6756
rect 13172 6722 13207 6756
rect 13241 6722 13276 6756
rect 13310 6722 13345 6756
rect 13379 6722 13414 6756
rect 13448 6722 13483 6756
rect 13517 6722 13552 6756
rect 13586 6722 13621 6756
rect 13655 6722 13690 6756
rect 13724 6722 13759 6756
rect 13793 6722 13828 6756
rect 13862 6722 13897 6756
rect 13931 6722 13966 6756
rect 14000 6722 14035 6756
rect 14069 6722 14104 6756
rect 14138 6722 14173 6756
rect 14207 6722 14242 6756
rect 14276 6722 14311 6756
rect 14345 6722 14380 6756
rect 14414 6722 14449 6756
rect 14483 6722 14518 6756
rect 14552 6722 14587 6756
rect 14621 6722 14655 6756
rect 14689 6722 14723 6756
rect 14757 6722 14791 6756
rect 14825 6722 14859 6756
rect 14893 6731 15117 6756
rect 14893 6722 14932 6731
rect 12493 6697 14932 6722
rect 14966 6697 15000 6731
rect 15034 6697 15068 6731
rect 15102 6697 15117 6731
rect 12493 6669 15117 6697
rect 12493 6635 12517 6669
rect 12551 6635 12586 6669
rect 12620 6635 12655 6669
rect 12689 6635 12724 6669
rect 12758 6635 12793 6669
rect 12827 6635 12862 6669
rect 12896 6635 12931 6669
rect 12965 6635 13000 6669
rect 13034 6635 13069 6669
rect 13103 6635 13138 6669
rect 13172 6635 13207 6669
rect 13241 6635 13276 6669
rect 13310 6635 13345 6669
rect 13379 6635 13414 6669
rect 13448 6635 13483 6669
rect 13517 6635 13552 6669
rect 13586 6635 13621 6669
rect 13655 6635 13690 6669
rect 13724 6635 13759 6669
rect 13793 6635 13828 6669
rect 13862 6635 13897 6669
rect 13931 6635 13966 6669
rect 14000 6635 14035 6669
rect 14069 6635 14104 6669
rect 14138 6635 14173 6669
rect 14207 6635 14242 6669
rect 14276 6635 14311 6669
rect 14345 6635 14380 6669
rect 14414 6635 14449 6669
rect 14483 6635 14518 6669
rect 14552 6635 14587 6669
rect 14621 6635 14655 6669
rect 14689 6635 14723 6669
rect 14757 6635 14791 6669
rect 14825 6635 14859 6669
rect 14893 6657 15117 6669
rect 14893 6635 14932 6657
rect 44 6623 14932 6635
rect 14966 6623 15000 6657
rect 15034 6623 15068 6657
rect 15102 6623 15117 6657
rect 44 6583 15117 6623
rect 44 6582 14932 6583
rect 44 6548 68 6582
rect 102 6548 137 6582
rect 171 6548 206 6582
rect 240 6548 275 6582
rect 309 6548 344 6582
rect 378 6548 413 6582
rect 447 6548 482 6582
rect 516 6548 551 6582
rect 585 6548 620 6582
rect 654 6548 689 6582
rect 723 6548 758 6582
rect 792 6548 827 6582
rect 861 6548 896 6582
rect 930 6548 965 6582
rect 999 6548 1034 6582
rect 1068 6548 1103 6582
rect 1137 6548 1172 6582
rect 1206 6548 1241 6582
rect 1275 6548 1310 6582
rect 1344 6548 1379 6582
rect 1413 6548 1448 6582
rect 1482 6548 1517 6582
rect 1551 6548 1586 6582
rect 1620 6548 1655 6582
rect 1689 6548 1724 6582
rect 1758 6548 1793 6582
rect 1827 6548 1862 6582
rect 1896 6548 1931 6582
rect 1965 6548 2000 6582
rect 2034 6548 2069 6582
rect 2103 6548 2138 6582
rect 2172 6548 2207 6582
rect 2241 6548 2276 6582
rect 2310 6548 2345 6582
rect 2379 6548 2414 6582
rect 2448 6548 2483 6582
rect 2517 6548 2551 6582
rect 2585 6548 2619 6582
rect 2653 6548 2687 6582
rect 2721 6548 2755 6582
rect 2789 6548 2823 6582
rect 2857 6548 2891 6582
rect 2925 6548 2959 6582
rect 2993 6548 3027 6582
rect 3061 6548 3095 6582
rect 3129 6548 3163 6582
rect 3197 6548 3231 6582
rect 3265 6548 3299 6582
rect 3333 6548 3367 6582
rect 3401 6548 3435 6582
rect 3469 6548 3503 6582
rect 3537 6548 3571 6582
rect 3605 6548 3639 6582
rect 3673 6548 3707 6582
rect 3741 6548 3775 6582
rect 3809 6548 3843 6582
rect 3877 6548 3911 6582
rect 3945 6548 3979 6582
rect 4013 6548 4047 6582
rect 4081 6548 4115 6582
rect 4149 6548 4183 6582
rect 4217 6548 4251 6582
rect 4285 6548 4319 6582
rect 4353 6548 4387 6582
rect 4421 6548 4455 6582
rect 4489 6548 4523 6582
rect 4557 6548 4591 6582
rect 4625 6548 4659 6582
rect 4693 6548 4727 6582
rect 4761 6548 4795 6582
rect 4829 6548 4863 6582
rect 4897 6548 4931 6582
rect 4965 6548 4999 6582
rect 5033 6548 5067 6582
rect 5101 6548 5135 6582
rect 5169 6548 5203 6582
rect 5237 6548 5271 6582
rect 5305 6548 5339 6582
rect 5373 6548 5407 6582
rect 5441 6548 5475 6582
rect 5509 6548 5543 6582
rect 5577 6548 5611 6582
rect 5645 6548 5679 6582
rect 5713 6548 5747 6582
rect 5781 6548 5815 6582
rect 5849 6548 5883 6582
rect 5917 6548 5951 6582
rect 5985 6548 6019 6582
rect 6053 6548 6087 6582
rect 6121 6548 6155 6582
rect 6189 6548 6223 6582
rect 6257 6548 6291 6582
rect 6325 6548 6359 6582
rect 6393 6548 6427 6582
rect 6461 6548 6495 6582
rect 6529 6548 6563 6582
rect 6597 6548 6631 6582
rect 6665 6548 6699 6582
rect 6733 6548 6767 6582
rect 6801 6548 6835 6582
rect 6869 6548 6903 6582
rect 6937 6548 6971 6582
rect 7005 6548 7039 6582
rect 7073 6548 7107 6582
rect 7141 6548 7175 6582
rect 7209 6548 7243 6582
rect 7277 6548 7311 6582
rect 7345 6548 7379 6582
rect 7413 6548 7447 6582
rect 7481 6548 7515 6582
rect 7549 6548 7583 6582
rect 7617 6548 7651 6582
rect 7685 6548 7719 6582
rect 7753 6548 7787 6582
rect 7821 6548 7855 6582
rect 7889 6548 7923 6582
rect 7957 6548 7991 6582
rect 8025 6548 8059 6582
rect 8093 6548 8127 6582
rect 8161 6548 8195 6582
rect 8229 6548 8263 6582
rect 8297 6548 8331 6582
rect 8365 6548 8399 6582
rect 8433 6548 8467 6582
rect 8501 6548 8535 6582
rect 8569 6548 8603 6582
rect 8637 6548 8671 6582
rect 8705 6548 8739 6582
rect 8773 6548 8807 6582
rect 8841 6548 8875 6582
rect 8909 6548 8943 6582
rect 8977 6548 9011 6582
rect 9045 6548 9079 6582
rect 9113 6548 9147 6582
rect 9181 6548 9215 6582
rect 9249 6548 9283 6582
rect 9317 6548 9351 6582
rect 9385 6548 9419 6582
rect 9453 6548 9487 6582
rect 9521 6548 9555 6582
rect 9589 6548 9623 6582
rect 9657 6548 9691 6582
rect 9725 6548 9759 6582
rect 9793 6548 9827 6582
rect 9861 6548 9895 6582
rect 9929 6548 9963 6582
rect 9997 6548 10031 6582
rect 10065 6548 10099 6582
rect 10133 6548 10167 6582
rect 10201 6548 10235 6582
rect 10269 6548 10303 6582
rect 10337 6548 10371 6582
rect 10405 6548 10439 6582
rect 10473 6548 10507 6582
rect 10541 6548 10575 6582
rect 10609 6548 10643 6582
rect 10677 6548 10711 6582
rect 10745 6548 10779 6582
rect 10813 6548 10847 6582
rect 10881 6548 10915 6582
rect 10949 6548 10983 6582
rect 11017 6548 11051 6582
rect 11085 6548 11119 6582
rect 11153 6548 11187 6582
rect 11221 6548 11255 6582
rect 11289 6548 11323 6582
rect 11357 6548 11391 6582
rect 11425 6548 11459 6582
rect 11493 6548 11527 6582
rect 11561 6548 11595 6582
rect 11629 6548 11663 6582
rect 11697 6548 11731 6582
rect 11765 6548 11799 6582
rect 11833 6548 11867 6582
rect 11901 6548 11935 6582
rect 11969 6548 12003 6582
rect 12037 6548 12071 6582
rect 12105 6548 12139 6582
rect 12173 6548 12207 6582
rect 12241 6548 12275 6582
rect 12309 6548 12343 6582
rect 12377 6548 12411 6582
rect 12445 6548 12479 6582
rect 12513 6548 12547 6582
rect 12581 6548 12615 6582
rect 12649 6548 12683 6582
rect 12717 6548 12751 6582
rect 12785 6548 12819 6582
rect 12853 6548 12887 6582
rect 12921 6548 12955 6582
rect 12989 6548 13023 6582
rect 13057 6548 13091 6582
rect 13125 6548 13159 6582
rect 13193 6548 13227 6582
rect 13261 6548 13295 6582
rect 13329 6548 13363 6582
rect 13397 6548 13431 6582
rect 13465 6548 13499 6582
rect 13533 6548 13567 6582
rect 13601 6548 13635 6582
rect 13669 6548 13703 6582
rect 13737 6548 13771 6582
rect 13805 6548 13839 6582
rect 13873 6548 13907 6582
rect 13941 6548 13975 6582
rect 14009 6548 14043 6582
rect 14077 6548 14111 6582
rect 14145 6548 14179 6582
rect 14213 6548 14247 6582
rect 14281 6548 14315 6582
rect 14349 6548 14383 6582
rect 14417 6548 14451 6582
rect 14485 6548 14519 6582
rect 14553 6548 14587 6582
rect 14621 6548 14655 6582
rect 14689 6548 14723 6582
rect 14757 6548 14791 6582
rect 14825 6548 14859 6582
rect 14893 6549 14932 6582
rect 14966 6549 15000 6583
rect 15034 6549 15068 6583
rect 15102 6549 15117 6583
rect 14893 6548 15117 6549
rect 44 6509 15117 6548
rect 44 6508 14932 6509
rect 44 6474 68 6508
rect 102 6474 137 6508
rect 171 6474 206 6508
rect 240 6474 275 6508
rect 309 6474 344 6508
rect 378 6474 413 6508
rect 447 6474 482 6508
rect 516 6474 551 6508
rect 585 6474 620 6508
rect 654 6474 689 6508
rect 723 6474 758 6508
rect 792 6474 827 6508
rect 861 6474 896 6508
rect 930 6474 965 6508
rect 999 6474 1034 6508
rect 1068 6474 1103 6508
rect 1137 6474 1172 6508
rect 1206 6474 1241 6508
rect 1275 6474 1310 6508
rect 1344 6474 1379 6508
rect 1413 6474 1448 6508
rect 1482 6474 1517 6508
rect 1551 6474 1586 6508
rect 1620 6474 1655 6508
rect 1689 6474 1724 6508
rect 1758 6474 1793 6508
rect 1827 6474 1862 6508
rect 1896 6474 1931 6508
rect 1965 6474 2000 6508
rect 2034 6474 2069 6508
rect 2103 6474 2138 6508
rect 2172 6474 2207 6508
rect 2241 6474 2276 6508
rect 2310 6474 2345 6508
rect 2379 6474 2414 6508
rect 2448 6474 2483 6508
rect 2517 6474 2551 6508
rect 2585 6474 2619 6508
rect 2653 6474 2687 6508
rect 2721 6474 2755 6508
rect 2789 6474 2823 6508
rect 2857 6474 2891 6508
rect 2925 6474 2959 6508
rect 2993 6474 3027 6508
rect 3061 6474 3095 6508
rect 3129 6474 3163 6508
rect 3197 6474 3231 6508
rect 3265 6474 3299 6508
rect 3333 6474 3367 6508
rect 3401 6474 3435 6508
rect 3469 6474 3503 6508
rect 3537 6474 3571 6508
rect 3605 6474 3639 6508
rect 3673 6474 3707 6508
rect 3741 6474 3775 6508
rect 3809 6474 3843 6508
rect 3877 6474 3911 6508
rect 3945 6474 3979 6508
rect 4013 6474 4047 6508
rect 4081 6474 4115 6508
rect 4149 6474 4183 6508
rect 4217 6474 4251 6508
rect 4285 6474 4319 6508
rect 4353 6474 4387 6508
rect 4421 6474 4455 6508
rect 4489 6474 4523 6508
rect 4557 6474 4591 6508
rect 4625 6474 4659 6508
rect 4693 6474 4727 6508
rect 4761 6474 4795 6508
rect 4829 6474 4863 6508
rect 4897 6474 4931 6508
rect 4965 6474 4999 6508
rect 5033 6474 5067 6508
rect 5101 6474 5135 6508
rect 5169 6474 5203 6508
rect 5237 6474 5271 6508
rect 5305 6474 5339 6508
rect 5373 6474 5407 6508
rect 5441 6474 5475 6508
rect 5509 6474 5543 6508
rect 5577 6474 5611 6508
rect 5645 6474 5679 6508
rect 5713 6474 5747 6508
rect 5781 6474 5815 6508
rect 5849 6474 5883 6508
rect 5917 6474 5951 6508
rect 5985 6474 6019 6508
rect 6053 6474 6087 6508
rect 6121 6474 6155 6508
rect 6189 6474 6223 6508
rect 6257 6474 6291 6508
rect 6325 6474 6359 6508
rect 6393 6474 6427 6508
rect 6461 6474 6495 6508
rect 6529 6474 6563 6508
rect 6597 6474 6631 6508
rect 6665 6474 6699 6508
rect 6733 6474 6767 6508
rect 6801 6474 6835 6508
rect 6869 6474 6903 6508
rect 6937 6474 6971 6508
rect 7005 6474 7039 6508
rect 7073 6474 7107 6508
rect 7141 6474 7175 6508
rect 7209 6474 7243 6508
rect 7277 6474 7311 6508
rect 7345 6474 7379 6508
rect 7413 6474 7447 6508
rect 7481 6474 7515 6508
rect 7549 6474 7583 6508
rect 7617 6474 7651 6508
rect 7685 6474 7719 6508
rect 7753 6474 7787 6508
rect 7821 6474 7855 6508
rect 7889 6474 7923 6508
rect 7957 6474 7991 6508
rect 8025 6474 8059 6508
rect 8093 6474 8127 6508
rect 8161 6474 8195 6508
rect 8229 6474 8263 6508
rect 8297 6474 8331 6508
rect 8365 6474 8399 6508
rect 8433 6474 8467 6508
rect 8501 6474 8535 6508
rect 8569 6474 8603 6508
rect 8637 6474 8671 6508
rect 8705 6474 8739 6508
rect 8773 6474 8807 6508
rect 8841 6474 8875 6508
rect 8909 6474 8943 6508
rect 8977 6474 9011 6508
rect 9045 6474 9079 6508
rect 9113 6474 9147 6508
rect 9181 6474 9215 6508
rect 9249 6474 9283 6508
rect 9317 6474 9351 6508
rect 9385 6474 9419 6508
rect 9453 6474 9487 6508
rect 9521 6474 9555 6508
rect 9589 6474 9623 6508
rect 9657 6474 9691 6508
rect 9725 6474 9759 6508
rect 9793 6474 9827 6508
rect 9861 6474 9895 6508
rect 9929 6474 9963 6508
rect 9997 6474 10031 6508
rect 10065 6474 10099 6508
rect 10133 6474 10167 6508
rect 10201 6474 10235 6508
rect 10269 6474 10303 6508
rect 10337 6474 10371 6508
rect 10405 6474 10439 6508
rect 10473 6474 10507 6508
rect 10541 6474 10575 6508
rect 10609 6474 10643 6508
rect 10677 6474 10711 6508
rect 10745 6474 10779 6508
rect 10813 6474 10847 6508
rect 10881 6474 10915 6508
rect 10949 6474 10983 6508
rect 11017 6474 11051 6508
rect 11085 6474 11119 6508
rect 11153 6474 11187 6508
rect 11221 6474 11255 6508
rect 11289 6474 11323 6508
rect 11357 6474 11391 6508
rect 11425 6474 11459 6508
rect 11493 6474 11527 6508
rect 11561 6474 11595 6508
rect 11629 6474 11663 6508
rect 11697 6474 11731 6508
rect 11765 6474 11799 6508
rect 11833 6474 11867 6508
rect 11901 6474 11935 6508
rect 11969 6474 12003 6508
rect 12037 6474 12071 6508
rect 12105 6474 12139 6508
rect 12173 6474 12207 6508
rect 12241 6474 12275 6508
rect 12309 6474 12343 6508
rect 12377 6474 12411 6508
rect 12445 6474 12479 6508
rect 12513 6474 12547 6508
rect 12581 6474 12615 6508
rect 12649 6474 12683 6508
rect 12717 6474 12751 6508
rect 12785 6474 12819 6508
rect 12853 6474 12887 6508
rect 12921 6474 12955 6508
rect 12989 6474 13023 6508
rect 13057 6474 13091 6508
rect 13125 6474 13159 6508
rect 13193 6474 13227 6508
rect 13261 6474 13295 6508
rect 13329 6474 13363 6508
rect 13397 6474 13431 6508
rect 13465 6474 13499 6508
rect 13533 6474 13567 6508
rect 13601 6474 13635 6508
rect 13669 6474 13703 6508
rect 13737 6474 13771 6508
rect 13805 6474 13839 6508
rect 13873 6474 13907 6508
rect 13941 6474 13975 6508
rect 14009 6474 14043 6508
rect 14077 6474 14111 6508
rect 14145 6474 14179 6508
rect 14213 6474 14247 6508
rect 14281 6474 14315 6508
rect 14349 6474 14383 6508
rect 14417 6474 14451 6508
rect 14485 6474 14519 6508
rect 14553 6474 14587 6508
rect 14621 6474 14655 6508
rect 14689 6474 14723 6508
rect 14757 6474 14791 6508
rect 14825 6474 14859 6508
rect 14893 6475 14932 6508
rect 14966 6475 15000 6509
rect 15034 6475 15068 6509
rect 15102 6475 15117 6509
rect 14893 6474 15117 6475
rect 44 6435 15117 6474
rect 44 6434 14932 6435
rect 44 6400 68 6434
rect 102 6400 137 6434
rect 171 6400 206 6434
rect 240 6400 275 6434
rect 309 6400 344 6434
rect 378 6400 413 6434
rect 447 6400 482 6434
rect 516 6400 551 6434
rect 585 6400 620 6434
rect 654 6400 689 6434
rect 723 6400 758 6434
rect 792 6400 827 6434
rect 861 6400 896 6434
rect 930 6400 965 6434
rect 999 6400 1034 6434
rect 1068 6400 1103 6434
rect 1137 6400 1172 6434
rect 1206 6400 1241 6434
rect 1275 6400 1310 6434
rect 1344 6400 1379 6434
rect 1413 6400 1448 6434
rect 1482 6400 1517 6434
rect 1551 6400 1586 6434
rect 1620 6400 1655 6434
rect 1689 6400 1724 6434
rect 1758 6400 1793 6434
rect 1827 6400 1862 6434
rect 1896 6400 1931 6434
rect 1965 6400 2000 6434
rect 2034 6400 2069 6434
rect 2103 6400 2138 6434
rect 2172 6400 2207 6434
rect 2241 6400 2276 6434
rect 2310 6400 2345 6434
rect 2379 6400 2414 6434
rect 2448 6400 2483 6434
rect 2517 6400 2551 6434
rect 2585 6400 2619 6434
rect 2653 6400 2687 6434
rect 2721 6400 2755 6434
rect 2789 6400 2823 6434
rect 2857 6400 2891 6434
rect 2925 6400 2959 6434
rect 2993 6400 3027 6434
rect 3061 6400 3095 6434
rect 3129 6400 3163 6434
rect 3197 6400 3231 6434
rect 3265 6400 3299 6434
rect 3333 6400 3367 6434
rect 3401 6400 3435 6434
rect 3469 6400 3503 6434
rect 3537 6400 3571 6434
rect 3605 6400 3639 6434
rect 3673 6400 3707 6434
rect 3741 6400 3775 6434
rect 3809 6400 3843 6434
rect 3877 6400 3911 6434
rect 3945 6400 3979 6434
rect 4013 6400 4047 6434
rect 4081 6400 4115 6434
rect 4149 6400 4183 6434
rect 4217 6400 4251 6434
rect 4285 6400 4319 6434
rect 4353 6400 4387 6434
rect 4421 6400 4455 6434
rect 4489 6400 4523 6434
rect 4557 6400 4591 6434
rect 4625 6400 4659 6434
rect 4693 6400 4727 6434
rect 4761 6400 4795 6434
rect 4829 6400 4863 6434
rect 4897 6400 4931 6434
rect 4965 6400 4999 6434
rect 5033 6400 5067 6434
rect 5101 6400 5135 6434
rect 5169 6400 5203 6434
rect 5237 6400 5271 6434
rect 5305 6400 5339 6434
rect 5373 6400 5407 6434
rect 5441 6400 5475 6434
rect 5509 6400 5543 6434
rect 5577 6400 5611 6434
rect 5645 6400 5679 6434
rect 5713 6400 5747 6434
rect 5781 6400 5815 6434
rect 5849 6400 5883 6434
rect 5917 6400 5951 6434
rect 5985 6400 6019 6434
rect 6053 6400 6087 6434
rect 6121 6400 6155 6434
rect 6189 6400 6223 6434
rect 6257 6400 6291 6434
rect 6325 6400 6359 6434
rect 6393 6400 6427 6434
rect 6461 6400 6495 6434
rect 6529 6400 6563 6434
rect 6597 6400 6631 6434
rect 6665 6400 6699 6434
rect 6733 6400 6767 6434
rect 6801 6400 6835 6434
rect 6869 6400 6903 6434
rect 6937 6400 6971 6434
rect 7005 6400 7039 6434
rect 7073 6400 7107 6434
rect 7141 6400 7175 6434
rect 7209 6400 7243 6434
rect 7277 6400 7311 6434
rect 7345 6400 7379 6434
rect 7413 6400 7447 6434
rect 7481 6400 7515 6434
rect 7549 6400 7583 6434
rect 7617 6400 7651 6434
rect 7685 6400 7719 6434
rect 7753 6400 7787 6434
rect 7821 6400 7855 6434
rect 7889 6400 7923 6434
rect 7957 6400 7991 6434
rect 8025 6400 8059 6434
rect 8093 6400 8127 6434
rect 8161 6400 8195 6434
rect 8229 6400 8263 6434
rect 8297 6400 8331 6434
rect 8365 6400 8399 6434
rect 8433 6400 8467 6434
rect 8501 6400 8535 6434
rect 8569 6400 8603 6434
rect 8637 6400 8671 6434
rect 8705 6400 8739 6434
rect 8773 6400 8807 6434
rect 8841 6400 8875 6434
rect 8909 6400 8943 6434
rect 8977 6400 9011 6434
rect 9045 6400 9079 6434
rect 9113 6400 9147 6434
rect 9181 6400 9215 6434
rect 9249 6400 9283 6434
rect 9317 6400 9351 6434
rect 9385 6400 9419 6434
rect 9453 6400 9487 6434
rect 9521 6400 9555 6434
rect 9589 6400 9623 6434
rect 9657 6400 9691 6434
rect 9725 6400 9759 6434
rect 9793 6400 9827 6434
rect 9861 6400 9895 6434
rect 9929 6400 9963 6434
rect 9997 6400 10031 6434
rect 10065 6400 10099 6434
rect 10133 6400 10167 6434
rect 10201 6400 10235 6434
rect 10269 6400 10303 6434
rect 10337 6400 10371 6434
rect 10405 6400 10439 6434
rect 10473 6400 10507 6434
rect 10541 6400 10575 6434
rect 10609 6400 10643 6434
rect 10677 6400 10711 6434
rect 10745 6400 10779 6434
rect 10813 6400 10847 6434
rect 10881 6400 10915 6434
rect 10949 6400 10983 6434
rect 11017 6400 11051 6434
rect 11085 6400 11119 6434
rect 11153 6400 11187 6434
rect 11221 6400 11255 6434
rect 11289 6400 11323 6434
rect 11357 6400 11391 6434
rect 11425 6400 11459 6434
rect 11493 6400 11527 6434
rect 11561 6400 11595 6434
rect 11629 6400 11663 6434
rect 11697 6400 11731 6434
rect 11765 6400 11799 6434
rect 11833 6400 11867 6434
rect 11901 6400 11935 6434
rect 11969 6400 12003 6434
rect 12037 6400 12071 6434
rect 12105 6400 12139 6434
rect 12173 6400 12207 6434
rect 12241 6400 12275 6434
rect 12309 6400 12343 6434
rect 12377 6400 12411 6434
rect 12445 6400 12479 6434
rect 12513 6400 12547 6434
rect 12581 6400 12615 6434
rect 12649 6400 12683 6434
rect 12717 6400 12751 6434
rect 12785 6400 12819 6434
rect 12853 6400 12887 6434
rect 12921 6400 12955 6434
rect 12989 6400 13023 6434
rect 13057 6400 13091 6434
rect 13125 6400 13159 6434
rect 13193 6400 13227 6434
rect 13261 6400 13295 6434
rect 13329 6400 13363 6434
rect 13397 6400 13431 6434
rect 13465 6400 13499 6434
rect 13533 6400 13567 6434
rect 13601 6400 13635 6434
rect 13669 6400 13703 6434
rect 13737 6400 13771 6434
rect 13805 6400 13839 6434
rect 13873 6400 13907 6434
rect 13941 6400 13975 6434
rect 14009 6400 14043 6434
rect 14077 6400 14111 6434
rect 14145 6400 14179 6434
rect 14213 6400 14247 6434
rect 14281 6400 14315 6434
rect 14349 6400 14383 6434
rect 14417 6400 14451 6434
rect 14485 6400 14519 6434
rect 14553 6400 14587 6434
rect 14621 6400 14655 6434
rect 14689 6400 14723 6434
rect 14757 6400 14791 6434
rect 14825 6400 14859 6434
rect 14893 6401 14932 6434
rect 14966 6401 15000 6435
rect 15034 6401 15068 6435
rect 15102 6401 15117 6435
rect 14893 6400 15117 6401
rect 44 6360 15117 6400
rect 44 6326 68 6360
rect 102 6326 137 6360
rect 171 6326 206 6360
rect 240 6326 275 6360
rect 309 6326 344 6360
rect 378 6326 413 6360
rect 447 6326 482 6360
rect 516 6326 551 6360
rect 585 6326 620 6360
rect 654 6326 689 6360
rect 723 6326 758 6360
rect 792 6326 827 6360
rect 861 6326 896 6360
rect 930 6326 965 6360
rect 999 6326 1034 6360
rect 1068 6326 1103 6360
rect 1137 6326 1172 6360
rect 1206 6326 1241 6360
rect 1275 6326 1310 6360
rect 1344 6326 1379 6360
rect 1413 6326 1448 6360
rect 1482 6326 1517 6360
rect 1551 6326 1586 6360
rect 1620 6326 1655 6360
rect 1689 6326 1724 6360
rect 1758 6326 1793 6360
rect 1827 6326 1862 6360
rect 1896 6326 1931 6360
rect 1965 6326 2000 6360
rect 2034 6326 2069 6360
rect 2103 6326 2138 6360
rect 2172 6326 2207 6360
rect 2241 6326 2276 6360
rect 2310 6326 2345 6360
rect 2379 6326 2414 6360
rect 2448 6326 2483 6360
rect 2517 6326 2551 6360
rect 2585 6326 2619 6360
rect 2653 6326 2687 6360
rect 2721 6326 2755 6360
rect 2789 6326 2823 6360
rect 2857 6326 2891 6360
rect 2925 6326 2959 6360
rect 2993 6326 3027 6360
rect 3061 6326 3095 6360
rect 3129 6326 3163 6360
rect 3197 6326 3231 6360
rect 3265 6326 3299 6360
rect 3333 6326 3367 6360
rect 3401 6326 3435 6360
rect 3469 6326 3503 6360
rect 3537 6326 3571 6360
rect 3605 6326 3639 6360
rect 3673 6326 3707 6360
rect 3741 6326 3775 6360
rect 3809 6326 3843 6360
rect 3877 6326 3911 6360
rect 3945 6326 3979 6360
rect 4013 6326 4047 6360
rect 4081 6326 4115 6360
rect 4149 6326 4183 6360
rect 4217 6326 4251 6360
rect 4285 6326 4319 6360
rect 4353 6326 4387 6360
rect 4421 6326 4455 6360
rect 4489 6326 4523 6360
rect 4557 6326 4591 6360
rect 4625 6326 4659 6360
rect 4693 6326 4727 6360
rect 4761 6326 4795 6360
rect 4829 6326 4863 6360
rect 4897 6326 4931 6360
rect 4965 6326 4999 6360
rect 5033 6326 5067 6360
rect 5101 6326 5135 6360
rect 5169 6326 5203 6360
rect 5237 6326 5271 6360
rect 5305 6326 5339 6360
rect 5373 6326 5407 6360
rect 5441 6326 5475 6360
rect 5509 6326 5543 6360
rect 5577 6326 5611 6360
rect 5645 6326 5679 6360
rect 5713 6326 5747 6360
rect 5781 6326 5815 6360
rect 5849 6326 5883 6360
rect 5917 6326 5951 6360
rect 5985 6326 6019 6360
rect 6053 6326 6087 6360
rect 6121 6326 6155 6360
rect 6189 6326 6223 6360
rect 6257 6326 6291 6360
rect 6325 6326 6359 6360
rect 6393 6326 6427 6360
rect 6461 6326 6495 6360
rect 6529 6326 6563 6360
rect 6597 6326 6631 6360
rect 6665 6326 6699 6360
rect 6733 6326 6767 6360
rect 6801 6326 6835 6360
rect 6869 6326 6903 6360
rect 6937 6326 6971 6360
rect 7005 6326 7039 6360
rect 7073 6326 7107 6360
rect 7141 6326 7175 6360
rect 7209 6326 7243 6360
rect 7277 6326 7311 6360
rect 7345 6326 7379 6360
rect 7413 6326 7447 6360
rect 7481 6326 7515 6360
rect 7549 6326 7583 6360
rect 7617 6326 7651 6360
rect 7685 6326 7719 6360
rect 7753 6326 7787 6360
rect 7821 6326 7855 6360
rect 7889 6326 7923 6360
rect 7957 6326 7991 6360
rect 8025 6326 8059 6360
rect 8093 6326 8127 6360
rect 8161 6326 8195 6360
rect 8229 6326 8263 6360
rect 8297 6326 8331 6360
rect 8365 6326 8399 6360
rect 8433 6326 8467 6360
rect 8501 6326 8535 6360
rect 8569 6326 8603 6360
rect 8637 6326 8671 6360
rect 8705 6326 8739 6360
rect 8773 6326 8807 6360
rect 8841 6326 8875 6360
rect 8909 6326 8943 6360
rect 8977 6326 9011 6360
rect 9045 6326 9079 6360
rect 9113 6326 9147 6360
rect 9181 6326 9215 6360
rect 9249 6326 9283 6360
rect 9317 6326 9351 6360
rect 9385 6326 9419 6360
rect 9453 6326 9487 6360
rect 9521 6326 9555 6360
rect 9589 6326 9623 6360
rect 9657 6326 9691 6360
rect 9725 6326 9759 6360
rect 9793 6326 9827 6360
rect 9861 6326 9895 6360
rect 9929 6326 9963 6360
rect 9997 6326 10031 6360
rect 10065 6326 10099 6360
rect 10133 6326 10167 6360
rect 10201 6326 10235 6360
rect 10269 6326 10303 6360
rect 10337 6326 10371 6360
rect 10405 6326 10439 6360
rect 10473 6326 10507 6360
rect 10541 6326 10575 6360
rect 10609 6326 10643 6360
rect 10677 6326 10711 6360
rect 10745 6326 10779 6360
rect 10813 6326 10847 6360
rect 10881 6326 10915 6360
rect 10949 6326 10983 6360
rect 11017 6326 11051 6360
rect 11085 6326 11119 6360
rect 11153 6326 11187 6360
rect 11221 6326 11255 6360
rect 11289 6326 11323 6360
rect 11357 6326 11391 6360
rect 11425 6326 11459 6360
rect 11493 6326 11527 6360
rect 11561 6326 11595 6360
rect 11629 6326 11663 6360
rect 11697 6326 11731 6360
rect 11765 6326 11799 6360
rect 11833 6326 11867 6360
rect 11901 6326 11935 6360
rect 11969 6326 12003 6360
rect 12037 6326 12071 6360
rect 12105 6326 12139 6360
rect 12173 6326 12207 6360
rect 12241 6326 12275 6360
rect 12309 6326 12343 6360
rect 12377 6326 12411 6360
rect 12445 6326 12479 6360
rect 12513 6326 12547 6360
rect 12581 6326 12615 6360
rect 12649 6326 12683 6360
rect 12717 6326 12751 6360
rect 12785 6326 12819 6360
rect 12853 6326 12887 6360
rect 12921 6326 12955 6360
rect 12989 6326 13023 6360
rect 13057 6326 13091 6360
rect 13125 6326 13159 6360
rect 13193 6326 13227 6360
rect 13261 6326 13295 6360
rect 13329 6326 13363 6360
rect 13397 6326 13431 6360
rect 13465 6326 13499 6360
rect 13533 6326 13567 6360
rect 13601 6326 13635 6360
rect 13669 6326 13703 6360
rect 13737 6326 13771 6360
rect 13805 6326 13839 6360
rect 13873 6326 13907 6360
rect 13941 6326 13975 6360
rect 14009 6326 14043 6360
rect 14077 6326 14111 6360
rect 14145 6326 14179 6360
rect 14213 6326 14247 6360
rect 14281 6326 14315 6360
rect 14349 6326 14383 6360
rect 14417 6326 14451 6360
rect 14485 6326 14519 6360
rect 14553 6326 14587 6360
rect 14621 6326 14655 6360
rect 14689 6326 14723 6360
rect 14757 6326 14791 6360
rect 14825 6326 14859 6360
rect 14893 6326 14932 6360
rect 14966 6326 15000 6360
rect 15034 6326 15068 6360
rect 15102 6326 15117 6360
rect 44 6286 15117 6326
rect 44 6252 68 6286
rect 102 6252 137 6286
rect 171 6252 206 6286
rect 240 6252 275 6286
rect 309 6252 344 6286
rect 378 6252 413 6286
rect 447 6252 482 6286
rect 516 6252 551 6286
rect 585 6252 620 6286
rect 654 6252 689 6286
rect 723 6252 758 6286
rect 792 6252 827 6286
rect 861 6252 896 6286
rect 930 6252 965 6286
rect 999 6252 1034 6286
rect 1068 6252 1103 6286
rect 1137 6252 1172 6286
rect 1206 6252 1241 6286
rect 1275 6252 1310 6286
rect 1344 6252 1379 6286
rect 1413 6252 1448 6286
rect 1482 6252 1517 6286
rect 1551 6252 1586 6286
rect 1620 6252 1655 6286
rect 1689 6252 1724 6286
rect 1758 6252 1793 6286
rect 1827 6252 1862 6286
rect 1896 6252 1931 6286
rect 1965 6252 2000 6286
rect 2034 6252 2069 6286
rect 2103 6252 2138 6286
rect 2172 6252 2207 6286
rect 2241 6252 2276 6286
rect 2310 6252 2345 6286
rect 2379 6252 2414 6286
rect 2448 6252 2483 6286
rect 2517 6252 2551 6286
rect 2585 6252 2619 6286
rect 2653 6252 2687 6286
rect 2721 6252 2755 6286
rect 2789 6252 2823 6286
rect 2857 6252 2891 6286
rect 2925 6252 2959 6286
rect 2993 6252 3027 6286
rect 3061 6252 3095 6286
rect 3129 6252 3163 6286
rect 3197 6252 3231 6286
rect 3265 6252 3299 6286
rect 3333 6252 3367 6286
rect 3401 6252 3435 6286
rect 3469 6252 3503 6286
rect 3537 6252 3571 6286
rect 3605 6252 3639 6286
rect 3673 6252 3707 6286
rect 3741 6252 3775 6286
rect 3809 6252 3843 6286
rect 3877 6252 3911 6286
rect 3945 6252 3979 6286
rect 4013 6252 4047 6286
rect 4081 6252 4115 6286
rect 4149 6252 4183 6286
rect 4217 6252 4251 6286
rect 4285 6252 4319 6286
rect 4353 6252 4387 6286
rect 4421 6252 4455 6286
rect 4489 6252 4523 6286
rect 4557 6252 4591 6286
rect 4625 6252 4659 6286
rect 4693 6252 4727 6286
rect 4761 6252 4795 6286
rect 4829 6252 4863 6286
rect 4897 6252 4931 6286
rect 4965 6252 4999 6286
rect 5033 6252 5067 6286
rect 5101 6252 5135 6286
rect 5169 6252 5203 6286
rect 5237 6252 5271 6286
rect 5305 6252 5339 6286
rect 5373 6252 5407 6286
rect 5441 6252 5475 6286
rect 5509 6252 5543 6286
rect 5577 6252 5611 6286
rect 5645 6252 5679 6286
rect 5713 6252 5747 6286
rect 5781 6252 5815 6286
rect 5849 6252 5883 6286
rect 5917 6252 5951 6286
rect 5985 6252 6019 6286
rect 6053 6252 6087 6286
rect 6121 6252 6155 6286
rect 6189 6252 6223 6286
rect 6257 6252 6291 6286
rect 6325 6252 6359 6286
rect 6393 6252 6427 6286
rect 6461 6252 6495 6286
rect 6529 6252 6563 6286
rect 6597 6252 6631 6286
rect 6665 6252 6699 6286
rect 6733 6252 6767 6286
rect 6801 6252 6835 6286
rect 6869 6252 6903 6286
rect 6937 6252 6971 6286
rect 7005 6252 7039 6286
rect 7073 6252 7107 6286
rect 7141 6252 7175 6286
rect 7209 6252 7243 6286
rect 7277 6252 7311 6286
rect 7345 6252 7379 6286
rect 7413 6252 7447 6286
rect 7481 6252 7515 6286
rect 7549 6252 7583 6286
rect 7617 6252 7651 6286
rect 7685 6252 7719 6286
rect 7753 6252 7787 6286
rect 7821 6252 7855 6286
rect 7889 6252 7923 6286
rect 7957 6252 7991 6286
rect 8025 6252 8059 6286
rect 8093 6252 8127 6286
rect 8161 6252 8195 6286
rect 8229 6252 8263 6286
rect 8297 6252 8331 6286
rect 8365 6252 8399 6286
rect 8433 6252 8467 6286
rect 8501 6252 8535 6286
rect 8569 6252 8603 6286
rect 8637 6252 8671 6286
rect 8705 6252 8739 6286
rect 8773 6252 8807 6286
rect 8841 6252 8875 6286
rect 8909 6252 8943 6286
rect 8977 6252 9011 6286
rect 9045 6252 9079 6286
rect 9113 6252 9147 6286
rect 9181 6252 9215 6286
rect 9249 6252 9283 6286
rect 9317 6252 9351 6286
rect 9385 6252 9419 6286
rect 9453 6252 9487 6286
rect 9521 6252 9555 6286
rect 9589 6252 9623 6286
rect 9657 6252 9691 6286
rect 9725 6252 9759 6286
rect 9793 6252 9827 6286
rect 9861 6252 9895 6286
rect 9929 6252 9963 6286
rect 9997 6252 10031 6286
rect 10065 6252 10099 6286
rect 10133 6252 10167 6286
rect 10201 6252 10235 6286
rect 10269 6252 10303 6286
rect 10337 6252 10371 6286
rect 10405 6252 10439 6286
rect 10473 6252 10507 6286
rect 10541 6252 10575 6286
rect 10609 6252 10643 6286
rect 10677 6252 10711 6286
rect 10745 6252 10779 6286
rect 10813 6252 10847 6286
rect 10881 6252 10915 6286
rect 10949 6252 10983 6286
rect 11017 6252 11051 6286
rect 11085 6252 11119 6286
rect 11153 6252 11187 6286
rect 11221 6252 11255 6286
rect 11289 6252 11323 6286
rect 11357 6252 11391 6286
rect 11425 6252 11459 6286
rect 11493 6252 11527 6286
rect 11561 6252 11595 6286
rect 11629 6252 11663 6286
rect 11697 6252 11731 6286
rect 11765 6252 11799 6286
rect 11833 6252 11867 6286
rect 11901 6252 11935 6286
rect 11969 6252 12003 6286
rect 12037 6252 12071 6286
rect 12105 6252 12139 6286
rect 12173 6252 12207 6286
rect 12241 6252 12275 6286
rect 12309 6252 12343 6286
rect 12377 6252 12411 6286
rect 12445 6252 12479 6286
rect 12513 6252 12547 6286
rect 12581 6252 12615 6286
rect 12649 6252 12683 6286
rect 12717 6252 12751 6286
rect 12785 6252 12819 6286
rect 12853 6252 12887 6286
rect 12921 6252 12955 6286
rect 12989 6252 13023 6286
rect 13057 6252 13091 6286
rect 13125 6252 13159 6286
rect 13193 6252 13227 6286
rect 13261 6252 13295 6286
rect 13329 6252 13363 6286
rect 13397 6252 13431 6286
rect 13465 6252 13499 6286
rect 13533 6252 13567 6286
rect 13601 6252 13635 6286
rect 13669 6252 13703 6286
rect 13737 6252 13771 6286
rect 13805 6252 13839 6286
rect 13873 6252 13907 6286
rect 13941 6252 13975 6286
rect 14009 6252 14043 6286
rect 14077 6252 14111 6286
rect 14145 6252 14179 6286
rect 14213 6252 14247 6286
rect 14281 6252 14315 6286
rect 14349 6252 14383 6286
rect 14417 6252 14451 6286
rect 14485 6252 14519 6286
rect 14553 6252 14587 6286
rect 14621 6252 14655 6286
rect 14689 6252 14723 6286
rect 14757 6252 14791 6286
rect 14825 6252 14859 6286
rect 14893 6285 15117 6286
rect 14893 6252 14932 6285
rect 44 6251 14932 6252
rect 14966 6251 15000 6285
rect 15034 6251 15068 6285
rect 15102 6251 15117 6285
rect 44 6212 15117 6251
rect 44 6178 68 6212
rect 102 6178 137 6212
rect 171 6178 206 6212
rect 240 6178 275 6212
rect 309 6178 344 6212
rect 378 6178 413 6212
rect 447 6178 482 6212
rect 516 6178 551 6212
rect 585 6178 620 6212
rect 654 6178 689 6212
rect 723 6178 758 6212
rect 792 6178 827 6212
rect 861 6178 896 6212
rect 930 6178 965 6212
rect 999 6178 1034 6212
rect 1068 6178 1103 6212
rect 1137 6178 1172 6212
rect 1206 6178 1241 6212
rect 1275 6178 1310 6212
rect 1344 6178 1379 6212
rect 1413 6178 1448 6212
rect 1482 6178 1517 6212
rect 1551 6178 1586 6212
rect 1620 6178 1655 6212
rect 1689 6178 1724 6212
rect 1758 6178 1793 6212
rect 1827 6178 1862 6212
rect 1896 6178 1931 6212
rect 1965 6178 2000 6212
rect 2034 6178 2069 6212
rect 2103 6178 2138 6212
rect 2172 6178 2207 6212
rect 2241 6178 2276 6212
rect 2310 6178 2345 6212
rect 2379 6178 2414 6212
rect 2448 6178 2483 6212
rect 2517 6178 2551 6212
rect 2585 6178 2619 6212
rect 2653 6178 2687 6212
rect 2721 6178 2755 6212
rect 2789 6178 2823 6212
rect 2857 6178 2891 6212
rect 2925 6178 2959 6212
rect 2993 6178 3027 6212
rect 3061 6178 3095 6212
rect 3129 6178 3163 6212
rect 3197 6178 3231 6212
rect 3265 6178 3299 6212
rect 3333 6178 3367 6212
rect 3401 6178 3435 6212
rect 3469 6178 3503 6212
rect 3537 6178 3571 6212
rect 3605 6178 3639 6212
rect 3673 6178 3707 6212
rect 3741 6178 3775 6212
rect 3809 6178 3843 6212
rect 3877 6178 3911 6212
rect 3945 6178 3979 6212
rect 4013 6178 4047 6212
rect 4081 6178 4115 6212
rect 4149 6178 4183 6212
rect 4217 6178 4251 6212
rect 4285 6178 4319 6212
rect 4353 6178 4387 6212
rect 4421 6178 4455 6212
rect 4489 6178 4523 6212
rect 4557 6178 4591 6212
rect 4625 6178 4659 6212
rect 4693 6178 4727 6212
rect 4761 6178 4795 6212
rect 4829 6178 4863 6212
rect 4897 6178 4931 6212
rect 4965 6178 4999 6212
rect 5033 6178 5067 6212
rect 5101 6178 5135 6212
rect 5169 6178 5203 6212
rect 5237 6178 5271 6212
rect 5305 6178 5339 6212
rect 5373 6178 5407 6212
rect 5441 6178 5475 6212
rect 5509 6178 5543 6212
rect 5577 6178 5611 6212
rect 5645 6178 5679 6212
rect 5713 6178 5747 6212
rect 5781 6178 5815 6212
rect 5849 6178 5883 6212
rect 5917 6178 5951 6212
rect 5985 6178 6019 6212
rect 6053 6178 6087 6212
rect 6121 6178 6155 6212
rect 6189 6178 6223 6212
rect 6257 6178 6291 6212
rect 6325 6178 6359 6212
rect 6393 6178 6427 6212
rect 6461 6178 6495 6212
rect 6529 6178 6563 6212
rect 6597 6178 6631 6212
rect 6665 6178 6699 6212
rect 6733 6178 6767 6212
rect 6801 6178 6835 6212
rect 6869 6178 6903 6212
rect 6937 6178 6971 6212
rect 7005 6178 7039 6212
rect 7073 6178 7107 6212
rect 7141 6178 7175 6212
rect 7209 6178 7243 6212
rect 7277 6178 7311 6212
rect 7345 6178 7379 6212
rect 7413 6178 7447 6212
rect 7481 6178 7515 6212
rect 7549 6178 7583 6212
rect 7617 6178 7651 6212
rect 7685 6178 7719 6212
rect 7753 6178 7787 6212
rect 7821 6178 7855 6212
rect 7889 6178 7923 6212
rect 7957 6178 7991 6212
rect 8025 6178 8059 6212
rect 8093 6178 8127 6212
rect 8161 6178 8195 6212
rect 8229 6178 8263 6212
rect 8297 6178 8331 6212
rect 8365 6178 8399 6212
rect 8433 6178 8467 6212
rect 8501 6178 8535 6212
rect 8569 6178 8603 6212
rect 8637 6178 8671 6212
rect 8705 6178 8739 6212
rect 8773 6178 8807 6212
rect 8841 6178 8875 6212
rect 8909 6178 8943 6212
rect 8977 6178 9011 6212
rect 9045 6178 9079 6212
rect 9113 6178 9147 6212
rect 9181 6178 9215 6212
rect 9249 6178 9283 6212
rect 9317 6178 9351 6212
rect 9385 6178 9419 6212
rect 9453 6178 9487 6212
rect 9521 6178 9555 6212
rect 9589 6178 9623 6212
rect 9657 6178 9691 6212
rect 9725 6178 9759 6212
rect 9793 6178 9827 6212
rect 9861 6178 9895 6212
rect 9929 6178 9963 6212
rect 9997 6178 10031 6212
rect 10065 6178 10099 6212
rect 10133 6178 10167 6212
rect 10201 6178 10235 6212
rect 10269 6178 10303 6212
rect 10337 6178 10371 6212
rect 10405 6178 10439 6212
rect 10473 6178 10507 6212
rect 10541 6178 10575 6212
rect 10609 6178 10643 6212
rect 10677 6178 10711 6212
rect 10745 6178 10779 6212
rect 10813 6178 10847 6212
rect 10881 6178 10915 6212
rect 10949 6178 10983 6212
rect 11017 6178 11051 6212
rect 11085 6178 11119 6212
rect 11153 6178 11187 6212
rect 11221 6178 11255 6212
rect 11289 6178 11323 6212
rect 11357 6178 11391 6212
rect 11425 6178 11459 6212
rect 11493 6178 11527 6212
rect 11561 6178 11595 6212
rect 11629 6178 11663 6212
rect 11697 6178 11731 6212
rect 11765 6178 11799 6212
rect 11833 6178 11867 6212
rect 11901 6178 11935 6212
rect 11969 6178 12003 6212
rect 12037 6178 12071 6212
rect 12105 6178 12139 6212
rect 12173 6178 12207 6212
rect 12241 6178 12275 6212
rect 12309 6178 12343 6212
rect 12377 6178 12411 6212
rect 12445 6178 12479 6212
rect 12513 6178 12547 6212
rect 12581 6178 12615 6212
rect 12649 6178 12683 6212
rect 12717 6178 12751 6212
rect 12785 6178 12819 6212
rect 12853 6178 12887 6212
rect 12921 6178 12955 6212
rect 12989 6178 13023 6212
rect 13057 6178 13091 6212
rect 13125 6178 13159 6212
rect 13193 6178 13227 6212
rect 13261 6178 13295 6212
rect 13329 6178 13363 6212
rect 13397 6178 13431 6212
rect 13465 6178 13499 6212
rect 13533 6178 13567 6212
rect 13601 6178 13635 6212
rect 13669 6178 13703 6212
rect 13737 6178 13771 6212
rect 13805 6178 13839 6212
rect 13873 6178 13907 6212
rect 13941 6178 13975 6212
rect 14009 6178 14043 6212
rect 14077 6178 14111 6212
rect 14145 6178 14179 6212
rect 14213 6178 14247 6212
rect 14281 6178 14315 6212
rect 14349 6178 14383 6212
rect 14417 6178 14451 6212
rect 14485 6178 14519 6212
rect 14553 6178 14587 6212
rect 14621 6178 14655 6212
rect 14689 6178 14723 6212
rect 14757 6178 14791 6212
rect 14825 6178 14859 6212
rect 14893 6210 15117 6212
rect 14893 6178 14932 6210
rect 44 6176 14932 6178
rect 14966 6176 15000 6210
rect 15034 6176 15068 6210
rect 15102 6176 15117 6210
rect 44 6138 15117 6176
rect 44 6104 68 6138
rect 102 6104 137 6138
rect 171 6104 206 6138
rect 240 6104 275 6138
rect 309 6104 344 6138
rect 378 6104 413 6138
rect 447 6104 482 6138
rect 516 6104 551 6138
rect 585 6104 620 6138
rect 654 6104 689 6138
rect 723 6104 758 6138
rect 792 6104 827 6138
rect 861 6104 896 6138
rect 930 6104 965 6138
rect 999 6104 1034 6138
rect 1068 6104 1103 6138
rect 1137 6104 1172 6138
rect 1206 6104 1241 6138
rect 1275 6104 1310 6138
rect 1344 6104 1379 6138
rect 1413 6104 1448 6138
rect 1482 6104 1517 6138
rect 1551 6104 1586 6138
rect 1620 6104 1655 6138
rect 1689 6104 1724 6138
rect 1758 6104 1793 6138
rect 1827 6104 1862 6138
rect 1896 6104 1931 6138
rect 1965 6104 2000 6138
rect 2034 6104 2069 6138
rect 2103 6104 2138 6138
rect 2172 6104 2207 6138
rect 2241 6104 2276 6138
rect 2310 6104 2345 6138
rect 2379 6104 2414 6138
rect 2448 6104 2483 6138
rect 2517 6104 2551 6138
rect 2585 6104 2619 6138
rect 2653 6104 2687 6138
rect 2721 6104 2755 6138
rect 2789 6104 2823 6138
rect 2857 6104 2891 6138
rect 2925 6104 2959 6138
rect 2993 6104 3027 6138
rect 3061 6104 3095 6138
rect 3129 6104 3163 6138
rect 3197 6104 3231 6138
rect 3265 6104 3299 6138
rect 3333 6104 3367 6138
rect 3401 6104 3435 6138
rect 3469 6104 3503 6138
rect 3537 6104 3571 6138
rect 3605 6104 3639 6138
rect 3673 6104 3707 6138
rect 3741 6104 3775 6138
rect 3809 6104 3843 6138
rect 3877 6104 3911 6138
rect 3945 6104 3979 6138
rect 4013 6104 4047 6138
rect 4081 6104 4115 6138
rect 4149 6104 4183 6138
rect 4217 6104 4251 6138
rect 4285 6104 4319 6138
rect 4353 6104 4387 6138
rect 4421 6104 4455 6138
rect 4489 6104 4523 6138
rect 4557 6104 4591 6138
rect 4625 6104 4659 6138
rect 4693 6104 4727 6138
rect 4761 6104 4795 6138
rect 4829 6104 4863 6138
rect 4897 6104 4931 6138
rect 4965 6104 4999 6138
rect 5033 6104 5067 6138
rect 5101 6104 5135 6138
rect 5169 6104 5203 6138
rect 5237 6104 5271 6138
rect 5305 6104 5339 6138
rect 5373 6104 5407 6138
rect 5441 6104 5475 6138
rect 5509 6104 5543 6138
rect 5577 6104 5611 6138
rect 5645 6104 5679 6138
rect 5713 6104 5747 6138
rect 5781 6104 5815 6138
rect 5849 6104 5883 6138
rect 5917 6104 5951 6138
rect 5985 6104 6019 6138
rect 6053 6104 6087 6138
rect 6121 6104 6155 6138
rect 6189 6104 6223 6138
rect 6257 6104 6291 6138
rect 6325 6104 6359 6138
rect 6393 6104 6427 6138
rect 6461 6104 6495 6138
rect 6529 6104 6563 6138
rect 6597 6104 6631 6138
rect 6665 6104 6699 6138
rect 6733 6104 6767 6138
rect 6801 6104 6835 6138
rect 6869 6104 6903 6138
rect 6937 6104 6971 6138
rect 7005 6104 7039 6138
rect 7073 6104 7107 6138
rect 7141 6104 7175 6138
rect 7209 6104 7243 6138
rect 7277 6104 7311 6138
rect 7345 6104 7379 6138
rect 7413 6104 7447 6138
rect 7481 6104 7515 6138
rect 7549 6104 7583 6138
rect 7617 6104 7651 6138
rect 7685 6104 7719 6138
rect 7753 6104 7787 6138
rect 7821 6104 7855 6138
rect 7889 6104 7923 6138
rect 7957 6104 7991 6138
rect 8025 6104 8059 6138
rect 8093 6104 8127 6138
rect 8161 6104 8195 6138
rect 8229 6104 8263 6138
rect 8297 6104 8331 6138
rect 8365 6104 8399 6138
rect 8433 6104 8467 6138
rect 8501 6104 8535 6138
rect 8569 6104 8603 6138
rect 8637 6104 8671 6138
rect 8705 6104 8739 6138
rect 8773 6104 8807 6138
rect 8841 6104 8875 6138
rect 8909 6104 8943 6138
rect 8977 6104 9011 6138
rect 9045 6104 9079 6138
rect 9113 6104 9147 6138
rect 9181 6104 9215 6138
rect 9249 6104 9283 6138
rect 9317 6104 9351 6138
rect 9385 6104 9419 6138
rect 9453 6104 9487 6138
rect 9521 6104 9555 6138
rect 9589 6104 9623 6138
rect 9657 6104 9691 6138
rect 9725 6104 9759 6138
rect 9793 6104 9827 6138
rect 9861 6104 9895 6138
rect 9929 6104 9963 6138
rect 9997 6104 10031 6138
rect 10065 6104 10099 6138
rect 10133 6104 10167 6138
rect 10201 6104 10235 6138
rect 10269 6104 10303 6138
rect 10337 6104 10371 6138
rect 10405 6104 10439 6138
rect 10473 6104 10507 6138
rect 10541 6104 10575 6138
rect 10609 6104 10643 6138
rect 10677 6104 10711 6138
rect 10745 6104 10779 6138
rect 10813 6104 10847 6138
rect 10881 6104 10915 6138
rect 10949 6104 10983 6138
rect 11017 6104 11051 6138
rect 11085 6104 11119 6138
rect 11153 6104 11187 6138
rect 11221 6104 11255 6138
rect 11289 6104 11323 6138
rect 11357 6104 11391 6138
rect 11425 6104 11459 6138
rect 11493 6104 11527 6138
rect 11561 6104 11595 6138
rect 11629 6104 11663 6138
rect 11697 6104 11731 6138
rect 11765 6104 11799 6138
rect 11833 6104 11867 6138
rect 11901 6104 11935 6138
rect 11969 6104 12003 6138
rect 12037 6104 12071 6138
rect 12105 6104 12139 6138
rect 12173 6104 12207 6138
rect 12241 6104 12275 6138
rect 12309 6104 12343 6138
rect 12377 6104 12411 6138
rect 12445 6104 12479 6138
rect 12513 6104 12547 6138
rect 12581 6104 12615 6138
rect 12649 6104 12683 6138
rect 12717 6104 12751 6138
rect 12785 6104 12819 6138
rect 12853 6104 12887 6138
rect 12921 6104 12955 6138
rect 12989 6104 13023 6138
rect 13057 6104 13091 6138
rect 13125 6104 13159 6138
rect 13193 6104 13227 6138
rect 13261 6104 13295 6138
rect 13329 6104 13363 6138
rect 13397 6104 13431 6138
rect 13465 6104 13499 6138
rect 13533 6104 13567 6138
rect 13601 6104 13635 6138
rect 13669 6104 13703 6138
rect 13737 6104 13771 6138
rect 13805 6104 13839 6138
rect 13873 6104 13907 6138
rect 13941 6104 13975 6138
rect 14009 6104 14043 6138
rect 14077 6104 14111 6138
rect 14145 6104 14179 6138
rect 14213 6104 14247 6138
rect 14281 6104 14315 6138
rect 14349 6104 14383 6138
rect 14417 6104 14451 6138
rect 14485 6104 14519 6138
rect 14553 6104 14587 6138
rect 14621 6104 14655 6138
rect 14689 6104 14723 6138
rect 14757 6104 14791 6138
rect 14825 6104 14859 6138
rect 14893 6135 15117 6138
rect 14893 6104 14932 6135
rect 44 6101 14932 6104
rect 14966 6101 15000 6135
rect 15034 6101 15068 6135
rect 15102 6101 15117 6135
rect 44 6060 15117 6101
rect 44 6051 14932 6060
rect 14917 6026 14932 6051
rect 14966 6026 15000 6060
rect 15034 6026 15068 6060
rect 15102 6026 15117 6060
rect 14917 5988 15117 6026
rect 14977 5954 15117 5988
rect 14977 4628 15000 5954
rect 15102 4628 15117 5954
rect 14977 4593 15117 4628
rect 14977 4559 15000 4593
rect 15034 4559 15068 4593
rect 15102 4559 15117 4593
rect 14977 4524 15117 4559
rect 14977 4490 15000 4524
rect 15034 4490 15068 4524
rect 15102 4490 15117 4524
rect 14977 4455 15117 4490
rect 14977 4421 15000 4455
rect 15034 4421 15068 4455
rect 15102 4421 15117 4455
rect 14977 4386 15117 4421
rect 14977 4352 15000 4386
rect 15034 4352 15068 4386
rect 15102 4352 15117 4386
rect 14977 4317 15117 4352
rect 14977 4283 15000 4317
rect 15034 4283 15068 4317
rect 15102 4283 15117 4317
rect 14977 4248 15117 4283
rect 14977 4214 15000 4248
rect 15034 4214 15068 4248
rect 15102 4214 15117 4248
rect 14977 4179 15117 4214
rect 14977 4145 15000 4179
rect 15034 4145 15068 4179
rect 15102 4145 15117 4179
rect 14977 4110 15117 4145
rect 14977 4076 15000 4110
rect 15034 4076 15068 4110
rect 15102 4076 15117 4110
rect 14977 4041 15117 4076
rect 14977 4007 15000 4041
rect 15034 4007 15068 4041
rect 15102 4007 15117 4041
rect 14977 3972 15117 4007
rect 14977 3938 15000 3972
rect 15034 3938 15068 3972
rect 15102 3938 15117 3972
rect 14977 3903 15117 3938
rect 14977 3869 15000 3903
rect 15034 3869 15068 3903
rect 15102 3869 15117 3903
rect 14977 3834 15117 3869
rect 14977 3800 15000 3834
rect 15034 3800 15068 3834
rect 15102 3800 15117 3834
rect 14977 3765 15117 3800
rect 14977 3731 15000 3765
rect 15034 3731 15068 3765
rect 15102 3731 15117 3765
rect 14977 3696 15117 3731
rect 14977 3662 15000 3696
rect 15034 3662 15068 3696
rect 15102 3662 15117 3696
rect 14977 3627 15117 3662
rect 14977 3593 15000 3627
rect 15034 3593 15068 3627
rect 15102 3593 15117 3627
rect 14977 3558 15117 3593
rect 14977 3524 15000 3558
rect 15034 3524 15068 3558
rect 15102 3524 15117 3558
rect 14977 3489 15117 3524
rect 14977 3455 15000 3489
rect 15034 3455 15068 3489
rect 15102 3455 15117 3489
rect 14977 3420 15117 3455
rect 14977 3386 15000 3420
rect 15034 3386 15068 3420
rect 15102 3386 15117 3420
rect 14977 3351 15117 3386
rect 14977 3317 15000 3351
rect 15034 3317 15068 3351
rect 15102 3317 15117 3351
rect 14977 3282 15117 3317
rect 14977 3248 15000 3282
rect 15034 3248 15068 3282
rect 15102 3248 15117 3282
rect 14977 3213 15117 3248
rect 14977 3179 15000 3213
rect 15034 3179 15068 3213
rect 15102 3179 15117 3213
rect 14977 3144 15117 3179
rect 14977 3110 15000 3144
rect 15034 3110 15068 3144
rect 15102 3110 15117 3144
rect 14977 3075 15117 3110
rect 14977 3041 15000 3075
rect 15034 3041 15068 3075
rect 15102 3041 15117 3075
rect 14977 3006 15117 3041
rect 14977 2972 15000 3006
rect 15034 2972 15068 3006
rect 15102 2972 15117 3006
rect 14977 2937 15117 2972
rect 14977 2903 15000 2937
rect 15034 2903 15068 2937
rect 15102 2903 15117 2937
rect 14977 2868 15117 2903
rect 14977 2834 15000 2868
rect 15034 2834 15068 2868
rect 15102 2834 15117 2868
rect 14977 2799 15117 2834
rect 14977 2765 15000 2799
rect 15034 2765 15068 2799
rect 15102 2765 15117 2799
rect 14977 2730 15117 2765
rect 14977 2696 15000 2730
rect 15034 2696 15068 2730
rect 15102 2696 15117 2730
rect 14977 2661 15117 2696
rect 14977 2627 15000 2661
rect 15034 2627 15068 2661
rect 15102 2627 15117 2661
rect 14977 2592 15117 2627
rect 14977 2558 15000 2592
rect 15034 2558 15068 2592
rect 15102 2558 15117 2592
rect 14977 2523 15117 2558
rect 14977 2489 15000 2523
rect 15034 2489 15068 2523
rect 15102 2489 15117 2523
rect 14977 2454 15117 2489
rect 14977 2420 15000 2454
rect 15034 2420 15068 2454
rect 15102 2420 15117 2454
rect 14977 2385 15117 2420
rect 14977 2351 15000 2385
rect 15034 2351 15068 2385
rect 15102 2351 15117 2385
rect 14977 2316 15117 2351
rect 14977 2282 15000 2316
rect 15034 2282 15068 2316
rect 15102 2282 15117 2316
rect 14977 2247 15117 2282
rect 14977 2213 15000 2247
rect 15034 2213 15068 2247
rect 15102 2213 15117 2247
rect 14977 2178 15117 2213
rect 14977 2144 15000 2178
rect 15034 2144 15068 2178
rect 15102 2144 15117 2178
rect 14977 2109 15117 2144
rect 14977 2075 15000 2109
rect 15034 2075 15068 2109
rect 15102 2075 15117 2109
rect 14977 2040 15117 2075
rect 14977 2006 15000 2040
rect 15034 2006 15068 2040
rect 15102 2006 15117 2040
rect 14977 1971 15117 2006
rect 14977 1937 15000 1971
rect 15034 1937 15068 1971
rect 15102 1937 15117 1971
rect 14977 1902 15117 1937
rect 14977 1868 15000 1902
rect 15034 1868 15068 1902
rect 15102 1868 15117 1902
rect 14977 1833 15117 1868
rect 14977 1799 15000 1833
rect 15034 1799 15068 1833
rect 15102 1799 15117 1833
rect 14977 1764 15117 1799
rect 14977 1730 15000 1764
rect 15034 1730 15068 1764
rect 15102 1730 15117 1764
rect 14977 1695 15117 1730
rect 14977 1661 15000 1695
rect 15034 1661 15068 1695
rect 15102 1661 15117 1695
rect 14977 1626 15117 1661
rect 14977 1592 15000 1626
rect 15034 1592 15068 1626
rect 15102 1592 15117 1626
rect 14977 1557 15117 1592
rect 14977 1523 15000 1557
rect 15034 1523 15068 1557
rect 15102 1523 15117 1557
rect 14977 1488 15117 1523
rect 14977 1454 15000 1488
rect 15034 1454 15068 1488
rect 15102 1454 15117 1488
rect 14977 1419 15117 1454
rect 14977 1385 15000 1419
rect 15034 1385 15068 1419
rect 15102 1385 15117 1419
rect 14977 1350 15117 1385
rect 14977 1316 15000 1350
rect 15034 1316 15068 1350
rect 15102 1316 15117 1350
rect 7044 1282 14917 1288
rect 14977 1282 15117 1316
rect 3427 1257 15117 1282
rect 3427 1251 7068 1257
rect 3537 1217 3577 1251
rect 3611 1217 3645 1251
rect 3679 1217 3713 1251
rect 3747 1217 3781 1251
rect 3815 1217 3849 1251
rect 3883 1217 3917 1251
rect 3951 1217 3985 1251
rect 4019 1217 4053 1251
rect 4087 1217 4121 1251
rect 4155 1217 4189 1251
rect 4223 1217 4257 1251
rect 4291 1217 4325 1251
rect 4359 1217 4393 1251
rect 4427 1217 4461 1251
rect 4495 1217 4529 1251
rect 4563 1217 4597 1251
rect 4631 1217 4665 1251
rect 4699 1217 4733 1251
rect 4767 1217 4801 1251
rect 4835 1217 4869 1251
rect 4903 1217 4937 1251
rect 4971 1217 5005 1251
rect 5039 1217 5073 1251
rect 5107 1217 5141 1251
rect 5175 1217 5209 1251
rect 5243 1217 5277 1251
rect 5311 1217 5345 1251
rect 5379 1217 5413 1251
rect 5447 1217 5481 1251
rect 5515 1217 5549 1251
rect 5583 1217 5617 1251
rect 5651 1217 5685 1251
rect 5719 1217 5753 1251
rect 5787 1217 5821 1251
rect 5855 1217 5889 1251
rect 5923 1217 5957 1251
rect 5991 1217 6025 1251
rect 6059 1217 6093 1251
rect 6127 1217 6161 1251
rect 6195 1217 6229 1251
rect 6263 1217 6297 1251
rect 6331 1217 6365 1251
rect 6399 1217 6433 1251
rect 6467 1217 6501 1251
rect 6535 1217 6569 1251
rect 6603 1217 6637 1251
rect 6671 1217 6705 1251
rect 6739 1217 6773 1251
rect 6807 1217 6841 1251
rect 6875 1217 6909 1251
rect 6943 1227 7068 1251
rect 6943 1217 6988 1227
rect 7022 1223 7068 1227
rect 7102 1223 7137 1257
rect 7171 1223 7206 1257
rect 7240 1223 7275 1257
rect 7309 1223 7344 1257
rect 7378 1223 7413 1257
rect 7447 1223 7482 1257
rect 7516 1223 7551 1257
rect 7585 1223 7620 1257
rect 7654 1223 7689 1257
rect 7723 1223 7758 1257
rect 7792 1223 7827 1257
rect 7861 1223 7896 1257
rect 7930 1223 7965 1257
rect 7999 1223 8034 1257
rect 8068 1223 8103 1257
rect 8137 1223 8172 1257
rect 8206 1223 8241 1257
rect 8275 1223 8310 1257
rect 8344 1223 8379 1257
rect 8413 1223 8448 1257
rect 8482 1223 8517 1257
rect 8551 1223 8586 1257
rect 8620 1223 8655 1257
rect 8689 1223 8724 1257
rect 8758 1223 8793 1257
rect 8827 1223 8862 1257
rect 8896 1223 8931 1257
rect 8965 1223 9000 1257
rect 9034 1223 9069 1257
rect 9103 1223 9138 1257
rect 9172 1223 9207 1257
rect 9241 1223 9276 1257
rect 9310 1223 9345 1257
rect 9379 1223 9414 1257
rect 9448 1223 9483 1257
rect 9517 1223 9552 1257
rect 9586 1223 9621 1257
rect 9655 1223 9690 1257
rect 9724 1223 9759 1257
rect 7022 1193 9759 1223
rect 6988 1189 9759 1193
rect 6988 1159 7068 1189
rect 7022 1155 7068 1159
rect 7102 1155 7137 1189
rect 7171 1155 7206 1189
rect 7240 1155 7275 1189
rect 7309 1155 7344 1189
rect 7378 1155 7413 1189
rect 7447 1155 7482 1189
rect 7516 1155 7551 1189
rect 7585 1155 7620 1189
rect 7654 1155 7689 1189
rect 7723 1155 7758 1189
rect 7792 1155 7827 1189
rect 7861 1155 7896 1189
rect 7930 1155 7965 1189
rect 7999 1155 8034 1189
rect 8068 1155 8103 1189
rect 8137 1155 8172 1189
rect 8206 1155 8241 1189
rect 8275 1155 8310 1189
rect 8344 1155 8379 1189
rect 8413 1155 8448 1189
rect 8482 1155 8517 1189
rect 8551 1155 8586 1189
rect 8620 1155 8655 1189
rect 8689 1155 8724 1189
rect 8758 1155 8793 1189
rect 8827 1155 8862 1189
rect 8896 1155 8931 1189
rect 8965 1155 9000 1189
rect 9034 1155 9069 1189
rect 9103 1155 9138 1189
rect 9172 1155 9207 1189
rect 9241 1155 9276 1189
rect 9310 1155 9345 1189
rect 9379 1155 9414 1189
rect 9448 1155 9483 1189
rect 9517 1155 9552 1189
rect 9586 1155 9621 1189
rect 9655 1155 9690 1189
rect 9724 1155 9759 1189
rect 7022 1125 9759 1155
rect 6988 1121 9759 1125
rect 6988 1091 7068 1121
rect 7022 1087 7068 1091
rect 7102 1087 7137 1121
rect 7171 1087 7206 1121
rect 7240 1087 7275 1121
rect 7309 1087 7344 1121
rect 7378 1087 7413 1121
rect 7447 1087 7482 1121
rect 7516 1087 7551 1121
rect 7585 1087 7620 1121
rect 7654 1087 7689 1121
rect 7723 1087 7758 1121
rect 7792 1087 7827 1121
rect 7861 1087 7896 1121
rect 7930 1087 7965 1121
rect 7999 1087 8034 1121
rect 8068 1087 8103 1121
rect 8137 1087 8172 1121
rect 8206 1087 8241 1121
rect 8275 1087 8310 1121
rect 8344 1087 8379 1121
rect 8413 1087 8448 1121
rect 8482 1087 8517 1121
rect 8551 1087 8586 1121
rect 8620 1087 8655 1121
rect 8689 1087 8724 1121
rect 8758 1087 8793 1121
rect 8827 1087 8862 1121
rect 8896 1087 8931 1121
rect 8965 1087 9000 1121
rect 9034 1087 9069 1121
rect 9103 1087 9138 1121
rect 9172 1087 9207 1121
rect 9241 1087 9276 1121
rect 9310 1087 9345 1121
rect 9379 1087 9414 1121
rect 9448 1087 9483 1121
rect 9517 1087 9552 1121
rect 9586 1087 9621 1121
rect 9655 1087 9690 1121
rect 9724 1087 9759 1121
rect 7022 1057 9759 1087
rect 6988 1053 9759 1057
rect 6988 1023 7068 1053
rect 7022 1019 7068 1023
rect 7102 1019 7137 1053
rect 7171 1019 7206 1053
rect 7240 1019 7275 1053
rect 7309 1019 7344 1053
rect 7378 1019 7413 1053
rect 7447 1019 7482 1053
rect 7516 1019 7551 1053
rect 7585 1019 7620 1053
rect 7654 1019 7689 1053
rect 7723 1019 7758 1053
rect 7792 1019 7827 1053
rect 7861 1019 7896 1053
rect 7930 1019 7965 1053
rect 7999 1019 8034 1053
rect 8068 1019 8103 1053
rect 8137 1019 8172 1053
rect 8206 1019 8241 1053
rect 8275 1019 8310 1053
rect 8344 1019 8379 1053
rect 8413 1019 8448 1053
rect 8482 1019 8517 1053
rect 8551 1019 8586 1053
rect 8620 1019 8655 1053
rect 8689 1019 8724 1053
rect 8758 1019 8793 1053
rect 8827 1019 8862 1053
rect 8896 1019 8931 1053
rect 8965 1019 9000 1053
rect 9034 1019 9069 1053
rect 9103 1019 9138 1053
rect 9172 1019 9207 1053
rect 9241 1019 9276 1053
rect 9310 1019 9345 1053
rect 9379 1019 9414 1053
rect 9448 1019 9483 1053
rect 9517 1019 9552 1053
rect 9586 1019 9621 1053
rect 9655 1019 9690 1053
rect 9724 1019 9759 1053
rect 14893 1244 15117 1257
rect 14893 1210 14932 1244
rect 14966 1210 15000 1244
rect 15034 1210 15068 1244
rect 15102 1210 15117 1244
rect 14893 1172 15117 1210
rect 14893 1138 14932 1172
rect 14966 1138 15000 1172
rect 15034 1138 15068 1172
rect 15102 1138 15117 1172
rect 14893 1100 15117 1138
rect 14893 1066 14932 1100
rect 14966 1066 15000 1100
rect 15034 1066 15068 1100
rect 15102 1066 15117 1100
rect 14893 1028 15117 1066
rect 14893 1019 14932 1028
rect 7022 994 14932 1019
rect 14966 994 15000 1028
rect 15034 994 15068 1028
rect 15102 994 15117 1028
rect 7022 989 15117 994
rect 6988 988 15117 989
rect 6988 955 7754 988
rect 7022 947 7754 955
rect 7022 921 7067 947
rect 6988 913 7067 921
rect 7101 913 7137 947
rect 7171 913 7207 947
rect 7241 913 7277 947
rect 7311 913 7347 947
rect 7381 913 7417 947
rect 7451 913 7487 947
rect 7521 913 7557 947
rect 7591 913 7627 947
rect 7661 913 7696 947
rect 7730 913 7754 947
rect 6988 887 7754 913
rect 7022 875 7754 887
rect 7022 853 7067 875
rect 6988 841 7067 853
rect 7101 841 7137 875
rect 7171 841 7207 875
rect 7241 841 7277 875
rect 7311 841 7347 875
rect 7381 841 7417 875
rect 7451 841 7487 875
rect 7521 841 7557 875
rect 7591 841 7627 875
rect 7661 841 7696 875
rect 7730 841 7754 875
rect 6988 819 7754 841
rect 7022 803 7754 819
rect 7022 785 7067 803
rect 6988 769 7067 785
rect 7101 769 7137 803
rect 7171 769 7207 803
rect 7241 769 7277 803
rect 7311 769 7347 803
rect 7381 769 7417 803
rect 7451 769 7487 803
rect 7521 769 7557 803
rect 7591 769 7627 803
rect 7661 769 7696 803
rect 7730 769 7754 803
rect 6988 751 7754 769
rect 7022 731 7754 751
rect 7022 717 7067 731
rect 6988 697 7067 717
rect 7101 697 7137 731
rect 7171 697 7207 731
rect 7241 697 7277 731
rect 7311 697 7347 731
rect 7381 697 7417 731
rect 7451 697 7487 731
rect 7521 697 7557 731
rect 7591 697 7627 731
rect 7661 697 7696 731
rect 7730 697 7754 731
rect 6988 683 7754 697
rect 7022 659 7754 683
rect 7022 649 7067 659
rect 6988 625 7067 649
rect 7101 625 7137 659
rect 7171 625 7207 659
rect 7241 625 7277 659
rect 7311 625 7347 659
rect 7381 625 7417 659
rect 7451 625 7487 659
rect 7521 625 7557 659
rect 7591 625 7627 659
rect 7661 625 7696 659
rect 7730 625 7754 659
rect 6988 615 7754 625
rect 7022 587 7754 615
rect 7022 581 7067 587
rect 6988 553 7067 581
rect 7101 553 7137 587
rect 7171 553 7207 587
rect 7241 553 7277 587
rect 7311 553 7347 587
rect 7381 553 7417 587
rect 7451 553 7487 587
rect 7521 553 7557 587
rect 7591 553 7627 587
rect 7661 553 7696 587
rect 7730 553 7754 587
rect 6988 547 7754 553
rect 7022 515 7754 547
rect 7022 513 7067 515
rect 6988 481 7067 513
rect 7101 481 7137 515
rect 7171 481 7207 515
rect 7241 481 7277 515
rect 7311 481 7347 515
rect 7381 481 7417 515
rect 7451 481 7487 515
rect 7521 481 7557 515
rect 7591 481 7627 515
rect 7661 481 7696 515
rect 7730 481 7754 515
rect 6988 479 7754 481
rect 7022 445 7754 479
rect 6988 443 7754 445
rect 6988 411 7067 443
rect 7022 409 7067 411
rect 7101 409 7137 443
rect 7171 409 7207 443
rect 7241 409 7277 443
rect 7311 409 7347 443
rect 7381 409 7417 443
rect 7451 409 7487 443
rect 7521 409 7557 443
rect 7591 409 7627 443
rect 7661 409 7696 443
rect 7730 409 7754 443
rect 7022 377 7754 409
rect 6988 369 7754 377
rect 9687 956 15117 988
rect 9687 955 14932 956
rect 9687 947 11680 955
rect 9687 913 9711 947
rect 9745 913 9781 947
rect 9815 913 9851 947
rect 9885 913 9921 947
rect 9955 913 9991 947
rect 10025 913 10061 947
rect 10095 913 10131 947
rect 10165 913 10201 947
rect 10235 913 10271 947
rect 10305 913 10341 947
rect 10375 913 10411 947
rect 10445 913 10481 947
rect 10515 913 10551 947
rect 10585 913 10621 947
rect 10655 913 10691 947
rect 10725 913 10761 947
rect 10795 913 10831 947
rect 10865 913 10901 947
rect 10935 913 10971 947
rect 11005 913 11041 947
rect 11075 913 11111 947
rect 11145 913 11181 947
rect 11215 913 11251 947
rect 11285 913 11321 947
rect 11355 913 11391 947
rect 11425 913 11460 947
rect 11494 913 11529 947
rect 11563 913 11598 947
rect 11632 921 11680 947
rect 11714 921 11750 955
rect 11784 921 11820 955
rect 11854 921 11890 955
rect 11924 921 11960 955
rect 11994 921 12030 955
rect 12064 921 12099 955
rect 12133 921 12168 955
rect 12202 921 12237 955
rect 12271 921 12306 955
rect 12340 921 12375 955
rect 12409 921 12444 955
rect 12478 921 12513 955
rect 12547 921 12582 955
rect 12616 921 12651 955
rect 12685 921 12720 955
rect 12754 921 12789 955
rect 12823 921 12858 955
rect 12892 921 12927 955
rect 12961 921 12996 955
rect 13030 921 13065 955
rect 13099 921 13134 955
rect 13168 921 13203 955
rect 13237 921 13272 955
rect 13306 921 13341 955
rect 13375 921 13410 955
rect 13444 921 13479 955
rect 13513 921 13548 955
rect 13582 921 13617 955
rect 13651 921 13686 955
rect 13720 921 13755 955
rect 13789 921 13824 955
rect 13858 921 13893 955
rect 13927 921 13962 955
rect 13996 921 14031 955
rect 14065 921 14100 955
rect 14134 921 14169 955
rect 14203 921 14238 955
rect 14272 921 14307 955
rect 14341 921 14376 955
rect 14410 921 14445 955
rect 14479 921 14514 955
rect 14548 921 14583 955
rect 14617 921 14652 955
rect 14686 921 14721 955
rect 14755 921 14790 955
rect 14824 921 14859 955
rect 14893 922 14932 955
rect 14966 922 15000 956
rect 15034 922 15068 956
rect 15102 922 15117 956
rect 14893 921 15117 922
rect 11632 913 15117 921
rect 9687 884 15117 913
rect 9687 875 14932 884
rect 9687 841 9711 875
rect 9745 841 9781 875
rect 9815 841 9851 875
rect 9885 841 9921 875
rect 9955 841 9991 875
rect 10025 841 10061 875
rect 10095 841 10131 875
rect 10165 841 10201 875
rect 10235 841 10271 875
rect 10305 841 10341 875
rect 10375 841 10411 875
rect 10445 841 10481 875
rect 10515 841 10551 875
rect 10585 841 10621 875
rect 10655 841 10691 875
rect 10725 841 10761 875
rect 10795 841 10831 875
rect 10865 841 10901 875
rect 10935 841 10971 875
rect 11005 841 11041 875
rect 11075 841 11111 875
rect 11145 841 11181 875
rect 11215 841 11251 875
rect 11285 841 11321 875
rect 11355 841 11391 875
rect 11425 841 11460 875
rect 11494 841 11529 875
rect 11563 841 11598 875
rect 11632 841 11680 875
rect 11714 841 11750 875
rect 11784 841 11820 875
rect 11854 841 11890 875
rect 11924 841 11960 875
rect 11994 841 12030 875
rect 12064 841 12099 875
rect 12133 841 12168 875
rect 12202 841 12237 875
rect 12271 841 12306 875
rect 12340 841 12375 875
rect 12409 841 12444 875
rect 12478 841 12513 875
rect 12547 841 12582 875
rect 12616 841 12651 875
rect 12685 841 12720 875
rect 12754 841 12789 875
rect 12823 841 12858 875
rect 12892 841 12927 875
rect 12961 841 12996 875
rect 13030 841 13065 875
rect 13099 841 13134 875
rect 13168 841 13203 875
rect 13237 841 13272 875
rect 13306 841 13341 875
rect 13375 841 13410 875
rect 13444 841 13479 875
rect 13513 841 13548 875
rect 13582 841 13617 875
rect 13651 841 13686 875
rect 13720 841 13755 875
rect 13789 841 13824 875
rect 13858 841 13893 875
rect 13927 841 13962 875
rect 13996 841 14031 875
rect 14065 841 14100 875
rect 14134 841 14169 875
rect 14203 841 14238 875
rect 14272 841 14307 875
rect 14341 841 14376 875
rect 14410 841 14445 875
rect 14479 841 14514 875
rect 14548 841 14583 875
rect 14617 841 14652 875
rect 14686 841 14721 875
rect 14755 841 14790 875
rect 14824 841 14859 875
rect 14893 850 14932 875
rect 14966 850 15000 884
rect 15034 850 15068 884
rect 15102 850 15117 884
rect 14893 841 15117 850
rect 9687 812 15117 841
rect 9687 803 14932 812
rect 9687 769 9711 803
rect 9745 769 9781 803
rect 9815 769 9851 803
rect 9885 769 9921 803
rect 9955 769 9991 803
rect 10025 769 10061 803
rect 10095 769 10131 803
rect 10165 769 10201 803
rect 10235 769 10271 803
rect 10305 769 10341 803
rect 10375 769 10411 803
rect 10445 769 10481 803
rect 10515 769 10551 803
rect 10585 769 10621 803
rect 10655 769 10691 803
rect 10725 769 10761 803
rect 10795 769 10831 803
rect 10865 769 10901 803
rect 10935 769 10971 803
rect 11005 769 11041 803
rect 11075 769 11111 803
rect 11145 769 11181 803
rect 11215 769 11251 803
rect 11285 769 11321 803
rect 11355 769 11391 803
rect 11425 769 11460 803
rect 11494 769 11529 803
rect 11563 769 11598 803
rect 11632 795 14932 803
rect 11632 769 11680 795
rect 9687 761 11680 769
rect 11714 761 11750 795
rect 11784 761 11820 795
rect 11854 761 11890 795
rect 11924 761 11960 795
rect 11994 761 12030 795
rect 12064 761 12099 795
rect 12133 761 12168 795
rect 12202 761 12237 795
rect 12271 761 12306 795
rect 12340 761 12375 795
rect 12409 761 12444 795
rect 12478 761 12513 795
rect 12547 761 12582 795
rect 12616 761 12651 795
rect 12685 761 12720 795
rect 12754 761 12789 795
rect 12823 761 12858 795
rect 12892 761 12927 795
rect 12961 761 12996 795
rect 13030 761 13065 795
rect 13099 761 13134 795
rect 13168 761 13203 795
rect 13237 761 13272 795
rect 13306 761 13341 795
rect 13375 761 13410 795
rect 13444 761 13479 795
rect 13513 761 13548 795
rect 13582 761 13617 795
rect 13651 761 13686 795
rect 13720 761 13755 795
rect 13789 761 13824 795
rect 13858 761 13893 795
rect 13927 761 13962 795
rect 13996 761 14031 795
rect 14065 761 14100 795
rect 14134 761 14169 795
rect 14203 761 14238 795
rect 14272 761 14307 795
rect 14341 761 14376 795
rect 14410 761 14445 795
rect 14479 761 14514 795
rect 14548 761 14583 795
rect 14617 761 14652 795
rect 14686 761 14721 795
rect 14755 761 14790 795
rect 14824 761 14859 795
rect 14893 778 14932 795
rect 14966 778 15000 812
rect 15034 778 15068 812
rect 15102 778 15117 812
rect 14893 761 15117 778
rect 9687 740 15117 761
rect 9687 731 14932 740
rect 9687 697 9711 731
rect 9745 697 9781 731
rect 9815 697 9851 731
rect 9885 697 9921 731
rect 9955 697 9991 731
rect 10025 697 10061 731
rect 10095 697 10131 731
rect 10165 697 10201 731
rect 10235 697 10271 731
rect 10305 697 10341 731
rect 10375 697 10411 731
rect 10445 697 10481 731
rect 10515 697 10551 731
rect 10585 697 10621 731
rect 10655 697 10691 731
rect 10725 697 10761 731
rect 10795 697 10831 731
rect 10865 697 10901 731
rect 10935 697 10971 731
rect 11005 697 11041 731
rect 11075 697 11111 731
rect 11145 697 11181 731
rect 11215 697 11251 731
rect 11285 697 11321 731
rect 11355 697 11391 731
rect 11425 697 11460 731
rect 11494 697 11529 731
rect 11563 697 11598 731
rect 11632 728 14932 731
rect 11632 697 11656 728
rect 9687 659 11656 697
rect 9687 625 9711 659
rect 9745 625 9781 659
rect 9815 625 9851 659
rect 9885 625 9921 659
rect 9955 625 9991 659
rect 10025 625 10061 659
rect 10095 625 10131 659
rect 10165 625 10201 659
rect 10235 625 10271 659
rect 10305 625 10341 659
rect 10375 625 10411 659
rect 10445 625 10481 659
rect 10515 625 10551 659
rect 10585 625 10621 659
rect 10655 625 10691 659
rect 10725 625 10761 659
rect 10795 625 10831 659
rect 10865 625 10901 659
rect 10935 625 10971 659
rect 11005 625 11041 659
rect 11075 625 11111 659
rect 11145 625 11181 659
rect 11215 625 11251 659
rect 11285 625 11321 659
rect 11355 625 11391 659
rect 11425 625 11460 659
rect 11494 625 11529 659
rect 11563 625 11598 659
rect 11632 625 11656 659
rect 9687 587 11656 625
rect 9687 553 9711 587
rect 9745 553 9781 587
rect 9815 553 9851 587
rect 9885 553 9921 587
rect 9955 553 9991 587
rect 10025 553 10061 587
rect 10095 553 10131 587
rect 10165 553 10201 587
rect 10235 553 10271 587
rect 10305 553 10341 587
rect 10375 553 10411 587
rect 10445 553 10481 587
rect 10515 553 10551 587
rect 10585 553 10621 587
rect 10655 553 10691 587
rect 10725 553 10761 587
rect 10795 553 10831 587
rect 10865 553 10901 587
rect 10935 553 10971 587
rect 11005 553 11041 587
rect 11075 553 11111 587
rect 11145 553 11181 587
rect 11215 553 11251 587
rect 11285 553 11321 587
rect 11355 553 11391 587
rect 11425 553 11460 587
rect 11494 553 11529 587
rect 11563 553 11598 587
rect 11632 553 11656 587
rect 9687 515 11656 553
rect 9687 481 9711 515
rect 9745 481 9781 515
rect 9815 481 9851 515
rect 9885 481 9921 515
rect 9955 481 9991 515
rect 10025 481 10061 515
rect 10095 481 10131 515
rect 10165 481 10201 515
rect 10235 481 10271 515
rect 10305 481 10341 515
rect 10375 481 10411 515
rect 10445 481 10481 515
rect 10515 481 10551 515
rect 10585 481 10621 515
rect 10655 481 10691 515
rect 10725 481 10761 515
rect 10795 481 10831 515
rect 10865 481 10901 515
rect 10935 481 10971 515
rect 11005 481 11041 515
rect 11075 481 11111 515
rect 11145 481 11181 515
rect 11215 481 11251 515
rect 11285 481 11321 515
rect 11355 481 11391 515
rect 11425 481 11460 515
rect 11494 481 11529 515
rect 11563 481 11598 515
rect 11632 481 11656 515
rect 9687 443 11656 481
rect 9687 409 9711 443
rect 9745 409 9781 443
rect 9815 409 9851 443
rect 9885 409 9921 443
rect 9955 409 9991 443
rect 10025 409 10061 443
rect 10095 409 10131 443
rect 10165 409 10201 443
rect 10235 409 10271 443
rect 10305 409 10341 443
rect 10375 409 10411 443
rect 10445 409 10481 443
rect 10515 409 10551 443
rect 10585 409 10621 443
rect 10655 409 10691 443
rect 10725 409 10761 443
rect 10795 409 10831 443
rect 10865 409 10901 443
rect 10935 409 10971 443
rect 11005 409 11041 443
rect 11075 409 11111 443
rect 11145 409 11181 443
rect 11215 409 11251 443
rect 11285 409 11321 443
rect 11355 409 11391 443
rect 11425 409 11460 443
rect 11494 409 11529 443
rect 11563 409 11598 443
rect 11632 409 11656 443
rect 9687 369 11656 409
rect 14465 706 14932 728
rect 14966 706 15000 740
rect 15034 706 15068 740
rect 15102 706 15117 740
rect 14465 695 15117 706
rect 14499 661 14543 695
rect 14577 661 14621 695
rect 14655 661 14698 695
rect 14732 661 14775 695
rect 14809 661 14852 695
rect 14886 668 15117 695
rect 14886 661 14932 668
rect 14465 634 14932 661
rect 14966 634 15000 668
rect 15034 634 15068 668
rect 15102 634 15117 668
rect 14465 609 15117 634
rect 14499 575 14543 609
rect 14577 575 14621 609
rect 14655 575 14698 609
rect 14732 575 14775 609
rect 14809 575 14852 609
rect 14886 596 15117 609
rect 14886 575 14932 596
rect 14465 562 14932 575
rect 14966 562 15000 596
rect 15034 562 15068 596
rect 15102 562 15117 596
rect 14465 524 15117 562
rect 14465 523 14932 524
rect 14499 489 14543 523
rect 14577 489 14621 523
rect 14655 489 14698 523
rect 14732 489 14775 523
rect 14809 489 14852 523
rect 14886 490 14932 523
rect 14966 490 15000 524
rect 15034 490 15068 524
rect 15102 490 15117 524
rect 14886 489 15117 490
rect 14465 452 15117 489
rect 14465 437 14932 452
rect 14499 403 14543 437
rect 14577 403 14621 437
rect 14655 403 14698 437
rect 14732 403 14775 437
rect 14809 403 14852 437
rect 14886 418 14932 437
rect 14966 418 15000 452
rect 15034 418 15068 452
rect 15102 418 15117 452
rect 14886 403 15117 418
rect 14465 380 15117 403
rect 14465 369 14932 380
rect 6988 367 14932 369
rect 6988 343 7056 367
rect 7022 333 7056 343
rect 7090 333 7125 367
rect 7159 333 7194 367
rect 7228 333 7263 367
rect 7297 333 7332 367
rect 7366 333 7401 367
rect 7435 333 7470 367
rect 7504 333 7539 367
rect 7573 333 7608 367
rect 7642 333 7677 367
rect 7711 333 7746 367
rect 7780 333 7815 367
rect 7849 333 7884 367
rect 7918 333 7953 367
rect 7987 333 8022 367
rect 8056 333 8091 367
rect 8125 333 8160 367
rect 8194 333 8229 367
rect 8263 333 8298 367
rect 8332 333 8367 367
rect 8401 333 8436 367
rect 8470 333 8505 367
rect 8539 333 8574 367
rect 8608 333 8643 367
rect 8677 333 8712 367
rect 8746 333 8781 367
rect 8815 333 8850 367
rect 8884 333 8919 367
rect 8953 333 8988 367
rect 9022 333 9057 367
rect 9091 333 9126 367
rect 9160 333 9195 367
rect 9229 333 9264 367
rect 9298 333 9333 367
rect 9367 333 9402 367
rect 9436 333 9471 367
rect 9505 333 9540 367
rect 9574 333 9609 367
rect 9643 333 9678 367
rect 9712 333 9747 367
rect 9781 333 9816 367
rect 9850 333 9885 367
rect 9919 333 9954 367
rect 9988 333 10023 367
rect 10057 333 10092 367
rect 10126 333 10161 367
rect 10195 333 10230 367
rect 10264 333 10299 367
rect 10333 333 10368 367
rect 10402 333 10437 367
rect 10471 333 10506 367
rect 10540 333 10575 367
rect 10609 333 10643 367
rect 10677 333 10711 367
rect 10745 333 10779 367
rect 10813 333 10847 367
rect 10881 333 10915 367
rect 10949 333 10983 367
rect 11017 333 11051 367
rect 11085 333 11119 367
rect 11153 333 11187 367
rect 11221 333 11255 367
rect 11289 333 11323 367
rect 11357 333 11391 367
rect 11425 333 11459 367
rect 11493 333 11527 367
rect 11561 333 11595 367
rect 11629 333 11663 367
rect 11697 333 11731 367
rect 11765 333 11799 367
rect 11833 333 11867 367
rect 11901 333 11935 367
rect 11969 333 12003 367
rect 12037 333 12071 367
rect 12105 333 12139 367
rect 12173 333 12207 367
rect 12241 333 12275 367
rect 12309 333 12343 367
rect 12377 333 12411 367
rect 12445 333 12479 367
rect 12513 333 12547 367
rect 12581 333 12615 367
rect 12649 333 12683 367
rect 12717 333 12751 367
rect 12785 333 12819 367
rect 12853 333 12887 367
rect 12921 333 12955 367
rect 12989 333 13023 367
rect 13057 333 13091 367
rect 13125 333 13159 367
rect 13193 333 13227 367
rect 13261 333 13295 367
rect 13329 333 13363 367
rect 13397 333 13431 367
rect 13465 333 13499 367
rect 13533 333 13567 367
rect 13601 333 13635 367
rect 13669 333 13703 367
rect 13737 333 13771 367
rect 13805 333 13839 367
rect 13873 333 13907 367
rect 13941 333 13975 367
rect 14009 333 14043 367
rect 14077 333 14111 367
rect 14145 333 14179 367
rect 14213 333 14247 367
rect 14281 333 14315 367
rect 14349 333 14383 367
rect 14417 333 14451 367
rect 14485 333 14519 367
rect 14553 333 14587 367
rect 14621 333 14655 367
rect 14689 333 14723 367
rect 14757 333 14791 367
rect 14825 333 14859 367
rect 14893 346 14932 367
rect 14966 346 15000 380
rect 15034 346 15068 380
rect 15102 346 15117 380
rect 14893 333 15117 346
rect 7022 309 15117 333
rect 6988 308 15117 309
rect 6988 289 14932 308
rect 6988 275 7056 289
rect 7022 255 7056 275
rect 7090 255 7125 289
rect 7159 255 7194 289
rect 7228 255 7263 289
rect 7297 255 7332 289
rect 7366 255 7401 289
rect 7435 255 7470 289
rect 7504 255 7539 289
rect 7573 255 7608 289
rect 7642 255 7677 289
rect 7711 255 7746 289
rect 7780 255 7815 289
rect 7849 255 7884 289
rect 7918 255 7953 289
rect 7987 255 8022 289
rect 8056 255 8091 289
rect 8125 255 8160 289
rect 8194 255 8229 289
rect 8263 255 8298 289
rect 8332 255 8367 289
rect 8401 255 8436 289
rect 8470 255 8505 289
rect 8539 255 8574 289
rect 8608 255 8643 289
rect 8677 255 8712 289
rect 8746 255 8781 289
rect 8815 255 8850 289
rect 8884 255 8919 289
rect 8953 255 8988 289
rect 9022 255 9057 289
rect 9091 255 9126 289
rect 9160 255 9195 289
rect 9229 255 9264 289
rect 9298 255 9333 289
rect 9367 255 9402 289
rect 9436 255 9471 289
rect 9505 255 9540 289
rect 9574 255 9609 289
rect 9643 255 9678 289
rect 9712 255 9747 289
rect 9781 255 9816 289
rect 9850 255 9885 289
rect 9919 255 9954 289
rect 9988 255 10023 289
rect 10057 255 10092 289
rect 10126 255 10161 289
rect 10195 255 10230 289
rect 10264 255 10299 289
rect 10333 255 10368 289
rect 10402 255 10437 289
rect 10471 255 10506 289
rect 10540 255 10575 289
rect 10609 255 10643 289
rect 10677 255 10711 289
rect 10745 255 10779 289
rect 10813 255 10847 289
rect 10881 255 10915 289
rect 10949 255 10983 289
rect 11017 255 11051 289
rect 11085 255 11119 289
rect 11153 255 11187 289
rect 11221 255 11255 289
rect 11289 255 11323 289
rect 11357 255 11391 289
rect 11425 255 11459 289
rect 11493 255 11527 289
rect 11561 255 11595 289
rect 11629 255 11663 289
rect 11697 255 11731 289
rect 11765 255 11799 289
rect 11833 255 11867 289
rect 11901 255 11935 289
rect 11969 255 12003 289
rect 12037 255 12071 289
rect 12105 255 12139 289
rect 12173 255 12207 289
rect 12241 255 12275 289
rect 12309 255 12343 289
rect 12377 255 12411 289
rect 12445 255 12479 289
rect 12513 255 12547 289
rect 12581 255 12615 289
rect 12649 255 12683 289
rect 12717 255 12751 289
rect 12785 255 12819 289
rect 12853 255 12887 289
rect 12921 255 12955 289
rect 12989 255 13023 289
rect 13057 255 13091 289
rect 13125 255 13159 289
rect 13193 255 13227 289
rect 13261 255 13295 289
rect 13329 255 13363 289
rect 13397 255 13431 289
rect 13465 255 13499 289
rect 13533 255 13567 289
rect 13601 255 13635 289
rect 13669 255 13703 289
rect 13737 255 13771 289
rect 13805 255 13839 289
rect 13873 255 13907 289
rect 13941 255 13975 289
rect 14009 255 14043 289
rect 14077 255 14111 289
rect 14145 255 14179 289
rect 14213 255 14247 289
rect 14281 255 14315 289
rect 14349 255 14383 289
rect 14417 255 14451 289
rect 14485 255 14519 289
rect 14553 255 14587 289
rect 14621 255 14655 289
rect 14689 255 14723 289
rect 14757 255 14791 289
rect 14825 255 14859 289
rect 14893 274 14932 289
rect 14966 274 15000 308
rect 15034 274 15068 308
rect 15102 274 15117 308
rect 14893 255 15117 274
rect 7022 241 15117 255
rect 6988 236 15117 241
rect 6988 211 14932 236
rect 6988 207 7056 211
rect 7022 177 7056 207
rect 7090 177 7125 211
rect 7159 177 7194 211
rect 7228 177 7263 211
rect 7297 177 7332 211
rect 7366 177 7401 211
rect 7435 177 7470 211
rect 7504 177 7539 211
rect 7573 177 7608 211
rect 7642 177 7677 211
rect 7711 177 7746 211
rect 7780 177 7815 211
rect 7849 177 7884 211
rect 7918 177 7953 211
rect 7987 177 8022 211
rect 8056 177 8091 211
rect 8125 177 8160 211
rect 8194 177 8229 211
rect 8263 177 8298 211
rect 8332 177 8367 211
rect 8401 177 8436 211
rect 8470 177 8505 211
rect 8539 177 8574 211
rect 8608 177 8643 211
rect 8677 177 8712 211
rect 8746 177 8781 211
rect 8815 177 8850 211
rect 8884 177 8919 211
rect 8953 177 8988 211
rect 9022 177 9057 211
rect 9091 177 9126 211
rect 9160 177 9195 211
rect 9229 177 9264 211
rect 9298 177 9333 211
rect 9367 177 9402 211
rect 9436 177 9471 211
rect 9505 177 9540 211
rect 9574 177 9609 211
rect 9643 177 9678 211
rect 9712 177 9747 211
rect 9781 177 9816 211
rect 9850 177 9885 211
rect 9919 177 9954 211
rect 9988 177 10023 211
rect 10057 177 10092 211
rect 10126 177 10161 211
rect 10195 177 10230 211
rect 10264 177 10299 211
rect 10333 177 10368 211
rect 10402 177 10437 211
rect 10471 177 10506 211
rect 10540 177 10575 211
rect 10609 177 10643 211
rect 10677 177 10711 211
rect 10745 177 10779 211
rect 10813 177 10847 211
rect 10881 177 10915 211
rect 10949 177 10983 211
rect 11017 177 11051 211
rect 11085 177 11119 211
rect 11153 177 11187 211
rect 11221 177 11255 211
rect 11289 177 11323 211
rect 11357 177 11391 211
rect 11425 177 11459 211
rect 11493 177 11527 211
rect 11561 177 11595 211
rect 11629 177 11663 211
rect 11697 177 11731 211
rect 11765 177 11799 211
rect 11833 177 11867 211
rect 11901 177 11935 211
rect 11969 177 12003 211
rect 12037 177 12071 211
rect 12105 177 12139 211
rect 12173 177 12207 211
rect 12241 177 12275 211
rect 12309 177 12343 211
rect 12377 177 12411 211
rect 12445 177 12479 211
rect 12513 177 12547 211
rect 12581 177 12615 211
rect 12649 177 12683 211
rect 12717 177 12751 211
rect 12785 177 12819 211
rect 12853 177 12887 211
rect 12921 177 12955 211
rect 12989 177 13023 211
rect 13057 177 13091 211
rect 13125 177 13159 211
rect 13193 177 13227 211
rect 13261 177 13295 211
rect 13329 177 13363 211
rect 13397 177 13431 211
rect 13465 177 13499 211
rect 13533 177 13567 211
rect 13601 177 13635 211
rect 13669 177 13703 211
rect 13737 177 13771 211
rect 13805 177 13839 211
rect 13873 177 13907 211
rect 13941 177 13975 211
rect 14009 177 14043 211
rect 14077 177 14111 211
rect 14145 177 14179 211
rect 14213 177 14247 211
rect 14281 177 14315 211
rect 14349 177 14383 211
rect 14417 177 14451 211
rect 14485 177 14519 211
rect 14553 177 14587 211
rect 14621 177 14655 211
rect 14689 177 14723 211
rect 14757 177 14791 211
rect 14825 177 14859 211
rect 14893 202 14932 211
rect 14966 202 15000 236
rect 15034 202 15068 236
rect 15102 202 15117 236
rect 14893 177 15117 202
rect 7022 173 15117 177
rect 6988 164 15117 173
rect 6988 139 14932 164
rect 7022 133 14932 139
rect 7022 105 7056 133
rect 6988 99 7056 105
rect 7090 99 7125 133
rect 7159 99 7194 133
rect 7228 99 7263 133
rect 7297 99 7332 133
rect 7366 99 7401 133
rect 7435 99 7470 133
rect 7504 99 7539 133
rect 7573 99 7608 133
rect 7642 99 7677 133
rect 7711 99 7746 133
rect 7780 99 7815 133
rect 7849 99 7884 133
rect 7918 99 7953 133
rect 7987 99 8022 133
rect 8056 99 8091 133
rect 8125 99 8160 133
rect 8194 99 8229 133
rect 8263 99 8298 133
rect 8332 99 8367 133
rect 8401 99 8436 133
rect 8470 99 8505 133
rect 8539 99 8574 133
rect 8608 99 8643 133
rect 8677 99 8712 133
rect 8746 99 8781 133
rect 8815 99 8850 133
rect 8884 99 8919 133
rect 8953 99 8988 133
rect 9022 99 9057 133
rect 9091 99 9126 133
rect 9160 99 9195 133
rect 9229 99 9264 133
rect 9298 99 9333 133
rect 9367 99 9402 133
rect 9436 99 9471 133
rect 9505 99 9540 133
rect 9574 99 9609 133
rect 9643 99 9678 133
rect 9712 99 9747 133
rect 9781 99 9816 133
rect 9850 99 9885 133
rect 9919 99 9954 133
rect 9988 99 10023 133
rect 10057 99 10092 133
rect 10126 99 10161 133
rect 10195 99 10230 133
rect 10264 99 10299 133
rect 10333 99 10368 133
rect 10402 99 10437 133
rect 10471 99 10506 133
rect 10540 99 10575 133
rect 10609 99 10643 133
rect 10677 99 10711 133
rect 10745 99 10779 133
rect 10813 99 10847 133
rect 10881 99 10915 133
rect 10949 99 10983 133
rect 11017 99 11051 133
rect 11085 99 11119 133
rect 11153 99 11187 133
rect 11221 99 11255 133
rect 11289 99 11323 133
rect 11357 99 11391 133
rect 11425 99 11459 133
rect 11493 99 11527 133
rect 11561 99 11595 133
rect 11629 99 11663 133
rect 11697 99 11731 133
rect 11765 99 11799 133
rect 11833 99 11867 133
rect 11901 99 11935 133
rect 11969 99 12003 133
rect 12037 99 12071 133
rect 12105 99 12139 133
rect 12173 99 12207 133
rect 12241 99 12275 133
rect 12309 99 12343 133
rect 12377 99 12411 133
rect 12445 99 12479 133
rect 12513 99 12547 133
rect 12581 99 12615 133
rect 12649 99 12683 133
rect 12717 99 12751 133
rect 12785 99 12819 133
rect 12853 99 12887 133
rect 12921 99 12955 133
rect 12989 99 13023 133
rect 13057 99 13091 133
rect 13125 99 13159 133
rect 13193 99 13227 133
rect 13261 99 13295 133
rect 13329 99 13363 133
rect 13397 99 13431 133
rect 13465 99 13499 133
rect 13533 99 13567 133
rect 13601 99 13635 133
rect 13669 99 13703 133
rect 13737 99 13771 133
rect 13805 99 13839 133
rect 13873 99 13907 133
rect 13941 99 13975 133
rect 14009 99 14043 133
rect 14077 99 14111 133
rect 14145 99 14179 133
rect 14213 99 14247 133
rect 14281 99 14315 133
rect 14349 99 14383 133
rect 14417 99 14451 133
rect 14485 99 14519 133
rect 14553 99 14587 133
rect 14621 99 14655 133
rect 14689 99 14723 133
rect 14757 99 14791 133
rect 14825 99 14859 133
rect 14893 130 14932 133
rect 14966 130 15000 164
rect 15034 130 15068 164
rect 15102 130 15117 164
rect 14893 99 15117 130
rect 6988 91 15117 99
rect 6988 57 14932 91
rect 14966 57 15000 91
rect 15034 57 15068 91
rect 15102 57 15117 91
rect 6988 55 15117 57
rect 6988 23 7056 55
rect 3545 -11 3632 23
rect 3666 -11 3700 23
rect 3734 -11 3768 23
rect 3802 -11 3836 23
rect 3870 -11 3904 23
rect 3938 -11 3972 23
rect 4006 -11 4040 23
rect 4074 -11 4108 23
rect 4142 -11 4176 23
rect 4210 -11 4244 23
rect 4278 -11 4312 23
rect 4346 -11 4380 23
rect 4414 -11 4448 23
rect 4482 -11 4516 23
rect 4550 -11 4584 23
rect 4618 -11 4652 23
rect 4686 -11 4720 23
rect 4754 -11 4788 23
rect 4822 -11 4856 23
rect 4890 -11 4924 23
rect 4958 -11 4992 23
rect 5026 -11 5060 23
rect 5094 -11 5128 23
rect 5162 -11 5196 23
rect 5230 -11 5264 23
rect 5298 -11 5332 23
rect 5366 -11 5400 23
rect 5434 -11 5468 23
rect 5502 -11 5536 23
rect 5570 -11 5604 23
rect 5638 -11 5672 23
rect 5706 -11 5740 23
rect 5774 -11 5808 23
rect 5842 -11 5876 23
rect 5910 -11 5944 23
rect 5978 -11 6012 23
rect 6046 -11 6080 23
rect 6114 -11 6148 23
rect 6182 -11 6216 23
rect 6250 -11 6284 23
rect 6318 -11 6352 23
rect 6386 -11 6420 23
rect 6454 -11 6488 23
rect 6522 -11 6556 23
rect 6590 -11 6624 23
rect 6658 -11 6692 23
rect 6726 -11 6760 23
rect 6794 -11 6828 23
rect 6862 -11 6896 23
rect 6930 -11 6964 23
rect 6998 21 7056 23
rect 7090 21 7125 55
rect 7159 21 7194 55
rect 7228 21 7263 55
rect 7297 21 7332 55
rect 7366 21 7401 55
rect 7435 21 7470 55
rect 7504 21 7539 55
rect 7573 21 7608 55
rect 7642 21 7677 55
rect 7711 21 7746 55
rect 7780 21 7815 55
rect 7849 21 7884 55
rect 7918 21 7953 55
rect 7987 21 8022 55
rect 8056 21 8091 55
rect 8125 21 8160 55
rect 8194 21 8229 55
rect 8263 21 8298 55
rect 8332 21 8367 55
rect 8401 21 8436 55
rect 8470 21 8505 55
rect 8539 21 8574 55
rect 8608 21 8643 55
rect 8677 21 8712 55
rect 8746 21 8781 55
rect 8815 21 8850 55
rect 8884 21 8919 55
rect 8953 21 8988 55
rect 9022 21 9057 55
rect 9091 21 9126 55
rect 9160 21 9195 55
rect 9229 21 9264 55
rect 9298 21 9333 55
rect 9367 21 9402 55
rect 9436 21 9471 55
rect 9505 21 9540 55
rect 9574 21 9609 55
rect 9643 21 9678 55
rect 9712 21 9747 55
rect 9781 21 9816 55
rect 9850 21 9885 55
rect 9919 21 9954 55
rect 9988 21 10023 55
rect 10057 21 10092 55
rect 10126 21 10161 55
rect 10195 21 10230 55
rect 10264 21 10299 55
rect 10333 21 10368 55
rect 10402 21 10437 55
rect 10471 21 10506 55
rect 10540 21 10575 55
rect 10609 21 10643 55
rect 10677 21 10711 55
rect 10745 21 10779 55
rect 10813 21 10847 55
rect 10881 21 10915 55
rect 10949 21 10983 55
rect 11017 21 11051 55
rect 11085 21 11119 55
rect 11153 21 11187 55
rect 11221 21 11255 55
rect 11289 21 11323 55
rect 11357 21 11391 55
rect 11425 21 11459 55
rect 11493 21 11527 55
rect 11561 21 11595 55
rect 11629 21 11663 55
rect 11697 21 11731 55
rect 11765 21 11799 55
rect 11833 21 11867 55
rect 11901 21 11935 55
rect 11969 21 12003 55
rect 12037 21 12071 55
rect 12105 21 12139 55
rect 12173 21 12207 55
rect 12241 21 12275 55
rect 12309 21 12343 55
rect 12377 21 12411 55
rect 12445 21 12479 55
rect 12513 21 12547 55
rect 12581 21 12615 55
rect 12649 21 12683 55
rect 12717 21 12751 55
rect 12785 21 12819 55
rect 12853 21 12887 55
rect 12921 21 12955 55
rect 12989 21 13023 55
rect 13057 21 13091 55
rect 13125 21 13159 55
rect 13193 21 13227 55
rect 13261 21 13295 55
rect 13329 21 13363 55
rect 13397 21 13431 55
rect 13465 21 13499 55
rect 13533 21 13567 55
rect 13601 21 13635 55
rect 13669 21 13703 55
rect 13737 21 13771 55
rect 13805 21 13839 55
rect 13873 21 13907 55
rect 13941 21 13975 55
rect 14009 21 14043 55
rect 14077 21 14111 55
rect 14145 21 14179 55
rect 14213 21 14247 55
rect 14281 21 14315 55
rect 14349 21 14383 55
rect 14417 21 14451 55
rect 14485 21 14519 55
rect 14553 21 14587 55
rect 14621 21 14655 55
rect 14689 21 14723 55
rect 14757 21 14791 55
rect 14825 21 14859 55
rect 14893 21 15117 55
rect 6998 19 15117 21
rect 6998 -11 7022 19
<< mvnsubdiff >>
rect 67 16503 15106 16527
rect 67 16493 14420 16503
rect 67 16459 68 16493
rect 102 16459 139 16493
rect 173 16459 210 16493
rect 244 16459 281 16493
rect 315 16459 352 16493
rect 386 16459 444 16493
rect 478 16459 513 16493
rect 547 16459 582 16493
rect 616 16459 651 16493
rect 685 16459 720 16493
rect 754 16459 789 16493
rect 823 16459 858 16493
rect 892 16459 927 16493
rect 961 16459 996 16493
rect 1030 16459 1065 16493
rect 1099 16459 1134 16493
rect 1168 16459 1203 16493
rect 1237 16459 1272 16493
rect 1306 16459 1341 16493
rect 1375 16459 1410 16493
rect 1444 16459 1479 16493
rect 1513 16459 1548 16493
rect 1582 16459 1617 16493
rect 1651 16459 1686 16493
rect 1720 16459 1755 16493
rect 1789 16459 1824 16493
rect 1858 16459 1893 16493
rect 1927 16459 1962 16493
rect 1996 16459 2031 16493
rect 2065 16459 2100 16493
rect 2134 16459 2169 16493
rect 2203 16459 2238 16493
rect 2272 16459 2307 16493
rect 2341 16459 2376 16493
rect 2410 16459 2445 16493
rect 2479 16459 2514 16493
rect 2548 16459 2583 16493
rect 2617 16459 2652 16493
rect 2686 16459 2721 16493
rect 2755 16459 2790 16493
rect 2824 16459 2859 16493
rect 2893 16459 2928 16493
rect 2962 16459 2996 16493
rect 3030 16459 3064 16493
rect 3098 16459 3132 16493
rect 3166 16459 3200 16493
rect 3234 16459 3268 16493
rect 3302 16459 3336 16493
rect 3370 16459 3404 16493
rect 3438 16459 3472 16493
rect 3506 16459 3540 16493
rect 3574 16459 3608 16493
rect 3642 16459 3676 16493
rect 3710 16459 3744 16493
rect 3778 16459 3812 16493
rect 3846 16459 3880 16493
rect 3914 16459 3948 16493
rect 3982 16459 4016 16493
rect 4050 16459 4084 16493
rect 4118 16459 4152 16493
rect 4186 16459 4220 16493
rect 4254 16459 4288 16493
rect 4322 16459 4356 16493
rect 4390 16459 4424 16493
rect 4458 16459 4492 16493
rect 4526 16459 4560 16493
rect 4594 16459 4628 16493
rect 4662 16459 4696 16493
rect 4730 16459 4764 16493
rect 4798 16459 4832 16493
rect 4866 16459 4900 16493
rect 4934 16459 4968 16493
rect 5002 16459 5036 16493
rect 5070 16459 5104 16493
rect 5138 16459 5172 16493
rect 5206 16459 5240 16493
rect 5274 16459 5308 16493
rect 5342 16459 5376 16493
rect 5410 16459 5444 16493
rect 5478 16459 5512 16493
rect 5546 16459 5580 16493
rect 5614 16459 5648 16493
rect 5682 16459 5716 16493
rect 5750 16459 5784 16493
rect 5818 16459 5852 16493
rect 5886 16459 5920 16493
rect 5954 16459 5988 16493
rect 6022 16459 6056 16493
rect 6090 16459 6124 16493
rect 6158 16459 6192 16493
rect 6226 16459 6260 16493
rect 6294 16459 6328 16493
rect 6362 16459 6396 16493
rect 6430 16459 6464 16493
rect 6498 16459 6532 16493
rect 6566 16459 6600 16493
rect 6634 16459 6668 16493
rect 6702 16459 6736 16493
rect 6770 16459 6804 16493
rect 6838 16459 6872 16493
rect 6906 16459 6940 16493
rect 6974 16459 7008 16493
rect 7042 16459 7076 16493
rect 7110 16459 7144 16493
rect 7178 16459 7212 16493
rect 7246 16459 7280 16493
rect 7314 16459 7348 16493
rect 7382 16459 7416 16493
rect 7450 16459 7484 16493
rect 7518 16459 7552 16493
rect 7586 16459 7620 16493
rect 7654 16459 7688 16493
rect 7722 16459 7756 16493
rect 7790 16459 7824 16493
rect 7858 16459 7892 16493
rect 7926 16459 7960 16493
rect 7994 16459 8028 16493
rect 8062 16459 8096 16493
rect 8130 16459 8164 16493
rect 8198 16459 8232 16493
rect 8266 16459 8300 16493
rect 8334 16459 8368 16493
rect 8402 16459 8436 16493
rect 8470 16459 8504 16493
rect 8538 16459 8572 16493
rect 8606 16459 8640 16493
rect 8674 16459 8708 16493
rect 8742 16459 8776 16493
rect 8810 16459 8844 16493
rect 8878 16459 8912 16493
rect 8946 16459 8980 16493
rect 9014 16459 9048 16493
rect 9082 16459 9116 16493
rect 9150 16459 9184 16493
rect 9218 16459 9252 16493
rect 9286 16459 9320 16493
rect 9354 16459 9388 16493
rect 9422 16459 9456 16493
rect 9490 16459 9524 16493
rect 9558 16459 9592 16493
rect 9626 16459 9660 16493
rect 9694 16459 9728 16493
rect 9762 16459 9796 16493
rect 9830 16459 9864 16493
rect 9898 16459 9932 16493
rect 9966 16459 10000 16493
rect 10034 16459 10068 16493
rect 10102 16459 10136 16493
rect 10170 16459 10204 16493
rect 10238 16459 10272 16493
rect 10306 16459 10340 16493
rect 10374 16459 10408 16493
rect 10442 16459 10476 16493
rect 10510 16459 10544 16493
rect 10578 16459 10612 16493
rect 10646 16459 10680 16493
rect 10714 16459 10748 16493
rect 10782 16459 10816 16493
rect 10850 16459 10884 16493
rect 10918 16459 10952 16493
rect 10986 16459 11020 16493
rect 11054 16459 11088 16493
rect 11122 16459 11156 16493
rect 11190 16459 11224 16493
rect 11258 16459 11292 16493
rect 11326 16459 11360 16493
rect 11394 16459 11428 16493
rect 11462 16459 11496 16493
rect 11530 16459 11564 16493
rect 11598 16459 11632 16493
rect 11666 16459 11700 16493
rect 11734 16459 11768 16493
rect 11802 16459 11836 16493
rect 11870 16459 11904 16493
rect 11938 16459 11972 16493
rect 12006 16459 12040 16493
rect 12074 16459 12108 16493
rect 12142 16459 12176 16493
rect 12210 16459 12244 16493
rect 12278 16459 12312 16493
rect 12346 16459 12380 16493
rect 12414 16459 12448 16493
rect 12482 16459 12516 16493
rect 12550 16459 12584 16493
rect 12618 16459 12652 16493
rect 12686 16459 12720 16493
rect 12754 16459 12788 16493
rect 12822 16459 12856 16493
rect 12890 16459 12924 16493
rect 12958 16459 12992 16493
rect 13026 16459 13060 16493
rect 13094 16459 13128 16493
rect 13162 16459 13196 16493
rect 13230 16459 13264 16493
rect 13298 16459 13332 16493
rect 13366 16459 13400 16493
rect 13434 16459 13468 16493
rect 13502 16459 13536 16493
rect 13570 16459 13604 16493
rect 13638 16459 13672 16493
rect 13706 16459 13740 16493
rect 13774 16459 13808 16493
rect 13842 16459 13876 16493
rect 13910 16459 13944 16493
rect 13978 16459 14012 16493
rect 14046 16459 14080 16493
rect 14114 16459 14148 16493
rect 14182 16459 14216 16493
rect 14250 16459 14284 16493
rect 14318 16459 14352 16493
rect 14386 16469 14420 16493
rect 14454 16469 14492 16503
rect 14526 16469 14564 16503
rect 14598 16469 14636 16503
rect 14670 16469 14708 16503
rect 14742 16469 14780 16503
rect 14814 16469 14852 16503
rect 14886 16469 14924 16503
rect 14958 16469 14996 16503
rect 15030 16469 15068 16503
rect 15102 16469 15106 16503
rect 14386 16459 15106 16469
rect 67 16434 15106 16459
rect 67 16425 14420 16434
rect 67 16391 68 16425
rect 102 16391 139 16425
rect 173 16391 210 16425
rect 244 16391 281 16425
rect 315 16391 352 16425
rect 386 16423 14420 16425
rect 386 16391 444 16423
rect 67 16389 444 16391
rect 478 16389 513 16423
rect 547 16389 582 16423
rect 616 16389 651 16423
rect 685 16389 720 16423
rect 754 16389 789 16423
rect 823 16389 858 16423
rect 892 16389 927 16423
rect 961 16389 996 16423
rect 1030 16389 1065 16423
rect 1099 16389 1134 16423
rect 1168 16389 1203 16423
rect 1237 16389 1272 16423
rect 1306 16389 1341 16423
rect 1375 16389 1410 16423
rect 1444 16389 1479 16423
rect 1513 16389 1548 16423
rect 1582 16389 1617 16423
rect 1651 16389 1686 16423
rect 1720 16389 1755 16423
rect 1789 16389 1824 16423
rect 1858 16389 1893 16423
rect 1927 16389 1962 16423
rect 1996 16389 2031 16423
rect 2065 16389 2100 16423
rect 2134 16389 2169 16423
rect 2203 16389 2238 16423
rect 2272 16389 2307 16423
rect 2341 16389 2376 16423
rect 2410 16389 2445 16423
rect 2479 16389 2514 16423
rect 2548 16389 2583 16423
rect 2617 16389 2652 16423
rect 2686 16389 2721 16423
rect 2755 16389 2790 16423
rect 2824 16389 2859 16423
rect 2893 16389 2928 16423
rect 2962 16389 2996 16423
rect 3030 16389 3064 16423
rect 3098 16389 3132 16423
rect 3166 16389 3200 16423
rect 3234 16389 3268 16423
rect 3302 16389 3336 16423
rect 3370 16389 3404 16423
rect 3438 16389 3472 16423
rect 3506 16389 3540 16423
rect 3574 16389 3608 16423
rect 3642 16389 3676 16423
rect 3710 16389 3744 16423
rect 3778 16389 3812 16423
rect 3846 16389 3880 16423
rect 3914 16389 3948 16423
rect 3982 16389 4016 16423
rect 4050 16389 4084 16423
rect 4118 16389 4152 16423
rect 4186 16389 4220 16423
rect 4254 16389 4288 16423
rect 4322 16389 4356 16423
rect 4390 16389 4424 16423
rect 4458 16389 4492 16423
rect 4526 16389 4560 16423
rect 4594 16389 4628 16423
rect 4662 16389 4696 16423
rect 4730 16389 4764 16423
rect 4798 16389 4832 16423
rect 4866 16389 4900 16423
rect 4934 16389 4968 16423
rect 5002 16389 5036 16423
rect 5070 16389 5104 16423
rect 5138 16389 5172 16423
rect 5206 16389 5240 16423
rect 5274 16389 5308 16423
rect 5342 16389 5376 16423
rect 5410 16389 5444 16423
rect 5478 16389 5512 16423
rect 5546 16389 5580 16423
rect 5614 16389 5648 16423
rect 5682 16389 5716 16423
rect 5750 16389 5784 16423
rect 5818 16389 5852 16423
rect 5886 16389 5920 16423
rect 5954 16389 5988 16423
rect 6022 16389 6056 16423
rect 6090 16389 6124 16423
rect 6158 16389 6192 16423
rect 6226 16389 6260 16423
rect 6294 16389 6328 16423
rect 6362 16389 6396 16423
rect 6430 16389 6464 16423
rect 6498 16389 6532 16423
rect 6566 16389 6600 16423
rect 6634 16389 6668 16423
rect 6702 16389 6736 16423
rect 6770 16389 6804 16423
rect 6838 16389 6872 16423
rect 6906 16389 6940 16423
rect 6974 16389 7008 16423
rect 7042 16389 7076 16423
rect 7110 16389 7144 16423
rect 7178 16389 7212 16423
rect 7246 16389 7280 16423
rect 7314 16389 7348 16423
rect 7382 16389 7416 16423
rect 7450 16389 7484 16423
rect 7518 16389 7552 16423
rect 7586 16389 7620 16423
rect 7654 16389 7688 16423
rect 7722 16389 7756 16423
rect 7790 16389 7824 16423
rect 7858 16389 7892 16423
rect 7926 16389 7960 16423
rect 7994 16389 8028 16423
rect 8062 16389 8096 16423
rect 8130 16389 8164 16423
rect 8198 16389 8232 16423
rect 8266 16389 8300 16423
rect 8334 16389 8368 16423
rect 8402 16389 8436 16423
rect 8470 16389 8504 16423
rect 8538 16389 8572 16423
rect 8606 16389 8640 16423
rect 8674 16389 8708 16423
rect 8742 16389 8776 16423
rect 8810 16389 8844 16423
rect 8878 16389 8912 16423
rect 8946 16389 8980 16423
rect 9014 16389 9048 16423
rect 9082 16389 9116 16423
rect 9150 16389 9184 16423
rect 9218 16389 9252 16423
rect 9286 16389 9320 16423
rect 9354 16389 9388 16423
rect 9422 16389 9456 16423
rect 9490 16389 9524 16423
rect 9558 16389 9592 16423
rect 9626 16389 9660 16423
rect 9694 16389 9728 16423
rect 9762 16389 9796 16423
rect 9830 16389 9864 16423
rect 9898 16389 9932 16423
rect 9966 16389 10000 16423
rect 10034 16389 10068 16423
rect 10102 16389 10136 16423
rect 10170 16389 10204 16423
rect 10238 16389 10272 16423
rect 10306 16389 10340 16423
rect 10374 16389 10408 16423
rect 10442 16389 10476 16423
rect 10510 16389 10544 16423
rect 10578 16389 10612 16423
rect 10646 16389 10680 16423
rect 10714 16389 10748 16423
rect 10782 16389 10816 16423
rect 10850 16389 10884 16423
rect 10918 16389 10952 16423
rect 10986 16389 11020 16423
rect 11054 16389 11088 16423
rect 11122 16389 11156 16423
rect 11190 16389 11224 16423
rect 11258 16389 11292 16423
rect 11326 16389 11360 16423
rect 11394 16389 11428 16423
rect 11462 16389 11496 16423
rect 11530 16389 11564 16423
rect 11598 16389 11632 16423
rect 11666 16389 11700 16423
rect 11734 16389 11768 16423
rect 11802 16389 11836 16423
rect 11870 16389 11904 16423
rect 11938 16389 11972 16423
rect 12006 16389 12040 16423
rect 12074 16389 12108 16423
rect 12142 16389 12176 16423
rect 12210 16389 12244 16423
rect 12278 16389 12312 16423
rect 12346 16389 12380 16423
rect 12414 16389 12448 16423
rect 12482 16389 12516 16423
rect 12550 16389 12584 16423
rect 12618 16389 12652 16423
rect 12686 16389 12720 16423
rect 12754 16389 12788 16423
rect 12822 16389 12856 16423
rect 12890 16389 12924 16423
rect 12958 16389 12992 16423
rect 13026 16389 13060 16423
rect 13094 16389 13128 16423
rect 13162 16389 13196 16423
rect 13230 16389 13264 16423
rect 13298 16389 13332 16423
rect 13366 16389 13400 16423
rect 13434 16389 13468 16423
rect 13502 16389 13536 16423
rect 13570 16389 13604 16423
rect 13638 16389 13672 16423
rect 13706 16389 13740 16423
rect 13774 16389 13808 16423
rect 13842 16389 13876 16423
rect 13910 16389 13944 16423
rect 13978 16389 14012 16423
rect 14046 16389 14080 16423
rect 14114 16389 14148 16423
rect 14182 16389 14216 16423
rect 14250 16389 14284 16423
rect 14318 16389 14352 16423
rect 14386 16400 14420 16423
rect 14454 16400 14492 16434
rect 14526 16400 14564 16434
rect 14598 16400 14636 16434
rect 14670 16400 14708 16434
rect 14742 16400 14780 16434
rect 14814 16400 14852 16434
rect 14886 16400 14924 16434
rect 14958 16400 14996 16434
rect 15030 16400 15068 16434
rect 15102 16400 15106 16434
rect 14386 16389 15106 16400
rect 67 16365 15106 16389
rect 67 16357 14420 16365
rect 67 16323 68 16357
rect 102 16323 139 16357
rect 173 16323 210 16357
rect 244 16323 281 16357
rect 315 16323 352 16357
rect 386 16353 14420 16357
rect 386 16323 444 16353
rect 67 16319 444 16323
rect 478 16319 513 16353
rect 547 16319 582 16353
rect 616 16319 651 16353
rect 685 16319 720 16353
rect 754 16319 789 16353
rect 823 16319 858 16353
rect 892 16319 927 16353
rect 961 16319 996 16353
rect 1030 16319 1065 16353
rect 1099 16319 1134 16353
rect 1168 16319 1203 16353
rect 1237 16319 1272 16353
rect 1306 16319 1341 16353
rect 1375 16319 1410 16353
rect 1444 16319 1479 16353
rect 1513 16319 1548 16353
rect 1582 16319 1617 16353
rect 1651 16319 1686 16353
rect 1720 16319 1755 16353
rect 1789 16319 1824 16353
rect 1858 16319 1893 16353
rect 1927 16319 1962 16353
rect 1996 16319 2031 16353
rect 2065 16319 2100 16353
rect 2134 16319 2169 16353
rect 2203 16319 2238 16353
rect 2272 16319 2307 16353
rect 2341 16319 2376 16353
rect 2410 16319 2445 16353
rect 2479 16319 2514 16353
rect 2548 16319 2583 16353
rect 2617 16319 2652 16353
rect 2686 16319 2721 16353
rect 2755 16319 2790 16353
rect 2824 16319 2859 16353
rect 2893 16319 2928 16353
rect 2962 16319 2996 16353
rect 3030 16319 3064 16353
rect 3098 16319 3132 16353
rect 3166 16319 3200 16353
rect 3234 16319 3268 16353
rect 3302 16319 3336 16353
rect 3370 16319 3404 16353
rect 3438 16319 3472 16353
rect 3506 16319 3540 16353
rect 3574 16319 3608 16353
rect 3642 16319 3676 16353
rect 3710 16319 3744 16353
rect 3778 16319 3812 16353
rect 3846 16319 3880 16353
rect 3914 16319 3948 16353
rect 3982 16319 4016 16353
rect 4050 16319 4084 16353
rect 4118 16319 4152 16353
rect 4186 16319 4220 16353
rect 4254 16319 4288 16353
rect 4322 16319 4356 16353
rect 4390 16319 4424 16353
rect 4458 16319 4492 16353
rect 4526 16319 4560 16353
rect 4594 16319 4628 16353
rect 4662 16319 4696 16353
rect 4730 16319 4764 16353
rect 4798 16319 4832 16353
rect 4866 16319 4900 16353
rect 4934 16319 4968 16353
rect 5002 16319 5036 16353
rect 5070 16319 5104 16353
rect 5138 16319 5172 16353
rect 5206 16319 5240 16353
rect 5274 16319 5308 16353
rect 5342 16319 5376 16353
rect 5410 16319 5444 16353
rect 5478 16319 5512 16353
rect 5546 16319 5580 16353
rect 5614 16319 5648 16353
rect 5682 16319 5716 16353
rect 5750 16319 5784 16353
rect 5818 16319 5852 16353
rect 5886 16319 5920 16353
rect 5954 16319 5988 16353
rect 6022 16319 6056 16353
rect 6090 16319 6124 16353
rect 6158 16319 6192 16353
rect 6226 16319 6260 16353
rect 6294 16319 6328 16353
rect 6362 16319 6396 16353
rect 6430 16319 6464 16353
rect 6498 16319 6532 16353
rect 6566 16319 6600 16353
rect 6634 16319 6668 16353
rect 6702 16319 6736 16353
rect 6770 16319 6804 16353
rect 6838 16319 6872 16353
rect 6906 16319 6940 16353
rect 6974 16319 7008 16353
rect 7042 16319 7076 16353
rect 7110 16319 7144 16353
rect 7178 16319 7212 16353
rect 7246 16319 7280 16353
rect 7314 16319 7348 16353
rect 7382 16319 7416 16353
rect 7450 16319 7484 16353
rect 7518 16319 7552 16353
rect 7586 16319 7620 16353
rect 7654 16319 7688 16353
rect 7722 16319 7756 16353
rect 7790 16319 7824 16353
rect 7858 16319 7892 16353
rect 7926 16319 7960 16353
rect 7994 16319 8028 16353
rect 8062 16319 8096 16353
rect 8130 16319 8164 16353
rect 8198 16319 8232 16353
rect 8266 16319 8300 16353
rect 8334 16319 8368 16353
rect 8402 16319 8436 16353
rect 8470 16319 8504 16353
rect 8538 16319 8572 16353
rect 8606 16319 8640 16353
rect 8674 16319 8708 16353
rect 8742 16319 8776 16353
rect 8810 16319 8844 16353
rect 8878 16319 8912 16353
rect 8946 16319 8980 16353
rect 9014 16319 9048 16353
rect 9082 16319 9116 16353
rect 9150 16319 9184 16353
rect 9218 16319 9252 16353
rect 9286 16319 9320 16353
rect 9354 16319 9388 16353
rect 9422 16319 9456 16353
rect 9490 16319 9524 16353
rect 9558 16319 9592 16353
rect 9626 16319 9660 16353
rect 9694 16319 9728 16353
rect 9762 16319 9796 16353
rect 9830 16319 9864 16353
rect 9898 16319 9932 16353
rect 9966 16319 10000 16353
rect 10034 16319 10068 16353
rect 10102 16319 10136 16353
rect 10170 16319 10204 16353
rect 10238 16319 10272 16353
rect 10306 16319 10340 16353
rect 10374 16319 10408 16353
rect 10442 16319 10476 16353
rect 10510 16319 10544 16353
rect 10578 16319 10612 16353
rect 10646 16319 10680 16353
rect 10714 16319 10748 16353
rect 10782 16319 10816 16353
rect 10850 16319 10884 16353
rect 10918 16319 10952 16353
rect 10986 16319 11020 16353
rect 11054 16319 11088 16353
rect 11122 16319 11156 16353
rect 11190 16319 11224 16353
rect 11258 16319 11292 16353
rect 11326 16319 11360 16353
rect 11394 16319 11428 16353
rect 11462 16319 11496 16353
rect 11530 16319 11564 16353
rect 11598 16319 11632 16353
rect 11666 16319 11700 16353
rect 11734 16319 11768 16353
rect 11802 16319 11836 16353
rect 11870 16319 11904 16353
rect 11938 16319 11972 16353
rect 12006 16319 12040 16353
rect 12074 16319 12108 16353
rect 12142 16319 12176 16353
rect 12210 16319 12244 16353
rect 12278 16319 12312 16353
rect 12346 16319 12380 16353
rect 12414 16319 12448 16353
rect 12482 16319 12516 16353
rect 12550 16319 12584 16353
rect 12618 16319 12652 16353
rect 12686 16319 12720 16353
rect 12754 16319 12788 16353
rect 12822 16319 12856 16353
rect 12890 16319 12924 16353
rect 12958 16319 12992 16353
rect 13026 16319 13060 16353
rect 13094 16319 13128 16353
rect 13162 16319 13196 16353
rect 13230 16319 13264 16353
rect 13298 16319 13332 16353
rect 13366 16319 13400 16353
rect 13434 16319 13468 16353
rect 13502 16319 13536 16353
rect 13570 16319 13604 16353
rect 13638 16319 13672 16353
rect 13706 16319 13740 16353
rect 13774 16319 13808 16353
rect 13842 16319 13876 16353
rect 13910 16319 13944 16353
rect 13978 16319 14012 16353
rect 14046 16319 14080 16353
rect 14114 16319 14148 16353
rect 14182 16319 14216 16353
rect 14250 16319 14284 16353
rect 14318 16319 14352 16353
rect 14386 16331 14420 16353
rect 14454 16331 14492 16365
rect 14526 16331 14564 16365
rect 14598 16331 14636 16365
rect 14670 16331 14708 16365
rect 14742 16331 14780 16365
rect 14814 16331 14852 16365
rect 14886 16331 14924 16365
rect 14958 16331 14996 16365
rect 15030 16331 15068 16365
rect 15102 16331 15106 16365
rect 14386 16319 15106 16331
rect 67 16296 15106 16319
rect 67 16289 14420 16296
rect 67 16255 68 16289
rect 102 16255 139 16289
rect 173 16255 210 16289
rect 244 16255 281 16289
rect 315 16255 352 16289
rect 386 16283 14420 16289
rect 386 16255 444 16283
rect 67 16249 444 16255
rect 478 16249 513 16283
rect 547 16249 582 16283
rect 616 16249 651 16283
rect 685 16249 720 16283
rect 754 16249 789 16283
rect 823 16249 858 16283
rect 892 16249 927 16283
rect 961 16249 996 16283
rect 1030 16249 1065 16283
rect 1099 16249 1134 16283
rect 1168 16249 1203 16283
rect 1237 16249 1272 16283
rect 1306 16249 1341 16283
rect 1375 16249 1410 16283
rect 1444 16249 1479 16283
rect 1513 16249 1548 16283
rect 1582 16249 1617 16283
rect 1651 16249 1686 16283
rect 1720 16249 1755 16283
rect 1789 16249 1824 16283
rect 1858 16249 1893 16283
rect 1927 16249 1962 16283
rect 1996 16249 2031 16283
rect 2065 16249 2100 16283
rect 2134 16249 2169 16283
rect 2203 16249 2238 16283
rect 2272 16249 2307 16283
rect 2341 16249 2376 16283
rect 2410 16249 2445 16283
rect 2479 16249 2514 16283
rect 2548 16249 2583 16283
rect 2617 16249 2652 16283
rect 2686 16249 2721 16283
rect 2755 16249 2790 16283
rect 2824 16249 2859 16283
rect 2893 16249 2928 16283
rect 2962 16249 2996 16283
rect 3030 16249 3064 16283
rect 3098 16249 3132 16283
rect 3166 16249 3200 16283
rect 3234 16249 3268 16283
rect 3302 16249 3336 16283
rect 3370 16249 3404 16283
rect 3438 16249 3472 16283
rect 3506 16249 3540 16283
rect 3574 16249 3608 16283
rect 3642 16249 3676 16283
rect 3710 16249 3744 16283
rect 3778 16249 3812 16283
rect 3846 16249 3880 16283
rect 3914 16249 3948 16283
rect 3982 16249 4016 16283
rect 4050 16249 4084 16283
rect 4118 16249 4152 16283
rect 4186 16249 4220 16283
rect 4254 16249 4288 16283
rect 4322 16249 4356 16283
rect 4390 16249 4424 16283
rect 4458 16249 4492 16283
rect 4526 16249 4560 16283
rect 4594 16249 4628 16283
rect 4662 16249 4696 16283
rect 4730 16249 4764 16283
rect 4798 16249 4832 16283
rect 4866 16249 4900 16283
rect 4934 16249 4968 16283
rect 5002 16249 5036 16283
rect 5070 16249 5104 16283
rect 5138 16249 5172 16283
rect 5206 16249 5240 16283
rect 5274 16249 5308 16283
rect 5342 16249 5376 16283
rect 5410 16249 5444 16283
rect 5478 16249 5512 16283
rect 5546 16249 5580 16283
rect 5614 16249 5648 16283
rect 5682 16249 5716 16283
rect 5750 16249 5784 16283
rect 5818 16249 5852 16283
rect 5886 16249 5920 16283
rect 5954 16249 5988 16283
rect 6022 16249 6056 16283
rect 6090 16249 6124 16283
rect 6158 16249 6192 16283
rect 6226 16249 6260 16283
rect 6294 16249 6328 16283
rect 6362 16249 6396 16283
rect 6430 16249 6464 16283
rect 6498 16249 6532 16283
rect 6566 16249 6600 16283
rect 6634 16249 6668 16283
rect 6702 16249 6736 16283
rect 6770 16249 6804 16283
rect 6838 16249 6872 16283
rect 6906 16249 6940 16283
rect 6974 16249 7008 16283
rect 7042 16249 7076 16283
rect 7110 16249 7144 16283
rect 7178 16249 7212 16283
rect 7246 16249 7280 16283
rect 7314 16249 7348 16283
rect 7382 16249 7416 16283
rect 7450 16249 7484 16283
rect 7518 16249 7552 16283
rect 7586 16249 7620 16283
rect 7654 16249 7688 16283
rect 7722 16249 7756 16283
rect 7790 16249 7824 16283
rect 7858 16249 7892 16283
rect 7926 16249 7960 16283
rect 7994 16249 8028 16283
rect 8062 16249 8096 16283
rect 8130 16249 8164 16283
rect 8198 16249 8232 16283
rect 8266 16249 8300 16283
rect 8334 16249 8368 16283
rect 8402 16249 8436 16283
rect 8470 16249 8504 16283
rect 8538 16249 8572 16283
rect 8606 16249 8640 16283
rect 8674 16249 8708 16283
rect 8742 16249 8776 16283
rect 8810 16249 8844 16283
rect 8878 16249 8912 16283
rect 8946 16249 8980 16283
rect 9014 16249 9048 16283
rect 9082 16249 9116 16283
rect 9150 16249 9184 16283
rect 9218 16249 9252 16283
rect 9286 16249 9320 16283
rect 9354 16249 9388 16283
rect 9422 16249 9456 16283
rect 9490 16249 9524 16283
rect 9558 16249 9592 16283
rect 9626 16249 9660 16283
rect 9694 16249 9728 16283
rect 9762 16249 9796 16283
rect 9830 16249 9864 16283
rect 9898 16249 9932 16283
rect 9966 16249 10000 16283
rect 10034 16249 10068 16283
rect 10102 16249 10136 16283
rect 10170 16249 10204 16283
rect 10238 16249 10272 16283
rect 10306 16249 10340 16283
rect 10374 16249 10408 16283
rect 10442 16249 10476 16283
rect 10510 16249 10544 16283
rect 10578 16249 10612 16283
rect 10646 16249 10680 16283
rect 10714 16249 10748 16283
rect 10782 16249 10816 16283
rect 10850 16249 10884 16283
rect 10918 16249 10952 16283
rect 10986 16249 11020 16283
rect 11054 16249 11088 16283
rect 11122 16249 11156 16283
rect 11190 16249 11224 16283
rect 11258 16249 11292 16283
rect 11326 16249 11360 16283
rect 11394 16249 11428 16283
rect 11462 16249 11496 16283
rect 11530 16249 11564 16283
rect 11598 16249 11632 16283
rect 11666 16249 11700 16283
rect 11734 16249 11768 16283
rect 11802 16249 11836 16283
rect 11870 16249 11904 16283
rect 11938 16249 11972 16283
rect 12006 16249 12040 16283
rect 12074 16249 12108 16283
rect 12142 16249 12176 16283
rect 12210 16249 12244 16283
rect 12278 16249 12312 16283
rect 12346 16249 12380 16283
rect 12414 16249 12448 16283
rect 12482 16249 12516 16283
rect 12550 16249 12584 16283
rect 12618 16249 12652 16283
rect 12686 16249 12720 16283
rect 12754 16249 12788 16283
rect 12822 16249 12856 16283
rect 12890 16249 12924 16283
rect 12958 16249 12992 16283
rect 13026 16249 13060 16283
rect 13094 16249 13128 16283
rect 13162 16249 13196 16283
rect 13230 16249 13264 16283
rect 13298 16249 13332 16283
rect 13366 16249 13400 16283
rect 13434 16249 13468 16283
rect 13502 16249 13536 16283
rect 13570 16249 13604 16283
rect 13638 16249 13672 16283
rect 13706 16249 13740 16283
rect 13774 16249 13808 16283
rect 13842 16249 13876 16283
rect 13910 16249 13944 16283
rect 13978 16249 14012 16283
rect 14046 16249 14080 16283
rect 14114 16249 14148 16283
rect 14182 16249 14216 16283
rect 14250 16249 14284 16283
rect 14318 16249 14352 16283
rect 14386 16262 14420 16283
rect 14454 16262 14492 16296
rect 14526 16262 14564 16296
rect 14598 16262 14636 16296
rect 14670 16262 14708 16296
rect 14742 16262 14780 16296
rect 14814 16262 14852 16296
rect 14886 16262 14924 16296
rect 14958 16262 14996 16296
rect 15030 16262 15068 16296
rect 15102 16262 15106 16296
rect 14386 16249 15106 16262
rect 67 16227 15106 16249
rect 67 16221 14420 16227
rect 67 16187 68 16221
rect 102 16187 139 16221
rect 173 16187 210 16221
rect 244 16187 281 16221
rect 315 16187 352 16221
rect 386 16213 14420 16221
rect 386 16187 444 16213
rect 67 16179 444 16187
rect 478 16179 513 16213
rect 547 16179 582 16213
rect 616 16179 651 16213
rect 685 16179 720 16213
rect 754 16179 789 16213
rect 823 16179 858 16213
rect 892 16179 927 16213
rect 961 16179 996 16213
rect 1030 16179 1065 16213
rect 1099 16179 1134 16213
rect 1168 16179 1203 16213
rect 1237 16179 1272 16213
rect 1306 16179 1341 16213
rect 1375 16179 1410 16213
rect 1444 16179 1479 16213
rect 1513 16179 1548 16213
rect 1582 16179 1617 16213
rect 1651 16179 1686 16213
rect 1720 16179 1755 16213
rect 1789 16179 1824 16213
rect 1858 16179 1893 16213
rect 1927 16179 1962 16213
rect 1996 16179 2031 16213
rect 2065 16179 2100 16213
rect 2134 16179 2169 16213
rect 2203 16179 2238 16213
rect 2272 16179 2307 16213
rect 2341 16179 2376 16213
rect 2410 16179 2445 16213
rect 2479 16179 2514 16213
rect 2548 16179 2583 16213
rect 2617 16179 2652 16213
rect 2686 16179 2721 16213
rect 2755 16179 2790 16213
rect 2824 16179 2859 16213
rect 2893 16179 2928 16213
rect 2962 16179 2996 16213
rect 3030 16179 3064 16213
rect 3098 16179 3132 16213
rect 3166 16179 3200 16213
rect 3234 16179 3268 16213
rect 3302 16179 3336 16213
rect 3370 16179 3404 16213
rect 3438 16179 3472 16213
rect 3506 16179 3540 16213
rect 3574 16179 3608 16213
rect 3642 16179 3676 16213
rect 3710 16179 3744 16213
rect 3778 16179 3812 16213
rect 3846 16179 3880 16213
rect 3914 16179 3948 16213
rect 3982 16179 4016 16213
rect 4050 16179 4084 16213
rect 4118 16179 4152 16213
rect 4186 16179 4220 16213
rect 4254 16179 4288 16213
rect 4322 16179 4356 16213
rect 4390 16179 4424 16213
rect 4458 16179 4492 16213
rect 4526 16179 4560 16213
rect 4594 16179 4628 16213
rect 4662 16179 4696 16213
rect 4730 16179 4764 16213
rect 4798 16179 4832 16213
rect 4866 16179 4900 16213
rect 4934 16179 4968 16213
rect 5002 16179 5036 16213
rect 5070 16179 5104 16213
rect 5138 16179 5172 16213
rect 5206 16179 5240 16213
rect 5274 16179 5308 16213
rect 5342 16179 5376 16213
rect 5410 16179 5444 16213
rect 5478 16179 5512 16213
rect 5546 16179 5580 16213
rect 5614 16179 5648 16213
rect 5682 16179 5716 16213
rect 5750 16179 5784 16213
rect 5818 16179 5852 16213
rect 5886 16179 5920 16213
rect 5954 16179 5988 16213
rect 6022 16179 6056 16213
rect 6090 16179 6124 16213
rect 6158 16179 6192 16213
rect 6226 16179 6260 16213
rect 6294 16179 6328 16213
rect 6362 16179 6396 16213
rect 6430 16179 6464 16213
rect 6498 16179 6532 16213
rect 6566 16179 6600 16213
rect 6634 16179 6668 16213
rect 6702 16179 6736 16213
rect 6770 16179 6804 16213
rect 6838 16179 6872 16213
rect 6906 16179 6940 16213
rect 6974 16179 7008 16213
rect 7042 16179 7076 16213
rect 7110 16179 7144 16213
rect 7178 16179 7212 16213
rect 7246 16179 7280 16213
rect 7314 16179 7348 16213
rect 7382 16179 7416 16213
rect 7450 16179 7484 16213
rect 7518 16179 7552 16213
rect 7586 16179 7620 16213
rect 7654 16179 7688 16213
rect 7722 16179 7756 16213
rect 7790 16179 7824 16213
rect 7858 16179 7892 16213
rect 7926 16179 7960 16213
rect 7994 16179 8028 16213
rect 8062 16179 8096 16213
rect 8130 16179 8164 16213
rect 8198 16179 8232 16213
rect 8266 16179 8300 16213
rect 8334 16179 8368 16213
rect 8402 16179 8436 16213
rect 8470 16179 8504 16213
rect 8538 16179 8572 16213
rect 8606 16179 8640 16213
rect 8674 16179 8708 16213
rect 8742 16179 8776 16213
rect 8810 16179 8844 16213
rect 8878 16179 8912 16213
rect 8946 16179 8980 16213
rect 9014 16179 9048 16213
rect 9082 16179 9116 16213
rect 9150 16179 9184 16213
rect 9218 16179 9252 16213
rect 9286 16179 9320 16213
rect 9354 16179 9388 16213
rect 9422 16179 9456 16213
rect 9490 16179 9524 16213
rect 9558 16179 9592 16213
rect 9626 16179 9660 16213
rect 9694 16179 9728 16213
rect 9762 16179 9796 16213
rect 9830 16179 9864 16213
rect 9898 16179 9932 16213
rect 9966 16179 10000 16213
rect 10034 16179 10068 16213
rect 10102 16179 10136 16213
rect 10170 16179 10204 16213
rect 10238 16179 10272 16213
rect 10306 16179 10340 16213
rect 10374 16179 10408 16213
rect 10442 16179 10476 16213
rect 10510 16179 10544 16213
rect 10578 16179 10612 16213
rect 10646 16179 10680 16213
rect 10714 16179 10748 16213
rect 10782 16179 10816 16213
rect 10850 16179 10884 16213
rect 10918 16179 10952 16213
rect 10986 16179 11020 16213
rect 11054 16179 11088 16213
rect 11122 16179 11156 16213
rect 11190 16179 11224 16213
rect 11258 16179 11292 16213
rect 11326 16179 11360 16213
rect 11394 16179 11428 16213
rect 11462 16179 11496 16213
rect 11530 16179 11564 16213
rect 11598 16179 11632 16213
rect 11666 16179 11700 16213
rect 11734 16179 11768 16213
rect 11802 16179 11836 16213
rect 11870 16179 11904 16213
rect 11938 16179 11972 16213
rect 12006 16179 12040 16213
rect 12074 16179 12108 16213
rect 12142 16179 12176 16213
rect 12210 16179 12244 16213
rect 12278 16179 12312 16213
rect 12346 16179 12380 16213
rect 12414 16179 12448 16213
rect 12482 16179 12516 16213
rect 12550 16179 12584 16213
rect 12618 16179 12652 16213
rect 12686 16179 12720 16213
rect 12754 16179 12788 16213
rect 12822 16179 12856 16213
rect 12890 16179 12924 16213
rect 12958 16179 12992 16213
rect 13026 16179 13060 16213
rect 13094 16179 13128 16213
rect 13162 16179 13196 16213
rect 13230 16179 13264 16213
rect 13298 16179 13332 16213
rect 13366 16179 13400 16213
rect 13434 16179 13468 16213
rect 13502 16179 13536 16213
rect 13570 16179 13604 16213
rect 13638 16179 13672 16213
rect 13706 16179 13740 16213
rect 13774 16179 13808 16213
rect 13842 16179 13876 16213
rect 13910 16179 13944 16213
rect 13978 16179 14012 16213
rect 14046 16179 14080 16213
rect 14114 16179 14148 16213
rect 14182 16179 14216 16213
rect 14250 16179 14284 16213
rect 14318 16179 14352 16213
rect 14386 16193 14420 16213
rect 14454 16193 14492 16227
rect 14526 16193 14564 16227
rect 14598 16193 14636 16227
rect 14670 16193 14708 16227
rect 14742 16193 14780 16227
rect 14814 16193 14852 16227
rect 14886 16193 14924 16227
rect 14958 16193 14996 16227
rect 15030 16193 15068 16227
rect 15102 16193 15106 16227
rect 14386 16179 15106 16193
rect 67 16158 15106 16179
rect 67 16153 14420 16158
rect 67 16119 68 16153
rect 102 16119 139 16153
rect 173 16119 210 16153
rect 244 16119 281 16153
rect 315 16119 352 16153
rect 386 16143 14420 16153
rect 386 16119 444 16143
rect 67 16109 444 16119
rect 478 16109 513 16143
rect 547 16109 582 16143
rect 616 16109 651 16143
rect 685 16109 720 16143
rect 754 16109 789 16143
rect 823 16109 858 16143
rect 892 16109 927 16143
rect 961 16109 996 16143
rect 1030 16109 1065 16143
rect 1099 16109 1134 16143
rect 1168 16109 1203 16143
rect 1237 16109 1272 16143
rect 1306 16109 1341 16143
rect 1375 16109 1410 16143
rect 1444 16109 1479 16143
rect 1513 16109 1548 16143
rect 1582 16109 1617 16143
rect 1651 16109 1686 16143
rect 1720 16109 1755 16143
rect 1789 16109 1824 16143
rect 1858 16109 1893 16143
rect 1927 16109 1962 16143
rect 1996 16109 2031 16143
rect 2065 16109 2100 16143
rect 2134 16109 2169 16143
rect 2203 16109 2238 16143
rect 2272 16109 2307 16143
rect 2341 16109 2376 16143
rect 2410 16109 2445 16143
rect 2479 16109 2514 16143
rect 2548 16109 2583 16143
rect 2617 16109 2652 16143
rect 2686 16109 2721 16143
rect 2755 16109 2790 16143
rect 2824 16109 2859 16143
rect 2893 16109 2928 16143
rect 2962 16109 2996 16143
rect 3030 16109 3064 16143
rect 3098 16109 3132 16143
rect 3166 16109 3200 16143
rect 3234 16109 3268 16143
rect 3302 16109 3336 16143
rect 3370 16109 3404 16143
rect 3438 16109 3472 16143
rect 3506 16109 3540 16143
rect 3574 16109 3608 16143
rect 3642 16109 3676 16143
rect 3710 16109 3744 16143
rect 3778 16109 3812 16143
rect 3846 16109 3880 16143
rect 3914 16109 3948 16143
rect 3982 16109 4016 16143
rect 4050 16109 4084 16143
rect 4118 16109 4152 16143
rect 4186 16109 4220 16143
rect 4254 16109 4288 16143
rect 4322 16109 4356 16143
rect 4390 16109 4424 16143
rect 4458 16109 4492 16143
rect 4526 16109 4560 16143
rect 4594 16109 4628 16143
rect 4662 16109 4696 16143
rect 4730 16109 4764 16143
rect 4798 16109 4832 16143
rect 4866 16109 4900 16143
rect 4934 16109 4968 16143
rect 5002 16109 5036 16143
rect 5070 16109 5104 16143
rect 5138 16109 5172 16143
rect 5206 16109 5240 16143
rect 5274 16109 5308 16143
rect 5342 16109 5376 16143
rect 5410 16109 5444 16143
rect 5478 16109 5512 16143
rect 5546 16109 5580 16143
rect 5614 16109 5648 16143
rect 5682 16109 5716 16143
rect 5750 16109 5784 16143
rect 5818 16109 5852 16143
rect 5886 16109 5920 16143
rect 5954 16109 5988 16143
rect 6022 16109 6056 16143
rect 6090 16109 6124 16143
rect 6158 16109 6192 16143
rect 6226 16109 6260 16143
rect 6294 16109 6328 16143
rect 6362 16109 6396 16143
rect 6430 16109 6464 16143
rect 6498 16109 6532 16143
rect 6566 16109 6600 16143
rect 6634 16109 6668 16143
rect 6702 16109 6736 16143
rect 6770 16109 6804 16143
rect 6838 16109 6872 16143
rect 6906 16109 6940 16143
rect 6974 16109 7008 16143
rect 7042 16109 7076 16143
rect 7110 16109 7144 16143
rect 7178 16109 7212 16143
rect 7246 16109 7280 16143
rect 7314 16109 7348 16143
rect 7382 16109 7416 16143
rect 7450 16109 7484 16143
rect 7518 16109 7552 16143
rect 7586 16109 7620 16143
rect 7654 16109 7688 16143
rect 7722 16109 7756 16143
rect 7790 16109 7824 16143
rect 7858 16109 7892 16143
rect 7926 16109 7960 16143
rect 7994 16109 8028 16143
rect 8062 16109 8096 16143
rect 8130 16109 8164 16143
rect 8198 16109 8232 16143
rect 8266 16109 8300 16143
rect 8334 16109 8368 16143
rect 8402 16109 8436 16143
rect 8470 16109 8504 16143
rect 8538 16109 8572 16143
rect 8606 16109 8640 16143
rect 8674 16109 8708 16143
rect 8742 16109 8776 16143
rect 8810 16109 8844 16143
rect 8878 16109 8912 16143
rect 8946 16109 8980 16143
rect 9014 16109 9048 16143
rect 9082 16109 9116 16143
rect 9150 16109 9184 16143
rect 9218 16109 9252 16143
rect 9286 16109 9320 16143
rect 9354 16109 9388 16143
rect 9422 16109 9456 16143
rect 9490 16109 9524 16143
rect 9558 16109 9592 16143
rect 9626 16109 9660 16143
rect 9694 16109 9728 16143
rect 9762 16109 9796 16143
rect 9830 16109 9864 16143
rect 9898 16109 9932 16143
rect 9966 16109 10000 16143
rect 10034 16109 10068 16143
rect 10102 16109 10136 16143
rect 10170 16109 10204 16143
rect 10238 16109 10272 16143
rect 10306 16109 10340 16143
rect 10374 16109 10408 16143
rect 10442 16109 10476 16143
rect 10510 16109 10544 16143
rect 10578 16109 10612 16143
rect 10646 16109 10680 16143
rect 10714 16109 10748 16143
rect 10782 16109 10816 16143
rect 10850 16109 10884 16143
rect 10918 16109 10952 16143
rect 10986 16109 11020 16143
rect 11054 16109 11088 16143
rect 11122 16109 11156 16143
rect 11190 16109 11224 16143
rect 11258 16109 11292 16143
rect 11326 16109 11360 16143
rect 11394 16109 11428 16143
rect 11462 16109 11496 16143
rect 11530 16109 11564 16143
rect 11598 16109 11632 16143
rect 11666 16109 11700 16143
rect 11734 16109 11768 16143
rect 11802 16109 11836 16143
rect 11870 16109 11904 16143
rect 11938 16109 11972 16143
rect 12006 16109 12040 16143
rect 12074 16109 12108 16143
rect 12142 16109 12176 16143
rect 12210 16109 12244 16143
rect 12278 16109 12312 16143
rect 12346 16109 12380 16143
rect 12414 16109 12448 16143
rect 12482 16109 12516 16143
rect 12550 16109 12584 16143
rect 12618 16109 12652 16143
rect 12686 16109 12720 16143
rect 12754 16109 12788 16143
rect 12822 16109 12856 16143
rect 12890 16109 12924 16143
rect 12958 16109 12992 16143
rect 13026 16109 13060 16143
rect 13094 16109 13128 16143
rect 13162 16109 13196 16143
rect 13230 16109 13264 16143
rect 13298 16109 13332 16143
rect 13366 16109 13400 16143
rect 13434 16109 13468 16143
rect 13502 16109 13536 16143
rect 13570 16109 13604 16143
rect 13638 16109 13672 16143
rect 13706 16109 13740 16143
rect 13774 16109 13808 16143
rect 13842 16109 13876 16143
rect 13910 16109 13944 16143
rect 13978 16109 14012 16143
rect 14046 16109 14080 16143
rect 14114 16109 14148 16143
rect 14182 16109 14216 16143
rect 14250 16109 14284 16143
rect 14318 16109 14352 16143
rect 14386 16124 14420 16143
rect 14454 16124 14492 16158
rect 14526 16124 14564 16158
rect 14598 16124 14636 16158
rect 14670 16124 14708 16158
rect 14742 16124 14780 16158
rect 14814 16124 14852 16158
rect 14886 16124 14924 16158
rect 14958 16124 14996 16158
rect 15030 16124 15068 16158
rect 15102 16124 15106 16158
rect 14386 16109 15106 16124
rect 67 16089 15106 16109
rect 67 16085 14420 16089
rect 67 16051 68 16085
rect 102 16051 139 16085
rect 173 16051 210 16085
rect 244 16051 281 16085
rect 315 16051 352 16085
rect 386 16073 14420 16085
rect 386 16051 444 16073
rect 67 16039 444 16051
rect 478 16039 513 16073
rect 547 16039 582 16073
rect 616 16039 651 16073
rect 685 16039 720 16073
rect 754 16039 789 16073
rect 823 16039 858 16073
rect 892 16039 927 16073
rect 961 16039 996 16073
rect 1030 16039 1065 16073
rect 1099 16039 1134 16073
rect 1168 16039 1203 16073
rect 1237 16039 1272 16073
rect 1306 16039 1341 16073
rect 1375 16039 1410 16073
rect 1444 16039 1479 16073
rect 1513 16039 1548 16073
rect 1582 16039 1617 16073
rect 1651 16039 1686 16073
rect 1720 16039 1755 16073
rect 1789 16039 1824 16073
rect 1858 16039 1893 16073
rect 1927 16039 1962 16073
rect 1996 16039 2031 16073
rect 2065 16039 2100 16073
rect 2134 16039 2169 16073
rect 2203 16039 2238 16073
rect 2272 16039 2307 16073
rect 2341 16039 2376 16073
rect 2410 16039 2445 16073
rect 2479 16039 2514 16073
rect 2548 16039 2583 16073
rect 2617 16039 2652 16073
rect 2686 16039 2721 16073
rect 2755 16039 2790 16073
rect 2824 16039 2859 16073
rect 2893 16039 2928 16073
rect 2962 16039 2996 16073
rect 3030 16039 3064 16073
rect 3098 16039 3132 16073
rect 3166 16039 3200 16073
rect 3234 16039 3268 16073
rect 3302 16039 3336 16073
rect 3370 16039 3404 16073
rect 3438 16039 3472 16073
rect 3506 16039 3540 16073
rect 3574 16039 3608 16073
rect 3642 16039 3676 16073
rect 3710 16039 3744 16073
rect 3778 16039 3812 16073
rect 3846 16039 3880 16073
rect 3914 16039 3948 16073
rect 3982 16039 4016 16073
rect 4050 16039 4084 16073
rect 4118 16039 4152 16073
rect 4186 16039 4220 16073
rect 4254 16039 4288 16073
rect 4322 16039 4356 16073
rect 4390 16039 4424 16073
rect 4458 16039 4492 16073
rect 4526 16039 4560 16073
rect 4594 16039 4628 16073
rect 4662 16039 4696 16073
rect 4730 16039 4764 16073
rect 4798 16039 4832 16073
rect 4866 16039 4900 16073
rect 4934 16039 4968 16073
rect 5002 16039 5036 16073
rect 5070 16039 5104 16073
rect 5138 16039 5172 16073
rect 5206 16039 5240 16073
rect 5274 16039 5308 16073
rect 5342 16039 5376 16073
rect 5410 16039 5444 16073
rect 5478 16039 5512 16073
rect 5546 16039 5580 16073
rect 5614 16039 5648 16073
rect 5682 16039 5716 16073
rect 5750 16039 5784 16073
rect 5818 16039 5852 16073
rect 5886 16039 5920 16073
rect 5954 16039 5988 16073
rect 6022 16039 6056 16073
rect 6090 16039 6124 16073
rect 6158 16039 6192 16073
rect 6226 16039 6260 16073
rect 6294 16039 6328 16073
rect 6362 16039 6396 16073
rect 6430 16039 6464 16073
rect 6498 16039 6532 16073
rect 6566 16039 6600 16073
rect 6634 16039 6668 16073
rect 6702 16039 6736 16073
rect 6770 16039 6804 16073
rect 6838 16039 6872 16073
rect 6906 16039 6940 16073
rect 6974 16039 7008 16073
rect 7042 16039 7076 16073
rect 7110 16039 7144 16073
rect 7178 16039 7212 16073
rect 7246 16039 7280 16073
rect 7314 16039 7348 16073
rect 7382 16039 7416 16073
rect 7450 16039 7484 16073
rect 7518 16039 7552 16073
rect 7586 16039 7620 16073
rect 7654 16039 7688 16073
rect 7722 16039 7756 16073
rect 7790 16039 7824 16073
rect 7858 16039 7892 16073
rect 7926 16039 7960 16073
rect 7994 16039 8028 16073
rect 8062 16039 8096 16073
rect 8130 16039 8164 16073
rect 8198 16039 8232 16073
rect 8266 16039 8300 16073
rect 8334 16039 8368 16073
rect 8402 16039 8436 16073
rect 8470 16039 8504 16073
rect 8538 16039 8572 16073
rect 8606 16039 8640 16073
rect 8674 16039 8708 16073
rect 8742 16039 8776 16073
rect 8810 16039 8844 16073
rect 8878 16039 8912 16073
rect 8946 16039 8980 16073
rect 9014 16039 9048 16073
rect 9082 16039 9116 16073
rect 9150 16039 9184 16073
rect 9218 16039 9252 16073
rect 9286 16039 9320 16073
rect 9354 16039 9388 16073
rect 9422 16039 9456 16073
rect 9490 16039 9524 16073
rect 9558 16039 9592 16073
rect 9626 16039 9660 16073
rect 9694 16039 9728 16073
rect 9762 16039 9796 16073
rect 9830 16039 9864 16073
rect 9898 16039 9932 16073
rect 9966 16039 10000 16073
rect 10034 16039 10068 16073
rect 10102 16039 10136 16073
rect 10170 16039 10204 16073
rect 10238 16039 10272 16073
rect 10306 16039 10340 16073
rect 10374 16039 10408 16073
rect 10442 16039 10476 16073
rect 10510 16039 10544 16073
rect 10578 16039 10612 16073
rect 10646 16039 10680 16073
rect 10714 16039 10748 16073
rect 10782 16039 10816 16073
rect 10850 16039 10884 16073
rect 10918 16039 10952 16073
rect 10986 16039 11020 16073
rect 11054 16039 11088 16073
rect 11122 16039 11156 16073
rect 11190 16039 11224 16073
rect 11258 16039 11292 16073
rect 11326 16039 11360 16073
rect 11394 16039 11428 16073
rect 11462 16039 11496 16073
rect 11530 16039 11564 16073
rect 11598 16039 11632 16073
rect 11666 16039 11700 16073
rect 11734 16039 11768 16073
rect 11802 16039 11836 16073
rect 11870 16039 11904 16073
rect 11938 16039 11972 16073
rect 12006 16039 12040 16073
rect 12074 16039 12108 16073
rect 12142 16039 12176 16073
rect 12210 16039 12244 16073
rect 12278 16039 12312 16073
rect 12346 16039 12380 16073
rect 12414 16039 12448 16073
rect 12482 16039 12516 16073
rect 12550 16039 12584 16073
rect 12618 16039 12652 16073
rect 12686 16039 12720 16073
rect 12754 16039 12788 16073
rect 12822 16039 12856 16073
rect 12890 16039 12924 16073
rect 12958 16039 12992 16073
rect 13026 16039 13060 16073
rect 13094 16039 13128 16073
rect 13162 16039 13196 16073
rect 13230 16039 13264 16073
rect 13298 16039 13332 16073
rect 13366 16039 13400 16073
rect 13434 16039 13468 16073
rect 13502 16039 13536 16073
rect 13570 16039 13604 16073
rect 13638 16039 13672 16073
rect 13706 16039 13740 16073
rect 13774 16039 13808 16073
rect 13842 16039 13876 16073
rect 13910 16039 13944 16073
rect 13978 16039 14012 16073
rect 14046 16039 14080 16073
rect 14114 16039 14148 16073
rect 14182 16039 14216 16073
rect 14250 16039 14284 16073
rect 14318 16039 14352 16073
rect 14386 16055 14420 16073
rect 14454 16055 14492 16089
rect 14526 16055 14564 16089
rect 14598 16055 14636 16089
rect 14670 16055 14708 16089
rect 14742 16055 14780 16089
rect 14814 16055 14852 16089
rect 14886 16055 14924 16089
rect 14958 16055 14996 16089
rect 15030 16055 15068 16089
rect 15102 16055 15106 16089
rect 14386 16039 15106 16055
rect 67 16020 15106 16039
rect 67 16017 14420 16020
rect 67 15983 68 16017
rect 102 15983 139 16017
rect 173 15983 210 16017
rect 244 15983 281 16017
rect 315 15983 352 16017
rect 386 16003 14420 16017
rect 386 15983 444 16003
rect 67 15969 444 15983
rect 478 15969 513 16003
rect 547 15969 582 16003
rect 616 15969 651 16003
rect 685 15969 720 16003
rect 754 15969 789 16003
rect 823 15969 858 16003
rect 892 15969 927 16003
rect 961 15969 996 16003
rect 1030 15969 1065 16003
rect 1099 15969 1134 16003
rect 1168 15969 1203 16003
rect 1237 15969 1272 16003
rect 1306 15969 1341 16003
rect 1375 15969 1410 16003
rect 1444 15969 1479 16003
rect 1513 15969 1548 16003
rect 1582 15969 1617 16003
rect 1651 15969 1686 16003
rect 1720 15969 1755 16003
rect 1789 15969 1824 16003
rect 1858 15969 1893 16003
rect 1927 15969 1962 16003
rect 1996 15969 2031 16003
rect 2065 15969 2100 16003
rect 2134 15969 2169 16003
rect 2203 15969 2238 16003
rect 2272 15969 2307 16003
rect 2341 15969 2376 16003
rect 2410 15969 2445 16003
rect 2479 15969 2514 16003
rect 2548 15969 2583 16003
rect 2617 15969 2652 16003
rect 2686 15969 2721 16003
rect 2755 15969 2790 16003
rect 2824 15969 2859 16003
rect 2893 15969 2928 16003
rect 2962 15969 2996 16003
rect 3030 15969 3064 16003
rect 3098 15969 3132 16003
rect 3166 15969 3200 16003
rect 3234 15969 3268 16003
rect 3302 15969 3336 16003
rect 3370 15969 3404 16003
rect 3438 15969 3472 16003
rect 3506 15969 3540 16003
rect 3574 15969 3608 16003
rect 3642 15969 3676 16003
rect 3710 15969 3744 16003
rect 3778 15969 3812 16003
rect 3846 15969 3880 16003
rect 3914 15969 3948 16003
rect 3982 15969 4016 16003
rect 4050 15969 4084 16003
rect 4118 15969 4152 16003
rect 4186 15969 4220 16003
rect 4254 15969 4288 16003
rect 4322 15969 4356 16003
rect 4390 15969 4424 16003
rect 4458 15969 4492 16003
rect 4526 15969 4560 16003
rect 4594 15969 4628 16003
rect 4662 15969 4696 16003
rect 4730 15969 4764 16003
rect 4798 15969 4832 16003
rect 4866 15969 4900 16003
rect 4934 15969 4968 16003
rect 5002 15969 5036 16003
rect 5070 15969 5104 16003
rect 5138 15969 5172 16003
rect 5206 15969 5240 16003
rect 5274 15969 5308 16003
rect 5342 15969 5376 16003
rect 5410 15969 5444 16003
rect 5478 15969 5512 16003
rect 5546 15969 5580 16003
rect 5614 15969 5648 16003
rect 5682 15969 5716 16003
rect 5750 15969 5784 16003
rect 5818 15969 5852 16003
rect 5886 15969 5920 16003
rect 5954 15969 5988 16003
rect 6022 15969 6056 16003
rect 6090 15969 6124 16003
rect 6158 15969 6192 16003
rect 6226 15969 6260 16003
rect 6294 15969 6328 16003
rect 6362 15969 6396 16003
rect 6430 15969 6464 16003
rect 6498 15969 6532 16003
rect 6566 15969 6600 16003
rect 6634 15969 6668 16003
rect 6702 15969 6736 16003
rect 6770 15969 6804 16003
rect 6838 15969 6872 16003
rect 6906 15969 6940 16003
rect 6974 15969 7008 16003
rect 7042 15969 7076 16003
rect 7110 15969 7144 16003
rect 7178 15969 7212 16003
rect 7246 15969 7280 16003
rect 7314 15969 7348 16003
rect 7382 15969 7416 16003
rect 7450 15969 7484 16003
rect 7518 15969 7552 16003
rect 7586 15969 7620 16003
rect 7654 15969 7688 16003
rect 7722 15969 7756 16003
rect 7790 15969 7824 16003
rect 7858 15969 7892 16003
rect 7926 15969 7960 16003
rect 7994 15969 8028 16003
rect 8062 15969 8096 16003
rect 8130 15969 8164 16003
rect 8198 15969 8232 16003
rect 8266 15969 8300 16003
rect 8334 15969 8368 16003
rect 8402 15969 8436 16003
rect 8470 15969 8504 16003
rect 8538 15969 8572 16003
rect 8606 15969 8640 16003
rect 8674 15969 8708 16003
rect 8742 15969 8776 16003
rect 8810 15969 8844 16003
rect 8878 15969 8912 16003
rect 8946 15969 8980 16003
rect 9014 15969 9048 16003
rect 9082 15969 9116 16003
rect 9150 15969 9184 16003
rect 9218 15969 9252 16003
rect 9286 15969 9320 16003
rect 9354 15969 9388 16003
rect 9422 15969 9456 16003
rect 9490 15969 9524 16003
rect 9558 15969 9592 16003
rect 9626 15969 9660 16003
rect 9694 15969 9728 16003
rect 9762 15969 9796 16003
rect 9830 15969 9864 16003
rect 9898 15969 9932 16003
rect 9966 15969 10000 16003
rect 10034 15969 10068 16003
rect 10102 15969 10136 16003
rect 10170 15969 10204 16003
rect 10238 15969 10272 16003
rect 10306 15969 10340 16003
rect 10374 15969 10408 16003
rect 10442 15969 10476 16003
rect 10510 15969 10544 16003
rect 10578 15969 10612 16003
rect 10646 15969 10680 16003
rect 10714 15969 10748 16003
rect 10782 15969 10816 16003
rect 10850 15969 10884 16003
rect 10918 15969 10952 16003
rect 10986 15969 11020 16003
rect 11054 15969 11088 16003
rect 11122 15969 11156 16003
rect 11190 15969 11224 16003
rect 11258 15969 11292 16003
rect 11326 15969 11360 16003
rect 11394 15969 11428 16003
rect 11462 15969 11496 16003
rect 11530 15969 11564 16003
rect 11598 15969 11632 16003
rect 11666 15969 11700 16003
rect 11734 15969 11768 16003
rect 11802 15969 11836 16003
rect 11870 15969 11904 16003
rect 11938 15969 11972 16003
rect 12006 15969 12040 16003
rect 12074 15969 12108 16003
rect 12142 15969 12176 16003
rect 12210 15969 12244 16003
rect 12278 15969 12312 16003
rect 12346 15969 12380 16003
rect 12414 15969 12448 16003
rect 12482 15969 12516 16003
rect 12550 15969 12584 16003
rect 12618 15969 12652 16003
rect 12686 15969 12720 16003
rect 12754 15969 12788 16003
rect 12822 15969 12856 16003
rect 12890 15969 12924 16003
rect 12958 15969 12992 16003
rect 13026 15969 13060 16003
rect 13094 15969 13128 16003
rect 13162 15969 13196 16003
rect 13230 15969 13264 16003
rect 13298 15969 13332 16003
rect 13366 15969 13400 16003
rect 13434 15969 13468 16003
rect 13502 15969 13536 16003
rect 13570 15969 13604 16003
rect 13638 15969 13672 16003
rect 13706 15969 13740 16003
rect 13774 15969 13808 16003
rect 13842 15969 13876 16003
rect 13910 15969 13944 16003
rect 13978 15969 14012 16003
rect 14046 15969 14080 16003
rect 14114 15969 14148 16003
rect 14182 15969 14216 16003
rect 14250 15969 14284 16003
rect 14318 15969 14352 16003
rect 14386 15986 14420 16003
rect 14454 15986 14492 16020
rect 14526 15986 14564 16020
rect 14598 15986 14636 16020
rect 14670 15986 14708 16020
rect 14742 15986 14780 16020
rect 14814 15986 14852 16020
rect 14886 15986 14924 16020
rect 14958 15986 14996 16020
rect 15030 15986 15068 16020
rect 15102 15986 15106 16020
rect 14386 15969 15106 15986
rect 67 15951 15106 15969
rect 67 15949 14420 15951
rect 67 15915 68 15949
rect 102 15915 139 15949
rect 173 15915 210 15949
rect 244 15915 281 15949
rect 315 15915 352 15949
rect 386 15933 14420 15949
rect 386 15915 444 15933
rect 67 15899 444 15915
rect 478 15899 513 15933
rect 547 15899 582 15933
rect 616 15899 651 15933
rect 685 15899 720 15933
rect 754 15899 789 15933
rect 823 15899 858 15933
rect 892 15899 927 15933
rect 961 15899 996 15933
rect 1030 15899 1065 15933
rect 1099 15899 1134 15933
rect 1168 15899 1203 15933
rect 1237 15899 1272 15933
rect 1306 15899 1341 15933
rect 1375 15899 1410 15933
rect 1444 15899 1479 15933
rect 1513 15899 1548 15933
rect 1582 15899 1617 15933
rect 1651 15899 1686 15933
rect 1720 15899 1755 15933
rect 1789 15899 1824 15933
rect 1858 15899 1893 15933
rect 1927 15899 1962 15933
rect 1996 15899 2031 15933
rect 2065 15899 2100 15933
rect 2134 15899 2169 15933
rect 2203 15899 2238 15933
rect 2272 15899 2307 15933
rect 2341 15899 2376 15933
rect 2410 15899 2445 15933
rect 2479 15899 2514 15933
rect 2548 15899 2583 15933
rect 2617 15899 2652 15933
rect 2686 15899 2721 15933
rect 2755 15899 2790 15933
rect 2824 15899 2859 15933
rect 2893 15899 2928 15933
rect 2962 15899 2996 15933
rect 3030 15899 3064 15933
rect 3098 15899 3132 15933
rect 3166 15899 3200 15933
rect 3234 15899 3268 15933
rect 3302 15899 3336 15933
rect 3370 15899 3404 15933
rect 3438 15899 3472 15933
rect 3506 15899 3540 15933
rect 3574 15899 3608 15933
rect 3642 15899 3676 15933
rect 3710 15899 3744 15933
rect 3778 15899 3812 15933
rect 3846 15899 3880 15933
rect 3914 15899 3948 15933
rect 3982 15899 4016 15933
rect 4050 15899 4084 15933
rect 4118 15899 4152 15933
rect 4186 15899 4220 15933
rect 4254 15899 4288 15933
rect 4322 15899 4356 15933
rect 4390 15899 4424 15933
rect 4458 15899 4492 15933
rect 4526 15899 4560 15933
rect 4594 15899 4628 15933
rect 4662 15899 4696 15933
rect 4730 15899 4764 15933
rect 4798 15899 4832 15933
rect 4866 15899 4900 15933
rect 4934 15899 4968 15933
rect 5002 15899 5036 15933
rect 5070 15899 5104 15933
rect 5138 15899 5172 15933
rect 5206 15899 5240 15933
rect 5274 15899 5308 15933
rect 5342 15899 5376 15933
rect 5410 15899 5444 15933
rect 5478 15899 5512 15933
rect 5546 15899 5580 15933
rect 5614 15899 5648 15933
rect 5682 15899 5716 15933
rect 5750 15899 5784 15933
rect 5818 15899 5852 15933
rect 5886 15899 5920 15933
rect 5954 15899 5988 15933
rect 6022 15899 6056 15933
rect 6090 15899 6124 15933
rect 6158 15899 6192 15933
rect 6226 15899 6260 15933
rect 6294 15899 6328 15933
rect 6362 15899 6396 15933
rect 6430 15899 6464 15933
rect 6498 15899 6532 15933
rect 6566 15899 6600 15933
rect 6634 15899 6668 15933
rect 6702 15899 6736 15933
rect 6770 15899 6804 15933
rect 6838 15899 6872 15933
rect 6906 15899 6940 15933
rect 6974 15899 7008 15933
rect 7042 15899 7076 15933
rect 7110 15899 7144 15933
rect 7178 15899 7212 15933
rect 7246 15899 7280 15933
rect 7314 15899 7348 15933
rect 7382 15899 7416 15933
rect 7450 15899 7484 15933
rect 7518 15899 7552 15933
rect 7586 15899 7620 15933
rect 7654 15899 7688 15933
rect 7722 15899 7756 15933
rect 7790 15899 7824 15933
rect 7858 15899 7892 15933
rect 7926 15899 7960 15933
rect 7994 15899 8028 15933
rect 8062 15899 8096 15933
rect 8130 15899 8164 15933
rect 8198 15899 8232 15933
rect 8266 15899 8300 15933
rect 8334 15899 8368 15933
rect 8402 15899 8436 15933
rect 8470 15899 8504 15933
rect 8538 15899 8572 15933
rect 8606 15899 8640 15933
rect 8674 15899 8708 15933
rect 8742 15899 8776 15933
rect 8810 15899 8844 15933
rect 8878 15899 8912 15933
rect 8946 15899 8980 15933
rect 9014 15899 9048 15933
rect 9082 15899 9116 15933
rect 9150 15899 9184 15933
rect 9218 15899 9252 15933
rect 9286 15899 9320 15933
rect 9354 15899 9388 15933
rect 9422 15899 9456 15933
rect 9490 15899 9524 15933
rect 9558 15899 9592 15933
rect 9626 15899 9660 15933
rect 9694 15899 9728 15933
rect 9762 15899 9796 15933
rect 9830 15899 9864 15933
rect 9898 15899 9932 15933
rect 9966 15899 10000 15933
rect 10034 15899 10068 15933
rect 10102 15899 10136 15933
rect 10170 15899 10204 15933
rect 10238 15899 10272 15933
rect 10306 15899 10340 15933
rect 10374 15899 10408 15933
rect 10442 15899 10476 15933
rect 10510 15899 10544 15933
rect 10578 15899 10612 15933
rect 10646 15899 10680 15933
rect 10714 15899 10748 15933
rect 10782 15899 10816 15933
rect 10850 15899 10884 15933
rect 10918 15899 10952 15933
rect 10986 15899 11020 15933
rect 11054 15899 11088 15933
rect 11122 15899 11156 15933
rect 11190 15899 11224 15933
rect 11258 15899 11292 15933
rect 11326 15899 11360 15933
rect 11394 15899 11428 15933
rect 11462 15899 11496 15933
rect 11530 15899 11564 15933
rect 11598 15899 11632 15933
rect 11666 15899 11700 15933
rect 11734 15899 11768 15933
rect 11802 15899 11836 15933
rect 11870 15899 11904 15933
rect 11938 15899 11972 15933
rect 12006 15899 12040 15933
rect 12074 15899 12108 15933
rect 12142 15899 12176 15933
rect 12210 15899 12244 15933
rect 12278 15899 12312 15933
rect 12346 15899 12380 15933
rect 12414 15899 12448 15933
rect 12482 15899 12516 15933
rect 12550 15899 12584 15933
rect 12618 15899 12652 15933
rect 12686 15899 12720 15933
rect 12754 15899 12788 15933
rect 12822 15899 12856 15933
rect 12890 15899 12924 15933
rect 12958 15899 12992 15933
rect 13026 15899 13060 15933
rect 13094 15899 13128 15933
rect 13162 15899 13196 15933
rect 13230 15899 13264 15933
rect 13298 15899 13332 15933
rect 13366 15899 13400 15933
rect 13434 15899 13468 15933
rect 13502 15899 13536 15933
rect 13570 15899 13604 15933
rect 13638 15899 13672 15933
rect 13706 15899 13740 15933
rect 13774 15899 13808 15933
rect 13842 15899 13876 15933
rect 13910 15899 13944 15933
rect 13978 15899 14012 15933
rect 14046 15899 14080 15933
rect 14114 15899 14148 15933
rect 14182 15899 14216 15933
rect 14250 15899 14284 15933
rect 14318 15899 14352 15933
rect 14386 15917 14420 15933
rect 14454 15917 14492 15951
rect 14526 15917 14564 15951
rect 14598 15917 14636 15951
rect 14670 15917 14708 15951
rect 14742 15917 14780 15951
rect 14814 15917 14852 15951
rect 14886 15917 14924 15951
rect 14958 15917 14996 15951
rect 15030 15917 15068 15951
rect 15102 15917 15106 15951
rect 14386 15899 15106 15917
rect 67 15882 15106 15899
rect 67 15880 14420 15882
rect 67 15846 68 15880
rect 102 15846 139 15880
rect 173 15846 210 15880
rect 244 15846 281 15880
rect 315 15846 352 15880
rect 386 15863 14420 15880
rect 386 15846 444 15863
rect 67 15829 444 15846
rect 478 15829 513 15863
rect 547 15829 582 15863
rect 616 15829 651 15863
rect 685 15829 720 15863
rect 754 15829 789 15863
rect 823 15829 858 15863
rect 892 15829 927 15863
rect 961 15829 996 15863
rect 1030 15829 1065 15863
rect 1099 15829 1134 15863
rect 1168 15829 1203 15863
rect 1237 15829 1272 15863
rect 1306 15829 1341 15863
rect 1375 15829 1410 15863
rect 1444 15829 1479 15863
rect 1513 15829 1548 15863
rect 1582 15829 1617 15863
rect 1651 15829 1686 15863
rect 1720 15829 1755 15863
rect 1789 15829 1824 15863
rect 1858 15829 1893 15863
rect 1927 15829 1962 15863
rect 1996 15829 2031 15863
rect 2065 15829 2100 15863
rect 2134 15829 2169 15863
rect 2203 15829 2238 15863
rect 2272 15829 2307 15863
rect 2341 15829 2376 15863
rect 2410 15829 2445 15863
rect 2479 15829 2514 15863
rect 2548 15829 2583 15863
rect 2617 15829 2652 15863
rect 2686 15829 2721 15863
rect 2755 15829 2790 15863
rect 2824 15829 2859 15863
rect 2893 15829 2928 15863
rect 2962 15829 2996 15863
rect 3030 15829 3064 15863
rect 3098 15829 3132 15863
rect 3166 15829 3200 15863
rect 3234 15829 3268 15863
rect 3302 15829 3336 15863
rect 3370 15829 3404 15863
rect 3438 15829 3472 15863
rect 3506 15829 3540 15863
rect 3574 15829 3608 15863
rect 3642 15829 3676 15863
rect 3710 15829 3744 15863
rect 3778 15829 3812 15863
rect 3846 15829 3880 15863
rect 3914 15829 3948 15863
rect 3982 15829 4016 15863
rect 4050 15829 4084 15863
rect 4118 15829 4152 15863
rect 4186 15829 4220 15863
rect 4254 15829 4288 15863
rect 4322 15829 4356 15863
rect 4390 15829 4424 15863
rect 4458 15829 4492 15863
rect 4526 15829 4560 15863
rect 4594 15829 4628 15863
rect 4662 15829 4696 15863
rect 4730 15829 4764 15863
rect 4798 15829 4832 15863
rect 4866 15829 4900 15863
rect 4934 15829 4968 15863
rect 5002 15829 5036 15863
rect 5070 15829 5104 15863
rect 5138 15829 5172 15863
rect 5206 15829 5240 15863
rect 5274 15829 5308 15863
rect 5342 15829 5376 15863
rect 5410 15829 5444 15863
rect 5478 15829 5512 15863
rect 5546 15829 5580 15863
rect 5614 15829 5648 15863
rect 5682 15829 5716 15863
rect 5750 15829 5784 15863
rect 5818 15829 5852 15863
rect 5886 15829 5920 15863
rect 5954 15829 5988 15863
rect 6022 15829 6056 15863
rect 6090 15829 6124 15863
rect 6158 15829 6192 15863
rect 6226 15829 6260 15863
rect 6294 15829 6328 15863
rect 6362 15829 6396 15863
rect 6430 15829 6464 15863
rect 6498 15829 6532 15863
rect 6566 15829 6600 15863
rect 6634 15829 6668 15863
rect 6702 15829 6736 15863
rect 6770 15829 6804 15863
rect 6838 15829 6872 15863
rect 6906 15829 6940 15863
rect 6974 15829 7008 15863
rect 7042 15829 7076 15863
rect 7110 15829 7144 15863
rect 7178 15829 7212 15863
rect 7246 15829 7280 15863
rect 7314 15829 7348 15863
rect 7382 15829 7416 15863
rect 7450 15829 7484 15863
rect 7518 15829 7552 15863
rect 7586 15829 7620 15863
rect 7654 15829 7688 15863
rect 7722 15829 7756 15863
rect 7790 15829 7824 15863
rect 7858 15829 7892 15863
rect 7926 15829 7960 15863
rect 7994 15829 8028 15863
rect 8062 15829 8096 15863
rect 8130 15829 8164 15863
rect 8198 15829 8232 15863
rect 8266 15829 8300 15863
rect 8334 15829 8368 15863
rect 8402 15829 8436 15863
rect 8470 15829 8504 15863
rect 8538 15829 8572 15863
rect 8606 15829 8640 15863
rect 8674 15829 8708 15863
rect 8742 15829 8776 15863
rect 8810 15829 8844 15863
rect 8878 15829 8912 15863
rect 8946 15829 8980 15863
rect 9014 15829 9048 15863
rect 9082 15829 9116 15863
rect 9150 15829 9184 15863
rect 9218 15829 9252 15863
rect 9286 15829 9320 15863
rect 9354 15829 9388 15863
rect 9422 15829 9456 15863
rect 9490 15829 9524 15863
rect 9558 15829 9592 15863
rect 9626 15829 9660 15863
rect 9694 15829 9728 15863
rect 9762 15829 9796 15863
rect 9830 15829 9864 15863
rect 9898 15829 9932 15863
rect 9966 15829 10000 15863
rect 10034 15829 10068 15863
rect 10102 15829 10136 15863
rect 10170 15829 10204 15863
rect 10238 15829 10272 15863
rect 10306 15829 10340 15863
rect 10374 15829 10408 15863
rect 10442 15829 10476 15863
rect 10510 15829 10544 15863
rect 10578 15829 10612 15863
rect 10646 15829 10680 15863
rect 10714 15829 10748 15863
rect 10782 15829 10816 15863
rect 10850 15829 10884 15863
rect 10918 15829 10952 15863
rect 10986 15829 11020 15863
rect 11054 15829 11088 15863
rect 11122 15829 11156 15863
rect 11190 15829 11224 15863
rect 11258 15829 11292 15863
rect 11326 15829 11360 15863
rect 11394 15829 11428 15863
rect 11462 15829 11496 15863
rect 11530 15829 11564 15863
rect 11598 15829 11632 15863
rect 11666 15829 11700 15863
rect 11734 15829 11768 15863
rect 11802 15829 11836 15863
rect 11870 15829 11904 15863
rect 11938 15829 11972 15863
rect 12006 15829 12040 15863
rect 12074 15829 12108 15863
rect 12142 15829 12176 15863
rect 12210 15829 12244 15863
rect 12278 15829 12312 15863
rect 12346 15829 12380 15863
rect 12414 15829 12448 15863
rect 12482 15829 12516 15863
rect 12550 15829 12584 15863
rect 12618 15829 12652 15863
rect 12686 15829 12720 15863
rect 12754 15829 12788 15863
rect 12822 15829 12856 15863
rect 12890 15829 12924 15863
rect 12958 15829 12992 15863
rect 13026 15829 13060 15863
rect 13094 15829 13128 15863
rect 13162 15829 13196 15863
rect 13230 15829 13264 15863
rect 13298 15829 13332 15863
rect 13366 15829 13400 15863
rect 13434 15829 13468 15863
rect 13502 15829 13536 15863
rect 13570 15829 13604 15863
rect 13638 15829 13672 15863
rect 13706 15829 13740 15863
rect 13774 15829 13808 15863
rect 13842 15829 13876 15863
rect 13910 15829 13944 15863
rect 13978 15829 14012 15863
rect 14046 15829 14080 15863
rect 14114 15829 14148 15863
rect 14182 15829 14216 15863
rect 14250 15829 14284 15863
rect 14318 15829 14352 15863
rect 14386 15848 14420 15863
rect 14454 15848 14492 15882
rect 14526 15848 14564 15882
rect 14598 15848 14636 15882
rect 14670 15848 14708 15882
rect 14742 15848 14780 15882
rect 14814 15848 14852 15882
rect 14886 15848 14924 15882
rect 14958 15848 14996 15882
rect 15030 15848 15068 15882
rect 15102 15848 15106 15882
rect 14386 15829 15106 15848
rect 67 15813 15106 15829
rect 67 15811 14420 15813
rect 67 15777 68 15811
rect 102 15777 139 15811
rect 173 15777 210 15811
rect 244 15777 281 15811
rect 315 15777 352 15811
rect 386 15793 14420 15811
rect 386 15777 444 15793
rect 67 15759 444 15777
rect 478 15759 513 15793
rect 547 15759 582 15793
rect 616 15759 651 15793
rect 685 15759 720 15793
rect 754 15759 789 15793
rect 823 15759 858 15793
rect 892 15759 927 15793
rect 961 15759 996 15793
rect 1030 15759 1065 15793
rect 1099 15759 1134 15793
rect 1168 15759 1203 15793
rect 1237 15759 1272 15793
rect 1306 15759 1341 15793
rect 1375 15759 1410 15793
rect 1444 15759 1479 15793
rect 1513 15759 1548 15793
rect 1582 15759 1617 15793
rect 1651 15759 1686 15793
rect 1720 15759 1755 15793
rect 1789 15759 1824 15793
rect 1858 15759 1893 15793
rect 1927 15759 1962 15793
rect 1996 15759 2031 15793
rect 2065 15759 2100 15793
rect 2134 15759 2169 15793
rect 2203 15759 2238 15793
rect 2272 15759 2307 15793
rect 2341 15759 2376 15793
rect 2410 15759 2445 15793
rect 2479 15759 2514 15793
rect 2548 15759 2583 15793
rect 2617 15759 2652 15793
rect 2686 15759 2721 15793
rect 2755 15759 2790 15793
rect 2824 15759 2859 15793
rect 2893 15759 2928 15793
rect 2962 15759 2996 15793
rect 3030 15759 3064 15793
rect 3098 15759 3132 15793
rect 3166 15759 3200 15793
rect 3234 15759 3268 15793
rect 3302 15759 3336 15793
rect 3370 15759 3404 15793
rect 3438 15759 3472 15793
rect 3506 15759 3540 15793
rect 3574 15759 3608 15793
rect 3642 15759 3676 15793
rect 3710 15759 3744 15793
rect 3778 15759 3812 15793
rect 3846 15759 3880 15793
rect 3914 15759 3948 15793
rect 3982 15759 4016 15793
rect 4050 15759 4084 15793
rect 4118 15759 4152 15793
rect 4186 15759 4220 15793
rect 4254 15759 4288 15793
rect 4322 15759 4356 15793
rect 4390 15759 4424 15793
rect 4458 15759 4492 15793
rect 4526 15759 4560 15793
rect 4594 15759 4628 15793
rect 4662 15759 4696 15793
rect 4730 15759 4764 15793
rect 4798 15759 4832 15793
rect 4866 15759 4900 15793
rect 4934 15759 4968 15793
rect 5002 15759 5036 15793
rect 5070 15759 5104 15793
rect 5138 15759 5172 15793
rect 5206 15759 5240 15793
rect 5274 15759 5308 15793
rect 5342 15759 5376 15793
rect 5410 15759 5444 15793
rect 5478 15759 5512 15793
rect 5546 15759 5580 15793
rect 5614 15759 5648 15793
rect 5682 15759 5716 15793
rect 5750 15759 5784 15793
rect 5818 15759 5852 15793
rect 5886 15759 5920 15793
rect 5954 15759 5988 15793
rect 6022 15759 6056 15793
rect 6090 15759 6124 15793
rect 6158 15759 6192 15793
rect 6226 15759 6260 15793
rect 6294 15759 6328 15793
rect 6362 15759 6396 15793
rect 6430 15759 6464 15793
rect 6498 15759 6532 15793
rect 6566 15759 6600 15793
rect 6634 15759 6668 15793
rect 6702 15759 6736 15793
rect 6770 15759 6804 15793
rect 6838 15759 6872 15793
rect 6906 15759 6940 15793
rect 6974 15759 7008 15793
rect 7042 15759 7076 15793
rect 7110 15759 7144 15793
rect 7178 15759 7212 15793
rect 7246 15759 7280 15793
rect 7314 15759 7348 15793
rect 7382 15759 7416 15793
rect 7450 15759 7484 15793
rect 7518 15759 7552 15793
rect 7586 15759 7620 15793
rect 7654 15759 7688 15793
rect 7722 15759 7756 15793
rect 7790 15759 7824 15793
rect 7858 15759 7892 15793
rect 7926 15759 7960 15793
rect 7994 15759 8028 15793
rect 8062 15759 8096 15793
rect 8130 15759 8164 15793
rect 8198 15759 8232 15793
rect 8266 15759 8300 15793
rect 8334 15759 8368 15793
rect 8402 15759 8436 15793
rect 8470 15759 8504 15793
rect 8538 15759 8572 15793
rect 8606 15759 8640 15793
rect 8674 15759 8708 15793
rect 8742 15759 8776 15793
rect 8810 15759 8844 15793
rect 8878 15759 8912 15793
rect 8946 15759 8980 15793
rect 9014 15759 9048 15793
rect 9082 15759 9116 15793
rect 9150 15759 9184 15793
rect 9218 15759 9252 15793
rect 9286 15759 9320 15793
rect 9354 15759 9388 15793
rect 9422 15759 9456 15793
rect 9490 15759 9524 15793
rect 9558 15759 9592 15793
rect 9626 15759 9660 15793
rect 9694 15759 9728 15793
rect 9762 15759 9796 15793
rect 9830 15759 9864 15793
rect 9898 15759 9932 15793
rect 9966 15759 10000 15793
rect 10034 15759 10068 15793
rect 10102 15759 10136 15793
rect 10170 15759 10204 15793
rect 10238 15759 10272 15793
rect 10306 15759 10340 15793
rect 10374 15759 10408 15793
rect 10442 15759 10476 15793
rect 10510 15759 10544 15793
rect 10578 15759 10612 15793
rect 10646 15759 10680 15793
rect 10714 15759 10748 15793
rect 10782 15759 10816 15793
rect 10850 15759 10884 15793
rect 10918 15759 10952 15793
rect 10986 15759 11020 15793
rect 11054 15759 11088 15793
rect 11122 15759 11156 15793
rect 11190 15759 11224 15793
rect 11258 15759 11292 15793
rect 11326 15759 11360 15793
rect 11394 15759 11428 15793
rect 11462 15759 11496 15793
rect 11530 15759 11564 15793
rect 11598 15759 11632 15793
rect 11666 15759 11700 15793
rect 11734 15759 11768 15793
rect 11802 15759 11836 15793
rect 11870 15759 11904 15793
rect 11938 15759 11972 15793
rect 12006 15759 12040 15793
rect 12074 15759 12108 15793
rect 12142 15759 12176 15793
rect 12210 15759 12244 15793
rect 12278 15759 12312 15793
rect 12346 15759 12380 15793
rect 12414 15759 12448 15793
rect 12482 15759 12516 15793
rect 12550 15759 12584 15793
rect 12618 15759 12652 15793
rect 12686 15759 12720 15793
rect 12754 15759 12788 15793
rect 12822 15759 12856 15793
rect 12890 15759 12924 15793
rect 12958 15759 12992 15793
rect 13026 15759 13060 15793
rect 13094 15759 13128 15793
rect 13162 15759 13196 15793
rect 13230 15759 13264 15793
rect 13298 15759 13332 15793
rect 13366 15759 13400 15793
rect 13434 15759 13468 15793
rect 13502 15759 13536 15793
rect 13570 15759 13604 15793
rect 13638 15759 13672 15793
rect 13706 15759 13740 15793
rect 13774 15759 13808 15793
rect 13842 15759 13876 15793
rect 13910 15759 13944 15793
rect 13978 15759 14012 15793
rect 14046 15759 14080 15793
rect 14114 15759 14148 15793
rect 14182 15759 14216 15793
rect 14250 15759 14284 15793
rect 14318 15759 14352 15793
rect 14386 15779 14420 15793
rect 14454 15779 14492 15813
rect 14526 15779 14564 15813
rect 14598 15779 14636 15813
rect 14670 15779 14708 15813
rect 14742 15779 14780 15813
rect 14814 15779 14852 15813
rect 14886 15779 14924 15813
rect 14958 15779 14996 15813
rect 15030 15779 15068 15813
rect 15102 15779 15106 15813
rect 14386 15759 15106 15779
rect 67 15744 15106 15759
rect 67 15742 14420 15744
rect 67 15708 68 15742
rect 102 15708 139 15742
rect 173 15708 210 15742
rect 244 15708 281 15742
rect 315 15708 352 15742
rect 386 15723 14420 15742
rect 386 15708 444 15723
rect 67 15689 444 15708
rect 478 15689 513 15723
rect 547 15689 582 15723
rect 616 15689 651 15723
rect 685 15689 720 15723
rect 754 15689 789 15723
rect 823 15689 858 15723
rect 892 15689 927 15723
rect 961 15689 996 15723
rect 1030 15689 1065 15723
rect 1099 15689 1134 15723
rect 1168 15689 1203 15723
rect 1237 15689 1272 15723
rect 1306 15689 1341 15723
rect 1375 15689 1410 15723
rect 1444 15689 1479 15723
rect 1513 15689 1548 15723
rect 1582 15689 1617 15723
rect 1651 15689 1686 15723
rect 1720 15689 1755 15723
rect 1789 15689 1824 15723
rect 1858 15689 1893 15723
rect 1927 15689 1962 15723
rect 1996 15689 2031 15723
rect 2065 15689 2100 15723
rect 2134 15689 2169 15723
rect 2203 15689 2238 15723
rect 2272 15689 2307 15723
rect 2341 15689 2376 15723
rect 2410 15689 2445 15723
rect 2479 15689 2514 15723
rect 2548 15689 2583 15723
rect 2617 15689 2652 15723
rect 2686 15689 2721 15723
rect 2755 15689 2790 15723
rect 2824 15689 2859 15723
rect 2893 15689 2928 15723
rect 2962 15689 2996 15723
rect 3030 15689 3064 15723
rect 3098 15689 3132 15723
rect 3166 15689 3200 15723
rect 3234 15689 3268 15723
rect 3302 15689 3336 15723
rect 3370 15689 3404 15723
rect 3438 15689 3472 15723
rect 3506 15689 3540 15723
rect 3574 15689 3608 15723
rect 3642 15689 3676 15723
rect 3710 15689 3744 15723
rect 3778 15689 3812 15723
rect 3846 15689 3880 15723
rect 3914 15689 3948 15723
rect 3982 15689 4016 15723
rect 4050 15689 4084 15723
rect 4118 15689 4152 15723
rect 4186 15689 4220 15723
rect 4254 15689 4288 15723
rect 4322 15689 4356 15723
rect 4390 15689 4424 15723
rect 4458 15689 4492 15723
rect 4526 15689 4560 15723
rect 4594 15689 4628 15723
rect 4662 15689 4696 15723
rect 4730 15689 4764 15723
rect 4798 15689 4832 15723
rect 4866 15689 4900 15723
rect 4934 15689 4968 15723
rect 5002 15689 5036 15723
rect 5070 15689 5104 15723
rect 5138 15689 5172 15723
rect 5206 15689 5240 15723
rect 5274 15689 5308 15723
rect 5342 15689 5376 15723
rect 5410 15689 5444 15723
rect 5478 15689 5512 15723
rect 5546 15689 5580 15723
rect 5614 15689 5648 15723
rect 5682 15689 5716 15723
rect 5750 15689 5784 15723
rect 5818 15689 5852 15723
rect 5886 15689 5920 15723
rect 5954 15689 5988 15723
rect 6022 15689 6056 15723
rect 6090 15689 6124 15723
rect 6158 15689 6192 15723
rect 6226 15689 6260 15723
rect 6294 15689 6328 15723
rect 6362 15689 6396 15723
rect 6430 15689 6464 15723
rect 6498 15689 6532 15723
rect 6566 15689 6600 15723
rect 6634 15689 6668 15723
rect 6702 15689 6736 15723
rect 6770 15689 6804 15723
rect 6838 15689 6872 15723
rect 6906 15689 6940 15723
rect 6974 15689 7008 15723
rect 7042 15689 7076 15723
rect 7110 15689 7144 15723
rect 7178 15689 7212 15723
rect 7246 15689 7280 15723
rect 7314 15689 7348 15723
rect 7382 15689 7416 15723
rect 7450 15689 7484 15723
rect 7518 15689 7552 15723
rect 7586 15689 7620 15723
rect 7654 15689 7688 15723
rect 7722 15689 7756 15723
rect 7790 15689 7824 15723
rect 7858 15689 7892 15723
rect 7926 15689 7960 15723
rect 7994 15689 8028 15723
rect 8062 15689 8096 15723
rect 8130 15689 8164 15723
rect 8198 15689 8232 15723
rect 8266 15689 8300 15723
rect 8334 15689 8368 15723
rect 8402 15689 8436 15723
rect 8470 15689 8504 15723
rect 8538 15689 8572 15723
rect 8606 15689 8640 15723
rect 8674 15689 8708 15723
rect 8742 15689 8776 15723
rect 8810 15689 8844 15723
rect 8878 15689 8912 15723
rect 8946 15689 8980 15723
rect 9014 15689 9048 15723
rect 9082 15689 9116 15723
rect 9150 15689 9184 15723
rect 9218 15689 9252 15723
rect 9286 15689 9320 15723
rect 9354 15689 9388 15723
rect 9422 15689 9456 15723
rect 9490 15689 9524 15723
rect 9558 15689 9592 15723
rect 9626 15689 9660 15723
rect 9694 15689 9728 15723
rect 9762 15689 9796 15723
rect 9830 15689 9864 15723
rect 9898 15689 9932 15723
rect 9966 15689 10000 15723
rect 10034 15689 10068 15723
rect 10102 15689 10136 15723
rect 10170 15689 10204 15723
rect 10238 15689 10272 15723
rect 10306 15689 10340 15723
rect 10374 15689 10408 15723
rect 10442 15689 10476 15723
rect 10510 15689 10544 15723
rect 10578 15689 10612 15723
rect 10646 15689 10680 15723
rect 10714 15689 10748 15723
rect 10782 15689 10816 15723
rect 10850 15689 10884 15723
rect 10918 15689 10952 15723
rect 10986 15689 11020 15723
rect 11054 15689 11088 15723
rect 11122 15689 11156 15723
rect 11190 15689 11224 15723
rect 11258 15689 11292 15723
rect 11326 15689 11360 15723
rect 11394 15689 11428 15723
rect 11462 15689 11496 15723
rect 11530 15689 11564 15723
rect 11598 15689 11632 15723
rect 11666 15689 11700 15723
rect 11734 15689 11768 15723
rect 11802 15689 11836 15723
rect 11870 15689 11904 15723
rect 11938 15689 11972 15723
rect 12006 15689 12040 15723
rect 12074 15689 12108 15723
rect 12142 15689 12176 15723
rect 12210 15689 12244 15723
rect 12278 15689 12312 15723
rect 12346 15689 12380 15723
rect 12414 15689 12448 15723
rect 12482 15689 12516 15723
rect 12550 15689 12584 15723
rect 12618 15689 12652 15723
rect 12686 15689 12720 15723
rect 12754 15689 12788 15723
rect 12822 15689 12856 15723
rect 12890 15689 12924 15723
rect 12958 15689 12992 15723
rect 13026 15689 13060 15723
rect 13094 15689 13128 15723
rect 13162 15689 13196 15723
rect 13230 15689 13264 15723
rect 13298 15689 13332 15723
rect 13366 15689 13400 15723
rect 13434 15689 13468 15723
rect 13502 15689 13536 15723
rect 13570 15689 13604 15723
rect 13638 15689 13672 15723
rect 13706 15689 13740 15723
rect 13774 15689 13808 15723
rect 13842 15689 13876 15723
rect 13910 15689 13944 15723
rect 13978 15689 14012 15723
rect 14046 15689 14080 15723
rect 14114 15689 14148 15723
rect 14182 15689 14216 15723
rect 14250 15689 14284 15723
rect 14318 15689 14352 15723
rect 14386 15710 14420 15723
rect 14454 15710 14492 15744
rect 14526 15710 14564 15744
rect 14598 15710 14636 15744
rect 14670 15710 14708 15744
rect 14742 15710 14780 15744
rect 14814 15710 14852 15744
rect 14886 15710 14924 15744
rect 14958 15710 14996 15744
rect 15030 15710 15068 15744
rect 15102 15710 15106 15744
rect 14386 15689 15106 15710
rect 67 15675 15106 15689
rect 67 15673 14420 15675
rect 67 15639 68 15673
rect 102 15639 139 15673
rect 173 15639 210 15673
rect 244 15639 281 15673
rect 315 15639 352 15673
rect 386 15651 14420 15673
rect 386 15639 12660 15651
rect 67 15617 12660 15639
rect 12694 15617 12730 15651
rect 12764 15617 12800 15651
rect 12834 15617 12869 15651
rect 12903 15617 12938 15651
rect 12972 15617 13007 15651
rect 13041 15617 13076 15651
rect 13110 15617 13145 15651
rect 13179 15617 13214 15651
rect 13248 15617 13283 15651
rect 13317 15617 13352 15651
rect 13386 15617 13421 15651
rect 13455 15617 13490 15651
rect 13524 15617 13559 15651
rect 13593 15617 13628 15651
rect 13662 15617 13697 15651
rect 13731 15617 13766 15651
rect 13800 15617 13835 15651
rect 13869 15617 13904 15651
rect 13938 15617 13973 15651
rect 14007 15617 14042 15651
rect 14076 15617 14111 15651
rect 14145 15617 14180 15651
rect 14214 15617 14249 15651
rect 14283 15617 14318 15651
rect 14352 15641 14420 15651
rect 14454 15641 14492 15675
rect 14526 15641 14564 15675
rect 14598 15641 14636 15675
rect 14670 15641 14708 15675
rect 14742 15641 14780 15675
rect 14814 15641 14852 15675
rect 14886 15641 14924 15675
rect 14958 15641 14996 15675
rect 15030 15641 15068 15675
rect 15102 15641 15106 15675
rect 14352 15617 15106 15641
rect 67 15607 15106 15617
rect 67 15604 594 15607
rect 67 15570 68 15604
rect 102 15570 139 15604
rect 173 15570 210 15604
rect 244 15570 281 15604
rect 315 15570 352 15604
rect 386 15583 594 15604
rect 386 15570 420 15583
rect 67 15549 420 15570
rect 454 15549 488 15583
rect 522 15573 594 15583
rect 628 15573 663 15607
rect 697 15573 732 15607
rect 766 15573 801 15607
rect 835 15573 870 15607
rect 904 15573 939 15607
rect 973 15573 1008 15607
rect 1042 15573 1077 15607
rect 1111 15573 1146 15607
rect 1180 15573 1215 15607
rect 1249 15573 1284 15607
rect 1318 15573 1353 15607
rect 1387 15573 1422 15607
rect 1456 15573 1491 15607
rect 1525 15573 1560 15607
rect 1594 15573 1629 15607
rect 1663 15573 1698 15607
rect 1732 15573 1767 15607
rect 1801 15573 1836 15607
rect 1870 15573 1904 15607
rect 1938 15573 1972 15607
rect 2006 15573 2040 15607
rect 2074 15573 2108 15607
rect 2142 15573 2176 15607
rect 2210 15573 2244 15607
rect 2278 15573 2312 15607
rect 2346 15573 2380 15607
rect 2414 15573 2448 15607
rect 2482 15573 2516 15607
rect 2550 15573 2584 15607
rect 2618 15573 2652 15607
rect 2686 15573 2720 15607
rect 2754 15573 2788 15607
rect 2822 15573 2856 15607
rect 2890 15573 2924 15607
rect 2958 15573 2992 15607
rect 3026 15573 3060 15607
rect 3094 15573 3128 15607
rect 3162 15573 3196 15607
rect 3230 15573 3264 15607
rect 3298 15573 3332 15607
rect 3366 15573 3400 15607
rect 3434 15573 3468 15607
rect 3502 15573 3536 15607
rect 3570 15573 3604 15607
rect 3638 15573 3672 15607
rect 3706 15573 3740 15607
rect 3774 15573 3808 15607
rect 3842 15573 3876 15607
rect 3910 15573 3944 15607
rect 3978 15573 4012 15607
rect 4046 15573 4080 15607
rect 4114 15573 4148 15607
rect 4182 15573 4216 15607
rect 4250 15573 4284 15607
rect 4318 15573 4352 15607
rect 4386 15573 4420 15607
rect 4454 15573 4488 15607
rect 4522 15573 4556 15607
rect 4590 15573 4624 15607
rect 4658 15573 4692 15607
rect 4726 15573 4760 15607
rect 4794 15573 4828 15607
rect 4862 15573 4896 15607
rect 4930 15573 4964 15607
rect 4998 15573 5032 15607
rect 5066 15573 5100 15607
rect 5134 15573 5168 15607
rect 5202 15573 5236 15607
rect 5270 15573 5304 15607
rect 5338 15573 5372 15607
rect 5406 15573 5430 15607
rect 67 15535 522 15549
rect 67 15501 68 15535
rect 102 15501 139 15535
rect 173 15501 210 15535
rect 244 15501 281 15535
rect 315 15501 352 15535
rect 386 15514 522 15535
rect 386 15501 420 15514
rect 67 15480 420 15501
rect 454 15480 488 15514
rect 67 15466 522 15480
rect 67 15432 68 15466
rect 102 15432 139 15466
rect 173 15432 210 15466
rect 244 15432 281 15466
rect 315 15432 352 15466
rect 386 15445 522 15466
rect 386 15432 420 15445
rect 67 15411 420 15432
rect 454 15411 488 15445
rect 67 15397 522 15411
rect 67 15363 68 15397
rect 102 15363 139 15397
rect 173 15363 210 15397
rect 244 15363 281 15397
rect 315 15363 352 15397
rect 386 15375 522 15397
rect 386 15363 420 15375
rect 67 15341 420 15363
rect 454 15341 488 15375
rect 67 15328 522 15341
rect 67 15294 68 15328
rect 102 15294 139 15328
rect 173 15294 210 15328
rect 244 15294 281 15328
rect 315 15294 352 15328
rect 386 15305 522 15328
rect 386 15294 420 15305
rect 67 15271 420 15294
rect 454 15271 488 15305
rect 67 15259 522 15271
rect 67 15225 68 15259
rect 102 15225 139 15259
rect 173 15225 210 15259
rect 244 15225 281 15259
rect 315 15225 352 15259
rect 386 15235 522 15259
rect 386 15225 420 15235
rect 67 15201 420 15225
rect 454 15201 488 15235
rect 67 15190 522 15201
rect 67 15156 68 15190
rect 102 15156 139 15190
rect 173 15156 210 15190
rect 244 15156 281 15190
rect 315 15156 352 15190
rect 386 15165 522 15190
rect 386 15156 420 15165
rect 67 15131 420 15156
rect 454 15131 488 15165
rect 67 15121 522 15131
rect 67 15087 68 15121
rect 102 15087 139 15121
rect 173 15087 210 15121
rect 244 15087 281 15121
rect 315 15087 352 15121
rect 386 15095 522 15121
rect 386 15087 420 15095
rect 67 15061 420 15087
rect 454 15061 488 15095
rect 67 15052 522 15061
rect 67 15018 68 15052
rect 102 15018 139 15052
rect 173 15018 210 15052
rect 244 15018 281 15052
rect 315 15018 352 15052
rect 386 15025 522 15052
rect 386 15018 420 15025
rect 67 14991 420 15018
rect 454 14991 488 15025
rect 67 14983 522 14991
rect 67 14949 68 14983
rect 102 14949 139 14983
rect 173 14949 210 14983
rect 244 14949 281 14983
rect 315 14949 352 14983
rect 386 14955 522 14983
rect 386 14949 420 14955
rect 67 14921 420 14949
rect 454 14921 488 14955
rect 67 14914 522 14921
rect 67 14880 68 14914
rect 102 14880 139 14914
rect 173 14880 210 14914
rect 244 14880 281 14914
rect 315 14880 352 14914
rect 386 14885 522 14914
rect 386 14880 420 14885
rect 67 14851 420 14880
rect 454 14851 488 14885
rect 67 14845 522 14851
rect 67 14811 68 14845
rect 102 14811 139 14845
rect 173 14811 210 14845
rect 244 14811 281 14845
rect 315 14811 352 14845
rect 386 14827 522 14845
rect 5396 14827 5430 15573
rect 386 14811 5430 14827
rect 67 14793 5430 14811
rect 12580 15606 15106 15607
rect 12580 15581 14420 15606
rect 12580 15547 12660 15581
rect 12694 15547 12730 15581
rect 12764 15547 12800 15581
rect 12834 15547 12869 15581
rect 12903 15547 12938 15581
rect 12972 15547 13007 15581
rect 13041 15547 13076 15581
rect 13110 15547 13145 15581
rect 13179 15547 13214 15581
rect 13248 15547 13283 15581
rect 13317 15547 13352 15581
rect 13386 15547 13421 15581
rect 13455 15547 13490 15581
rect 13524 15547 13559 15581
rect 13593 15547 13628 15581
rect 13662 15547 13697 15581
rect 13731 15547 13766 15581
rect 13800 15547 13835 15581
rect 13869 15547 13904 15581
rect 13938 15547 13973 15581
rect 14007 15547 14042 15581
rect 14076 15547 14111 15581
rect 14145 15547 14180 15581
rect 14214 15547 14249 15581
rect 14283 15547 14318 15581
rect 14352 15572 14420 15581
rect 14454 15572 14492 15606
rect 14526 15572 14564 15606
rect 14598 15572 14636 15606
rect 14670 15572 14708 15606
rect 14742 15572 14780 15606
rect 14814 15572 14852 15606
rect 14886 15572 14924 15606
rect 14958 15572 14996 15606
rect 15030 15572 15068 15606
rect 15102 15572 15106 15606
rect 14352 15547 15106 15572
rect 12580 15537 15106 15547
rect 12580 15511 14420 15537
rect 12580 15477 12660 15511
rect 12694 15477 12730 15511
rect 12764 15477 12800 15511
rect 12834 15477 12869 15511
rect 12903 15477 12938 15511
rect 12972 15477 13007 15511
rect 13041 15477 13076 15511
rect 13110 15477 13145 15511
rect 13179 15477 13214 15511
rect 13248 15477 13283 15511
rect 13317 15477 13352 15511
rect 13386 15477 13421 15511
rect 13455 15477 13490 15511
rect 13524 15477 13559 15511
rect 13593 15477 13628 15511
rect 13662 15477 13697 15511
rect 13731 15477 13766 15511
rect 13800 15477 13835 15511
rect 13869 15477 13904 15511
rect 13938 15477 13973 15511
rect 14007 15477 14042 15511
rect 14076 15477 14111 15511
rect 14145 15477 14180 15511
rect 14214 15477 14249 15511
rect 14283 15477 14318 15511
rect 14352 15503 14420 15511
rect 14454 15503 14492 15537
rect 14526 15503 14564 15537
rect 14598 15503 14636 15537
rect 14670 15503 14708 15537
rect 14742 15503 14780 15537
rect 14814 15503 14852 15537
rect 14886 15503 14924 15537
rect 14958 15503 14996 15537
rect 15030 15503 15068 15537
rect 15102 15503 15106 15537
rect 14352 15477 15106 15503
rect 12580 15468 15106 15477
rect 12580 15441 14420 15468
rect 12580 15407 12660 15441
rect 12694 15407 12730 15441
rect 12764 15407 12800 15441
rect 12834 15407 12869 15441
rect 12903 15407 12938 15441
rect 12972 15407 13007 15441
rect 13041 15407 13076 15441
rect 13110 15407 13145 15441
rect 13179 15407 13214 15441
rect 13248 15407 13283 15441
rect 13317 15407 13352 15441
rect 13386 15407 13421 15441
rect 13455 15407 13490 15441
rect 13524 15407 13559 15441
rect 13593 15407 13628 15441
rect 13662 15407 13697 15441
rect 13731 15407 13766 15441
rect 13800 15407 13835 15441
rect 13869 15407 13904 15441
rect 13938 15407 13973 15441
rect 14007 15407 14042 15441
rect 14076 15407 14111 15441
rect 14145 15407 14180 15441
rect 14214 15407 14249 15441
rect 14283 15407 14318 15441
rect 14352 15434 14420 15441
rect 14454 15434 14492 15468
rect 14526 15434 14564 15468
rect 14598 15434 14636 15468
rect 14670 15434 14708 15468
rect 14742 15434 14780 15468
rect 14814 15434 14852 15468
rect 14886 15434 14924 15468
rect 14958 15434 14996 15468
rect 15030 15434 15068 15468
rect 15102 15434 15106 15468
rect 14352 15407 15106 15434
rect 12580 15399 15106 15407
rect 12580 15371 14420 15399
rect 12580 15337 12660 15371
rect 12694 15337 12730 15371
rect 12764 15337 12800 15371
rect 12834 15337 12869 15371
rect 12903 15337 12938 15371
rect 12972 15337 13007 15371
rect 13041 15337 13076 15371
rect 13110 15337 13145 15371
rect 13179 15337 13214 15371
rect 13248 15337 13283 15371
rect 13317 15337 13352 15371
rect 13386 15337 13421 15371
rect 13455 15337 13490 15371
rect 13524 15337 13559 15371
rect 13593 15337 13628 15371
rect 13662 15337 13697 15371
rect 13731 15337 13766 15371
rect 13800 15337 13835 15371
rect 13869 15337 13904 15371
rect 13938 15337 13973 15371
rect 14007 15337 14042 15371
rect 14076 15337 14111 15371
rect 14145 15337 14180 15371
rect 14214 15337 14249 15371
rect 14283 15337 14318 15371
rect 14352 15365 14420 15371
rect 14454 15365 14492 15399
rect 14526 15365 14564 15399
rect 14598 15365 14636 15399
rect 14670 15365 14708 15399
rect 14742 15365 14780 15399
rect 14814 15365 14852 15399
rect 14886 15365 14924 15399
rect 14958 15365 14996 15399
rect 15030 15365 15068 15399
rect 15102 15365 15106 15399
rect 14352 15337 15106 15365
rect 12580 15330 15106 15337
rect 12580 15301 14420 15330
rect 12580 15267 12660 15301
rect 12694 15267 12730 15301
rect 12764 15267 12800 15301
rect 12834 15267 12869 15301
rect 12903 15267 12938 15301
rect 12972 15267 13007 15301
rect 13041 15267 13076 15301
rect 13110 15267 13145 15301
rect 13179 15267 13214 15301
rect 13248 15267 13283 15301
rect 13317 15267 13352 15301
rect 13386 15267 13421 15301
rect 13455 15267 13490 15301
rect 13524 15267 13559 15301
rect 13593 15267 13628 15301
rect 13662 15267 13697 15301
rect 13731 15267 13766 15301
rect 13800 15267 13835 15301
rect 13869 15267 13904 15301
rect 13938 15267 13973 15301
rect 14007 15267 14042 15301
rect 14076 15267 14111 15301
rect 14145 15267 14180 15301
rect 14214 15267 14249 15301
rect 14283 15267 14318 15301
rect 14352 15296 14420 15301
rect 14454 15296 14492 15330
rect 14526 15296 14564 15330
rect 14598 15296 14636 15330
rect 14670 15296 14708 15330
rect 14742 15296 14780 15330
rect 14814 15296 14852 15330
rect 14886 15296 14924 15330
rect 14958 15296 14996 15330
rect 15030 15296 15068 15330
rect 15102 15296 15106 15330
rect 14352 15267 15106 15296
rect 12580 15261 15106 15267
rect 12580 15231 14420 15261
rect 12580 15197 12660 15231
rect 12694 15197 12730 15231
rect 12764 15197 12800 15231
rect 12834 15197 12869 15231
rect 12903 15197 12938 15231
rect 12972 15197 13007 15231
rect 13041 15197 13076 15231
rect 13110 15197 13145 15231
rect 13179 15197 13214 15231
rect 13248 15197 13283 15231
rect 13317 15197 13352 15231
rect 13386 15197 13421 15231
rect 13455 15197 13490 15231
rect 13524 15197 13559 15231
rect 13593 15197 13628 15231
rect 13662 15197 13697 15231
rect 13731 15197 13766 15231
rect 13800 15197 13835 15231
rect 13869 15197 13904 15231
rect 13938 15197 13973 15231
rect 14007 15197 14042 15231
rect 14076 15197 14111 15231
rect 14145 15197 14180 15231
rect 14214 15197 14249 15231
rect 14283 15197 14318 15231
rect 14352 15227 14420 15231
rect 14454 15227 14492 15261
rect 14526 15227 14564 15261
rect 14598 15227 14636 15261
rect 14670 15227 14708 15261
rect 14742 15227 14780 15261
rect 14814 15227 14852 15261
rect 14886 15227 14924 15261
rect 14958 15227 14996 15261
rect 15030 15227 15068 15261
rect 15102 15227 15106 15261
rect 14352 15197 15106 15227
rect 12580 15192 15106 15197
rect 12580 15161 14420 15192
rect 12580 15127 12660 15161
rect 12694 15127 12730 15161
rect 12764 15127 12800 15161
rect 12834 15127 12869 15161
rect 12903 15127 12938 15161
rect 12972 15127 13007 15161
rect 13041 15127 13076 15161
rect 13110 15127 13145 15161
rect 13179 15127 13214 15161
rect 13248 15127 13283 15161
rect 13317 15127 13352 15161
rect 13386 15127 13421 15161
rect 13455 15127 13490 15161
rect 13524 15127 13559 15161
rect 13593 15127 13628 15161
rect 13662 15127 13697 15161
rect 13731 15127 13766 15161
rect 13800 15127 13835 15161
rect 13869 15127 13904 15161
rect 13938 15127 13973 15161
rect 14007 15127 14042 15161
rect 14076 15127 14111 15161
rect 14145 15127 14180 15161
rect 14214 15127 14249 15161
rect 14283 15127 14318 15161
rect 14352 15158 14420 15161
rect 14454 15158 14492 15192
rect 14526 15158 14564 15192
rect 14598 15158 14636 15192
rect 14670 15158 14708 15192
rect 14742 15158 14780 15192
rect 14814 15158 14852 15192
rect 14886 15158 14924 15192
rect 14958 15158 14996 15192
rect 15030 15158 15068 15192
rect 15102 15158 15106 15192
rect 14352 15127 15106 15158
rect 12580 15123 15106 15127
rect 12580 15091 14420 15123
rect 12580 15057 12660 15091
rect 12694 15057 12730 15091
rect 12764 15057 12800 15091
rect 12834 15057 12869 15091
rect 12903 15057 12938 15091
rect 12972 15057 13007 15091
rect 13041 15057 13076 15091
rect 13110 15057 13145 15091
rect 13179 15057 13214 15091
rect 13248 15057 13283 15091
rect 13317 15057 13352 15091
rect 13386 15057 13421 15091
rect 13455 15057 13490 15091
rect 13524 15057 13559 15091
rect 13593 15057 13628 15091
rect 13662 15057 13697 15091
rect 13731 15057 13766 15091
rect 13800 15057 13835 15091
rect 13869 15057 13904 15091
rect 13938 15057 13973 15091
rect 14007 15057 14042 15091
rect 14076 15057 14111 15091
rect 14145 15057 14180 15091
rect 14214 15057 14249 15091
rect 14283 15057 14318 15091
rect 14352 15089 14420 15091
rect 14454 15089 14492 15123
rect 14526 15089 14564 15123
rect 14598 15089 14636 15123
rect 14670 15089 14708 15123
rect 14742 15089 14780 15123
rect 14814 15089 14852 15123
rect 14886 15089 14924 15123
rect 14958 15089 14996 15123
rect 15030 15089 15068 15123
rect 15102 15089 15106 15123
rect 14352 15057 15106 15089
rect 12580 15054 15106 15057
rect 12580 15021 14420 15054
rect 12580 14987 12660 15021
rect 12694 14987 12730 15021
rect 12764 14987 12800 15021
rect 12834 14987 12869 15021
rect 12903 14987 12938 15021
rect 12972 14987 13007 15021
rect 13041 14987 13076 15021
rect 13110 14987 13145 15021
rect 13179 14987 13214 15021
rect 13248 14987 13283 15021
rect 13317 14987 13352 15021
rect 13386 14987 13421 15021
rect 13455 14987 13490 15021
rect 13524 14987 13559 15021
rect 13593 14987 13628 15021
rect 13662 14987 13697 15021
rect 13731 14987 13766 15021
rect 13800 14987 13835 15021
rect 13869 14987 13904 15021
rect 13938 14987 13973 15021
rect 14007 14987 14042 15021
rect 14076 14987 14111 15021
rect 14145 14987 14180 15021
rect 14214 14987 14249 15021
rect 14283 14987 14318 15021
rect 14352 15020 14420 15021
rect 14454 15020 14492 15054
rect 14526 15020 14564 15054
rect 14598 15020 14636 15054
rect 14670 15020 14708 15054
rect 14742 15020 14780 15054
rect 14814 15020 14852 15054
rect 14886 15020 14924 15054
rect 14958 15020 14996 15054
rect 15030 15020 15068 15054
rect 15102 15020 15106 15054
rect 14352 14987 15106 15020
rect 12580 14985 15106 14987
rect 12580 14951 14420 14985
rect 14454 14951 14492 14985
rect 14526 14951 14564 14985
rect 14598 14951 14636 14985
rect 14670 14951 14708 14985
rect 14742 14951 14780 14985
rect 14814 14951 14852 14985
rect 14886 14951 14924 14985
rect 14958 14951 14996 14985
rect 15030 14951 15068 14985
rect 15102 14951 15106 14985
rect 12580 14917 12660 14951
rect 12694 14917 12730 14951
rect 12764 14917 12800 14951
rect 12834 14917 12869 14951
rect 12903 14917 12938 14951
rect 12972 14917 13007 14951
rect 13041 14917 13076 14951
rect 13110 14917 13145 14951
rect 13179 14917 13214 14951
rect 13248 14917 13283 14951
rect 13317 14917 13352 14951
rect 13386 14917 13421 14951
rect 13455 14917 13490 14951
rect 13524 14917 13559 14951
rect 13593 14917 13628 14951
rect 13662 14917 13697 14951
rect 13731 14917 13766 14951
rect 13800 14917 13835 14951
rect 13869 14917 13904 14951
rect 13938 14917 13973 14951
rect 14007 14917 14042 14951
rect 14076 14917 14111 14951
rect 14145 14917 14180 14951
rect 14214 14917 14249 14951
rect 14283 14917 14318 14951
rect 14352 14917 15106 14951
rect 12580 14916 15106 14917
rect 12580 14882 14420 14916
rect 14454 14882 14492 14916
rect 14526 14882 14564 14916
rect 14598 14882 14636 14916
rect 14670 14882 14708 14916
rect 14742 14882 14780 14916
rect 14814 14882 14852 14916
rect 14886 14882 14924 14916
rect 14958 14882 14996 14916
rect 15030 14882 15068 14916
rect 15102 14882 15106 14916
rect 12580 14881 15106 14882
rect 12580 14847 12660 14881
rect 12694 14847 12730 14881
rect 12764 14847 12800 14881
rect 12834 14847 12869 14881
rect 12903 14847 12938 14881
rect 12972 14847 13007 14881
rect 13041 14847 13076 14881
rect 13110 14847 13145 14881
rect 13179 14847 13214 14881
rect 13248 14847 13283 14881
rect 13317 14847 13352 14881
rect 13386 14847 13421 14881
rect 13455 14847 13490 14881
rect 13524 14847 13559 14881
rect 13593 14847 13628 14881
rect 13662 14847 13697 14881
rect 13731 14847 13766 14881
rect 13800 14847 13835 14881
rect 13869 14847 13904 14881
rect 13938 14847 13973 14881
rect 14007 14847 14042 14881
rect 14076 14847 14111 14881
rect 14145 14847 14180 14881
rect 14214 14847 14249 14881
rect 14283 14847 14318 14881
rect 14352 14847 15106 14881
rect 12580 14813 14420 14847
rect 14454 14813 14492 14847
rect 14526 14813 14564 14847
rect 14598 14813 14636 14847
rect 14670 14813 14708 14847
rect 14742 14813 14780 14847
rect 14814 14813 14852 14847
rect 14886 14813 14924 14847
rect 14958 14813 14996 14847
rect 15030 14813 15068 14847
rect 15102 14813 15106 14847
rect 12580 14793 15106 14813
rect 67 14777 5556 14793
rect 12467 14777 15106 14793
rect 8359 8808 15102 8809
rect 34 8774 15102 8808
rect 34 8740 68 8774
rect 102 8740 138 8774
rect 172 8740 208 8774
rect 242 8740 278 8774
rect 312 8740 348 8774
rect 382 8740 418 8774
rect 452 8740 488 8774
rect 522 8740 558 8774
rect 592 8740 628 8774
rect 662 8740 698 8774
rect 732 8740 768 8774
rect 802 8740 838 8774
rect 872 8740 908 8774
rect 942 8740 978 8774
rect 1012 8740 1048 8774
rect 1082 8740 1118 8774
rect 1152 8740 1188 8774
rect 1222 8740 1258 8774
rect 1292 8740 1328 8774
rect 1362 8740 1398 8774
rect 1432 8740 1467 8774
rect 1501 8740 1536 8774
rect 1570 8740 1605 8774
rect 1639 8740 1674 8774
rect 1708 8740 1743 8774
rect 1777 8740 1812 8774
rect 1846 8740 1881 8774
rect 1915 8740 1950 8774
rect 1984 8740 2019 8774
rect 2053 8740 2088 8774
rect 2122 8740 2157 8774
rect 2191 8740 2226 8774
rect 2260 8740 2295 8774
rect 2329 8740 2364 8774
rect 2398 8740 2433 8774
rect 2467 8740 2502 8774
rect 2536 8740 2571 8774
rect 2605 8740 2640 8774
rect 2674 8740 2709 8774
rect 2743 8740 2778 8774
rect 2812 8740 2847 8774
rect 2881 8773 15102 8774
rect 2881 8770 8393 8773
rect 2881 8740 2933 8770
rect 34 8736 2933 8740
rect 2967 8736 3002 8770
rect 3036 8736 3071 8770
rect 3105 8736 3139 8770
rect 3173 8736 3207 8770
rect 3241 8736 3275 8770
rect 3309 8736 3343 8770
rect 3377 8736 3411 8770
rect 3445 8736 3479 8770
rect 3513 8736 3547 8770
rect 3581 8736 3615 8770
rect 3649 8736 3683 8770
rect 3717 8736 3751 8770
rect 3785 8736 3819 8770
rect 3853 8736 3887 8770
rect 3921 8736 3955 8770
rect 3989 8736 4023 8770
rect 4057 8736 4091 8770
rect 4125 8736 4159 8770
rect 4193 8736 4227 8770
rect 4261 8736 4295 8770
rect 4329 8736 4363 8770
rect 4397 8736 4431 8770
rect 4465 8736 4499 8770
rect 4533 8736 4567 8770
rect 4601 8736 4635 8770
rect 4669 8736 4703 8770
rect 4737 8736 4771 8770
rect 4805 8736 4839 8770
rect 4873 8736 4907 8770
rect 4941 8736 4975 8770
rect 5009 8736 5043 8770
rect 5077 8736 5111 8770
rect 5145 8736 5179 8770
rect 5213 8736 5247 8770
rect 5281 8736 5315 8770
rect 5349 8736 5383 8770
rect 5417 8736 5451 8770
rect 5485 8736 5519 8770
rect 5553 8736 5587 8770
rect 5621 8736 5655 8770
rect 5689 8736 5723 8770
rect 5757 8736 5791 8770
rect 5825 8736 5859 8770
rect 5893 8736 5927 8770
rect 5961 8736 5995 8770
rect 6029 8736 6063 8770
rect 6097 8736 6131 8770
rect 6165 8736 6199 8770
rect 6233 8736 6267 8770
rect 6301 8736 6335 8770
rect 6369 8736 6403 8770
rect 6437 8736 6471 8770
rect 6505 8736 6539 8770
rect 6573 8736 6607 8770
rect 6641 8736 6675 8770
rect 6709 8736 6743 8770
rect 6777 8736 6811 8770
rect 6845 8736 6879 8770
rect 6913 8736 6947 8770
rect 6981 8736 7015 8770
rect 7049 8736 7083 8770
rect 7117 8736 7151 8770
rect 7185 8736 7219 8770
rect 7253 8736 7287 8770
rect 7321 8736 7355 8770
rect 7389 8736 7423 8770
rect 7457 8736 7491 8770
rect 7525 8736 7559 8770
rect 7593 8736 7627 8770
rect 7661 8736 7695 8770
rect 7729 8736 7763 8770
rect 7797 8736 7831 8770
rect 7865 8736 7899 8770
rect 7933 8736 7967 8770
rect 8001 8736 8035 8770
rect 8069 8736 8103 8770
rect 8137 8736 8171 8770
rect 8205 8736 8239 8770
rect 8273 8736 8307 8770
rect 8341 8739 8393 8770
rect 8427 8739 8462 8773
rect 8496 8739 8531 8773
rect 8565 8739 8600 8773
rect 8634 8739 8669 8773
rect 8703 8739 8738 8773
rect 8772 8739 8807 8773
rect 8841 8739 8876 8773
rect 8910 8739 8945 8773
rect 8979 8739 9014 8773
rect 9048 8739 9083 8773
rect 9117 8739 9152 8773
rect 9186 8739 9220 8773
rect 9254 8739 9288 8773
rect 9322 8739 9356 8773
rect 9390 8739 9424 8773
rect 9458 8739 9492 8773
rect 9526 8739 9560 8773
rect 9594 8739 9628 8773
rect 9662 8739 9696 8773
rect 9730 8739 9764 8773
rect 9798 8739 9832 8773
rect 9866 8739 9900 8773
rect 9934 8739 9968 8773
rect 10002 8739 10036 8773
rect 10070 8739 10104 8773
rect 10138 8739 10172 8773
rect 10206 8739 10240 8773
rect 10274 8739 10308 8773
rect 10342 8739 10376 8773
rect 10410 8739 10444 8773
rect 10478 8739 10512 8773
rect 10546 8739 10580 8773
rect 10614 8739 10648 8773
rect 10682 8739 10716 8773
rect 10750 8739 10784 8773
rect 10818 8739 10852 8773
rect 10886 8739 10920 8773
rect 10954 8739 10988 8773
rect 11022 8739 11056 8773
rect 11090 8739 11124 8773
rect 11158 8739 11192 8773
rect 11226 8739 11260 8773
rect 11294 8739 11328 8773
rect 11362 8739 11396 8773
rect 11430 8739 11464 8773
rect 11498 8739 11532 8773
rect 11566 8739 11600 8773
rect 11634 8739 11668 8773
rect 11702 8739 11736 8773
rect 11770 8739 11804 8773
rect 11838 8739 11872 8773
rect 11906 8739 11940 8773
rect 11974 8739 12008 8773
rect 12042 8739 12076 8773
rect 12110 8739 12144 8773
rect 12178 8739 12212 8773
rect 12246 8739 12280 8773
rect 12314 8739 12348 8773
rect 12382 8739 12416 8773
rect 12450 8739 12484 8773
rect 12518 8739 12552 8773
rect 12586 8739 12620 8773
rect 12654 8739 12688 8773
rect 12722 8739 12756 8773
rect 12790 8739 12824 8773
rect 12858 8739 12892 8773
rect 12926 8739 12960 8773
rect 12994 8739 13028 8773
rect 13062 8739 13096 8773
rect 13130 8739 13164 8773
rect 13198 8739 13232 8773
rect 13266 8739 13300 8773
rect 13334 8739 13368 8773
rect 13402 8739 13436 8773
rect 13470 8739 13504 8773
rect 13538 8739 13572 8773
rect 13606 8739 13640 8773
rect 13674 8739 13708 8773
rect 13742 8739 13776 8773
rect 13810 8739 13844 8773
rect 13878 8739 13912 8773
rect 13946 8739 13980 8773
rect 14014 8739 14048 8773
rect 14082 8739 14116 8773
rect 14150 8739 14184 8773
rect 14218 8739 14252 8773
rect 14286 8739 14320 8773
rect 14354 8739 14388 8773
rect 14422 8739 14456 8773
rect 14490 8739 14524 8773
rect 14558 8739 14592 8773
rect 14626 8739 14660 8773
rect 14694 8739 14728 8773
rect 14762 8739 14796 8773
rect 14830 8739 14864 8773
rect 14898 8739 15102 8773
rect 8341 8736 15102 8739
rect 34 8721 15102 8736
rect 34 8700 14932 8721
rect 34 8666 68 8700
rect 102 8666 138 8700
rect 172 8666 208 8700
rect 242 8666 278 8700
rect 312 8666 348 8700
rect 382 8666 418 8700
rect 452 8666 488 8700
rect 522 8666 558 8700
rect 592 8666 628 8700
rect 662 8666 698 8700
rect 732 8666 768 8700
rect 802 8666 838 8700
rect 872 8666 908 8700
rect 942 8666 978 8700
rect 1012 8666 1048 8700
rect 1082 8666 1118 8700
rect 1152 8666 1188 8700
rect 1222 8666 1258 8700
rect 1292 8666 1328 8700
rect 1362 8666 1398 8700
rect 1432 8666 1467 8700
rect 1501 8666 1536 8700
rect 1570 8666 1605 8700
rect 1639 8666 1674 8700
rect 1708 8666 1743 8700
rect 1777 8666 1812 8700
rect 1846 8666 1881 8700
rect 1915 8666 1950 8700
rect 1984 8666 2019 8700
rect 2053 8666 2088 8700
rect 2122 8666 2157 8700
rect 2191 8666 2226 8700
rect 2260 8666 2295 8700
rect 2329 8666 2364 8700
rect 2398 8666 2433 8700
rect 2467 8666 2502 8700
rect 2536 8666 2571 8700
rect 2605 8666 2640 8700
rect 2674 8666 2709 8700
rect 2743 8666 2778 8700
rect 2812 8666 2847 8700
rect 2881 8666 2933 8700
rect 2967 8666 3002 8700
rect 3036 8666 3071 8700
rect 3105 8666 3139 8700
rect 3173 8666 3207 8700
rect 3241 8666 3275 8700
rect 3309 8666 3343 8700
rect 3377 8666 3411 8700
rect 3445 8666 3479 8700
rect 3513 8666 3547 8700
rect 3581 8666 3615 8700
rect 3649 8666 3683 8700
rect 3717 8666 3751 8700
rect 3785 8666 3819 8700
rect 3853 8666 3887 8700
rect 3921 8666 3955 8700
rect 3989 8666 4023 8700
rect 4057 8666 4091 8700
rect 4125 8666 4159 8700
rect 4193 8666 4227 8700
rect 4261 8666 4295 8700
rect 4329 8666 4363 8700
rect 4397 8666 4431 8700
rect 4465 8666 4499 8700
rect 4533 8666 4567 8700
rect 4601 8666 4635 8700
rect 4669 8666 4703 8700
rect 4737 8666 4771 8700
rect 4805 8666 4839 8700
rect 4873 8666 4907 8700
rect 4941 8666 4975 8700
rect 5009 8666 5043 8700
rect 5077 8666 5111 8700
rect 5145 8666 5179 8700
rect 5213 8666 5247 8700
rect 5281 8666 5315 8700
rect 5349 8666 5383 8700
rect 5417 8666 5451 8700
rect 5485 8666 5519 8700
rect 5553 8666 5587 8700
rect 5621 8666 5655 8700
rect 5689 8666 5723 8700
rect 5757 8666 5791 8700
rect 5825 8666 5859 8700
rect 5893 8666 5927 8700
rect 5961 8666 5995 8700
rect 6029 8666 6063 8700
rect 6097 8666 6131 8700
rect 6165 8666 6199 8700
rect 6233 8666 6267 8700
rect 6301 8666 6335 8700
rect 6369 8666 6403 8700
rect 6437 8666 6471 8700
rect 6505 8666 6539 8700
rect 6573 8666 6607 8700
rect 6641 8666 6675 8700
rect 6709 8666 6743 8700
rect 6777 8666 6811 8700
rect 6845 8666 6879 8700
rect 6913 8666 6947 8700
rect 6981 8666 7015 8700
rect 7049 8666 7083 8700
rect 7117 8666 7151 8700
rect 7185 8666 7219 8700
rect 7253 8666 7287 8700
rect 7321 8666 7355 8700
rect 7389 8666 7423 8700
rect 7457 8666 7491 8700
rect 7525 8666 7559 8700
rect 7593 8666 7627 8700
rect 7661 8666 7695 8700
rect 7729 8666 7763 8700
rect 7797 8666 7831 8700
rect 7865 8666 7899 8700
rect 7933 8666 7967 8700
rect 8001 8666 8035 8700
rect 8069 8666 8103 8700
rect 8137 8666 8171 8700
rect 8205 8666 8239 8700
rect 8273 8666 8307 8700
rect 8341 8693 14932 8700
rect 8341 8666 8393 8693
rect 34 8659 8393 8666
rect 8427 8659 8462 8693
rect 8496 8659 8531 8693
rect 8565 8659 8600 8693
rect 8634 8659 8669 8693
rect 8703 8659 8738 8693
rect 8772 8659 8807 8693
rect 8841 8659 8876 8693
rect 8910 8659 8945 8693
rect 8979 8659 9014 8693
rect 9048 8659 9083 8693
rect 9117 8659 9152 8693
rect 9186 8659 9220 8693
rect 9254 8659 9288 8693
rect 9322 8659 9356 8693
rect 9390 8659 9424 8693
rect 9458 8659 9492 8693
rect 9526 8659 9560 8693
rect 9594 8659 9628 8693
rect 9662 8659 9696 8693
rect 9730 8659 9764 8693
rect 9798 8659 9832 8693
rect 9866 8659 9900 8693
rect 9934 8659 9968 8693
rect 10002 8659 10036 8693
rect 10070 8659 10104 8693
rect 10138 8659 10172 8693
rect 10206 8659 10240 8693
rect 10274 8659 10308 8693
rect 10342 8659 10376 8693
rect 10410 8659 10444 8693
rect 10478 8659 10512 8693
rect 10546 8659 10580 8693
rect 10614 8659 10648 8693
rect 10682 8659 10716 8693
rect 10750 8659 10784 8693
rect 10818 8659 10852 8693
rect 10886 8659 10920 8693
rect 10954 8659 10988 8693
rect 11022 8659 11056 8693
rect 11090 8659 11124 8693
rect 11158 8659 11192 8693
rect 11226 8659 11260 8693
rect 11294 8659 11328 8693
rect 11362 8659 11396 8693
rect 11430 8659 11464 8693
rect 11498 8659 11532 8693
rect 11566 8659 11600 8693
rect 11634 8659 11668 8693
rect 11702 8659 11736 8693
rect 11770 8659 11804 8693
rect 11838 8659 11872 8693
rect 11906 8659 11940 8693
rect 11974 8659 12008 8693
rect 12042 8659 12076 8693
rect 12110 8659 12144 8693
rect 12178 8659 12212 8693
rect 12246 8659 12280 8693
rect 12314 8659 12348 8693
rect 12382 8659 12416 8693
rect 12450 8659 12484 8693
rect 12518 8659 12552 8693
rect 12586 8659 12620 8693
rect 12654 8659 12688 8693
rect 12722 8659 12756 8693
rect 12790 8659 12824 8693
rect 12858 8659 12892 8693
rect 12926 8659 12960 8693
rect 12994 8659 13028 8693
rect 13062 8659 13096 8693
rect 13130 8659 13164 8693
rect 13198 8659 13232 8693
rect 13266 8659 13300 8693
rect 13334 8659 13368 8693
rect 13402 8659 13436 8693
rect 13470 8659 13504 8693
rect 13538 8659 13572 8693
rect 13606 8659 13640 8693
rect 13674 8659 13708 8693
rect 13742 8659 13776 8693
rect 13810 8659 13844 8693
rect 13878 8659 13912 8693
rect 13946 8659 13980 8693
rect 14014 8659 14048 8693
rect 14082 8659 14116 8693
rect 14150 8659 14184 8693
rect 14218 8659 14252 8693
rect 14286 8659 14320 8693
rect 14354 8659 14388 8693
rect 14422 8659 14456 8693
rect 14490 8659 14524 8693
rect 14558 8659 14592 8693
rect 14626 8659 14660 8693
rect 14694 8659 14728 8693
rect 14762 8659 14796 8693
rect 14830 8659 14864 8693
rect 14898 8687 14932 8693
rect 14966 8687 15000 8721
rect 15034 8687 15068 8721
rect 14898 8659 15102 8687
rect 34 8649 15102 8659
rect 34 8630 14932 8649
rect 34 8626 2933 8630
rect 34 8592 68 8626
rect 102 8592 138 8626
rect 172 8592 208 8626
rect 242 8592 278 8626
rect 312 8592 348 8626
rect 382 8592 418 8626
rect 452 8592 488 8626
rect 522 8592 558 8626
rect 592 8592 628 8626
rect 662 8592 698 8626
rect 732 8592 768 8626
rect 802 8592 838 8626
rect 872 8592 908 8626
rect 942 8592 978 8626
rect 1012 8592 1048 8626
rect 1082 8592 1118 8626
rect 1152 8592 1188 8626
rect 1222 8592 1258 8626
rect 1292 8592 1328 8626
rect 1362 8592 1398 8626
rect 1432 8592 1467 8626
rect 1501 8592 1536 8626
rect 1570 8592 1605 8626
rect 1639 8592 1674 8626
rect 1708 8592 1743 8626
rect 1777 8592 1812 8626
rect 1846 8592 1881 8626
rect 1915 8592 1950 8626
rect 1984 8592 2019 8626
rect 2053 8592 2088 8626
rect 2122 8592 2157 8626
rect 2191 8592 2226 8626
rect 2260 8592 2295 8626
rect 2329 8592 2364 8626
rect 2398 8592 2433 8626
rect 2467 8592 2502 8626
rect 2536 8592 2571 8626
rect 2605 8592 2640 8626
rect 2674 8592 2709 8626
rect 2743 8592 2778 8626
rect 2812 8592 2847 8626
rect 2881 8596 2933 8626
rect 2967 8596 3002 8630
rect 3036 8596 3071 8630
rect 3105 8596 3139 8630
rect 3173 8596 3207 8630
rect 3241 8596 3275 8630
rect 3309 8596 3343 8630
rect 3377 8596 3411 8630
rect 3445 8596 3479 8630
rect 3513 8596 3547 8630
rect 3581 8596 3615 8630
rect 3649 8596 3683 8630
rect 3717 8596 3751 8630
rect 3785 8596 3819 8630
rect 3853 8596 3887 8630
rect 3921 8596 3955 8630
rect 3989 8596 4023 8630
rect 4057 8596 4091 8630
rect 4125 8596 4159 8630
rect 4193 8596 4227 8630
rect 4261 8596 4295 8630
rect 4329 8596 4363 8630
rect 4397 8596 4431 8630
rect 4465 8596 4499 8630
rect 4533 8596 4567 8630
rect 4601 8596 4635 8630
rect 4669 8596 4703 8630
rect 4737 8596 4771 8630
rect 4805 8596 4839 8630
rect 4873 8596 4907 8630
rect 4941 8596 4975 8630
rect 5009 8596 5043 8630
rect 5077 8596 5111 8630
rect 5145 8596 5179 8630
rect 5213 8596 5247 8630
rect 5281 8596 5315 8630
rect 5349 8596 5383 8630
rect 5417 8596 5451 8630
rect 5485 8596 5519 8630
rect 5553 8596 5587 8630
rect 5621 8596 5655 8630
rect 5689 8596 5723 8630
rect 5757 8596 5791 8630
rect 5825 8596 5859 8630
rect 5893 8596 5927 8630
rect 5961 8596 5995 8630
rect 6029 8596 6063 8630
rect 6097 8596 6131 8630
rect 6165 8596 6199 8630
rect 6233 8596 6267 8630
rect 6301 8596 6335 8630
rect 6369 8596 6403 8630
rect 6437 8596 6471 8630
rect 6505 8596 6539 8630
rect 6573 8596 6607 8630
rect 6641 8596 6675 8630
rect 6709 8596 6743 8630
rect 6777 8596 6811 8630
rect 6845 8596 6879 8630
rect 6913 8596 6947 8630
rect 6981 8596 7015 8630
rect 7049 8596 7083 8630
rect 7117 8596 7151 8630
rect 7185 8596 7219 8630
rect 7253 8596 7287 8630
rect 7321 8596 7355 8630
rect 7389 8596 7423 8630
rect 7457 8596 7491 8630
rect 7525 8596 7559 8630
rect 7593 8596 7627 8630
rect 7661 8596 7695 8630
rect 7729 8596 7763 8630
rect 7797 8596 7831 8630
rect 7865 8596 7899 8630
rect 7933 8596 7967 8630
rect 8001 8596 8035 8630
rect 8069 8596 8103 8630
rect 8137 8596 8171 8630
rect 8205 8596 8239 8630
rect 8273 8596 8307 8630
rect 8341 8615 14932 8630
rect 14966 8615 15000 8649
rect 15034 8615 15068 8649
rect 8341 8613 15102 8615
rect 8341 8596 8393 8613
rect 2881 8592 8393 8596
rect 34 8579 8393 8592
rect 8427 8579 8462 8613
rect 8496 8579 8531 8613
rect 8565 8579 8600 8613
rect 8634 8579 8669 8613
rect 8703 8579 8738 8613
rect 8772 8579 8807 8613
rect 8841 8579 8876 8613
rect 8910 8579 8945 8613
rect 8979 8579 9014 8613
rect 9048 8579 9083 8613
rect 9117 8579 9152 8613
rect 9186 8579 9220 8613
rect 9254 8579 9288 8613
rect 9322 8579 9356 8613
rect 9390 8579 9424 8613
rect 9458 8579 9492 8613
rect 9526 8579 9560 8613
rect 9594 8579 9628 8613
rect 9662 8579 9696 8613
rect 9730 8579 9764 8613
rect 9798 8579 9832 8613
rect 9866 8579 9900 8613
rect 9934 8579 9968 8613
rect 10002 8579 10036 8613
rect 10070 8579 10104 8613
rect 10138 8579 10172 8613
rect 10206 8579 10240 8613
rect 10274 8579 10308 8613
rect 10342 8579 10376 8613
rect 10410 8579 10444 8613
rect 10478 8579 10512 8613
rect 10546 8579 10580 8613
rect 10614 8579 10648 8613
rect 10682 8579 10716 8613
rect 10750 8579 10784 8613
rect 10818 8579 10852 8613
rect 10886 8579 10920 8613
rect 10954 8579 10988 8613
rect 11022 8579 11056 8613
rect 11090 8579 11124 8613
rect 11158 8579 11192 8613
rect 11226 8579 11260 8613
rect 11294 8579 11328 8613
rect 11362 8579 11396 8613
rect 11430 8579 11464 8613
rect 11498 8579 11532 8613
rect 11566 8579 11600 8613
rect 11634 8579 11668 8613
rect 11702 8579 11736 8613
rect 11770 8579 11804 8613
rect 11838 8579 11872 8613
rect 11906 8579 11940 8613
rect 11974 8579 12008 8613
rect 12042 8579 12076 8613
rect 12110 8579 12144 8613
rect 12178 8579 12212 8613
rect 12246 8579 12280 8613
rect 12314 8579 12348 8613
rect 12382 8579 12416 8613
rect 12450 8579 12484 8613
rect 12518 8579 12552 8613
rect 12586 8579 12620 8613
rect 12654 8579 12688 8613
rect 12722 8579 12756 8613
rect 12790 8579 12824 8613
rect 12858 8579 12892 8613
rect 12926 8579 12960 8613
rect 12994 8579 13028 8613
rect 13062 8579 13096 8613
rect 13130 8579 13164 8613
rect 13198 8579 13232 8613
rect 13266 8579 13300 8613
rect 13334 8579 13368 8613
rect 13402 8579 13436 8613
rect 13470 8579 13504 8613
rect 13538 8579 13572 8613
rect 13606 8579 13640 8613
rect 13674 8579 13708 8613
rect 13742 8579 13776 8613
rect 13810 8579 13844 8613
rect 13878 8579 13912 8613
rect 13946 8579 13980 8613
rect 14014 8579 14048 8613
rect 14082 8579 14116 8613
rect 14150 8579 14184 8613
rect 14218 8579 14252 8613
rect 14286 8579 14320 8613
rect 14354 8579 14388 8613
rect 14422 8579 14456 8613
rect 14490 8579 14524 8613
rect 14558 8579 14592 8613
rect 14626 8579 14660 8613
rect 14694 8579 14728 8613
rect 14762 8579 14796 8613
rect 14830 8579 14864 8613
rect 14898 8579 15102 8613
rect 34 8577 15102 8579
rect 34 8560 14932 8577
rect 34 8552 2933 8560
rect 34 8518 68 8552
rect 102 8518 138 8552
rect 172 8518 208 8552
rect 242 8518 278 8552
rect 312 8518 348 8552
rect 382 8518 418 8552
rect 452 8518 488 8552
rect 522 8518 558 8552
rect 592 8518 628 8552
rect 662 8518 698 8552
rect 732 8518 768 8552
rect 802 8518 838 8552
rect 872 8518 908 8552
rect 942 8518 978 8552
rect 1012 8518 1048 8552
rect 1082 8518 1118 8552
rect 1152 8518 1188 8552
rect 1222 8518 1258 8552
rect 1292 8518 1328 8552
rect 1362 8518 1398 8552
rect 1432 8518 1467 8552
rect 1501 8518 1536 8552
rect 1570 8518 1605 8552
rect 1639 8518 1674 8552
rect 1708 8518 1743 8552
rect 1777 8518 1812 8552
rect 1846 8518 1881 8552
rect 1915 8518 1950 8552
rect 1984 8518 2019 8552
rect 2053 8518 2088 8552
rect 2122 8518 2157 8552
rect 2191 8518 2226 8552
rect 2260 8518 2295 8552
rect 2329 8518 2364 8552
rect 2398 8518 2433 8552
rect 2467 8518 2502 8552
rect 2536 8518 2571 8552
rect 2605 8518 2640 8552
rect 2674 8518 2709 8552
rect 2743 8518 2778 8552
rect 2812 8518 2847 8552
rect 2881 8526 2933 8552
rect 2967 8526 3002 8560
rect 3036 8526 3071 8560
rect 3105 8526 3139 8560
rect 3173 8526 3207 8560
rect 3241 8526 3275 8560
rect 3309 8526 3343 8560
rect 3377 8526 3411 8560
rect 3445 8526 3479 8560
rect 3513 8526 3547 8560
rect 3581 8526 3615 8560
rect 3649 8526 3683 8560
rect 3717 8526 3751 8560
rect 3785 8526 3819 8560
rect 3853 8526 3887 8560
rect 3921 8526 3955 8560
rect 3989 8526 4023 8560
rect 4057 8526 4091 8560
rect 4125 8526 4159 8560
rect 4193 8526 4227 8560
rect 4261 8526 4295 8560
rect 4329 8526 4363 8560
rect 4397 8526 4431 8560
rect 4465 8526 4499 8560
rect 4533 8526 4567 8560
rect 4601 8526 4635 8560
rect 4669 8526 4703 8560
rect 4737 8526 4771 8560
rect 4805 8526 4839 8560
rect 4873 8526 4907 8560
rect 4941 8526 4975 8560
rect 5009 8526 5043 8560
rect 5077 8526 5111 8560
rect 5145 8526 5179 8560
rect 5213 8526 5247 8560
rect 5281 8526 5315 8560
rect 5349 8526 5383 8560
rect 5417 8526 5451 8560
rect 5485 8526 5519 8560
rect 5553 8526 5587 8560
rect 5621 8526 5655 8560
rect 5689 8526 5723 8560
rect 5757 8526 5791 8560
rect 5825 8526 5859 8560
rect 5893 8526 5927 8560
rect 5961 8526 5995 8560
rect 6029 8526 6063 8560
rect 6097 8526 6131 8560
rect 6165 8526 6199 8560
rect 6233 8526 6267 8560
rect 6301 8526 6335 8560
rect 6369 8526 6403 8560
rect 6437 8526 6471 8560
rect 6505 8526 6539 8560
rect 6573 8526 6607 8560
rect 6641 8526 6675 8560
rect 6709 8526 6743 8560
rect 6777 8526 6811 8560
rect 6845 8526 6879 8560
rect 6913 8526 6947 8560
rect 6981 8526 7015 8560
rect 7049 8526 7083 8560
rect 7117 8526 7151 8560
rect 7185 8526 7219 8560
rect 7253 8526 7287 8560
rect 7321 8526 7355 8560
rect 7389 8526 7423 8560
rect 7457 8526 7491 8560
rect 7525 8526 7559 8560
rect 7593 8526 7627 8560
rect 7661 8526 7695 8560
rect 7729 8526 7763 8560
rect 7797 8526 7831 8560
rect 7865 8526 7899 8560
rect 7933 8526 7967 8560
rect 8001 8526 8035 8560
rect 8069 8526 8103 8560
rect 8137 8526 8171 8560
rect 8205 8526 8239 8560
rect 8273 8526 8307 8560
rect 8341 8543 14932 8560
rect 14966 8543 15000 8577
rect 15034 8543 15068 8577
rect 8341 8533 15102 8543
rect 8341 8526 8393 8533
rect 2881 8518 8393 8526
rect 34 8499 8393 8518
rect 8427 8499 8462 8533
rect 8496 8499 8531 8533
rect 8565 8499 8600 8533
rect 8634 8499 8669 8533
rect 8703 8499 8738 8533
rect 8772 8499 8807 8533
rect 8841 8499 8876 8533
rect 8910 8499 8945 8533
rect 8979 8499 9014 8533
rect 9048 8499 9083 8533
rect 9117 8499 9152 8533
rect 9186 8499 9220 8533
rect 9254 8499 9288 8533
rect 9322 8499 9356 8533
rect 9390 8499 9424 8533
rect 9458 8499 9492 8533
rect 9526 8499 9560 8533
rect 9594 8499 9628 8533
rect 9662 8499 9696 8533
rect 9730 8499 9764 8533
rect 9798 8499 9832 8533
rect 9866 8499 9900 8533
rect 9934 8499 9968 8533
rect 10002 8499 10036 8533
rect 10070 8499 10104 8533
rect 10138 8499 10172 8533
rect 10206 8499 10240 8533
rect 10274 8499 10308 8533
rect 10342 8499 10376 8533
rect 10410 8499 10444 8533
rect 10478 8499 10512 8533
rect 10546 8499 10580 8533
rect 10614 8499 10648 8533
rect 10682 8499 10716 8533
rect 10750 8499 10784 8533
rect 10818 8499 10852 8533
rect 10886 8499 10920 8533
rect 10954 8499 10988 8533
rect 11022 8499 11056 8533
rect 11090 8499 11124 8533
rect 11158 8499 11192 8533
rect 11226 8499 11260 8533
rect 11294 8499 11328 8533
rect 11362 8499 11396 8533
rect 11430 8499 11464 8533
rect 11498 8499 11532 8533
rect 11566 8499 11600 8533
rect 11634 8499 11668 8533
rect 11702 8499 11736 8533
rect 11770 8499 11804 8533
rect 11838 8499 11872 8533
rect 11906 8499 11940 8533
rect 11974 8499 12008 8533
rect 12042 8499 12076 8533
rect 12110 8499 12144 8533
rect 12178 8499 12212 8533
rect 12246 8499 12280 8533
rect 12314 8499 12348 8533
rect 12382 8499 12416 8533
rect 12450 8499 12484 8533
rect 12518 8499 12552 8533
rect 12586 8499 12620 8533
rect 12654 8499 12688 8533
rect 12722 8499 12756 8533
rect 12790 8499 12824 8533
rect 12858 8499 12892 8533
rect 12926 8499 12960 8533
rect 12994 8499 13028 8533
rect 13062 8499 13096 8533
rect 13130 8499 13164 8533
rect 13198 8499 13232 8533
rect 13266 8499 13300 8533
rect 13334 8499 13368 8533
rect 13402 8499 13436 8533
rect 13470 8499 13504 8533
rect 13538 8499 13572 8533
rect 13606 8499 13640 8533
rect 13674 8499 13708 8533
rect 13742 8499 13776 8533
rect 13810 8499 13844 8533
rect 13878 8499 13912 8533
rect 13946 8499 13980 8533
rect 14014 8499 14048 8533
rect 14082 8499 14116 8533
rect 14150 8499 14184 8533
rect 14218 8499 14252 8533
rect 14286 8499 14320 8533
rect 14354 8499 14388 8533
rect 14422 8499 14456 8533
rect 14490 8499 14524 8533
rect 14558 8499 14592 8533
rect 14626 8499 14660 8533
rect 14694 8499 14728 8533
rect 14762 8499 14796 8533
rect 14830 8499 14864 8533
rect 14898 8505 15102 8533
rect 14898 8499 14932 8505
rect 34 8490 14932 8499
rect 34 8484 2933 8490
rect 34 8460 136 8484
rect 34 8426 68 8460
rect 102 8426 136 8460
rect 34 8392 136 8426
rect 34 8358 68 8392
rect 102 8358 136 8392
rect 2899 8456 2933 8484
rect 2967 8456 3002 8490
rect 3036 8456 3071 8490
rect 3105 8456 3139 8490
rect 3173 8456 3207 8490
rect 3241 8456 3275 8490
rect 3309 8456 3343 8490
rect 3377 8456 3411 8490
rect 3445 8456 3479 8490
rect 3513 8456 3547 8490
rect 3581 8456 3615 8490
rect 3649 8456 3683 8490
rect 3717 8456 3751 8490
rect 3785 8456 3819 8490
rect 3853 8456 3887 8490
rect 3921 8456 3955 8490
rect 3989 8456 4023 8490
rect 4057 8456 4091 8490
rect 4125 8456 4159 8490
rect 4193 8456 4227 8490
rect 4261 8456 4295 8490
rect 4329 8456 4363 8490
rect 4397 8456 4431 8490
rect 4465 8456 4499 8490
rect 4533 8456 4567 8490
rect 4601 8456 4635 8490
rect 4669 8456 4703 8490
rect 4737 8456 4771 8490
rect 4805 8456 4839 8490
rect 4873 8456 4907 8490
rect 4941 8456 4975 8490
rect 5009 8456 5043 8490
rect 5077 8456 5111 8490
rect 5145 8456 5179 8490
rect 5213 8456 5247 8490
rect 5281 8456 5315 8490
rect 5349 8456 5383 8490
rect 5417 8456 5451 8490
rect 5485 8456 5519 8490
rect 5553 8456 5587 8490
rect 5621 8456 5655 8490
rect 5689 8456 5723 8490
rect 5757 8456 5791 8490
rect 5825 8456 5859 8490
rect 5893 8456 5927 8490
rect 5961 8456 5995 8490
rect 6029 8456 6063 8490
rect 6097 8456 6131 8490
rect 6165 8456 6199 8490
rect 6233 8456 6267 8490
rect 6301 8456 6335 8490
rect 6369 8456 6403 8490
rect 6437 8456 6471 8490
rect 6505 8456 6539 8490
rect 6573 8456 6607 8490
rect 6641 8456 6675 8490
rect 6709 8456 6743 8490
rect 6777 8456 6811 8490
rect 6845 8456 6879 8490
rect 6913 8456 6947 8490
rect 6981 8456 7015 8490
rect 7049 8456 7083 8490
rect 7117 8456 7151 8490
rect 7185 8456 7219 8490
rect 7253 8456 7287 8490
rect 7321 8456 7355 8490
rect 7389 8456 7423 8490
rect 7457 8456 7491 8490
rect 7525 8456 7559 8490
rect 7593 8456 7627 8490
rect 7661 8456 7695 8490
rect 7729 8456 7763 8490
rect 7797 8456 7831 8490
rect 7865 8456 7899 8490
rect 7933 8456 7967 8490
rect 8001 8456 8035 8490
rect 8069 8456 8103 8490
rect 8137 8456 8171 8490
rect 8205 8456 8239 8490
rect 8273 8456 8307 8490
rect 8341 8471 14932 8490
rect 14966 8471 15000 8505
rect 15034 8471 15068 8505
rect 8341 8456 15102 8471
rect 2899 8453 15102 8456
rect 2899 8420 8393 8453
rect 34 8324 136 8358
rect 34 8290 68 8324
rect 102 8290 136 8324
rect 34 8256 136 8290
rect 2899 8386 2933 8420
rect 2967 8386 3002 8420
rect 3036 8386 3071 8420
rect 3105 8386 3139 8420
rect 3173 8386 3207 8420
rect 3241 8386 3275 8420
rect 3309 8386 3343 8420
rect 3377 8386 3411 8420
rect 3445 8386 3479 8420
rect 3513 8386 3547 8420
rect 3581 8386 3615 8420
rect 3649 8386 3683 8420
rect 3717 8386 3751 8420
rect 3785 8386 3819 8420
rect 3853 8386 3887 8420
rect 3921 8386 3955 8420
rect 3989 8386 4023 8420
rect 4057 8386 4091 8420
rect 4125 8386 4159 8420
rect 4193 8386 4227 8420
rect 4261 8386 4295 8420
rect 4329 8386 4363 8420
rect 4397 8386 4431 8420
rect 4465 8386 4499 8420
rect 4533 8386 4567 8420
rect 4601 8386 4635 8420
rect 4669 8386 4703 8420
rect 4737 8386 4771 8420
rect 4805 8386 4839 8420
rect 4873 8386 4907 8420
rect 4941 8386 4975 8420
rect 5009 8386 5043 8420
rect 5077 8386 5111 8420
rect 5145 8386 5179 8420
rect 5213 8386 5247 8420
rect 5281 8386 5315 8420
rect 5349 8386 5383 8420
rect 5417 8386 5451 8420
rect 5485 8386 5519 8420
rect 5553 8386 5587 8420
rect 5621 8386 5655 8420
rect 5689 8386 5723 8420
rect 5757 8386 5791 8420
rect 5825 8386 5859 8420
rect 5893 8386 5927 8420
rect 5961 8386 5995 8420
rect 6029 8386 6063 8420
rect 6097 8386 6131 8420
rect 6165 8386 6199 8420
rect 6233 8386 6267 8420
rect 6301 8386 6335 8420
rect 6369 8386 6403 8420
rect 6437 8386 6471 8420
rect 6505 8386 6539 8420
rect 6573 8386 6607 8420
rect 6641 8386 6675 8420
rect 6709 8386 6743 8420
rect 6777 8386 6811 8420
rect 6845 8386 6879 8420
rect 6913 8386 6947 8420
rect 6981 8386 7015 8420
rect 7049 8386 7083 8420
rect 7117 8386 7151 8420
rect 7185 8386 7219 8420
rect 7253 8386 7287 8420
rect 7321 8386 7355 8420
rect 7389 8386 7423 8420
rect 7457 8386 7491 8420
rect 7525 8386 7559 8420
rect 7593 8386 7627 8420
rect 7661 8386 7695 8420
rect 7729 8386 7763 8420
rect 7797 8386 7831 8420
rect 7865 8386 7899 8420
rect 7933 8386 7967 8420
rect 8001 8386 8035 8420
rect 8069 8386 8103 8420
rect 8137 8386 8171 8420
rect 8205 8386 8239 8420
rect 8273 8386 8307 8420
rect 8341 8419 8393 8420
rect 8427 8419 8462 8453
rect 8496 8419 8531 8453
rect 8565 8419 8600 8453
rect 8634 8419 8669 8453
rect 8703 8419 8738 8453
rect 8772 8419 8807 8453
rect 8841 8419 8876 8453
rect 8910 8419 8945 8453
rect 8979 8419 9014 8453
rect 9048 8419 9083 8453
rect 9117 8419 9152 8453
rect 9186 8419 9220 8453
rect 9254 8419 9288 8453
rect 9322 8419 9356 8453
rect 9390 8419 9424 8453
rect 9458 8419 9492 8453
rect 9526 8419 9560 8453
rect 9594 8419 9628 8453
rect 9662 8419 9696 8453
rect 9730 8419 9764 8453
rect 9798 8419 9832 8453
rect 9866 8419 9900 8453
rect 9934 8419 9968 8453
rect 10002 8419 10036 8453
rect 10070 8419 10104 8453
rect 10138 8419 10172 8453
rect 10206 8419 10240 8453
rect 10274 8419 10308 8453
rect 10342 8419 10376 8453
rect 10410 8419 10444 8453
rect 10478 8419 10512 8453
rect 10546 8419 10580 8453
rect 10614 8419 10648 8453
rect 10682 8419 10716 8453
rect 10750 8419 10784 8453
rect 10818 8419 10852 8453
rect 10886 8419 10920 8453
rect 10954 8419 10988 8453
rect 11022 8419 11056 8453
rect 11090 8419 11124 8453
rect 11158 8419 11192 8453
rect 11226 8419 11260 8453
rect 11294 8419 11328 8453
rect 11362 8419 11396 8453
rect 11430 8419 11464 8453
rect 11498 8419 11532 8453
rect 11566 8419 11600 8453
rect 11634 8419 11668 8453
rect 11702 8419 11736 8453
rect 11770 8419 11804 8453
rect 11838 8419 11872 8453
rect 11906 8419 11940 8453
rect 11974 8419 12008 8453
rect 12042 8419 12076 8453
rect 12110 8419 12144 8453
rect 12178 8419 12212 8453
rect 12246 8419 12280 8453
rect 12314 8419 12348 8453
rect 12382 8419 12416 8453
rect 12450 8419 12484 8453
rect 12518 8419 12552 8453
rect 12586 8419 12620 8453
rect 12654 8419 12688 8453
rect 12722 8419 12756 8453
rect 12790 8419 12824 8453
rect 12858 8419 12892 8453
rect 12926 8419 12960 8453
rect 12994 8419 13028 8453
rect 13062 8419 13096 8453
rect 13130 8419 13164 8453
rect 13198 8419 13232 8453
rect 13266 8419 13300 8453
rect 13334 8419 13368 8453
rect 13402 8419 13436 8453
rect 13470 8419 13504 8453
rect 13538 8419 13572 8453
rect 13606 8419 13640 8453
rect 13674 8419 13708 8453
rect 13742 8419 13776 8453
rect 13810 8419 13844 8453
rect 13878 8419 13912 8453
rect 13946 8419 13980 8453
rect 14014 8419 14048 8453
rect 14082 8419 14116 8453
rect 14150 8419 14184 8453
rect 14218 8419 14252 8453
rect 14286 8419 14320 8453
rect 14354 8419 14388 8453
rect 14422 8419 14456 8453
rect 14490 8419 14524 8453
rect 14558 8419 14592 8453
rect 14626 8419 14660 8453
rect 14694 8419 14728 8453
rect 14762 8419 14796 8453
rect 14830 8419 14864 8453
rect 14898 8433 15102 8453
rect 14898 8419 14932 8433
rect 8341 8399 14932 8419
rect 14966 8399 15000 8433
rect 15034 8399 15068 8433
rect 8341 8386 15102 8399
rect 2899 8383 15102 8386
rect 2899 8350 8375 8383
rect 2899 8316 2933 8350
rect 2967 8316 3002 8350
rect 3036 8316 3071 8350
rect 3105 8316 3139 8350
rect 3173 8316 3207 8350
rect 3241 8316 3275 8350
rect 3309 8316 3343 8350
rect 3377 8316 3411 8350
rect 3445 8316 3479 8350
rect 3513 8316 3547 8350
rect 3581 8316 3615 8350
rect 3649 8316 3683 8350
rect 3717 8316 3751 8350
rect 3785 8316 3819 8350
rect 3853 8316 3887 8350
rect 3921 8316 3955 8350
rect 3989 8316 4023 8350
rect 4057 8316 4091 8350
rect 4125 8316 4159 8350
rect 4193 8316 4227 8350
rect 4261 8316 4295 8350
rect 4329 8316 4363 8350
rect 4397 8316 4431 8350
rect 4465 8316 4499 8350
rect 4533 8316 4567 8350
rect 4601 8316 4635 8350
rect 4669 8316 4703 8350
rect 4737 8316 4771 8350
rect 4805 8316 4839 8350
rect 4873 8316 4907 8350
rect 4941 8316 4975 8350
rect 5009 8316 5043 8350
rect 5077 8316 5111 8350
rect 5145 8316 5179 8350
rect 5213 8316 5247 8350
rect 5281 8316 5315 8350
rect 5349 8316 5383 8350
rect 5417 8316 5451 8350
rect 5485 8316 5519 8350
rect 5553 8316 5587 8350
rect 5621 8316 5655 8350
rect 5689 8316 5723 8350
rect 5757 8316 5791 8350
rect 5825 8316 5859 8350
rect 5893 8316 5927 8350
rect 5961 8316 5995 8350
rect 6029 8316 6063 8350
rect 6097 8316 6131 8350
rect 6165 8316 6199 8350
rect 6233 8316 6267 8350
rect 6301 8316 6335 8350
rect 6369 8316 6403 8350
rect 6437 8316 6471 8350
rect 6505 8316 6539 8350
rect 6573 8316 6607 8350
rect 6641 8316 6675 8350
rect 6709 8316 6743 8350
rect 6777 8316 6811 8350
rect 6845 8316 6879 8350
rect 6913 8316 6947 8350
rect 6981 8316 7015 8350
rect 7049 8316 7083 8350
rect 7117 8316 7151 8350
rect 7185 8316 7219 8350
rect 7253 8316 7287 8350
rect 7321 8316 7355 8350
rect 7389 8316 7423 8350
rect 7457 8316 7491 8350
rect 7525 8316 7559 8350
rect 7593 8316 7627 8350
rect 7661 8316 7695 8350
rect 7729 8316 7763 8350
rect 7797 8316 7831 8350
rect 7865 8316 7899 8350
rect 7933 8316 7967 8350
rect 8001 8316 8035 8350
rect 8069 8316 8103 8350
rect 8137 8316 8171 8350
rect 8205 8316 8239 8350
rect 8273 8316 8307 8350
rect 8341 8316 8375 8350
rect 34 8222 68 8256
rect 102 8222 136 8256
rect 34 8192 136 8222
rect 2899 8280 8375 8316
rect 13498 8361 15102 8383
rect 13498 8357 14932 8361
rect 13498 8323 13532 8357
rect 13566 8323 13603 8357
rect 13637 8323 13674 8357
rect 13708 8323 13744 8357
rect 13778 8323 13814 8357
rect 13848 8323 13884 8357
rect 13918 8323 13954 8357
rect 13988 8323 14024 8357
rect 14058 8323 14094 8357
rect 14128 8323 14164 8357
rect 14198 8323 14234 8357
rect 14268 8323 14304 8357
rect 14338 8323 14374 8357
rect 14408 8323 14444 8357
rect 14478 8323 14514 8357
rect 14548 8323 14584 8357
rect 14618 8323 14654 8357
rect 14688 8323 14724 8357
rect 14758 8323 14794 8357
rect 14828 8323 14864 8357
rect 14898 8327 14932 8357
rect 14966 8327 15000 8361
rect 15034 8327 15068 8361
rect 14898 8323 15102 8327
rect 13498 8289 15102 8323
rect 2899 8246 2933 8280
rect 2967 8246 3002 8280
rect 3036 8246 3071 8280
rect 3105 8246 3139 8280
rect 3173 8246 3207 8280
rect 3241 8246 3275 8280
rect 3309 8246 3343 8280
rect 3377 8246 3411 8280
rect 3445 8246 3479 8280
rect 3513 8246 3547 8280
rect 3581 8246 3615 8280
rect 3649 8246 3683 8280
rect 3717 8246 3751 8280
rect 3785 8246 3819 8280
rect 3853 8246 3887 8280
rect 3921 8246 3955 8280
rect 3989 8246 4023 8280
rect 4057 8246 4091 8280
rect 4125 8246 4159 8280
rect 4193 8246 4227 8280
rect 4261 8246 4295 8280
rect 4329 8246 4363 8280
rect 4397 8246 4431 8280
rect 4465 8246 4499 8280
rect 4533 8246 4567 8280
rect 4601 8246 4635 8280
rect 4669 8246 4703 8280
rect 4737 8246 4771 8280
rect 4805 8246 4839 8280
rect 4873 8246 4907 8280
rect 4941 8246 4975 8280
rect 5009 8246 5043 8280
rect 5077 8246 5111 8280
rect 5145 8246 5179 8280
rect 5213 8246 5247 8280
rect 5281 8246 5315 8280
rect 5349 8246 5383 8280
rect 5417 8246 5451 8280
rect 5485 8246 5519 8280
rect 5553 8246 5587 8280
rect 5621 8246 5655 8280
rect 5689 8246 5723 8280
rect 5757 8246 5791 8280
rect 5825 8246 5859 8280
rect 5893 8246 5927 8280
rect 5961 8246 5995 8280
rect 6029 8246 6063 8280
rect 6097 8246 6131 8280
rect 6165 8246 6199 8280
rect 6233 8246 6267 8280
rect 6301 8246 6335 8280
rect 6369 8246 6403 8280
rect 6437 8246 6471 8280
rect 6505 8246 6539 8280
rect 6573 8246 6607 8280
rect 6641 8246 6675 8280
rect 6709 8246 6743 8280
rect 6777 8246 6811 8280
rect 6845 8246 6879 8280
rect 6913 8246 6947 8280
rect 6981 8246 7015 8280
rect 7049 8246 7083 8280
rect 7117 8246 7151 8280
rect 7185 8246 7219 8280
rect 7253 8246 7287 8280
rect 7321 8246 7355 8280
rect 7389 8246 7423 8280
rect 7457 8246 7491 8280
rect 7525 8246 7559 8280
rect 7593 8246 7627 8280
rect 7661 8246 7695 8280
rect 7729 8246 7763 8280
rect 7797 8246 7831 8280
rect 7865 8246 7899 8280
rect 7933 8246 7967 8280
rect 8001 8246 8035 8280
rect 8069 8246 8103 8280
rect 8137 8246 8171 8280
rect 8205 8246 8239 8280
rect 8273 8246 8307 8280
rect 8341 8246 8375 8280
rect 2899 8210 8375 8246
rect 2899 8192 2933 8210
rect 34 8176 2933 8192
rect 2967 8176 3002 8210
rect 3036 8176 3071 8210
rect 3105 8176 3139 8210
rect 3173 8176 3207 8210
rect 3241 8176 3275 8210
rect 3309 8176 3343 8210
rect 3377 8176 3411 8210
rect 3445 8176 3479 8210
rect 3513 8176 3547 8210
rect 3581 8176 3615 8210
rect 3649 8176 3683 8210
rect 3717 8176 3751 8210
rect 3785 8176 3819 8210
rect 3853 8176 3887 8210
rect 3921 8176 3955 8210
rect 3989 8176 4023 8210
rect 4057 8176 4091 8210
rect 4125 8176 4159 8210
rect 4193 8176 4227 8210
rect 4261 8176 4295 8210
rect 4329 8176 4363 8210
rect 4397 8176 4431 8210
rect 4465 8176 4499 8210
rect 4533 8176 4567 8210
rect 4601 8176 4635 8210
rect 4669 8176 4703 8210
rect 4737 8176 4771 8210
rect 4805 8176 4839 8210
rect 4873 8176 4907 8210
rect 4941 8176 4975 8210
rect 5009 8176 5043 8210
rect 5077 8176 5111 8210
rect 5145 8176 5179 8210
rect 5213 8176 5247 8210
rect 5281 8176 5315 8210
rect 5349 8176 5383 8210
rect 5417 8176 5451 8210
rect 5485 8176 5519 8210
rect 5553 8176 5587 8210
rect 5621 8176 5655 8210
rect 5689 8176 5723 8210
rect 5757 8176 5791 8210
rect 5825 8176 5859 8210
rect 5893 8176 5927 8210
rect 5961 8176 5995 8210
rect 6029 8176 6063 8210
rect 6097 8176 6131 8210
rect 6165 8176 6199 8210
rect 6233 8176 6267 8210
rect 6301 8176 6335 8210
rect 6369 8176 6403 8210
rect 6437 8176 6471 8210
rect 6505 8176 6539 8210
rect 6573 8176 6607 8210
rect 6641 8176 6675 8210
rect 6709 8176 6743 8210
rect 6777 8176 6811 8210
rect 6845 8176 6879 8210
rect 6913 8176 6947 8210
rect 6981 8176 7015 8210
rect 7049 8176 7083 8210
rect 7117 8176 7151 8210
rect 7185 8176 7219 8210
rect 7253 8176 7287 8210
rect 7321 8176 7355 8210
rect 7389 8176 7423 8210
rect 7457 8176 7491 8210
rect 7525 8176 7559 8210
rect 7593 8176 7627 8210
rect 7661 8176 7695 8210
rect 7729 8176 7763 8210
rect 7797 8176 7831 8210
rect 7865 8176 7899 8210
rect 7933 8176 7967 8210
rect 8001 8176 8035 8210
rect 8069 8176 8103 8210
rect 8137 8176 8171 8210
rect 8205 8176 8239 8210
rect 8273 8176 8307 8210
rect 8341 8176 8375 8210
rect 34 8157 8375 8176
rect 34 8123 68 8157
rect 102 8123 138 8157
rect 172 8123 208 8157
rect 242 8123 278 8157
rect 312 8123 348 8157
rect 382 8123 418 8157
rect 452 8123 488 8157
rect 522 8123 558 8157
rect 592 8123 628 8157
rect 662 8123 698 8157
rect 732 8123 768 8157
rect 802 8123 838 8157
rect 872 8123 908 8157
rect 942 8123 978 8157
rect 1012 8123 1048 8157
rect 1082 8123 1118 8157
rect 1152 8123 1188 8157
rect 1222 8123 1258 8157
rect 1292 8123 1328 8157
rect 1362 8123 1398 8157
rect 1432 8123 1467 8157
rect 1501 8123 1536 8157
rect 1570 8123 1605 8157
rect 1639 8123 1674 8157
rect 1708 8123 1743 8157
rect 1777 8123 1812 8157
rect 1846 8123 1881 8157
rect 1915 8123 1950 8157
rect 1984 8123 2019 8157
rect 2053 8123 2088 8157
rect 2122 8123 2157 8157
rect 2191 8123 2226 8157
rect 2260 8123 2295 8157
rect 2329 8123 2364 8157
rect 2398 8123 2433 8157
rect 2467 8123 2502 8157
rect 2536 8123 2571 8157
rect 2605 8123 2640 8157
rect 2674 8123 2709 8157
rect 2743 8123 2778 8157
rect 2812 8123 2847 8157
rect 2881 8140 8375 8157
rect 2881 8123 2933 8140
rect 34 8106 2933 8123
rect 2967 8106 3002 8140
rect 3036 8106 3071 8140
rect 3105 8106 3139 8140
rect 3173 8106 3207 8140
rect 3241 8106 3275 8140
rect 3309 8106 3343 8140
rect 3377 8106 3411 8140
rect 3445 8106 3479 8140
rect 3513 8106 3547 8140
rect 3581 8106 3615 8140
rect 3649 8106 3683 8140
rect 3717 8106 3751 8140
rect 3785 8106 3819 8140
rect 3853 8106 3887 8140
rect 3921 8106 3955 8140
rect 3989 8106 4023 8140
rect 4057 8106 4091 8140
rect 4125 8106 4159 8140
rect 4193 8106 4227 8140
rect 4261 8106 4295 8140
rect 4329 8106 4363 8140
rect 4397 8106 4431 8140
rect 4465 8106 4499 8140
rect 4533 8106 4567 8140
rect 4601 8106 4635 8140
rect 4669 8106 4703 8140
rect 4737 8106 4771 8140
rect 4805 8106 4839 8140
rect 4873 8106 4907 8140
rect 4941 8106 4975 8140
rect 5009 8106 5043 8140
rect 5077 8106 5111 8140
rect 5145 8106 5179 8140
rect 5213 8106 5247 8140
rect 5281 8106 5315 8140
rect 5349 8106 5383 8140
rect 5417 8106 5451 8140
rect 5485 8106 5519 8140
rect 5553 8106 5587 8140
rect 5621 8106 5655 8140
rect 5689 8106 5723 8140
rect 5757 8106 5791 8140
rect 5825 8106 5859 8140
rect 5893 8106 5927 8140
rect 5961 8106 5995 8140
rect 6029 8106 6063 8140
rect 6097 8106 6131 8140
rect 6165 8106 6199 8140
rect 6233 8106 6267 8140
rect 6301 8106 6335 8140
rect 6369 8106 6403 8140
rect 6437 8106 6471 8140
rect 6505 8106 6539 8140
rect 6573 8106 6607 8140
rect 6641 8106 6675 8140
rect 6709 8106 6743 8140
rect 6777 8106 6811 8140
rect 6845 8106 6879 8140
rect 6913 8106 6947 8140
rect 6981 8106 7015 8140
rect 7049 8106 7083 8140
rect 7117 8106 7151 8140
rect 7185 8106 7219 8140
rect 7253 8106 7287 8140
rect 7321 8106 7355 8140
rect 7389 8106 7423 8140
rect 7457 8106 7491 8140
rect 7525 8106 7559 8140
rect 7593 8106 7627 8140
rect 7661 8106 7695 8140
rect 7729 8106 7763 8140
rect 7797 8106 7831 8140
rect 7865 8106 7899 8140
rect 7933 8106 7967 8140
rect 8001 8106 8035 8140
rect 8069 8106 8103 8140
rect 8137 8106 8171 8140
rect 8205 8106 8239 8140
rect 8273 8106 8307 8140
rect 8341 8106 8375 8140
rect 34 8082 8375 8106
rect 34 8048 68 8082
rect 102 8048 138 8082
rect 172 8048 208 8082
rect 242 8048 278 8082
rect 312 8048 348 8082
rect 382 8048 418 8082
rect 452 8048 488 8082
rect 522 8048 558 8082
rect 592 8048 628 8082
rect 662 8048 698 8082
rect 732 8048 768 8082
rect 802 8048 838 8082
rect 872 8048 908 8082
rect 942 8048 978 8082
rect 1012 8048 1048 8082
rect 1082 8048 1118 8082
rect 1152 8048 1188 8082
rect 1222 8048 1258 8082
rect 1292 8048 1328 8082
rect 1362 8048 1398 8082
rect 1432 8048 1467 8082
rect 1501 8048 1536 8082
rect 1570 8048 1605 8082
rect 1639 8048 1674 8082
rect 1708 8048 1743 8082
rect 1777 8048 1812 8082
rect 1846 8048 1881 8082
rect 1915 8048 1950 8082
rect 1984 8048 2019 8082
rect 2053 8048 2088 8082
rect 2122 8048 2157 8082
rect 2191 8048 2226 8082
rect 2260 8048 2295 8082
rect 2329 8048 2364 8082
rect 2398 8048 2433 8082
rect 2467 8048 2502 8082
rect 2536 8048 2571 8082
rect 2605 8048 2640 8082
rect 2674 8048 2709 8082
rect 2743 8048 2778 8082
rect 2812 8048 2847 8082
rect 2881 8070 8375 8082
rect 2881 8048 2933 8070
rect 34 8036 2933 8048
rect 2967 8036 3002 8070
rect 3036 8036 3071 8070
rect 3105 8036 3139 8070
rect 3173 8036 3207 8070
rect 3241 8036 3275 8070
rect 3309 8036 3343 8070
rect 3377 8036 3411 8070
rect 3445 8036 3479 8070
rect 3513 8036 3547 8070
rect 3581 8036 3615 8070
rect 3649 8036 3683 8070
rect 3717 8036 3751 8070
rect 3785 8036 3819 8070
rect 3853 8036 3887 8070
rect 3921 8036 3955 8070
rect 3989 8036 4023 8070
rect 4057 8036 4091 8070
rect 4125 8036 4159 8070
rect 4193 8036 4227 8070
rect 4261 8036 4295 8070
rect 4329 8036 4363 8070
rect 4397 8036 4431 8070
rect 4465 8036 4499 8070
rect 4533 8036 4567 8070
rect 4601 8036 4635 8070
rect 4669 8036 4703 8070
rect 4737 8036 4771 8070
rect 4805 8036 4839 8070
rect 4873 8036 4907 8070
rect 4941 8036 4975 8070
rect 5009 8036 5043 8070
rect 5077 8036 5111 8070
rect 5145 8036 5179 8070
rect 5213 8036 5247 8070
rect 5281 8036 5315 8070
rect 5349 8036 5383 8070
rect 5417 8036 5451 8070
rect 5485 8036 5519 8070
rect 5553 8036 5587 8070
rect 5621 8036 5655 8070
rect 5689 8036 5723 8070
rect 5757 8036 5791 8070
rect 5825 8036 5859 8070
rect 5893 8036 5927 8070
rect 5961 8036 5995 8070
rect 6029 8036 6063 8070
rect 6097 8036 6131 8070
rect 6165 8036 6199 8070
rect 6233 8036 6267 8070
rect 6301 8036 6335 8070
rect 6369 8036 6403 8070
rect 6437 8036 6471 8070
rect 6505 8036 6539 8070
rect 6573 8036 6607 8070
rect 6641 8036 6675 8070
rect 6709 8036 6743 8070
rect 6777 8036 6811 8070
rect 6845 8036 6879 8070
rect 6913 8036 6947 8070
rect 6981 8036 7015 8070
rect 7049 8036 7083 8070
rect 7117 8036 7151 8070
rect 7185 8036 7219 8070
rect 7253 8036 7287 8070
rect 7321 8036 7355 8070
rect 7389 8036 7423 8070
rect 7457 8036 7491 8070
rect 7525 8036 7559 8070
rect 7593 8036 7627 8070
rect 7661 8036 7695 8070
rect 7729 8036 7763 8070
rect 7797 8036 7831 8070
rect 7865 8036 7899 8070
rect 7933 8036 7967 8070
rect 8001 8036 8035 8070
rect 8069 8036 8103 8070
rect 8137 8036 8171 8070
rect 8205 8036 8239 8070
rect 8273 8036 8307 8070
rect 8341 8036 8375 8070
rect 34 8007 8375 8036
rect 34 7973 68 8007
rect 102 7973 138 8007
rect 172 7973 208 8007
rect 242 7973 278 8007
rect 312 7973 348 8007
rect 382 7973 418 8007
rect 452 7973 488 8007
rect 522 7973 558 8007
rect 592 7973 628 8007
rect 662 7973 698 8007
rect 732 7973 768 8007
rect 802 7973 838 8007
rect 872 7973 908 8007
rect 942 7973 978 8007
rect 1012 7973 1048 8007
rect 1082 7973 1118 8007
rect 1152 7973 1188 8007
rect 1222 7973 1258 8007
rect 1292 7973 1328 8007
rect 1362 7973 1398 8007
rect 1432 7973 1467 8007
rect 1501 7973 1536 8007
rect 1570 7973 1605 8007
rect 1639 7973 1674 8007
rect 1708 7973 1743 8007
rect 1777 7973 1812 8007
rect 1846 7973 1881 8007
rect 1915 7973 1950 8007
rect 1984 7973 2019 8007
rect 2053 7973 2088 8007
rect 2122 7973 2157 8007
rect 2191 7973 2226 8007
rect 2260 7973 2295 8007
rect 2329 7973 2364 8007
rect 2398 7973 2433 8007
rect 2467 7973 2502 8007
rect 2536 7973 2571 8007
rect 2605 7973 2640 8007
rect 2674 7973 2709 8007
rect 2743 7973 2778 8007
rect 2812 7973 2847 8007
rect 2881 8000 8375 8007
rect 2881 7973 2933 8000
rect 34 7966 2933 7973
rect 2967 7966 3002 8000
rect 3036 7966 3071 8000
rect 3105 7966 3139 8000
rect 3173 7966 3207 8000
rect 3241 7966 3275 8000
rect 3309 7966 3343 8000
rect 3377 7966 3411 8000
rect 3445 7966 3479 8000
rect 3513 7966 3547 8000
rect 3581 7966 3615 8000
rect 3649 7966 3683 8000
rect 3717 7966 3751 8000
rect 3785 7966 3819 8000
rect 3853 7966 3887 8000
rect 3921 7966 3955 8000
rect 3989 7966 4023 8000
rect 4057 7966 4091 8000
rect 4125 7966 4159 8000
rect 4193 7966 4227 8000
rect 4261 7966 4295 8000
rect 4329 7966 4363 8000
rect 4397 7966 4431 8000
rect 4465 7966 4499 8000
rect 4533 7966 4567 8000
rect 4601 7966 4635 8000
rect 4669 7966 4703 8000
rect 4737 7966 4771 8000
rect 4805 7966 4839 8000
rect 4873 7966 4907 8000
rect 4941 7966 4975 8000
rect 5009 7966 5043 8000
rect 5077 7966 5111 8000
rect 5145 7966 5179 8000
rect 5213 7966 5247 8000
rect 5281 7966 5315 8000
rect 5349 7966 5383 8000
rect 5417 7966 5451 8000
rect 5485 7966 5519 8000
rect 5553 7966 5587 8000
rect 5621 7966 5655 8000
rect 5689 7966 5723 8000
rect 5757 7966 5791 8000
rect 5825 7966 5859 8000
rect 5893 7966 5927 8000
rect 5961 7966 5995 8000
rect 6029 7966 6063 8000
rect 6097 7966 6131 8000
rect 6165 7966 6199 8000
rect 6233 7966 6267 8000
rect 6301 7966 6335 8000
rect 6369 7966 6403 8000
rect 6437 7966 6471 8000
rect 6505 7966 6539 8000
rect 6573 7966 6607 8000
rect 6641 7966 6675 8000
rect 6709 7966 6743 8000
rect 6777 7966 6811 8000
rect 6845 7966 6879 8000
rect 6913 7966 6947 8000
rect 6981 7966 7015 8000
rect 7049 7966 7083 8000
rect 7117 7966 7151 8000
rect 7185 7966 7219 8000
rect 7253 7966 7287 8000
rect 7321 7966 7355 8000
rect 7389 7966 7423 8000
rect 7457 7966 7491 8000
rect 7525 7966 7559 8000
rect 7593 7966 7627 8000
rect 7661 7966 7695 8000
rect 7729 7966 7763 8000
rect 7797 7966 7831 8000
rect 7865 7966 7899 8000
rect 7933 7966 7967 8000
rect 8001 7966 8035 8000
rect 8069 7966 8103 8000
rect 8137 7966 8171 8000
rect 8205 7966 8239 8000
rect 8273 7966 8307 8000
rect 8341 7966 8375 8000
rect 34 7932 8375 7966
rect 34 7898 68 7932
rect 102 7898 138 7932
rect 172 7898 208 7932
rect 242 7898 278 7932
rect 312 7898 348 7932
rect 382 7898 418 7932
rect 452 7898 488 7932
rect 522 7898 558 7932
rect 592 7898 628 7932
rect 662 7898 698 7932
rect 732 7898 768 7932
rect 802 7898 838 7932
rect 872 7898 908 7932
rect 942 7898 978 7932
rect 1012 7898 1048 7932
rect 1082 7898 1118 7932
rect 1152 7898 1188 7932
rect 1222 7898 1258 7932
rect 1292 7898 1328 7932
rect 1362 7898 1398 7932
rect 1432 7898 1467 7932
rect 1501 7898 1536 7932
rect 1570 7898 1605 7932
rect 1639 7898 1674 7932
rect 1708 7898 1743 7932
rect 1777 7898 1812 7932
rect 1846 7898 1881 7932
rect 1915 7898 1950 7932
rect 1984 7898 2019 7932
rect 2053 7898 2088 7932
rect 2122 7898 2157 7932
rect 2191 7898 2226 7932
rect 2260 7898 2295 7932
rect 2329 7898 2364 7932
rect 2398 7898 2433 7932
rect 2467 7898 2502 7932
rect 2536 7898 2571 7932
rect 2605 7898 2640 7932
rect 2674 7898 2709 7932
rect 2743 7898 2778 7932
rect 2812 7898 2847 7932
rect 2881 7930 8375 7932
rect 2881 7898 2933 7930
rect 34 7896 2933 7898
rect 2967 7896 3002 7930
rect 3036 7896 3071 7930
rect 3105 7896 3139 7930
rect 3173 7896 3207 7930
rect 3241 7896 3275 7930
rect 3309 7896 3343 7930
rect 3377 7896 3411 7930
rect 3445 7896 3479 7930
rect 3513 7896 3547 7930
rect 3581 7896 3615 7930
rect 3649 7896 3683 7930
rect 3717 7896 3751 7930
rect 3785 7896 3819 7930
rect 3853 7896 3887 7930
rect 3921 7896 3955 7930
rect 3989 7896 4023 7930
rect 4057 7896 4091 7930
rect 4125 7896 4159 7930
rect 4193 7896 4227 7930
rect 4261 7896 4295 7930
rect 4329 7896 4363 7930
rect 4397 7896 4431 7930
rect 4465 7896 4499 7930
rect 4533 7896 4567 7930
rect 4601 7896 4635 7930
rect 4669 7896 4703 7930
rect 4737 7896 4771 7930
rect 4805 7896 4839 7930
rect 4873 7896 4907 7930
rect 4941 7896 4975 7930
rect 5009 7896 5043 7930
rect 5077 7896 5111 7930
rect 5145 7896 5179 7930
rect 5213 7896 5247 7930
rect 5281 7896 5315 7930
rect 5349 7896 5383 7930
rect 5417 7896 5451 7930
rect 5485 7896 5519 7930
rect 5553 7896 5587 7930
rect 5621 7896 5655 7930
rect 5689 7896 5723 7930
rect 5757 7896 5791 7930
rect 5825 7896 5859 7930
rect 5893 7896 5927 7930
rect 5961 7896 5995 7930
rect 6029 7896 6063 7930
rect 6097 7896 6131 7930
rect 6165 7896 6199 7930
rect 6233 7896 6267 7930
rect 6301 7896 6335 7930
rect 6369 7896 6403 7930
rect 6437 7896 6471 7930
rect 6505 7896 6539 7930
rect 6573 7896 6607 7930
rect 6641 7896 6675 7930
rect 6709 7896 6743 7930
rect 6777 7896 6811 7930
rect 6845 7896 6879 7930
rect 6913 7896 6947 7930
rect 6981 7896 7015 7930
rect 7049 7896 7083 7930
rect 7117 7896 7151 7930
rect 7185 7896 7219 7930
rect 7253 7896 7287 7930
rect 7321 7896 7355 7930
rect 7389 7896 7423 7930
rect 7457 7896 7491 7930
rect 7525 7896 7559 7930
rect 7593 7896 7627 7930
rect 7661 7896 7695 7930
rect 7729 7896 7763 7930
rect 7797 7896 7831 7930
rect 7865 7896 7899 7930
rect 7933 7896 7967 7930
rect 8001 7896 8035 7930
rect 8069 7896 8103 7930
rect 8137 7896 8171 7930
rect 8205 7896 8239 7930
rect 8273 7896 8307 7930
rect 8341 7896 8375 7930
rect 34 7860 8375 7896
rect 13498 8283 14932 8289
rect 13498 8249 13532 8283
rect 13566 8249 13603 8283
rect 13637 8249 13674 8283
rect 13708 8249 13744 8283
rect 13778 8249 13814 8283
rect 13848 8249 13884 8283
rect 13918 8249 13954 8283
rect 13988 8249 14024 8283
rect 14058 8249 14094 8283
rect 14128 8249 14164 8283
rect 14198 8249 14234 8283
rect 14268 8249 14304 8283
rect 14338 8249 14374 8283
rect 14408 8249 14444 8283
rect 14478 8249 14514 8283
rect 14548 8249 14584 8283
rect 14618 8249 14654 8283
rect 14688 8249 14724 8283
rect 14758 8249 14794 8283
rect 14828 8249 14864 8283
rect 14898 8255 14932 8283
rect 14966 8255 15000 8289
rect 15034 8255 15068 8289
rect 14898 8249 15102 8255
rect 13498 8217 15102 8249
rect 13498 8209 14932 8217
rect 13498 8175 13532 8209
rect 13566 8175 13603 8209
rect 13637 8175 13674 8209
rect 13708 8175 13744 8209
rect 13778 8175 13814 8209
rect 13848 8175 13884 8209
rect 13918 8175 13954 8209
rect 13988 8175 14024 8209
rect 14058 8175 14094 8209
rect 14128 8175 14164 8209
rect 14198 8175 14234 8209
rect 14268 8175 14304 8209
rect 14338 8175 14374 8209
rect 14408 8175 14444 8209
rect 14478 8175 14514 8209
rect 14548 8175 14584 8209
rect 14618 8175 14654 8209
rect 14688 8175 14724 8209
rect 14758 8175 14794 8209
rect 14828 8175 14864 8209
rect 14898 8183 14932 8209
rect 14966 8183 15000 8217
rect 15034 8183 15068 8217
rect 14898 8175 15102 8183
rect 13498 8145 15102 8175
rect 13498 8135 14932 8145
rect 13498 8101 13532 8135
rect 13566 8101 13603 8135
rect 13637 8101 13674 8135
rect 13708 8101 13744 8135
rect 13778 8101 13814 8135
rect 13848 8101 13884 8135
rect 13918 8101 13954 8135
rect 13988 8101 14024 8135
rect 14058 8101 14094 8135
rect 14128 8101 14164 8135
rect 14198 8101 14234 8135
rect 14268 8101 14304 8135
rect 14338 8101 14374 8135
rect 14408 8101 14444 8135
rect 14478 8101 14514 8135
rect 14548 8101 14584 8135
rect 14618 8101 14654 8135
rect 14688 8101 14724 8135
rect 14758 8101 14794 8135
rect 14828 8101 14864 8135
rect 14898 8111 14932 8135
rect 14966 8111 15000 8145
rect 15034 8111 15068 8145
rect 14898 8101 15102 8111
rect 13498 8073 15102 8101
rect 13498 8061 14932 8073
rect 13498 8027 13532 8061
rect 13566 8027 13603 8061
rect 13637 8027 13674 8061
rect 13708 8027 13744 8061
rect 13778 8027 13814 8061
rect 13848 8027 13884 8061
rect 13918 8027 13954 8061
rect 13988 8027 14024 8061
rect 14058 8027 14094 8061
rect 14128 8027 14164 8061
rect 14198 8027 14234 8061
rect 14268 8027 14304 8061
rect 14338 8027 14374 8061
rect 14408 8027 14444 8061
rect 14478 8027 14514 8061
rect 14548 8027 14584 8061
rect 14618 8027 14654 8061
rect 14688 8027 14724 8061
rect 14758 8027 14794 8061
rect 14828 8027 14864 8061
rect 14898 8039 14932 8061
rect 14966 8039 15000 8073
rect 15034 8039 15068 8073
rect 14898 8027 15102 8039
rect 13498 8001 15102 8027
rect 13498 7987 14932 8001
rect 13498 7953 13532 7987
rect 13566 7953 13603 7987
rect 13637 7953 13674 7987
rect 13708 7953 13744 7987
rect 13778 7953 13814 7987
rect 13848 7953 13884 7987
rect 13918 7953 13954 7987
rect 13988 7953 14024 7987
rect 14058 7953 14094 7987
rect 14128 7953 14164 7987
rect 14198 7953 14234 7987
rect 14268 7953 14304 7987
rect 14338 7953 14374 7987
rect 14408 7953 14444 7987
rect 14478 7953 14514 7987
rect 14548 7953 14584 7987
rect 14618 7953 14654 7987
rect 14688 7953 14724 7987
rect 14758 7953 14794 7987
rect 14828 7953 14864 7987
rect 14898 7967 14932 7987
rect 14966 7967 15000 8001
rect 15034 7967 15068 8001
rect 14898 7953 15102 7967
rect 13498 7929 15102 7953
rect 13498 7913 14932 7929
rect 34 7857 2933 7860
rect 34 7823 68 7857
rect 102 7823 138 7857
rect 172 7823 208 7857
rect 242 7823 278 7857
rect 312 7823 348 7857
rect 382 7823 418 7857
rect 452 7823 488 7857
rect 522 7823 558 7857
rect 592 7823 628 7857
rect 662 7823 698 7857
rect 732 7823 768 7857
rect 802 7823 838 7857
rect 872 7823 908 7857
rect 942 7823 978 7857
rect 1012 7823 1048 7857
rect 1082 7823 1118 7857
rect 1152 7823 1188 7857
rect 1222 7823 1258 7857
rect 1292 7823 1328 7857
rect 1362 7823 1398 7857
rect 1432 7823 1467 7857
rect 1501 7823 1536 7857
rect 1570 7823 1605 7857
rect 1639 7823 1674 7857
rect 1708 7823 1743 7857
rect 1777 7823 1812 7857
rect 1846 7823 1881 7857
rect 1915 7823 1950 7857
rect 1984 7823 2019 7857
rect 2053 7823 2088 7857
rect 2122 7823 2157 7857
rect 2191 7823 2226 7857
rect 2260 7823 2295 7857
rect 2329 7823 2364 7857
rect 2398 7823 2433 7857
rect 2467 7823 2502 7857
rect 2536 7823 2571 7857
rect 2605 7823 2640 7857
rect 2674 7823 2709 7857
rect 2743 7823 2778 7857
rect 2812 7823 2847 7857
rect 2881 7826 2933 7857
rect 2967 7826 3002 7860
rect 3036 7826 3071 7860
rect 3105 7826 3139 7860
rect 3173 7826 3207 7860
rect 3241 7826 3275 7860
rect 3309 7826 3343 7860
rect 3377 7826 3411 7860
rect 3445 7826 3479 7860
rect 3513 7826 3547 7860
rect 3581 7826 3615 7860
rect 3649 7826 3683 7860
rect 3717 7826 3751 7860
rect 3785 7826 3819 7860
rect 3853 7826 3887 7860
rect 3921 7826 3955 7860
rect 3989 7826 4023 7860
rect 4057 7826 4091 7860
rect 4125 7826 4159 7860
rect 4193 7826 4227 7860
rect 4261 7826 4295 7860
rect 4329 7826 4363 7860
rect 4397 7826 4431 7860
rect 4465 7826 4499 7860
rect 4533 7826 4567 7860
rect 4601 7826 4635 7860
rect 4669 7826 4703 7860
rect 4737 7826 4771 7860
rect 4805 7826 4839 7860
rect 4873 7826 4907 7860
rect 4941 7826 4975 7860
rect 5009 7826 5043 7860
rect 5077 7826 5111 7860
rect 5145 7826 5179 7860
rect 5213 7826 5247 7860
rect 5281 7826 5315 7860
rect 5349 7826 5383 7860
rect 5417 7826 5451 7860
rect 5485 7826 5519 7860
rect 5553 7826 5587 7860
rect 5621 7826 5655 7860
rect 5689 7826 5723 7860
rect 5757 7826 5791 7860
rect 5825 7826 5859 7860
rect 5893 7826 5927 7860
rect 5961 7826 5995 7860
rect 6029 7826 6063 7860
rect 6097 7826 6131 7860
rect 6165 7826 6199 7860
rect 6233 7826 6267 7860
rect 6301 7826 6335 7860
rect 6369 7826 6403 7860
rect 6437 7826 6471 7860
rect 6505 7826 6539 7860
rect 6573 7826 6607 7860
rect 6641 7826 6675 7860
rect 6709 7826 6743 7860
rect 6777 7826 6811 7860
rect 6845 7826 6879 7860
rect 6913 7826 6947 7860
rect 6981 7826 7015 7860
rect 7049 7826 7083 7860
rect 7117 7826 7151 7860
rect 7185 7826 7219 7860
rect 7253 7826 7287 7860
rect 7321 7826 7355 7860
rect 7389 7826 7423 7860
rect 7457 7826 7491 7860
rect 7525 7826 7559 7860
rect 7593 7826 7627 7860
rect 7661 7826 7695 7860
rect 7729 7826 7763 7860
rect 7797 7826 7831 7860
rect 7865 7826 7899 7860
rect 7933 7826 7967 7860
rect 8001 7826 8035 7860
rect 8069 7826 8103 7860
rect 8137 7826 8171 7860
rect 8205 7826 8239 7860
rect 8273 7826 8307 7860
rect 8341 7826 8375 7860
rect 2881 7823 8375 7826
rect 34 7788 8375 7823
rect 13498 7879 13532 7913
rect 13566 7879 13603 7913
rect 13637 7879 13674 7913
rect 13708 7879 13744 7913
rect 13778 7879 13814 7913
rect 13848 7879 13884 7913
rect 13918 7879 13954 7913
rect 13988 7879 14024 7913
rect 14058 7879 14094 7913
rect 14128 7879 14164 7913
rect 14198 7879 14234 7913
rect 14268 7879 14304 7913
rect 14338 7879 14374 7913
rect 14408 7879 14444 7913
rect 14478 7879 14514 7913
rect 14548 7879 14584 7913
rect 14618 7879 14654 7913
rect 14688 7879 14724 7913
rect 14758 7879 14794 7913
rect 14828 7879 14864 7913
rect 14898 7895 14932 7913
rect 14966 7895 15000 7929
rect 15034 7895 15068 7929
rect 14898 7879 15102 7895
rect 13498 7857 15102 7879
rect 13498 7839 14932 7857
rect 13498 7805 13532 7839
rect 13566 7805 13603 7839
rect 13637 7805 13674 7839
rect 13708 7805 13744 7839
rect 13778 7805 13814 7839
rect 13848 7805 13884 7839
rect 13918 7805 13954 7839
rect 13988 7805 14024 7839
rect 14058 7805 14094 7839
rect 14128 7805 14164 7839
rect 14198 7805 14234 7839
rect 14268 7805 14304 7839
rect 14338 7805 14374 7839
rect 14408 7805 14444 7839
rect 14478 7805 14514 7839
rect 14548 7805 14584 7839
rect 14618 7805 14654 7839
rect 14688 7805 14724 7839
rect 14758 7805 14794 7839
rect 14828 7805 14864 7839
rect 14898 7823 14932 7839
rect 14966 7823 15000 7857
rect 15034 7823 15068 7857
rect 14898 7805 15102 7823
rect 13498 7788 15102 7805
rect 34 7785 15102 7788
rect 34 7751 14932 7785
rect 14966 7751 15000 7785
rect 15034 7751 15068 7785
rect 34 7749 15102 7751
rect 34 7715 68 7749
rect 102 7715 137 7749
rect 171 7715 206 7749
rect 240 7715 275 7749
rect 309 7715 344 7749
rect 378 7715 413 7749
rect 447 7715 482 7749
rect 516 7715 551 7749
rect 585 7715 620 7749
rect 654 7715 689 7749
rect 723 7715 758 7749
rect 792 7715 827 7749
rect 861 7715 896 7749
rect 930 7715 965 7749
rect 999 7715 1034 7749
rect 1068 7715 1103 7749
rect 1137 7715 1172 7749
rect 1206 7715 1241 7749
rect 1275 7715 1310 7749
rect 1344 7715 1379 7749
rect 1413 7715 1448 7749
rect 1482 7715 1517 7749
rect 1551 7715 1586 7749
rect 1620 7715 1655 7749
rect 1689 7715 1724 7749
rect 1758 7715 1793 7749
rect 1827 7715 1862 7749
rect 1896 7715 1931 7749
rect 1965 7715 2000 7749
rect 2034 7715 2069 7749
rect 2103 7715 2138 7749
rect 2172 7715 2207 7749
rect 2241 7715 2276 7749
rect 2310 7715 2345 7749
rect 2379 7715 2414 7749
rect 2448 7715 2483 7749
rect 2517 7715 2552 7749
rect 2586 7715 2621 7749
rect 2655 7715 2690 7749
rect 2724 7715 2759 7749
rect 2793 7715 2828 7749
rect 2862 7715 2896 7749
rect 2930 7715 2964 7749
rect 2998 7715 3032 7749
rect 3066 7715 3100 7749
rect 3134 7715 3168 7749
rect 3202 7715 3236 7749
rect 3270 7715 3304 7749
rect 3338 7715 3372 7749
rect 3406 7715 3440 7749
rect 3474 7715 3508 7749
rect 3542 7715 3576 7749
rect 3610 7715 3644 7749
rect 3678 7715 3712 7749
rect 3746 7715 3780 7749
rect 3814 7715 3848 7749
rect 3882 7715 3916 7749
rect 3950 7715 3984 7749
rect 4018 7715 4052 7749
rect 4086 7715 4120 7749
rect 4154 7715 4188 7749
rect 4222 7715 4256 7749
rect 4290 7715 4324 7749
rect 4358 7715 4392 7749
rect 4426 7715 4460 7749
rect 4494 7715 4528 7749
rect 4562 7715 4596 7749
rect 4630 7715 4664 7749
rect 4698 7715 4732 7749
rect 4766 7715 4800 7749
rect 4834 7715 4868 7749
rect 4902 7715 4936 7749
rect 4970 7715 5004 7749
rect 5038 7715 5072 7749
rect 5106 7715 5140 7749
rect 5174 7715 5208 7749
rect 5242 7715 5276 7749
rect 5310 7715 5344 7749
rect 5378 7715 5412 7749
rect 5446 7715 5480 7749
rect 5514 7715 5548 7749
rect 5582 7715 5616 7749
rect 5650 7715 5684 7749
rect 5718 7715 5752 7749
rect 5786 7715 5820 7749
rect 5854 7715 5888 7749
rect 5922 7715 5956 7749
rect 5990 7715 6024 7749
rect 6058 7715 6092 7749
rect 6126 7715 6160 7749
rect 6194 7715 6228 7749
rect 6262 7715 6296 7749
rect 6330 7715 6364 7749
rect 6398 7715 6432 7749
rect 6466 7715 6500 7749
rect 6534 7715 6568 7749
rect 6602 7715 6636 7749
rect 6670 7715 6704 7749
rect 6738 7715 6772 7749
rect 6806 7715 6840 7749
rect 6874 7715 6908 7749
rect 6942 7715 6976 7749
rect 7010 7715 7044 7749
rect 7078 7715 7112 7749
rect 7146 7715 7180 7749
rect 7214 7715 7248 7749
rect 7282 7715 7316 7749
rect 7350 7715 7384 7749
rect 7418 7715 7452 7749
rect 7486 7715 7520 7749
rect 7554 7715 7588 7749
rect 7622 7715 7656 7749
rect 7690 7715 7724 7749
rect 7758 7715 7792 7749
rect 7826 7715 7860 7749
rect 7894 7715 7928 7749
rect 7962 7715 7996 7749
rect 8030 7715 8064 7749
rect 8098 7715 8132 7749
rect 8166 7715 8200 7749
rect 8234 7715 8268 7749
rect 8302 7715 8336 7749
rect 8370 7715 8404 7749
rect 8438 7715 8472 7749
rect 8506 7715 8540 7749
rect 8574 7715 8608 7749
rect 8642 7715 8676 7749
rect 8710 7715 8744 7749
rect 8778 7715 8812 7749
rect 8846 7715 8880 7749
rect 8914 7715 8948 7749
rect 8982 7715 9016 7749
rect 9050 7715 9084 7749
rect 9118 7715 9152 7749
rect 9186 7715 9220 7749
rect 9254 7715 9288 7749
rect 9322 7715 9356 7749
rect 9390 7715 9424 7749
rect 9458 7715 9492 7749
rect 9526 7715 9560 7749
rect 9594 7715 9628 7749
rect 9662 7715 9696 7749
rect 9730 7715 9764 7749
rect 9798 7715 9832 7749
rect 9866 7715 9900 7749
rect 9934 7715 9968 7749
rect 10002 7715 10036 7749
rect 10070 7715 10104 7749
rect 10138 7715 10172 7749
rect 10206 7715 10240 7749
rect 10274 7715 10308 7749
rect 10342 7715 10376 7749
rect 10410 7715 10444 7749
rect 10478 7715 10512 7749
rect 10546 7715 10580 7749
rect 10614 7715 10648 7749
rect 10682 7715 10716 7749
rect 10750 7715 10784 7749
rect 10818 7715 10852 7749
rect 10886 7715 10920 7749
rect 10954 7715 10988 7749
rect 11022 7715 11056 7749
rect 11090 7715 11124 7749
rect 11158 7715 11192 7749
rect 11226 7715 11260 7749
rect 11294 7715 11328 7749
rect 11362 7715 11396 7749
rect 11430 7715 11464 7749
rect 11498 7715 11532 7749
rect 11566 7715 11600 7749
rect 11634 7715 11668 7749
rect 11702 7715 11736 7749
rect 11770 7715 11804 7749
rect 11838 7715 11872 7749
rect 11906 7715 11940 7749
rect 11974 7715 12008 7749
rect 12042 7715 12076 7749
rect 12110 7715 12144 7749
rect 12178 7715 12212 7749
rect 12246 7715 12280 7749
rect 12314 7715 12348 7749
rect 12382 7715 12416 7749
rect 12450 7715 12484 7749
rect 12518 7715 12552 7749
rect 12586 7715 12620 7749
rect 12654 7715 12688 7749
rect 12722 7715 12756 7749
rect 12790 7715 12824 7749
rect 12858 7715 12892 7749
rect 12926 7715 12960 7749
rect 12994 7715 13028 7749
rect 13062 7715 13096 7749
rect 13130 7715 13164 7749
rect 13198 7715 13232 7749
rect 13266 7715 13300 7749
rect 13334 7715 13368 7749
rect 13402 7715 13436 7749
rect 13470 7715 13504 7749
rect 13538 7715 13572 7749
rect 13606 7715 13640 7749
rect 13674 7715 13708 7749
rect 13742 7715 13776 7749
rect 13810 7715 13844 7749
rect 13878 7715 13912 7749
rect 13946 7715 13980 7749
rect 14014 7715 14048 7749
rect 14082 7715 14116 7749
rect 14150 7715 14184 7749
rect 14218 7715 14252 7749
rect 14286 7715 14320 7749
rect 14354 7715 14388 7749
rect 14422 7715 14456 7749
rect 14490 7715 14524 7749
rect 14558 7715 14592 7749
rect 14626 7715 14660 7749
rect 14694 7715 14728 7749
rect 14762 7715 14796 7749
rect 14830 7715 14864 7749
rect 14898 7715 15102 7749
rect 34 7713 15102 7715
rect 34 7679 14932 7713
rect 14966 7679 15000 7713
rect 15034 7679 15068 7713
rect 34 7676 15102 7679
rect 34 7642 2733 7676
rect 34 7608 68 7642
rect 102 7608 137 7642
rect 171 7608 206 7642
rect 240 7608 275 7642
rect 309 7608 344 7642
rect 378 7608 413 7642
rect 447 7608 482 7642
rect 516 7608 551 7642
rect 585 7608 620 7642
rect 654 7608 689 7642
rect 723 7608 758 7642
rect 792 7608 827 7642
rect 861 7608 896 7642
rect 930 7608 965 7642
rect 999 7608 1033 7642
rect 1067 7608 1101 7642
rect 1135 7608 1169 7642
rect 1203 7608 1237 7642
rect 1271 7608 1305 7642
rect 1339 7608 1373 7642
rect 1407 7608 1441 7642
rect 1475 7608 1509 7642
rect 1543 7608 1577 7642
rect 1611 7608 1645 7642
rect 1679 7608 1713 7642
rect 1747 7608 1781 7642
rect 1815 7608 1849 7642
rect 1883 7608 1917 7642
rect 1951 7608 1985 7642
rect 2019 7608 2053 7642
rect 2087 7608 2121 7642
rect 2155 7608 2189 7642
rect 2223 7608 2257 7642
rect 2291 7608 2325 7642
rect 2359 7608 2393 7642
rect 2427 7608 2461 7642
rect 2495 7608 2529 7642
rect 2563 7608 2597 7642
rect 2631 7608 2665 7642
rect 2699 7608 2733 7642
rect 34 7570 2733 7608
rect 34 7536 68 7570
rect 102 7536 137 7570
rect 171 7536 206 7570
rect 240 7536 275 7570
rect 309 7536 344 7570
rect 378 7536 413 7570
rect 447 7536 482 7570
rect 516 7536 551 7570
rect 585 7536 620 7570
rect 654 7536 689 7570
rect 723 7536 758 7570
rect 792 7536 827 7570
rect 861 7536 896 7570
rect 930 7536 965 7570
rect 999 7536 1033 7570
rect 1067 7536 1101 7570
rect 1135 7536 1169 7570
rect 1203 7536 1237 7570
rect 1271 7536 1305 7570
rect 1339 7536 1373 7570
rect 1407 7536 1441 7570
rect 1475 7536 1509 7570
rect 1543 7536 1577 7570
rect 1611 7536 1645 7570
rect 1679 7536 1713 7570
rect 1747 7536 1781 7570
rect 1815 7536 1849 7570
rect 1883 7536 1917 7570
rect 1951 7536 1985 7570
rect 2019 7536 2053 7570
rect 2087 7536 2121 7570
rect 2155 7536 2189 7570
rect 2223 7536 2257 7570
rect 2291 7536 2325 7570
rect 2359 7536 2393 7570
rect 2427 7536 2461 7570
rect 2495 7536 2529 7570
rect 2563 7536 2597 7570
rect 2631 7536 2665 7570
rect 2699 7536 2733 7570
rect 34 7498 2733 7536
rect 34 7464 68 7498
rect 102 7464 137 7498
rect 171 7464 206 7498
rect 240 7464 275 7498
rect 309 7464 344 7498
rect 378 7464 413 7498
rect 447 7464 482 7498
rect 516 7464 551 7498
rect 585 7464 620 7498
rect 654 7464 689 7498
rect 723 7464 758 7498
rect 792 7464 827 7498
rect 861 7464 896 7498
rect 930 7464 965 7498
rect 999 7464 1033 7498
rect 1067 7464 1101 7498
rect 1135 7464 1169 7498
rect 1203 7464 1237 7498
rect 1271 7464 1305 7498
rect 1339 7464 1373 7498
rect 1407 7464 1441 7498
rect 1475 7464 1509 7498
rect 1543 7464 1577 7498
rect 1611 7464 1645 7498
rect 1679 7464 1713 7498
rect 1747 7464 1781 7498
rect 1815 7464 1849 7498
rect 1883 7464 1917 7498
rect 1951 7464 1985 7498
rect 2019 7464 2053 7498
rect 2087 7464 2121 7498
rect 2155 7464 2189 7498
rect 2223 7464 2257 7498
rect 2291 7464 2325 7498
rect 2359 7464 2393 7498
rect 2427 7464 2461 7498
rect 2495 7464 2529 7498
rect 2563 7464 2597 7498
rect 2631 7464 2665 7498
rect 2699 7464 2733 7498
rect 34 7426 2733 7464
rect 34 7392 68 7426
rect 102 7392 137 7426
rect 171 7392 206 7426
rect 240 7392 275 7426
rect 309 7392 344 7426
rect 378 7392 413 7426
rect 447 7392 482 7426
rect 516 7392 551 7426
rect 585 7392 620 7426
rect 654 7392 689 7426
rect 723 7392 758 7426
rect 792 7392 827 7426
rect 861 7392 896 7426
rect 930 7392 965 7426
rect 999 7392 1033 7426
rect 1067 7392 1101 7426
rect 1135 7392 1169 7426
rect 1203 7392 1237 7426
rect 1271 7392 1305 7426
rect 1339 7392 1373 7426
rect 1407 7392 1441 7426
rect 1475 7392 1509 7426
rect 1543 7392 1577 7426
rect 1611 7392 1645 7426
rect 1679 7392 1713 7426
rect 1747 7392 1781 7426
rect 1815 7392 1849 7426
rect 1883 7392 1917 7426
rect 1951 7392 1985 7426
rect 2019 7392 2053 7426
rect 2087 7392 2121 7426
rect 2155 7392 2189 7426
rect 2223 7392 2257 7426
rect 2291 7392 2325 7426
rect 2359 7392 2393 7426
rect 2427 7392 2461 7426
rect 2495 7392 2529 7426
rect 2563 7392 2597 7426
rect 2631 7392 2665 7426
rect 2699 7392 2733 7426
rect 34 7354 2733 7392
rect 34 7320 68 7354
rect 102 7320 137 7354
rect 171 7320 206 7354
rect 240 7320 275 7354
rect 309 7320 344 7354
rect 378 7320 413 7354
rect 447 7320 482 7354
rect 516 7320 551 7354
rect 585 7320 620 7354
rect 654 7320 689 7354
rect 723 7320 758 7354
rect 792 7320 827 7354
rect 861 7320 896 7354
rect 930 7320 965 7354
rect 999 7320 1033 7354
rect 1067 7320 1101 7354
rect 1135 7320 1169 7354
rect 1203 7320 1237 7354
rect 1271 7320 1305 7354
rect 1339 7320 1373 7354
rect 1407 7320 1441 7354
rect 1475 7320 1509 7354
rect 1543 7320 1577 7354
rect 1611 7320 1645 7354
rect 1679 7320 1713 7354
rect 1747 7320 1781 7354
rect 1815 7320 1849 7354
rect 1883 7320 1917 7354
rect 1951 7320 1985 7354
rect 2019 7320 2053 7354
rect 2087 7320 2121 7354
rect 2155 7320 2189 7354
rect 2223 7320 2257 7354
rect 2291 7320 2325 7354
rect 2359 7320 2393 7354
rect 2427 7320 2461 7354
rect 2495 7320 2529 7354
rect 2563 7320 2597 7354
rect 2631 7320 2665 7354
rect 2699 7320 2733 7354
rect 34 7282 2733 7320
rect 12490 7641 15102 7676
rect 12490 7640 14932 7641
rect 12490 7606 12524 7640
rect 12558 7606 12593 7640
rect 12627 7606 12662 7640
rect 12696 7606 12731 7640
rect 12765 7606 12800 7640
rect 12834 7606 12869 7640
rect 12903 7606 12938 7640
rect 12972 7606 13007 7640
rect 13041 7606 13076 7640
rect 13110 7606 13145 7640
rect 13179 7606 13214 7640
rect 13248 7606 13283 7640
rect 13317 7606 13352 7640
rect 13386 7606 13421 7640
rect 13455 7606 13490 7640
rect 13524 7606 13559 7640
rect 13593 7606 13628 7640
rect 13662 7606 13697 7640
rect 13731 7606 13766 7640
rect 13800 7606 13835 7640
rect 13869 7606 13904 7640
rect 13938 7606 13973 7640
rect 14007 7606 14042 7640
rect 14076 7606 14111 7640
rect 14145 7606 14180 7640
rect 14214 7606 14249 7640
rect 14283 7606 14318 7640
rect 14352 7606 14387 7640
rect 14421 7606 14456 7640
rect 14490 7606 14524 7640
rect 14558 7606 14592 7640
rect 14626 7606 14660 7640
rect 14694 7606 14728 7640
rect 14762 7606 14796 7640
rect 14830 7606 14864 7640
rect 14898 7607 14932 7640
rect 14966 7607 15000 7641
rect 15034 7607 15068 7641
rect 14898 7606 15102 7607
rect 12490 7569 15102 7606
rect 12490 7556 14932 7569
rect 12490 7522 12524 7556
rect 12558 7522 12593 7556
rect 12627 7522 12662 7556
rect 12696 7522 12731 7556
rect 12765 7522 12800 7556
rect 12834 7522 12869 7556
rect 12903 7522 12938 7556
rect 12972 7522 13007 7556
rect 13041 7522 13076 7556
rect 13110 7522 13145 7556
rect 13179 7522 13214 7556
rect 13248 7522 13283 7556
rect 13317 7522 13352 7556
rect 13386 7522 13421 7556
rect 13455 7522 13490 7556
rect 13524 7522 13559 7556
rect 13593 7522 13628 7556
rect 13662 7522 13697 7556
rect 13731 7522 13766 7556
rect 13800 7522 13835 7556
rect 13869 7522 13904 7556
rect 13938 7522 13973 7556
rect 14007 7522 14042 7556
rect 14076 7522 14111 7556
rect 14145 7522 14180 7556
rect 14214 7522 14249 7556
rect 14283 7522 14318 7556
rect 14352 7522 14387 7556
rect 14421 7522 14456 7556
rect 14490 7522 14524 7556
rect 14558 7522 14592 7556
rect 14626 7522 14660 7556
rect 14694 7522 14728 7556
rect 14762 7522 14796 7556
rect 14830 7522 14864 7556
rect 14898 7535 14932 7556
rect 14966 7535 15000 7569
rect 15034 7535 15068 7569
rect 14898 7522 15102 7535
rect 12490 7497 15102 7522
rect 12490 7472 14932 7497
rect 12490 7438 12524 7472
rect 12558 7438 12593 7472
rect 12627 7438 12662 7472
rect 12696 7438 12731 7472
rect 12765 7438 12800 7472
rect 12834 7438 12869 7472
rect 12903 7438 12938 7472
rect 12972 7438 13007 7472
rect 13041 7438 13076 7472
rect 13110 7438 13145 7472
rect 13179 7438 13214 7472
rect 13248 7438 13283 7472
rect 13317 7438 13352 7472
rect 13386 7438 13421 7472
rect 13455 7438 13490 7472
rect 13524 7438 13559 7472
rect 13593 7438 13628 7472
rect 13662 7438 13697 7472
rect 13731 7438 13766 7472
rect 13800 7438 13835 7472
rect 13869 7438 13904 7472
rect 13938 7438 13973 7472
rect 14007 7438 14042 7472
rect 14076 7438 14111 7472
rect 14145 7438 14180 7472
rect 14214 7438 14249 7472
rect 14283 7438 14318 7472
rect 14352 7438 14387 7472
rect 14421 7438 14456 7472
rect 14490 7438 14524 7472
rect 14558 7438 14592 7472
rect 14626 7438 14660 7472
rect 14694 7438 14728 7472
rect 14762 7438 14796 7472
rect 14830 7438 14864 7472
rect 14898 7463 14932 7472
rect 14966 7463 15000 7497
rect 15034 7463 15068 7497
rect 14898 7438 15102 7463
rect 12490 7425 15102 7438
rect 12490 7391 14932 7425
rect 14966 7391 15000 7425
rect 15034 7391 15068 7425
rect 12490 7388 15102 7391
rect 12490 7354 12524 7388
rect 12558 7354 12593 7388
rect 12627 7354 12662 7388
rect 12696 7354 12731 7388
rect 12765 7354 12800 7388
rect 12834 7354 12869 7388
rect 12903 7354 12938 7388
rect 12972 7354 13007 7388
rect 13041 7354 13076 7388
rect 13110 7354 13145 7388
rect 13179 7354 13214 7388
rect 13248 7354 13283 7388
rect 13317 7354 13352 7388
rect 13386 7354 13421 7388
rect 13455 7354 13490 7388
rect 13524 7354 13559 7388
rect 13593 7354 13628 7388
rect 13662 7354 13697 7388
rect 13731 7354 13766 7388
rect 13800 7354 13835 7388
rect 13869 7354 13904 7388
rect 13938 7354 13973 7388
rect 14007 7354 14042 7388
rect 14076 7354 14111 7388
rect 14145 7354 14180 7388
rect 14214 7354 14249 7388
rect 14283 7354 14318 7388
rect 14352 7354 14387 7388
rect 14421 7354 14456 7388
rect 14490 7354 14524 7388
rect 14558 7354 14592 7388
rect 14626 7354 14660 7388
rect 14694 7354 14728 7388
rect 14762 7354 14796 7388
rect 14830 7354 14864 7388
rect 14898 7354 15102 7388
rect 12490 7353 15102 7354
rect 12490 7319 14932 7353
rect 14966 7319 15000 7353
rect 15034 7319 15068 7353
rect 12490 7317 15102 7319
rect 34 7248 68 7282
rect 102 7248 137 7282
rect 171 7248 206 7282
rect 240 7248 275 7282
rect 309 7248 344 7282
rect 378 7248 413 7282
rect 447 7248 482 7282
rect 516 7248 551 7282
rect 585 7248 620 7282
rect 654 7248 689 7282
rect 723 7248 758 7282
rect 792 7248 827 7282
rect 861 7248 896 7282
rect 930 7248 965 7282
rect 999 7248 1033 7282
rect 1067 7248 1101 7282
rect 1135 7248 1169 7282
rect 1203 7248 1237 7282
rect 1271 7248 1305 7282
rect 1339 7248 1373 7282
rect 1407 7248 1441 7282
rect 1475 7248 1509 7282
rect 1543 7248 1577 7282
rect 1611 7248 1645 7282
rect 1679 7248 1713 7282
rect 1747 7248 1781 7282
rect 1815 7248 1849 7282
rect 1883 7248 1917 7282
rect 1951 7248 1985 7282
rect 2019 7248 2053 7282
rect 2087 7248 2121 7282
rect 2155 7248 2189 7282
rect 2223 7248 2257 7282
rect 2291 7248 2325 7282
rect 2359 7248 2393 7282
rect 2427 7248 2461 7282
rect 2495 7248 2529 7282
rect 2563 7248 2597 7282
rect 2631 7248 2665 7282
rect 2699 7248 2733 7282
rect 34 7210 2733 7248
rect 34 7176 68 7210
rect 102 7176 137 7210
rect 171 7176 206 7210
rect 240 7176 275 7210
rect 309 7176 344 7210
rect 378 7176 413 7210
rect 447 7176 482 7210
rect 516 7176 551 7210
rect 585 7176 620 7210
rect 654 7176 689 7210
rect 723 7176 758 7210
rect 792 7176 827 7210
rect 861 7176 896 7210
rect 930 7176 965 7210
rect 999 7176 1033 7210
rect 1067 7176 1101 7210
rect 1135 7176 1169 7210
rect 1203 7176 1237 7210
rect 1271 7176 1305 7210
rect 1339 7176 1373 7210
rect 1407 7176 1441 7210
rect 1475 7176 1509 7210
rect 1543 7176 1577 7210
rect 1611 7176 1645 7210
rect 1679 7176 1713 7210
rect 1747 7176 1781 7210
rect 1815 7176 1849 7210
rect 1883 7176 1917 7210
rect 1951 7176 1985 7210
rect 2019 7176 2053 7210
rect 2087 7176 2121 7210
rect 2155 7176 2189 7210
rect 2223 7176 2257 7210
rect 2291 7176 2325 7210
rect 2359 7176 2393 7210
rect 2427 7176 2461 7210
rect 2495 7176 2529 7210
rect 2563 7176 2597 7210
rect 2631 7176 2665 7210
rect 2699 7176 2733 7210
rect 34 7138 2733 7176
rect 34 7104 68 7138
rect 102 7104 137 7138
rect 171 7104 206 7138
rect 240 7104 275 7138
rect 309 7104 344 7138
rect 378 7104 413 7138
rect 447 7104 482 7138
rect 516 7104 551 7138
rect 585 7104 620 7138
rect 654 7104 689 7138
rect 723 7104 758 7138
rect 792 7104 827 7138
rect 861 7104 896 7138
rect 930 7104 965 7138
rect 999 7104 1033 7138
rect 1067 7104 1101 7138
rect 1135 7104 1169 7138
rect 1203 7104 1237 7138
rect 1271 7104 1305 7138
rect 1339 7104 1373 7138
rect 1407 7104 1441 7138
rect 1475 7104 1509 7138
rect 1543 7104 1577 7138
rect 1611 7104 1645 7138
rect 1679 7104 1713 7138
rect 1747 7104 1781 7138
rect 1815 7104 1849 7138
rect 1883 7104 1917 7138
rect 1951 7104 1985 7138
rect 2019 7104 2053 7138
rect 2087 7104 2121 7138
rect 2155 7104 2189 7138
rect 2223 7104 2257 7138
rect 2291 7104 2325 7138
rect 2359 7104 2393 7138
rect 2427 7104 2461 7138
rect 2495 7104 2529 7138
rect 2563 7104 2597 7138
rect 2631 7104 2665 7138
rect 2699 7104 2733 7138
rect 34 7066 2733 7104
rect 34 7032 68 7066
rect 102 7032 137 7066
rect 171 7032 206 7066
rect 240 7032 275 7066
rect 309 7032 344 7066
rect 378 7032 413 7066
rect 447 7032 482 7066
rect 516 7032 551 7066
rect 585 7032 620 7066
rect 654 7032 689 7066
rect 723 7032 758 7066
rect 792 7032 827 7066
rect 861 7032 896 7066
rect 930 7032 965 7066
rect 999 7032 1033 7066
rect 1067 7032 1101 7066
rect 1135 7032 1169 7066
rect 1203 7032 1237 7066
rect 1271 7032 1305 7066
rect 1339 7032 1373 7066
rect 1407 7032 1441 7066
rect 1475 7032 1509 7066
rect 1543 7032 1577 7066
rect 1611 7032 1645 7066
rect 1679 7032 1713 7066
rect 1747 7032 1781 7066
rect 1815 7032 1849 7066
rect 1883 7032 1917 7066
rect 1951 7032 1985 7066
rect 2019 7032 2053 7066
rect 2087 7032 2121 7066
rect 2155 7032 2189 7066
rect 2223 7032 2257 7066
rect 2291 7032 2325 7066
rect 2359 7032 2393 7066
rect 2427 7032 2461 7066
rect 2495 7032 2529 7066
rect 2563 7032 2597 7066
rect 2631 7032 2665 7066
rect 2699 7063 2733 7066
rect 8176 7282 15102 7317
rect 8176 7248 8210 7282
rect 8244 7248 8279 7282
rect 8313 7248 8348 7282
rect 8382 7248 8417 7282
rect 8451 7248 8486 7282
rect 8520 7248 8555 7282
rect 8589 7248 8624 7282
rect 8658 7248 8693 7282
rect 8727 7248 8762 7282
rect 8796 7248 8831 7282
rect 8865 7248 8900 7282
rect 8934 7248 8969 7282
rect 9003 7248 9038 7282
rect 9072 7248 9107 7282
rect 9141 7248 9176 7282
rect 9210 7248 9245 7282
rect 9279 7248 9314 7282
rect 9348 7248 9383 7282
rect 9417 7248 9452 7282
rect 9486 7248 9521 7282
rect 9555 7248 9590 7282
rect 9624 7248 9659 7282
rect 9693 7248 9728 7282
rect 9762 7248 9797 7282
rect 9831 7248 9866 7282
rect 9900 7248 9935 7282
rect 9969 7248 10004 7282
rect 10038 7248 10073 7282
rect 10107 7248 10142 7282
rect 10176 7248 10211 7282
rect 10245 7248 10280 7282
rect 10314 7248 10349 7282
rect 10383 7248 10418 7282
rect 10452 7248 10487 7282
rect 10521 7248 10556 7282
rect 10590 7248 10625 7282
rect 10659 7248 10694 7282
rect 10728 7248 10763 7282
rect 10797 7248 10832 7282
rect 10866 7248 10901 7282
rect 10935 7248 10970 7282
rect 11004 7248 11039 7282
rect 11073 7248 11108 7282
rect 11142 7248 11177 7282
rect 11211 7248 11246 7282
rect 11280 7248 11315 7282
rect 11349 7248 11384 7282
rect 11418 7248 11453 7282
rect 11487 7248 11522 7282
rect 11556 7248 11591 7282
rect 11625 7248 11660 7282
rect 11694 7248 11729 7282
rect 11763 7248 11798 7282
rect 11832 7248 11867 7282
rect 11901 7248 11936 7282
rect 11970 7248 12005 7282
rect 12039 7248 12074 7282
rect 12108 7248 12143 7282
rect 12177 7248 12212 7282
rect 12246 7248 12280 7282
rect 12314 7248 12348 7282
rect 12382 7248 12416 7282
rect 12450 7248 12484 7282
rect 12518 7248 12552 7282
rect 12586 7248 12620 7282
rect 12654 7248 12688 7282
rect 12722 7248 12756 7282
rect 12790 7248 12824 7282
rect 12858 7248 12892 7282
rect 12926 7248 12960 7282
rect 12994 7248 13028 7282
rect 13062 7248 13096 7282
rect 13130 7248 13164 7282
rect 13198 7248 13232 7282
rect 13266 7248 13300 7282
rect 13334 7248 13368 7282
rect 13402 7248 13436 7282
rect 13470 7248 13504 7282
rect 13538 7248 13572 7282
rect 13606 7248 13640 7282
rect 13674 7248 13708 7282
rect 13742 7248 13776 7282
rect 13810 7248 13844 7282
rect 13878 7248 13912 7282
rect 13946 7248 13980 7282
rect 14014 7248 14048 7282
rect 14082 7248 14116 7282
rect 14150 7248 14184 7282
rect 14218 7248 14252 7282
rect 14286 7248 14320 7282
rect 14354 7248 14388 7282
rect 14422 7248 14456 7282
rect 14490 7248 14524 7282
rect 14558 7248 14592 7282
rect 14626 7248 14660 7282
rect 14694 7248 14728 7282
rect 14762 7248 14796 7282
rect 14830 7248 14864 7282
rect 14898 7281 15102 7282
rect 14898 7248 14932 7281
rect 8176 7247 14932 7248
rect 14966 7247 15000 7281
rect 15034 7247 15068 7281
rect 8176 7210 15102 7247
rect 8176 7176 8210 7210
rect 8244 7176 8279 7210
rect 8313 7176 8348 7210
rect 8382 7176 8417 7210
rect 8451 7176 8486 7210
rect 8520 7176 8555 7210
rect 8589 7176 8624 7210
rect 8658 7176 8693 7210
rect 8727 7176 8762 7210
rect 8796 7176 8831 7210
rect 8865 7176 8900 7210
rect 8934 7176 8969 7210
rect 9003 7176 9038 7210
rect 9072 7176 9107 7210
rect 9141 7176 9176 7210
rect 9210 7176 9245 7210
rect 9279 7176 9314 7210
rect 9348 7176 9383 7210
rect 9417 7176 9452 7210
rect 9486 7176 9521 7210
rect 9555 7176 9590 7210
rect 9624 7176 9659 7210
rect 9693 7176 9728 7210
rect 9762 7176 9797 7210
rect 9831 7176 9866 7210
rect 9900 7176 9935 7210
rect 9969 7176 10004 7210
rect 10038 7176 10073 7210
rect 10107 7176 10142 7210
rect 10176 7176 10211 7210
rect 10245 7176 10280 7210
rect 10314 7176 10349 7210
rect 10383 7176 10418 7210
rect 10452 7176 10487 7210
rect 10521 7176 10556 7210
rect 10590 7176 10625 7210
rect 10659 7176 10694 7210
rect 10728 7176 10763 7210
rect 10797 7176 10832 7210
rect 10866 7176 10901 7210
rect 10935 7176 10970 7210
rect 11004 7176 11039 7210
rect 11073 7176 11108 7210
rect 11142 7176 11177 7210
rect 11211 7176 11246 7210
rect 11280 7176 11315 7210
rect 11349 7176 11384 7210
rect 11418 7176 11453 7210
rect 11487 7176 11522 7210
rect 11556 7176 11591 7210
rect 11625 7176 11660 7210
rect 11694 7176 11729 7210
rect 11763 7176 11798 7210
rect 11832 7176 11867 7210
rect 11901 7176 11936 7210
rect 11970 7176 12005 7210
rect 12039 7176 12074 7210
rect 12108 7176 12143 7210
rect 12177 7176 12212 7210
rect 12246 7176 12280 7210
rect 12314 7176 12348 7210
rect 12382 7176 12416 7210
rect 12450 7176 12484 7210
rect 12518 7176 12552 7210
rect 12586 7176 12620 7210
rect 12654 7176 12688 7210
rect 12722 7176 12756 7210
rect 12790 7176 12824 7210
rect 12858 7176 12892 7210
rect 12926 7176 12960 7210
rect 12994 7176 13028 7210
rect 13062 7176 13096 7210
rect 13130 7176 13164 7210
rect 13198 7176 13232 7210
rect 13266 7176 13300 7210
rect 13334 7176 13368 7210
rect 13402 7176 13436 7210
rect 13470 7176 13504 7210
rect 13538 7176 13572 7210
rect 13606 7176 13640 7210
rect 13674 7176 13708 7210
rect 13742 7176 13776 7210
rect 13810 7176 13844 7210
rect 13878 7176 13912 7210
rect 13946 7176 13980 7210
rect 14014 7176 14048 7210
rect 14082 7176 14116 7210
rect 14150 7176 14184 7210
rect 14218 7176 14252 7210
rect 14286 7176 14320 7210
rect 14354 7176 14388 7210
rect 14422 7176 14456 7210
rect 14490 7176 14524 7210
rect 14558 7176 14592 7210
rect 14626 7176 14660 7210
rect 14694 7176 14728 7210
rect 14762 7176 14796 7210
rect 14830 7176 14864 7210
rect 14898 7209 15102 7210
rect 14898 7176 14932 7209
rect 8176 7175 14932 7176
rect 14966 7175 15000 7209
rect 15034 7175 15068 7209
rect 8176 7138 15102 7175
rect 8176 7104 8210 7138
rect 8244 7104 8279 7138
rect 8313 7104 8348 7138
rect 8382 7104 8417 7138
rect 8451 7104 8486 7138
rect 8520 7104 8555 7138
rect 8589 7104 8624 7138
rect 8658 7104 8693 7138
rect 8727 7104 8762 7138
rect 8796 7104 8831 7138
rect 8865 7104 8900 7138
rect 8934 7104 8969 7138
rect 9003 7104 9038 7138
rect 9072 7104 9107 7138
rect 9141 7104 9176 7138
rect 9210 7104 9245 7138
rect 9279 7104 9314 7138
rect 9348 7104 9383 7138
rect 9417 7104 9452 7138
rect 9486 7104 9521 7138
rect 9555 7104 9590 7138
rect 9624 7104 9659 7138
rect 9693 7104 9728 7138
rect 9762 7104 9797 7138
rect 9831 7104 9866 7138
rect 9900 7104 9935 7138
rect 9969 7104 10004 7138
rect 10038 7104 10073 7138
rect 10107 7104 10142 7138
rect 10176 7104 10211 7138
rect 10245 7104 10280 7138
rect 10314 7104 10349 7138
rect 10383 7104 10418 7138
rect 10452 7104 10487 7138
rect 10521 7104 10556 7138
rect 10590 7104 10625 7138
rect 10659 7104 10694 7138
rect 10728 7104 10763 7138
rect 10797 7104 10832 7138
rect 10866 7104 10901 7138
rect 10935 7104 10970 7138
rect 11004 7104 11039 7138
rect 11073 7104 11108 7138
rect 11142 7104 11177 7138
rect 11211 7104 11246 7138
rect 11280 7104 11315 7138
rect 11349 7104 11384 7138
rect 11418 7104 11453 7138
rect 11487 7104 11522 7138
rect 11556 7104 11591 7138
rect 11625 7104 11660 7138
rect 11694 7104 11729 7138
rect 11763 7104 11798 7138
rect 11832 7104 11867 7138
rect 11901 7104 11936 7138
rect 11970 7104 12005 7138
rect 12039 7104 12074 7138
rect 12108 7104 12143 7138
rect 12177 7104 12212 7138
rect 12246 7104 12280 7138
rect 12314 7104 12348 7138
rect 12382 7104 12416 7138
rect 12450 7104 12484 7138
rect 12518 7104 12552 7138
rect 12586 7104 12620 7138
rect 12654 7104 12688 7138
rect 12722 7104 12756 7138
rect 12790 7104 12824 7138
rect 12858 7104 12892 7138
rect 12926 7104 12960 7138
rect 12994 7104 13028 7138
rect 13062 7104 13096 7138
rect 13130 7104 13164 7138
rect 13198 7104 13232 7138
rect 13266 7104 13300 7138
rect 13334 7104 13368 7138
rect 13402 7104 13436 7138
rect 13470 7104 13504 7138
rect 13538 7104 13572 7138
rect 13606 7104 13640 7138
rect 13674 7104 13708 7138
rect 13742 7104 13776 7138
rect 13810 7104 13844 7138
rect 13878 7104 13912 7138
rect 13946 7104 13980 7138
rect 14014 7104 14048 7138
rect 14082 7104 14116 7138
rect 14150 7104 14184 7138
rect 14218 7104 14252 7138
rect 14286 7104 14320 7138
rect 14354 7104 14388 7138
rect 14422 7104 14456 7138
rect 14490 7104 14524 7138
rect 14558 7104 14592 7138
rect 14626 7104 14660 7138
rect 14694 7104 14728 7138
rect 14762 7104 14796 7138
rect 14830 7104 14864 7138
rect 14898 7137 15102 7138
rect 14898 7104 14932 7137
rect 8176 7103 14932 7104
rect 14966 7103 15000 7137
rect 15034 7103 15068 7137
rect 8176 7066 15102 7103
rect 2699 7047 7756 7063
rect 2699 7032 2757 7047
rect 34 7013 2757 7032
rect 2791 7013 2825 7047
rect 2859 7013 2893 7047
rect 2927 7013 2961 7047
rect 2995 7013 3029 7047
rect 3063 7013 3097 7047
rect 3131 7013 3165 7047
rect 3199 7013 3233 7047
rect 3267 7013 3301 7047
rect 3335 7013 3369 7047
rect 3403 7013 3437 7047
rect 3471 7013 3505 7047
rect 3539 7013 3573 7047
rect 3607 7013 3641 7047
rect 3675 7013 3709 7047
rect 3743 7013 3777 7047
rect 3811 7013 3845 7047
rect 3879 7013 3913 7047
rect 3947 7013 3981 7047
rect 4015 7013 4049 7047
rect 4083 7013 4117 7047
rect 4151 7013 4185 7047
rect 4219 7013 4253 7047
rect 4287 7013 4321 7047
rect 4355 7013 4389 7047
rect 4423 7013 4457 7047
rect 4491 7013 4525 7047
rect 4559 7013 4593 7047
rect 4627 7013 4661 7047
rect 4695 7013 4729 7047
rect 4763 7013 4797 7047
rect 4831 7013 4865 7047
rect 4899 7013 4933 7047
rect 4967 7013 5001 7047
rect 5035 7013 5069 7047
rect 5103 7013 5137 7047
rect 5171 7013 5205 7047
rect 5239 7013 5273 7047
rect 5307 7013 5341 7047
rect 5375 7013 5409 7047
rect 5443 7013 5477 7047
rect 5511 7013 5545 7047
rect 5579 7013 5613 7047
rect 5647 7013 5681 7047
rect 5715 7013 5749 7047
rect 5783 7013 5817 7047
rect 5851 7013 5885 7047
rect 5919 7013 5953 7047
rect 5987 7013 6021 7047
rect 6055 7013 6089 7047
rect 6123 7013 6157 7047
rect 6191 7013 6225 7047
rect 6259 7013 6293 7047
rect 6327 7013 6361 7047
rect 6395 7013 6429 7047
rect 6463 7013 6497 7047
rect 6531 7013 6565 7047
rect 6599 7013 6633 7047
rect 6667 7013 6701 7047
rect 6735 7013 6769 7047
rect 6803 7013 6837 7047
rect 6871 7013 6905 7047
rect 6939 7013 6973 7047
rect 7007 7013 7041 7047
rect 7075 7013 7109 7047
rect 7143 7013 7177 7047
rect 7211 7013 7245 7047
rect 7279 7013 7313 7047
rect 7347 7013 7381 7047
rect 7415 7013 7449 7047
rect 7483 7013 7517 7047
rect 7551 7013 7585 7047
rect 7619 7013 7653 7047
rect 7687 7013 7756 7047
rect 34 6997 7756 7013
rect 8176 7032 8210 7066
rect 8244 7032 8279 7066
rect 8313 7032 8348 7066
rect 8382 7032 8417 7066
rect 8451 7032 8486 7066
rect 8520 7032 8555 7066
rect 8589 7032 8624 7066
rect 8658 7032 8693 7066
rect 8727 7032 8762 7066
rect 8796 7032 8831 7066
rect 8865 7032 8900 7066
rect 8934 7032 8969 7066
rect 9003 7032 9038 7066
rect 9072 7032 9107 7066
rect 9141 7032 9176 7066
rect 9210 7032 9245 7066
rect 9279 7032 9314 7066
rect 9348 7032 9383 7066
rect 9417 7032 9452 7066
rect 9486 7032 9521 7066
rect 9555 7032 9590 7066
rect 9624 7032 9659 7066
rect 9693 7032 9728 7066
rect 9762 7032 9797 7066
rect 9831 7032 9866 7066
rect 9900 7032 9935 7066
rect 9969 7032 10004 7066
rect 10038 7032 10073 7066
rect 10107 7032 10142 7066
rect 10176 7032 10211 7066
rect 10245 7032 10280 7066
rect 10314 7032 10349 7066
rect 10383 7032 10418 7066
rect 10452 7032 10487 7066
rect 10521 7032 10556 7066
rect 10590 7032 10625 7066
rect 10659 7032 10694 7066
rect 10728 7032 10763 7066
rect 10797 7032 10832 7066
rect 10866 7032 10901 7066
rect 10935 7032 10970 7066
rect 11004 7032 11039 7066
rect 11073 7032 11108 7066
rect 11142 7032 11177 7066
rect 11211 7032 11246 7066
rect 11280 7032 11315 7066
rect 11349 7032 11384 7066
rect 11418 7032 11453 7066
rect 11487 7032 11522 7066
rect 11556 7032 11591 7066
rect 11625 7032 11660 7066
rect 11694 7032 11729 7066
rect 11763 7032 11798 7066
rect 11832 7032 11867 7066
rect 11901 7032 11936 7066
rect 11970 7032 12005 7066
rect 12039 7032 12074 7066
rect 12108 7032 12143 7066
rect 12177 7032 12212 7066
rect 12246 7032 12280 7066
rect 12314 7032 12348 7066
rect 12382 7032 12416 7066
rect 12450 7032 12484 7066
rect 12518 7032 12552 7066
rect 12586 7032 12620 7066
rect 12654 7032 12688 7066
rect 12722 7032 12756 7066
rect 12790 7032 12824 7066
rect 12858 7032 12892 7066
rect 12926 7032 12960 7066
rect 12994 7032 13028 7066
rect 13062 7032 13096 7066
rect 13130 7032 13164 7066
rect 13198 7032 13232 7066
rect 13266 7032 13300 7066
rect 13334 7032 13368 7066
rect 13402 7032 13436 7066
rect 13470 7032 13504 7066
rect 13538 7032 13572 7066
rect 13606 7032 13640 7066
rect 13674 7032 13708 7066
rect 13742 7032 13776 7066
rect 13810 7032 13844 7066
rect 13878 7032 13912 7066
rect 13946 7032 13980 7066
rect 14014 7032 14048 7066
rect 14082 7032 14116 7066
rect 14150 7032 14184 7066
rect 14218 7032 14252 7066
rect 14286 7032 14320 7066
rect 14354 7032 14388 7066
rect 14422 7032 14456 7066
rect 14490 7032 14524 7066
rect 14558 7032 14592 7066
rect 14626 7032 14660 7066
rect 14694 7032 14728 7066
rect 14762 7032 14796 7066
rect 14830 7032 14864 7066
rect 14898 7065 15102 7066
rect 14898 7032 14932 7065
rect 8176 7031 14932 7032
rect 14966 7031 15000 7065
rect 15034 7031 15068 7065
rect 8176 6997 15102 7031
rect 3528 1031 3597 1065
rect 3631 1031 3666 1065
rect 3700 1031 3735 1065
rect 3769 1031 3804 1065
rect 3838 1031 3873 1065
rect 3907 1031 3942 1065
rect 3976 1031 4011 1065
rect 4045 1031 4080 1065
rect 4114 1031 4149 1065
rect 4183 1031 4218 1065
rect 4252 1031 4287 1065
rect 4321 1031 4356 1065
rect 4390 1031 4425 1065
rect 4459 1031 4494 1065
rect 4528 1031 4563 1065
rect 4597 1031 4632 1065
rect 4666 1031 4701 1065
rect 4735 1031 4770 1065
rect 4804 1031 4839 1065
rect 4873 1031 4908 1065
rect 4942 1031 4977 1065
rect 5011 1031 5046 1065
rect 5080 1031 5115 1065
rect 5149 1031 5184 1065
rect 5218 1031 5253 1065
rect 5287 1031 5322 1065
rect 5356 1031 5392 1065
rect 5426 1031 5462 1065
rect 5496 1031 5532 1065
rect 5566 1031 5602 1065
rect 5636 1031 5672 1065
rect 5706 1031 5742 1065
rect 5776 1031 5812 1065
rect 5846 1031 5882 1065
rect 5916 1031 5952 1065
rect 5986 1031 6022 1065
rect 6056 1031 6092 1065
rect 6126 1031 6162 1065
rect 6196 1031 6232 1065
rect 6266 1031 6302 1065
rect 6336 1031 6372 1065
rect 6406 1031 6442 1065
rect 6476 1031 6512 1065
rect 6546 1031 6582 1065
rect 6616 1031 6652 1065
rect 6686 1031 6722 1065
rect 6756 1031 6824 1065
rect 3528 209 3562 1031
rect 6790 966 6824 1031
rect 6790 845 6824 932
rect 6790 777 6824 811
rect 6790 709 6824 743
rect 6790 641 6824 675
rect 6790 573 6824 607
rect 6790 505 6824 539
rect 6790 437 6824 471
rect 6790 369 6824 403
rect 6790 301 6824 335
rect 6790 233 6824 267
rect 3528 175 3632 209
rect 3666 175 3700 209
rect 3734 175 3768 209
rect 3802 175 3836 209
rect 3870 175 3904 209
rect 3938 175 3972 209
rect 4006 175 4040 209
rect 4074 175 4108 209
rect 4142 175 4176 209
rect 4210 175 4244 209
rect 4278 175 4312 209
rect 4346 175 4380 209
rect 4414 175 4448 209
rect 4482 175 4516 209
rect 4550 175 4584 209
rect 4618 175 4652 209
rect 4686 175 4720 209
rect 4754 175 4788 209
rect 4822 175 4856 209
rect 4890 175 4924 209
rect 4958 175 4992 209
rect 5026 175 5060 209
rect 5094 175 5128 209
rect 5162 175 5196 209
rect 5230 175 5264 209
rect 5298 175 5332 209
rect 5366 175 5400 209
rect 5434 175 5468 209
rect 5502 175 5536 209
rect 5570 175 5604 209
rect 5638 175 5672 209
rect 5706 175 5740 209
rect 5774 175 5808 209
rect 5842 175 5876 209
rect 5910 175 5944 209
rect 5978 175 6012 209
rect 6046 175 6080 209
rect 6114 175 6148 209
rect 6182 175 6216 209
rect 6250 175 6284 209
rect 6318 175 6352 209
rect 6386 175 6420 209
rect 6454 175 6488 209
rect 6522 175 6556 209
rect 6590 175 6624 209
rect 6658 175 6692 209
rect 6726 199 6790 209
rect 6726 175 6824 199
<< mvpsubdiffcont >>
rect 698 15387 732 15421
rect 767 15387 801 15421
rect 836 15387 870 15421
rect 905 15387 939 15421
rect 974 15387 1008 15421
rect 1043 15387 1077 15421
rect 1112 15387 1146 15421
rect 1181 15387 1215 15421
rect 1250 15387 1284 15421
rect 1319 15387 1353 15421
rect 1388 15387 1422 15421
rect 1457 15387 1491 15421
rect 1526 15387 1560 15421
rect 1595 15387 1629 15421
rect 1664 15387 1698 15421
rect 1733 15387 1767 15421
rect 1802 15387 1836 15421
rect 1871 15387 1905 15421
rect 1940 15387 1974 15421
rect 2009 15387 2043 15421
rect 2078 15387 2112 15421
rect 2147 15387 2181 15421
rect 2216 15387 2250 15421
rect 2285 15387 2319 15421
rect 2354 15387 2388 15421
rect 2423 15387 2457 15421
rect 2492 15387 2526 15421
rect 2561 15387 2595 15421
rect 2630 15387 2664 15421
rect 2699 15387 2733 15421
rect 2768 15387 2802 15421
rect 2837 15387 2871 15421
rect 2906 15387 2940 15421
rect 2975 15387 3009 15421
rect 3044 15387 3078 15421
rect 3113 15387 3147 15421
rect 3182 15387 3216 15421
rect 3251 15387 3285 15421
rect 3320 15387 3354 15421
rect 3389 15387 3423 15421
rect 3458 15387 3492 15421
rect 3527 15387 3561 15421
rect 3596 15387 3630 15421
rect 3665 15387 3699 15421
rect 3734 15387 3768 15421
rect 3803 15387 3837 15421
rect 3872 15387 3906 15421
rect 3941 15387 3975 15421
rect 4010 15387 4044 15421
rect 4079 15387 4113 15421
rect 4148 15387 4182 15421
rect 4217 15387 4251 15421
rect 4286 15387 4320 15421
rect 4355 15387 4389 15421
rect 4424 15387 4458 15421
rect 4493 15387 4527 15421
rect 4562 15387 4596 15421
rect 4631 15387 4665 15421
rect 4700 15387 4734 15421
rect 4769 15387 4803 15421
rect 4838 15387 4872 15421
rect 4907 15387 4941 15421
rect 4976 15387 5010 15421
rect 5045 15387 5079 15421
rect 5114 15387 5148 15421
rect 674 15289 708 15323
rect 5208 15363 5242 15397
rect 674 15218 708 15252
rect 674 15147 708 15181
rect 5208 15250 5242 15284
rect 674 15075 708 15109
rect 5208 15116 5242 15150
rect 674 15003 708 15037
rect 768 14979 802 15013
rect 837 14979 871 15013
rect 906 14979 940 15013
rect 975 14979 1009 15013
rect 1044 14979 1078 15013
rect 1113 14979 1147 15013
rect 1182 14979 1216 15013
rect 1251 14979 1285 15013
rect 1320 14979 1354 15013
rect 1389 14979 1423 15013
rect 1458 14979 1492 15013
rect 1527 14979 1561 15013
rect 1596 14979 1630 15013
rect 1665 14979 1699 15013
rect 1734 14979 1768 15013
rect 1803 14979 1837 15013
rect 1872 14979 1906 15013
rect 1941 14979 1975 15013
rect 2010 14979 2044 15013
rect 2079 14979 2113 15013
rect 2148 14979 2182 15013
rect 2217 14979 2251 15013
rect 2286 14979 2320 15013
rect 2355 14979 2389 15013
rect 2424 14979 2458 15013
rect 2493 14979 2527 15013
rect 2562 14979 2596 15013
rect 2631 14979 2665 15013
rect 2700 14979 2734 15013
rect 2769 14979 2803 15013
rect 2838 14979 2872 15013
rect 2907 14979 2941 15013
rect 2976 14979 3010 15013
rect 3045 14979 3079 15013
rect 3114 14979 3148 15013
rect 3183 14979 3217 15013
rect 3252 14979 3286 15013
rect 3321 14979 3355 15013
rect 3390 14979 3424 15013
rect 3459 14979 3493 15013
rect 3528 14979 3562 15013
rect 3597 14979 3631 15013
rect 3666 14979 3700 15013
rect 3735 14979 3769 15013
rect 3804 14979 3838 15013
rect 3873 14979 3907 15013
rect 3942 14979 3976 15013
rect 4011 14979 4045 15013
rect 4080 14979 4114 15013
rect 4149 14979 4183 15013
rect 4218 14979 4252 15013
rect 4287 14979 4321 15013
rect 4356 14979 4390 15013
rect 4425 14979 4459 15013
rect 4494 14979 4528 15013
rect 4563 14979 4597 15013
rect 4632 14979 4666 15013
rect 4701 14979 4735 15013
rect 4770 14979 4804 15013
rect 4839 14979 4873 15013
rect 4908 14979 4942 15013
rect 4977 14979 5011 15013
rect 5046 14979 5080 15013
rect 5115 14979 5149 15013
rect 5184 14979 5218 15013
rect -932 9613 -898 9647
rect -864 9613 -830 9647
rect -796 9613 -762 9647
rect -723 9646 -689 9680
rect -654 9646 -620 9680
rect -585 9646 -551 9680
rect -516 9646 -482 9680
rect -447 9646 -413 9680
rect -378 9646 -344 9680
rect -309 9646 -275 9680
rect -240 9646 -206 9680
rect -171 9646 -137 9680
rect -102 9646 -68 9680
rect -723 9578 -689 9612
rect -654 9578 -620 9612
rect -585 9578 -551 9612
rect -516 9578 -482 9612
rect -447 9578 -413 9612
rect -378 9578 -344 9612
rect -309 9578 -275 9612
rect -240 9578 -206 9612
rect -171 9578 -137 9612
rect -102 9578 -68 9612
rect -932 9537 -898 9571
rect -864 9537 -830 9571
rect -796 9537 -762 9571
rect -723 9510 -689 9544
rect -654 9510 -620 9544
rect -585 9510 -551 9544
rect -516 9510 -482 9544
rect -447 9510 -413 9544
rect -378 9510 -344 9544
rect -309 9510 -275 9544
rect -240 9510 -206 9544
rect -171 9510 -137 9544
rect -102 9510 -68 9544
rect -932 9461 -898 9495
rect -864 9461 -830 9495
rect -796 9461 -762 9495
rect -723 9442 -689 9476
rect -654 9442 -620 9476
rect -585 9442 -551 9476
rect -516 9442 -482 9476
rect -447 9442 -413 9476
rect -378 9442 -344 9476
rect -309 9442 -275 9476
rect -240 9442 -206 9476
rect -171 9442 -137 9476
rect -102 9442 -68 9476
rect -932 9384 -898 9418
rect -864 9384 -830 9418
rect -796 9384 -762 9418
rect -723 9374 -689 9408
rect -654 9374 -620 9408
rect -585 9374 -551 9408
rect -516 9374 -482 9408
rect -447 9374 -413 9408
rect -378 9374 -344 9408
rect -309 9374 -275 9408
rect -240 9374 -206 9408
rect -171 9374 -137 9408
rect -102 9374 -68 9408
rect -932 9307 -898 9341
rect -864 9307 -830 9341
rect -796 9307 -762 9341
rect -723 9306 -689 9340
rect -654 9306 -620 9340
rect -585 9306 -551 9340
rect -516 9306 -482 9340
rect -447 9306 -413 9340
rect -378 9306 -344 9340
rect -309 9306 -275 9340
rect -240 9306 -206 9340
rect -171 9306 -137 9340
rect -102 9306 -68 9340
rect -932 9230 -898 9264
rect -864 9230 -830 9264
rect -796 9230 -762 9264
rect -723 9238 -689 9272
rect -654 9238 -620 9272
rect -585 9238 -551 9272
rect -516 9238 -482 9272
rect -447 9238 -413 9272
rect -378 9238 -344 9272
rect -309 9238 -275 9272
rect -240 9238 -206 9272
rect -171 9238 -137 9272
rect -102 9238 -68 9272
rect -932 9153 -898 9187
rect -864 9153 -830 9187
rect -796 9153 -762 9187
rect -723 9170 -689 9204
rect -654 9170 -620 9204
rect -585 9170 -551 9204
rect -516 9170 -482 9204
rect -447 9170 -413 9204
rect -378 9170 -344 9204
rect -309 9170 -275 9204
rect -240 9170 -206 9204
rect -171 9170 -137 9204
rect -102 9170 -68 9204
rect -932 9076 -898 9110
rect -864 9076 -830 9110
rect -796 9076 -762 9110
rect -723 9102 -689 9136
rect -654 9102 -620 9136
rect -585 9102 -551 9136
rect -516 9102 -482 9136
rect -447 9102 -413 9136
rect -378 9102 -344 9136
rect -309 9102 -275 9136
rect -240 9102 -206 9136
rect -171 9102 -137 9136
rect -102 9102 -68 9136
rect -723 9034 -689 9068
rect -654 9034 -620 9068
rect -585 9034 -551 9068
rect -516 9034 -482 9068
rect -447 9034 -413 9068
rect -378 9034 -344 9068
rect -309 9034 -275 9068
rect -240 9034 -206 9068
rect -171 9034 -137 9068
rect -102 9034 -68 9068
rect -932 8999 -898 9033
rect -864 8999 -830 9033
rect -796 8999 -762 9033
rect -723 8966 -689 9000
rect -654 8966 -620 9000
rect -585 8966 -551 9000
rect -516 8966 -482 9000
rect -447 8966 -413 9000
rect -378 8966 -344 9000
rect -309 8966 -275 9000
rect -240 8966 -206 9000
rect -171 8966 -137 9000
rect -102 8966 -68 9000
rect -33 8966 14893 9680
rect 14932 9613 14966 9647
rect 15000 9613 15034 9647
rect 15068 9613 15102 9647
rect 14932 9537 14966 9571
rect 15000 9537 15034 9571
rect 15068 9537 15102 9571
rect 14932 9461 14966 9495
rect 15000 9461 15034 9495
rect 15068 9461 15102 9495
rect 14932 9384 14966 9418
rect 15000 9384 15034 9418
rect 15068 9384 15102 9418
rect 14932 9307 14966 9341
rect 15000 9307 15034 9341
rect 15068 9307 15102 9341
rect 14932 9230 14966 9264
rect 15000 9230 15034 9264
rect 15068 9230 15102 9264
rect 14932 9153 14966 9187
rect 15000 9153 15034 9187
rect 15068 9153 15102 9187
rect 14932 9076 14966 9110
rect 15000 9076 15034 9110
rect 15068 9076 15102 9110
rect 14932 8999 14966 9033
rect 15000 8999 15034 9033
rect 15068 8999 15102 9033
rect 68 6809 102 6843
rect 137 6809 171 6843
rect 206 6809 240 6843
rect 275 6809 309 6843
rect 344 6809 378 6843
rect 413 6809 447 6843
rect 482 6809 516 6843
rect 551 6809 585 6843
rect 620 6809 654 6843
rect 689 6809 723 6843
rect 758 6809 792 6843
rect 827 6809 861 6843
rect 896 6809 930 6843
rect 965 6809 999 6843
rect 1034 6809 1068 6843
rect 1103 6809 1137 6843
rect 1172 6809 1206 6843
rect 1241 6809 1275 6843
rect 1310 6809 1344 6843
rect 1379 6809 1413 6843
rect 1448 6809 1482 6843
rect 1517 6809 1551 6843
rect 1586 6809 1620 6843
rect 1655 6809 1689 6843
rect 1724 6809 1758 6843
rect 1793 6809 1827 6843
rect 1862 6809 1896 6843
rect 1931 6809 1965 6843
rect 2000 6809 2034 6843
rect 2069 6809 2103 6843
rect 2138 6809 2172 6843
rect 2207 6809 2241 6843
rect 2276 6809 2310 6843
rect 2345 6809 2379 6843
rect 2414 6809 2448 6843
rect 2483 6809 2517 6843
rect 2552 6809 2586 6843
rect 2621 6809 2655 6843
rect 2690 6809 2724 6843
rect 2759 6809 2793 6843
rect 2828 6809 2862 6843
rect 2897 6809 2931 6843
rect 2966 6809 3000 6843
rect 3035 6809 3069 6843
rect 3104 6809 3138 6843
rect 3173 6809 3207 6843
rect 3242 6809 3276 6843
rect 3310 6809 3344 6843
rect 3378 6809 3412 6843
rect 3446 6809 3480 6843
rect 3514 6809 3548 6843
rect 3582 6809 3616 6843
rect 3650 6809 3684 6843
rect 3718 6809 3752 6843
rect 3786 6809 3820 6843
rect 3854 6809 3888 6843
rect 3922 6809 3956 6843
rect 3990 6809 4024 6843
rect 4058 6809 4092 6843
rect 4126 6809 4160 6843
rect 4194 6809 4228 6843
rect 4262 6809 4296 6843
rect 4330 6809 4364 6843
rect 4398 6809 4432 6843
rect 4466 6809 4500 6843
rect 4534 6809 4568 6843
rect 4602 6809 4636 6843
rect 4670 6809 4704 6843
rect 4738 6809 4772 6843
rect 4806 6809 4840 6843
rect 4874 6809 4908 6843
rect 4942 6809 4976 6843
rect 5010 6809 5044 6843
rect 5078 6809 5112 6843
rect 5146 6809 5180 6843
rect 5214 6809 5248 6843
rect 5282 6809 5316 6843
rect 5350 6809 5384 6843
rect 5418 6809 5452 6843
rect 5486 6809 5520 6843
rect 5554 6809 5588 6843
rect 5622 6809 5656 6843
rect 5690 6809 5724 6843
rect 5758 6809 5792 6843
rect 5826 6809 5860 6843
rect 5894 6809 5928 6843
rect 5962 6809 5996 6843
rect 6030 6809 6064 6843
rect 6098 6809 6132 6843
rect 6166 6809 6200 6843
rect 6234 6809 6268 6843
rect 6302 6809 6336 6843
rect 6370 6809 6404 6843
rect 6438 6809 6472 6843
rect 6506 6809 6540 6843
rect 6574 6809 6608 6843
rect 6642 6809 6676 6843
rect 6710 6809 6744 6843
rect 6778 6809 6812 6843
rect 6846 6809 6880 6843
rect 6914 6809 6948 6843
rect 6982 6809 7016 6843
rect 7050 6809 7084 6843
rect 68 6722 102 6756
rect 137 6722 171 6756
rect 206 6722 240 6756
rect 275 6722 309 6756
rect 344 6722 378 6756
rect 413 6722 447 6756
rect 482 6722 516 6756
rect 551 6722 585 6756
rect 620 6722 654 6756
rect 689 6722 723 6756
rect 758 6722 792 6756
rect 827 6722 861 6756
rect 896 6722 930 6756
rect 965 6722 999 6756
rect 1034 6722 1068 6756
rect 1103 6722 1137 6756
rect 1172 6722 1206 6756
rect 1241 6722 1275 6756
rect 1310 6722 1344 6756
rect 1379 6722 1413 6756
rect 1448 6722 1482 6756
rect 1517 6722 1551 6756
rect 1586 6722 1620 6756
rect 1655 6722 1689 6756
rect 1724 6722 1758 6756
rect 1793 6722 1827 6756
rect 1862 6722 1896 6756
rect 1931 6722 1965 6756
rect 2000 6722 2034 6756
rect 2069 6722 2103 6756
rect 2138 6722 2172 6756
rect 2207 6722 2241 6756
rect 2276 6722 2310 6756
rect 2345 6722 2379 6756
rect 2414 6722 2448 6756
rect 2483 6722 2517 6756
rect 2552 6722 2586 6756
rect 2621 6722 2655 6756
rect 2690 6722 2724 6756
rect 2759 6722 2793 6756
rect 2828 6722 2862 6756
rect 2897 6722 2931 6756
rect 2966 6722 3000 6756
rect 3035 6722 3069 6756
rect 3104 6722 3138 6756
rect 3173 6722 3207 6756
rect 3242 6722 3276 6756
rect 3310 6722 3344 6756
rect 3378 6722 3412 6756
rect 3446 6722 3480 6756
rect 3514 6722 3548 6756
rect 3582 6722 3616 6756
rect 3650 6722 3684 6756
rect 3718 6722 3752 6756
rect 3786 6722 3820 6756
rect 3854 6722 3888 6756
rect 3922 6722 3956 6756
rect 3990 6722 4024 6756
rect 4058 6722 4092 6756
rect 4126 6722 4160 6756
rect 4194 6722 4228 6756
rect 4262 6722 4296 6756
rect 4330 6722 4364 6756
rect 4398 6722 4432 6756
rect 4466 6722 4500 6756
rect 4534 6722 4568 6756
rect 4602 6722 4636 6756
rect 4670 6722 4704 6756
rect 4738 6722 4772 6756
rect 4806 6722 4840 6756
rect 4874 6722 4908 6756
rect 4942 6722 4976 6756
rect 5010 6722 5044 6756
rect 5078 6722 5112 6756
rect 5146 6722 5180 6756
rect 5214 6722 5248 6756
rect 5282 6722 5316 6756
rect 5350 6722 5384 6756
rect 5418 6722 5452 6756
rect 5486 6722 5520 6756
rect 5554 6722 5588 6756
rect 5622 6722 5656 6756
rect 5690 6722 5724 6756
rect 5758 6722 5792 6756
rect 5826 6722 5860 6756
rect 5894 6722 5928 6756
rect 5962 6722 5996 6756
rect 6030 6722 6064 6756
rect 6098 6722 6132 6756
rect 6166 6722 6200 6756
rect 6234 6722 6268 6756
rect 6302 6722 6336 6756
rect 6370 6722 6404 6756
rect 6438 6722 6472 6756
rect 6506 6722 6540 6756
rect 6574 6722 6608 6756
rect 6642 6722 6676 6756
rect 6710 6722 6744 6756
rect 6778 6722 6812 6756
rect 6846 6722 6880 6756
rect 6914 6722 6948 6756
rect 6982 6722 7016 6756
rect 7050 6722 7084 6756
rect 68 6635 102 6669
rect 137 6635 171 6669
rect 206 6635 240 6669
rect 275 6635 309 6669
rect 344 6635 378 6669
rect 413 6635 447 6669
rect 482 6635 516 6669
rect 551 6635 585 6669
rect 620 6635 654 6669
rect 689 6635 723 6669
rect 758 6635 792 6669
rect 827 6635 861 6669
rect 896 6635 930 6669
rect 965 6635 999 6669
rect 1034 6635 1068 6669
rect 1103 6635 1137 6669
rect 1172 6635 1206 6669
rect 1241 6635 1275 6669
rect 1310 6635 1344 6669
rect 1379 6635 1413 6669
rect 1448 6635 1482 6669
rect 1517 6635 1551 6669
rect 1586 6635 1620 6669
rect 1655 6635 1689 6669
rect 1724 6635 1758 6669
rect 1793 6635 1827 6669
rect 1862 6635 1896 6669
rect 1931 6635 1965 6669
rect 2000 6635 2034 6669
rect 2069 6635 2103 6669
rect 2138 6635 2172 6669
rect 2207 6635 2241 6669
rect 2276 6635 2310 6669
rect 2345 6635 2379 6669
rect 2414 6635 2448 6669
rect 2483 6635 2517 6669
rect 2552 6635 2586 6669
rect 2621 6635 2655 6669
rect 2690 6635 2724 6669
rect 2759 6635 2793 6669
rect 2828 6635 2862 6669
rect 2897 6635 2931 6669
rect 2966 6635 3000 6669
rect 3035 6635 3069 6669
rect 3104 6635 3138 6669
rect 3173 6635 3207 6669
rect 3242 6635 3276 6669
rect 3310 6635 3344 6669
rect 3378 6635 3412 6669
rect 3446 6635 3480 6669
rect 3514 6635 3548 6669
rect 3582 6635 3616 6669
rect 3650 6635 3684 6669
rect 3718 6635 3752 6669
rect 3786 6635 3820 6669
rect 3854 6635 3888 6669
rect 3922 6635 3956 6669
rect 3990 6635 4024 6669
rect 4058 6635 4092 6669
rect 4126 6635 4160 6669
rect 4194 6635 4228 6669
rect 4262 6635 4296 6669
rect 4330 6635 4364 6669
rect 4398 6635 4432 6669
rect 4466 6635 4500 6669
rect 4534 6635 4568 6669
rect 4602 6635 4636 6669
rect 4670 6635 4704 6669
rect 4738 6635 4772 6669
rect 4806 6635 4840 6669
rect 4874 6635 4908 6669
rect 4942 6635 4976 6669
rect 5010 6635 5044 6669
rect 5078 6635 5112 6669
rect 5146 6635 5180 6669
rect 5214 6635 5248 6669
rect 5282 6635 5316 6669
rect 5350 6635 5384 6669
rect 5418 6635 5452 6669
rect 5486 6635 5520 6669
rect 5554 6635 5588 6669
rect 5622 6635 5656 6669
rect 5690 6635 5724 6669
rect 5758 6635 5792 6669
rect 5826 6635 5860 6669
rect 5894 6635 5928 6669
rect 5962 6635 5996 6669
rect 6030 6635 6064 6669
rect 6098 6635 6132 6669
rect 6166 6635 6200 6669
rect 6234 6635 6268 6669
rect 6302 6635 6336 6669
rect 6370 6635 6404 6669
rect 6438 6635 6472 6669
rect 6506 6635 6540 6669
rect 6574 6635 6608 6669
rect 6642 6635 6676 6669
rect 6710 6635 6744 6669
rect 6778 6635 6812 6669
rect 6846 6635 6880 6669
rect 6914 6635 6948 6669
rect 6982 6635 7016 6669
rect 7050 6635 7084 6669
rect 12517 6809 12551 6843
rect 12586 6809 12620 6843
rect 12655 6809 12689 6843
rect 12724 6809 12758 6843
rect 12793 6809 12827 6843
rect 12862 6809 12896 6843
rect 12931 6809 12965 6843
rect 13000 6809 13034 6843
rect 13069 6809 13103 6843
rect 13138 6809 13172 6843
rect 13207 6809 13241 6843
rect 13276 6809 13310 6843
rect 13345 6809 13379 6843
rect 13414 6809 13448 6843
rect 13483 6809 13517 6843
rect 13552 6809 13586 6843
rect 13621 6809 13655 6843
rect 13690 6809 13724 6843
rect 13759 6809 13793 6843
rect 13828 6809 13862 6843
rect 13897 6809 13931 6843
rect 13966 6809 14000 6843
rect 14035 6809 14069 6843
rect 14104 6809 14138 6843
rect 14173 6809 14207 6843
rect 14242 6809 14276 6843
rect 14311 6809 14345 6843
rect 14380 6809 14414 6843
rect 14449 6809 14483 6843
rect 14518 6809 14552 6843
rect 14587 6809 14621 6843
rect 14655 6809 14689 6843
rect 14723 6809 14757 6843
rect 14791 6809 14825 6843
rect 14859 6809 14893 6843
rect 14932 6771 14966 6805
rect 15000 6771 15034 6805
rect 15068 6771 15102 6805
rect 12517 6722 12551 6756
rect 12586 6722 12620 6756
rect 12655 6722 12689 6756
rect 12724 6722 12758 6756
rect 12793 6722 12827 6756
rect 12862 6722 12896 6756
rect 12931 6722 12965 6756
rect 13000 6722 13034 6756
rect 13069 6722 13103 6756
rect 13138 6722 13172 6756
rect 13207 6722 13241 6756
rect 13276 6722 13310 6756
rect 13345 6722 13379 6756
rect 13414 6722 13448 6756
rect 13483 6722 13517 6756
rect 13552 6722 13586 6756
rect 13621 6722 13655 6756
rect 13690 6722 13724 6756
rect 13759 6722 13793 6756
rect 13828 6722 13862 6756
rect 13897 6722 13931 6756
rect 13966 6722 14000 6756
rect 14035 6722 14069 6756
rect 14104 6722 14138 6756
rect 14173 6722 14207 6756
rect 14242 6722 14276 6756
rect 14311 6722 14345 6756
rect 14380 6722 14414 6756
rect 14449 6722 14483 6756
rect 14518 6722 14552 6756
rect 14587 6722 14621 6756
rect 14655 6722 14689 6756
rect 14723 6722 14757 6756
rect 14791 6722 14825 6756
rect 14859 6722 14893 6756
rect 14932 6697 14966 6731
rect 15000 6697 15034 6731
rect 15068 6697 15102 6731
rect 12517 6635 12551 6669
rect 12586 6635 12620 6669
rect 12655 6635 12689 6669
rect 12724 6635 12758 6669
rect 12793 6635 12827 6669
rect 12862 6635 12896 6669
rect 12931 6635 12965 6669
rect 13000 6635 13034 6669
rect 13069 6635 13103 6669
rect 13138 6635 13172 6669
rect 13207 6635 13241 6669
rect 13276 6635 13310 6669
rect 13345 6635 13379 6669
rect 13414 6635 13448 6669
rect 13483 6635 13517 6669
rect 13552 6635 13586 6669
rect 13621 6635 13655 6669
rect 13690 6635 13724 6669
rect 13759 6635 13793 6669
rect 13828 6635 13862 6669
rect 13897 6635 13931 6669
rect 13966 6635 14000 6669
rect 14035 6635 14069 6669
rect 14104 6635 14138 6669
rect 14173 6635 14207 6669
rect 14242 6635 14276 6669
rect 14311 6635 14345 6669
rect 14380 6635 14414 6669
rect 14449 6635 14483 6669
rect 14518 6635 14552 6669
rect 14587 6635 14621 6669
rect 14655 6635 14689 6669
rect 14723 6635 14757 6669
rect 14791 6635 14825 6669
rect 14859 6635 14893 6669
rect 14932 6623 14966 6657
rect 15000 6623 15034 6657
rect 15068 6623 15102 6657
rect 68 6548 102 6582
rect 137 6548 171 6582
rect 206 6548 240 6582
rect 275 6548 309 6582
rect 344 6548 378 6582
rect 413 6548 447 6582
rect 482 6548 516 6582
rect 551 6548 585 6582
rect 620 6548 654 6582
rect 689 6548 723 6582
rect 758 6548 792 6582
rect 827 6548 861 6582
rect 896 6548 930 6582
rect 965 6548 999 6582
rect 1034 6548 1068 6582
rect 1103 6548 1137 6582
rect 1172 6548 1206 6582
rect 1241 6548 1275 6582
rect 1310 6548 1344 6582
rect 1379 6548 1413 6582
rect 1448 6548 1482 6582
rect 1517 6548 1551 6582
rect 1586 6548 1620 6582
rect 1655 6548 1689 6582
rect 1724 6548 1758 6582
rect 1793 6548 1827 6582
rect 1862 6548 1896 6582
rect 1931 6548 1965 6582
rect 2000 6548 2034 6582
rect 2069 6548 2103 6582
rect 2138 6548 2172 6582
rect 2207 6548 2241 6582
rect 2276 6548 2310 6582
rect 2345 6548 2379 6582
rect 2414 6548 2448 6582
rect 2483 6548 2517 6582
rect 2551 6548 2585 6582
rect 2619 6548 2653 6582
rect 2687 6548 2721 6582
rect 2755 6548 2789 6582
rect 2823 6548 2857 6582
rect 2891 6548 2925 6582
rect 2959 6548 2993 6582
rect 3027 6548 3061 6582
rect 3095 6548 3129 6582
rect 3163 6548 3197 6582
rect 3231 6548 3265 6582
rect 3299 6548 3333 6582
rect 3367 6548 3401 6582
rect 3435 6548 3469 6582
rect 3503 6548 3537 6582
rect 3571 6548 3605 6582
rect 3639 6548 3673 6582
rect 3707 6548 3741 6582
rect 3775 6548 3809 6582
rect 3843 6548 3877 6582
rect 3911 6548 3945 6582
rect 3979 6548 4013 6582
rect 4047 6548 4081 6582
rect 4115 6548 4149 6582
rect 4183 6548 4217 6582
rect 4251 6548 4285 6582
rect 4319 6548 4353 6582
rect 4387 6548 4421 6582
rect 4455 6548 4489 6582
rect 4523 6548 4557 6582
rect 4591 6548 4625 6582
rect 4659 6548 4693 6582
rect 4727 6548 4761 6582
rect 4795 6548 4829 6582
rect 4863 6548 4897 6582
rect 4931 6548 4965 6582
rect 4999 6548 5033 6582
rect 5067 6548 5101 6582
rect 5135 6548 5169 6582
rect 5203 6548 5237 6582
rect 5271 6548 5305 6582
rect 5339 6548 5373 6582
rect 5407 6548 5441 6582
rect 5475 6548 5509 6582
rect 5543 6548 5577 6582
rect 5611 6548 5645 6582
rect 5679 6548 5713 6582
rect 5747 6548 5781 6582
rect 5815 6548 5849 6582
rect 5883 6548 5917 6582
rect 5951 6548 5985 6582
rect 6019 6548 6053 6582
rect 6087 6548 6121 6582
rect 6155 6548 6189 6582
rect 6223 6548 6257 6582
rect 6291 6548 6325 6582
rect 6359 6548 6393 6582
rect 6427 6548 6461 6582
rect 6495 6548 6529 6582
rect 6563 6548 6597 6582
rect 6631 6548 6665 6582
rect 6699 6548 6733 6582
rect 6767 6548 6801 6582
rect 6835 6548 6869 6582
rect 6903 6548 6937 6582
rect 6971 6548 7005 6582
rect 7039 6548 7073 6582
rect 7107 6548 7141 6582
rect 7175 6548 7209 6582
rect 7243 6548 7277 6582
rect 7311 6548 7345 6582
rect 7379 6548 7413 6582
rect 7447 6548 7481 6582
rect 7515 6548 7549 6582
rect 7583 6548 7617 6582
rect 7651 6548 7685 6582
rect 7719 6548 7753 6582
rect 7787 6548 7821 6582
rect 7855 6548 7889 6582
rect 7923 6548 7957 6582
rect 7991 6548 8025 6582
rect 8059 6548 8093 6582
rect 8127 6548 8161 6582
rect 8195 6548 8229 6582
rect 8263 6548 8297 6582
rect 8331 6548 8365 6582
rect 8399 6548 8433 6582
rect 8467 6548 8501 6582
rect 8535 6548 8569 6582
rect 8603 6548 8637 6582
rect 8671 6548 8705 6582
rect 8739 6548 8773 6582
rect 8807 6548 8841 6582
rect 8875 6548 8909 6582
rect 8943 6548 8977 6582
rect 9011 6548 9045 6582
rect 9079 6548 9113 6582
rect 9147 6548 9181 6582
rect 9215 6548 9249 6582
rect 9283 6548 9317 6582
rect 9351 6548 9385 6582
rect 9419 6548 9453 6582
rect 9487 6548 9521 6582
rect 9555 6548 9589 6582
rect 9623 6548 9657 6582
rect 9691 6548 9725 6582
rect 9759 6548 9793 6582
rect 9827 6548 9861 6582
rect 9895 6548 9929 6582
rect 9963 6548 9997 6582
rect 10031 6548 10065 6582
rect 10099 6548 10133 6582
rect 10167 6548 10201 6582
rect 10235 6548 10269 6582
rect 10303 6548 10337 6582
rect 10371 6548 10405 6582
rect 10439 6548 10473 6582
rect 10507 6548 10541 6582
rect 10575 6548 10609 6582
rect 10643 6548 10677 6582
rect 10711 6548 10745 6582
rect 10779 6548 10813 6582
rect 10847 6548 10881 6582
rect 10915 6548 10949 6582
rect 10983 6548 11017 6582
rect 11051 6548 11085 6582
rect 11119 6548 11153 6582
rect 11187 6548 11221 6582
rect 11255 6548 11289 6582
rect 11323 6548 11357 6582
rect 11391 6548 11425 6582
rect 11459 6548 11493 6582
rect 11527 6548 11561 6582
rect 11595 6548 11629 6582
rect 11663 6548 11697 6582
rect 11731 6548 11765 6582
rect 11799 6548 11833 6582
rect 11867 6548 11901 6582
rect 11935 6548 11969 6582
rect 12003 6548 12037 6582
rect 12071 6548 12105 6582
rect 12139 6548 12173 6582
rect 12207 6548 12241 6582
rect 12275 6548 12309 6582
rect 12343 6548 12377 6582
rect 12411 6548 12445 6582
rect 12479 6548 12513 6582
rect 12547 6548 12581 6582
rect 12615 6548 12649 6582
rect 12683 6548 12717 6582
rect 12751 6548 12785 6582
rect 12819 6548 12853 6582
rect 12887 6548 12921 6582
rect 12955 6548 12989 6582
rect 13023 6548 13057 6582
rect 13091 6548 13125 6582
rect 13159 6548 13193 6582
rect 13227 6548 13261 6582
rect 13295 6548 13329 6582
rect 13363 6548 13397 6582
rect 13431 6548 13465 6582
rect 13499 6548 13533 6582
rect 13567 6548 13601 6582
rect 13635 6548 13669 6582
rect 13703 6548 13737 6582
rect 13771 6548 13805 6582
rect 13839 6548 13873 6582
rect 13907 6548 13941 6582
rect 13975 6548 14009 6582
rect 14043 6548 14077 6582
rect 14111 6548 14145 6582
rect 14179 6548 14213 6582
rect 14247 6548 14281 6582
rect 14315 6548 14349 6582
rect 14383 6548 14417 6582
rect 14451 6548 14485 6582
rect 14519 6548 14553 6582
rect 14587 6548 14621 6582
rect 14655 6548 14689 6582
rect 14723 6548 14757 6582
rect 14791 6548 14825 6582
rect 14859 6548 14893 6582
rect 14932 6549 14966 6583
rect 15000 6549 15034 6583
rect 15068 6549 15102 6583
rect 68 6474 102 6508
rect 137 6474 171 6508
rect 206 6474 240 6508
rect 275 6474 309 6508
rect 344 6474 378 6508
rect 413 6474 447 6508
rect 482 6474 516 6508
rect 551 6474 585 6508
rect 620 6474 654 6508
rect 689 6474 723 6508
rect 758 6474 792 6508
rect 827 6474 861 6508
rect 896 6474 930 6508
rect 965 6474 999 6508
rect 1034 6474 1068 6508
rect 1103 6474 1137 6508
rect 1172 6474 1206 6508
rect 1241 6474 1275 6508
rect 1310 6474 1344 6508
rect 1379 6474 1413 6508
rect 1448 6474 1482 6508
rect 1517 6474 1551 6508
rect 1586 6474 1620 6508
rect 1655 6474 1689 6508
rect 1724 6474 1758 6508
rect 1793 6474 1827 6508
rect 1862 6474 1896 6508
rect 1931 6474 1965 6508
rect 2000 6474 2034 6508
rect 2069 6474 2103 6508
rect 2138 6474 2172 6508
rect 2207 6474 2241 6508
rect 2276 6474 2310 6508
rect 2345 6474 2379 6508
rect 2414 6474 2448 6508
rect 2483 6474 2517 6508
rect 2551 6474 2585 6508
rect 2619 6474 2653 6508
rect 2687 6474 2721 6508
rect 2755 6474 2789 6508
rect 2823 6474 2857 6508
rect 2891 6474 2925 6508
rect 2959 6474 2993 6508
rect 3027 6474 3061 6508
rect 3095 6474 3129 6508
rect 3163 6474 3197 6508
rect 3231 6474 3265 6508
rect 3299 6474 3333 6508
rect 3367 6474 3401 6508
rect 3435 6474 3469 6508
rect 3503 6474 3537 6508
rect 3571 6474 3605 6508
rect 3639 6474 3673 6508
rect 3707 6474 3741 6508
rect 3775 6474 3809 6508
rect 3843 6474 3877 6508
rect 3911 6474 3945 6508
rect 3979 6474 4013 6508
rect 4047 6474 4081 6508
rect 4115 6474 4149 6508
rect 4183 6474 4217 6508
rect 4251 6474 4285 6508
rect 4319 6474 4353 6508
rect 4387 6474 4421 6508
rect 4455 6474 4489 6508
rect 4523 6474 4557 6508
rect 4591 6474 4625 6508
rect 4659 6474 4693 6508
rect 4727 6474 4761 6508
rect 4795 6474 4829 6508
rect 4863 6474 4897 6508
rect 4931 6474 4965 6508
rect 4999 6474 5033 6508
rect 5067 6474 5101 6508
rect 5135 6474 5169 6508
rect 5203 6474 5237 6508
rect 5271 6474 5305 6508
rect 5339 6474 5373 6508
rect 5407 6474 5441 6508
rect 5475 6474 5509 6508
rect 5543 6474 5577 6508
rect 5611 6474 5645 6508
rect 5679 6474 5713 6508
rect 5747 6474 5781 6508
rect 5815 6474 5849 6508
rect 5883 6474 5917 6508
rect 5951 6474 5985 6508
rect 6019 6474 6053 6508
rect 6087 6474 6121 6508
rect 6155 6474 6189 6508
rect 6223 6474 6257 6508
rect 6291 6474 6325 6508
rect 6359 6474 6393 6508
rect 6427 6474 6461 6508
rect 6495 6474 6529 6508
rect 6563 6474 6597 6508
rect 6631 6474 6665 6508
rect 6699 6474 6733 6508
rect 6767 6474 6801 6508
rect 6835 6474 6869 6508
rect 6903 6474 6937 6508
rect 6971 6474 7005 6508
rect 7039 6474 7073 6508
rect 7107 6474 7141 6508
rect 7175 6474 7209 6508
rect 7243 6474 7277 6508
rect 7311 6474 7345 6508
rect 7379 6474 7413 6508
rect 7447 6474 7481 6508
rect 7515 6474 7549 6508
rect 7583 6474 7617 6508
rect 7651 6474 7685 6508
rect 7719 6474 7753 6508
rect 7787 6474 7821 6508
rect 7855 6474 7889 6508
rect 7923 6474 7957 6508
rect 7991 6474 8025 6508
rect 8059 6474 8093 6508
rect 8127 6474 8161 6508
rect 8195 6474 8229 6508
rect 8263 6474 8297 6508
rect 8331 6474 8365 6508
rect 8399 6474 8433 6508
rect 8467 6474 8501 6508
rect 8535 6474 8569 6508
rect 8603 6474 8637 6508
rect 8671 6474 8705 6508
rect 8739 6474 8773 6508
rect 8807 6474 8841 6508
rect 8875 6474 8909 6508
rect 8943 6474 8977 6508
rect 9011 6474 9045 6508
rect 9079 6474 9113 6508
rect 9147 6474 9181 6508
rect 9215 6474 9249 6508
rect 9283 6474 9317 6508
rect 9351 6474 9385 6508
rect 9419 6474 9453 6508
rect 9487 6474 9521 6508
rect 9555 6474 9589 6508
rect 9623 6474 9657 6508
rect 9691 6474 9725 6508
rect 9759 6474 9793 6508
rect 9827 6474 9861 6508
rect 9895 6474 9929 6508
rect 9963 6474 9997 6508
rect 10031 6474 10065 6508
rect 10099 6474 10133 6508
rect 10167 6474 10201 6508
rect 10235 6474 10269 6508
rect 10303 6474 10337 6508
rect 10371 6474 10405 6508
rect 10439 6474 10473 6508
rect 10507 6474 10541 6508
rect 10575 6474 10609 6508
rect 10643 6474 10677 6508
rect 10711 6474 10745 6508
rect 10779 6474 10813 6508
rect 10847 6474 10881 6508
rect 10915 6474 10949 6508
rect 10983 6474 11017 6508
rect 11051 6474 11085 6508
rect 11119 6474 11153 6508
rect 11187 6474 11221 6508
rect 11255 6474 11289 6508
rect 11323 6474 11357 6508
rect 11391 6474 11425 6508
rect 11459 6474 11493 6508
rect 11527 6474 11561 6508
rect 11595 6474 11629 6508
rect 11663 6474 11697 6508
rect 11731 6474 11765 6508
rect 11799 6474 11833 6508
rect 11867 6474 11901 6508
rect 11935 6474 11969 6508
rect 12003 6474 12037 6508
rect 12071 6474 12105 6508
rect 12139 6474 12173 6508
rect 12207 6474 12241 6508
rect 12275 6474 12309 6508
rect 12343 6474 12377 6508
rect 12411 6474 12445 6508
rect 12479 6474 12513 6508
rect 12547 6474 12581 6508
rect 12615 6474 12649 6508
rect 12683 6474 12717 6508
rect 12751 6474 12785 6508
rect 12819 6474 12853 6508
rect 12887 6474 12921 6508
rect 12955 6474 12989 6508
rect 13023 6474 13057 6508
rect 13091 6474 13125 6508
rect 13159 6474 13193 6508
rect 13227 6474 13261 6508
rect 13295 6474 13329 6508
rect 13363 6474 13397 6508
rect 13431 6474 13465 6508
rect 13499 6474 13533 6508
rect 13567 6474 13601 6508
rect 13635 6474 13669 6508
rect 13703 6474 13737 6508
rect 13771 6474 13805 6508
rect 13839 6474 13873 6508
rect 13907 6474 13941 6508
rect 13975 6474 14009 6508
rect 14043 6474 14077 6508
rect 14111 6474 14145 6508
rect 14179 6474 14213 6508
rect 14247 6474 14281 6508
rect 14315 6474 14349 6508
rect 14383 6474 14417 6508
rect 14451 6474 14485 6508
rect 14519 6474 14553 6508
rect 14587 6474 14621 6508
rect 14655 6474 14689 6508
rect 14723 6474 14757 6508
rect 14791 6474 14825 6508
rect 14859 6474 14893 6508
rect 14932 6475 14966 6509
rect 15000 6475 15034 6509
rect 15068 6475 15102 6509
rect 68 6400 102 6434
rect 137 6400 171 6434
rect 206 6400 240 6434
rect 275 6400 309 6434
rect 344 6400 378 6434
rect 413 6400 447 6434
rect 482 6400 516 6434
rect 551 6400 585 6434
rect 620 6400 654 6434
rect 689 6400 723 6434
rect 758 6400 792 6434
rect 827 6400 861 6434
rect 896 6400 930 6434
rect 965 6400 999 6434
rect 1034 6400 1068 6434
rect 1103 6400 1137 6434
rect 1172 6400 1206 6434
rect 1241 6400 1275 6434
rect 1310 6400 1344 6434
rect 1379 6400 1413 6434
rect 1448 6400 1482 6434
rect 1517 6400 1551 6434
rect 1586 6400 1620 6434
rect 1655 6400 1689 6434
rect 1724 6400 1758 6434
rect 1793 6400 1827 6434
rect 1862 6400 1896 6434
rect 1931 6400 1965 6434
rect 2000 6400 2034 6434
rect 2069 6400 2103 6434
rect 2138 6400 2172 6434
rect 2207 6400 2241 6434
rect 2276 6400 2310 6434
rect 2345 6400 2379 6434
rect 2414 6400 2448 6434
rect 2483 6400 2517 6434
rect 2551 6400 2585 6434
rect 2619 6400 2653 6434
rect 2687 6400 2721 6434
rect 2755 6400 2789 6434
rect 2823 6400 2857 6434
rect 2891 6400 2925 6434
rect 2959 6400 2993 6434
rect 3027 6400 3061 6434
rect 3095 6400 3129 6434
rect 3163 6400 3197 6434
rect 3231 6400 3265 6434
rect 3299 6400 3333 6434
rect 3367 6400 3401 6434
rect 3435 6400 3469 6434
rect 3503 6400 3537 6434
rect 3571 6400 3605 6434
rect 3639 6400 3673 6434
rect 3707 6400 3741 6434
rect 3775 6400 3809 6434
rect 3843 6400 3877 6434
rect 3911 6400 3945 6434
rect 3979 6400 4013 6434
rect 4047 6400 4081 6434
rect 4115 6400 4149 6434
rect 4183 6400 4217 6434
rect 4251 6400 4285 6434
rect 4319 6400 4353 6434
rect 4387 6400 4421 6434
rect 4455 6400 4489 6434
rect 4523 6400 4557 6434
rect 4591 6400 4625 6434
rect 4659 6400 4693 6434
rect 4727 6400 4761 6434
rect 4795 6400 4829 6434
rect 4863 6400 4897 6434
rect 4931 6400 4965 6434
rect 4999 6400 5033 6434
rect 5067 6400 5101 6434
rect 5135 6400 5169 6434
rect 5203 6400 5237 6434
rect 5271 6400 5305 6434
rect 5339 6400 5373 6434
rect 5407 6400 5441 6434
rect 5475 6400 5509 6434
rect 5543 6400 5577 6434
rect 5611 6400 5645 6434
rect 5679 6400 5713 6434
rect 5747 6400 5781 6434
rect 5815 6400 5849 6434
rect 5883 6400 5917 6434
rect 5951 6400 5985 6434
rect 6019 6400 6053 6434
rect 6087 6400 6121 6434
rect 6155 6400 6189 6434
rect 6223 6400 6257 6434
rect 6291 6400 6325 6434
rect 6359 6400 6393 6434
rect 6427 6400 6461 6434
rect 6495 6400 6529 6434
rect 6563 6400 6597 6434
rect 6631 6400 6665 6434
rect 6699 6400 6733 6434
rect 6767 6400 6801 6434
rect 6835 6400 6869 6434
rect 6903 6400 6937 6434
rect 6971 6400 7005 6434
rect 7039 6400 7073 6434
rect 7107 6400 7141 6434
rect 7175 6400 7209 6434
rect 7243 6400 7277 6434
rect 7311 6400 7345 6434
rect 7379 6400 7413 6434
rect 7447 6400 7481 6434
rect 7515 6400 7549 6434
rect 7583 6400 7617 6434
rect 7651 6400 7685 6434
rect 7719 6400 7753 6434
rect 7787 6400 7821 6434
rect 7855 6400 7889 6434
rect 7923 6400 7957 6434
rect 7991 6400 8025 6434
rect 8059 6400 8093 6434
rect 8127 6400 8161 6434
rect 8195 6400 8229 6434
rect 8263 6400 8297 6434
rect 8331 6400 8365 6434
rect 8399 6400 8433 6434
rect 8467 6400 8501 6434
rect 8535 6400 8569 6434
rect 8603 6400 8637 6434
rect 8671 6400 8705 6434
rect 8739 6400 8773 6434
rect 8807 6400 8841 6434
rect 8875 6400 8909 6434
rect 8943 6400 8977 6434
rect 9011 6400 9045 6434
rect 9079 6400 9113 6434
rect 9147 6400 9181 6434
rect 9215 6400 9249 6434
rect 9283 6400 9317 6434
rect 9351 6400 9385 6434
rect 9419 6400 9453 6434
rect 9487 6400 9521 6434
rect 9555 6400 9589 6434
rect 9623 6400 9657 6434
rect 9691 6400 9725 6434
rect 9759 6400 9793 6434
rect 9827 6400 9861 6434
rect 9895 6400 9929 6434
rect 9963 6400 9997 6434
rect 10031 6400 10065 6434
rect 10099 6400 10133 6434
rect 10167 6400 10201 6434
rect 10235 6400 10269 6434
rect 10303 6400 10337 6434
rect 10371 6400 10405 6434
rect 10439 6400 10473 6434
rect 10507 6400 10541 6434
rect 10575 6400 10609 6434
rect 10643 6400 10677 6434
rect 10711 6400 10745 6434
rect 10779 6400 10813 6434
rect 10847 6400 10881 6434
rect 10915 6400 10949 6434
rect 10983 6400 11017 6434
rect 11051 6400 11085 6434
rect 11119 6400 11153 6434
rect 11187 6400 11221 6434
rect 11255 6400 11289 6434
rect 11323 6400 11357 6434
rect 11391 6400 11425 6434
rect 11459 6400 11493 6434
rect 11527 6400 11561 6434
rect 11595 6400 11629 6434
rect 11663 6400 11697 6434
rect 11731 6400 11765 6434
rect 11799 6400 11833 6434
rect 11867 6400 11901 6434
rect 11935 6400 11969 6434
rect 12003 6400 12037 6434
rect 12071 6400 12105 6434
rect 12139 6400 12173 6434
rect 12207 6400 12241 6434
rect 12275 6400 12309 6434
rect 12343 6400 12377 6434
rect 12411 6400 12445 6434
rect 12479 6400 12513 6434
rect 12547 6400 12581 6434
rect 12615 6400 12649 6434
rect 12683 6400 12717 6434
rect 12751 6400 12785 6434
rect 12819 6400 12853 6434
rect 12887 6400 12921 6434
rect 12955 6400 12989 6434
rect 13023 6400 13057 6434
rect 13091 6400 13125 6434
rect 13159 6400 13193 6434
rect 13227 6400 13261 6434
rect 13295 6400 13329 6434
rect 13363 6400 13397 6434
rect 13431 6400 13465 6434
rect 13499 6400 13533 6434
rect 13567 6400 13601 6434
rect 13635 6400 13669 6434
rect 13703 6400 13737 6434
rect 13771 6400 13805 6434
rect 13839 6400 13873 6434
rect 13907 6400 13941 6434
rect 13975 6400 14009 6434
rect 14043 6400 14077 6434
rect 14111 6400 14145 6434
rect 14179 6400 14213 6434
rect 14247 6400 14281 6434
rect 14315 6400 14349 6434
rect 14383 6400 14417 6434
rect 14451 6400 14485 6434
rect 14519 6400 14553 6434
rect 14587 6400 14621 6434
rect 14655 6400 14689 6434
rect 14723 6400 14757 6434
rect 14791 6400 14825 6434
rect 14859 6400 14893 6434
rect 14932 6401 14966 6435
rect 15000 6401 15034 6435
rect 15068 6401 15102 6435
rect 68 6326 102 6360
rect 137 6326 171 6360
rect 206 6326 240 6360
rect 275 6326 309 6360
rect 344 6326 378 6360
rect 413 6326 447 6360
rect 482 6326 516 6360
rect 551 6326 585 6360
rect 620 6326 654 6360
rect 689 6326 723 6360
rect 758 6326 792 6360
rect 827 6326 861 6360
rect 896 6326 930 6360
rect 965 6326 999 6360
rect 1034 6326 1068 6360
rect 1103 6326 1137 6360
rect 1172 6326 1206 6360
rect 1241 6326 1275 6360
rect 1310 6326 1344 6360
rect 1379 6326 1413 6360
rect 1448 6326 1482 6360
rect 1517 6326 1551 6360
rect 1586 6326 1620 6360
rect 1655 6326 1689 6360
rect 1724 6326 1758 6360
rect 1793 6326 1827 6360
rect 1862 6326 1896 6360
rect 1931 6326 1965 6360
rect 2000 6326 2034 6360
rect 2069 6326 2103 6360
rect 2138 6326 2172 6360
rect 2207 6326 2241 6360
rect 2276 6326 2310 6360
rect 2345 6326 2379 6360
rect 2414 6326 2448 6360
rect 2483 6326 2517 6360
rect 2551 6326 2585 6360
rect 2619 6326 2653 6360
rect 2687 6326 2721 6360
rect 2755 6326 2789 6360
rect 2823 6326 2857 6360
rect 2891 6326 2925 6360
rect 2959 6326 2993 6360
rect 3027 6326 3061 6360
rect 3095 6326 3129 6360
rect 3163 6326 3197 6360
rect 3231 6326 3265 6360
rect 3299 6326 3333 6360
rect 3367 6326 3401 6360
rect 3435 6326 3469 6360
rect 3503 6326 3537 6360
rect 3571 6326 3605 6360
rect 3639 6326 3673 6360
rect 3707 6326 3741 6360
rect 3775 6326 3809 6360
rect 3843 6326 3877 6360
rect 3911 6326 3945 6360
rect 3979 6326 4013 6360
rect 4047 6326 4081 6360
rect 4115 6326 4149 6360
rect 4183 6326 4217 6360
rect 4251 6326 4285 6360
rect 4319 6326 4353 6360
rect 4387 6326 4421 6360
rect 4455 6326 4489 6360
rect 4523 6326 4557 6360
rect 4591 6326 4625 6360
rect 4659 6326 4693 6360
rect 4727 6326 4761 6360
rect 4795 6326 4829 6360
rect 4863 6326 4897 6360
rect 4931 6326 4965 6360
rect 4999 6326 5033 6360
rect 5067 6326 5101 6360
rect 5135 6326 5169 6360
rect 5203 6326 5237 6360
rect 5271 6326 5305 6360
rect 5339 6326 5373 6360
rect 5407 6326 5441 6360
rect 5475 6326 5509 6360
rect 5543 6326 5577 6360
rect 5611 6326 5645 6360
rect 5679 6326 5713 6360
rect 5747 6326 5781 6360
rect 5815 6326 5849 6360
rect 5883 6326 5917 6360
rect 5951 6326 5985 6360
rect 6019 6326 6053 6360
rect 6087 6326 6121 6360
rect 6155 6326 6189 6360
rect 6223 6326 6257 6360
rect 6291 6326 6325 6360
rect 6359 6326 6393 6360
rect 6427 6326 6461 6360
rect 6495 6326 6529 6360
rect 6563 6326 6597 6360
rect 6631 6326 6665 6360
rect 6699 6326 6733 6360
rect 6767 6326 6801 6360
rect 6835 6326 6869 6360
rect 6903 6326 6937 6360
rect 6971 6326 7005 6360
rect 7039 6326 7073 6360
rect 7107 6326 7141 6360
rect 7175 6326 7209 6360
rect 7243 6326 7277 6360
rect 7311 6326 7345 6360
rect 7379 6326 7413 6360
rect 7447 6326 7481 6360
rect 7515 6326 7549 6360
rect 7583 6326 7617 6360
rect 7651 6326 7685 6360
rect 7719 6326 7753 6360
rect 7787 6326 7821 6360
rect 7855 6326 7889 6360
rect 7923 6326 7957 6360
rect 7991 6326 8025 6360
rect 8059 6326 8093 6360
rect 8127 6326 8161 6360
rect 8195 6326 8229 6360
rect 8263 6326 8297 6360
rect 8331 6326 8365 6360
rect 8399 6326 8433 6360
rect 8467 6326 8501 6360
rect 8535 6326 8569 6360
rect 8603 6326 8637 6360
rect 8671 6326 8705 6360
rect 8739 6326 8773 6360
rect 8807 6326 8841 6360
rect 8875 6326 8909 6360
rect 8943 6326 8977 6360
rect 9011 6326 9045 6360
rect 9079 6326 9113 6360
rect 9147 6326 9181 6360
rect 9215 6326 9249 6360
rect 9283 6326 9317 6360
rect 9351 6326 9385 6360
rect 9419 6326 9453 6360
rect 9487 6326 9521 6360
rect 9555 6326 9589 6360
rect 9623 6326 9657 6360
rect 9691 6326 9725 6360
rect 9759 6326 9793 6360
rect 9827 6326 9861 6360
rect 9895 6326 9929 6360
rect 9963 6326 9997 6360
rect 10031 6326 10065 6360
rect 10099 6326 10133 6360
rect 10167 6326 10201 6360
rect 10235 6326 10269 6360
rect 10303 6326 10337 6360
rect 10371 6326 10405 6360
rect 10439 6326 10473 6360
rect 10507 6326 10541 6360
rect 10575 6326 10609 6360
rect 10643 6326 10677 6360
rect 10711 6326 10745 6360
rect 10779 6326 10813 6360
rect 10847 6326 10881 6360
rect 10915 6326 10949 6360
rect 10983 6326 11017 6360
rect 11051 6326 11085 6360
rect 11119 6326 11153 6360
rect 11187 6326 11221 6360
rect 11255 6326 11289 6360
rect 11323 6326 11357 6360
rect 11391 6326 11425 6360
rect 11459 6326 11493 6360
rect 11527 6326 11561 6360
rect 11595 6326 11629 6360
rect 11663 6326 11697 6360
rect 11731 6326 11765 6360
rect 11799 6326 11833 6360
rect 11867 6326 11901 6360
rect 11935 6326 11969 6360
rect 12003 6326 12037 6360
rect 12071 6326 12105 6360
rect 12139 6326 12173 6360
rect 12207 6326 12241 6360
rect 12275 6326 12309 6360
rect 12343 6326 12377 6360
rect 12411 6326 12445 6360
rect 12479 6326 12513 6360
rect 12547 6326 12581 6360
rect 12615 6326 12649 6360
rect 12683 6326 12717 6360
rect 12751 6326 12785 6360
rect 12819 6326 12853 6360
rect 12887 6326 12921 6360
rect 12955 6326 12989 6360
rect 13023 6326 13057 6360
rect 13091 6326 13125 6360
rect 13159 6326 13193 6360
rect 13227 6326 13261 6360
rect 13295 6326 13329 6360
rect 13363 6326 13397 6360
rect 13431 6326 13465 6360
rect 13499 6326 13533 6360
rect 13567 6326 13601 6360
rect 13635 6326 13669 6360
rect 13703 6326 13737 6360
rect 13771 6326 13805 6360
rect 13839 6326 13873 6360
rect 13907 6326 13941 6360
rect 13975 6326 14009 6360
rect 14043 6326 14077 6360
rect 14111 6326 14145 6360
rect 14179 6326 14213 6360
rect 14247 6326 14281 6360
rect 14315 6326 14349 6360
rect 14383 6326 14417 6360
rect 14451 6326 14485 6360
rect 14519 6326 14553 6360
rect 14587 6326 14621 6360
rect 14655 6326 14689 6360
rect 14723 6326 14757 6360
rect 14791 6326 14825 6360
rect 14859 6326 14893 6360
rect 14932 6326 14966 6360
rect 15000 6326 15034 6360
rect 15068 6326 15102 6360
rect 68 6252 102 6286
rect 137 6252 171 6286
rect 206 6252 240 6286
rect 275 6252 309 6286
rect 344 6252 378 6286
rect 413 6252 447 6286
rect 482 6252 516 6286
rect 551 6252 585 6286
rect 620 6252 654 6286
rect 689 6252 723 6286
rect 758 6252 792 6286
rect 827 6252 861 6286
rect 896 6252 930 6286
rect 965 6252 999 6286
rect 1034 6252 1068 6286
rect 1103 6252 1137 6286
rect 1172 6252 1206 6286
rect 1241 6252 1275 6286
rect 1310 6252 1344 6286
rect 1379 6252 1413 6286
rect 1448 6252 1482 6286
rect 1517 6252 1551 6286
rect 1586 6252 1620 6286
rect 1655 6252 1689 6286
rect 1724 6252 1758 6286
rect 1793 6252 1827 6286
rect 1862 6252 1896 6286
rect 1931 6252 1965 6286
rect 2000 6252 2034 6286
rect 2069 6252 2103 6286
rect 2138 6252 2172 6286
rect 2207 6252 2241 6286
rect 2276 6252 2310 6286
rect 2345 6252 2379 6286
rect 2414 6252 2448 6286
rect 2483 6252 2517 6286
rect 2551 6252 2585 6286
rect 2619 6252 2653 6286
rect 2687 6252 2721 6286
rect 2755 6252 2789 6286
rect 2823 6252 2857 6286
rect 2891 6252 2925 6286
rect 2959 6252 2993 6286
rect 3027 6252 3061 6286
rect 3095 6252 3129 6286
rect 3163 6252 3197 6286
rect 3231 6252 3265 6286
rect 3299 6252 3333 6286
rect 3367 6252 3401 6286
rect 3435 6252 3469 6286
rect 3503 6252 3537 6286
rect 3571 6252 3605 6286
rect 3639 6252 3673 6286
rect 3707 6252 3741 6286
rect 3775 6252 3809 6286
rect 3843 6252 3877 6286
rect 3911 6252 3945 6286
rect 3979 6252 4013 6286
rect 4047 6252 4081 6286
rect 4115 6252 4149 6286
rect 4183 6252 4217 6286
rect 4251 6252 4285 6286
rect 4319 6252 4353 6286
rect 4387 6252 4421 6286
rect 4455 6252 4489 6286
rect 4523 6252 4557 6286
rect 4591 6252 4625 6286
rect 4659 6252 4693 6286
rect 4727 6252 4761 6286
rect 4795 6252 4829 6286
rect 4863 6252 4897 6286
rect 4931 6252 4965 6286
rect 4999 6252 5033 6286
rect 5067 6252 5101 6286
rect 5135 6252 5169 6286
rect 5203 6252 5237 6286
rect 5271 6252 5305 6286
rect 5339 6252 5373 6286
rect 5407 6252 5441 6286
rect 5475 6252 5509 6286
rect 5543 6252 5577 6286
rect 5611 6252 5645 6286
rect 5679 6252 5713 6286
rect 5747 6252 5781 6286
rect 5815 6252 5849 6286
rect 5883 6252 5917 6286
rect 5951 6252 5985 6286
rect 6019 6252 6053 6286
rect 6087 6252 6121 6286
rect 6155 6252 6189 6286
rect 6223 6252 6257 6286
rect 6291 6252 6325 6286
rect 6359 6252 6393 6286
rect 6427 6252 6461 6286
rect 6495 6252 6529 6286
rect 6563 6252 6597 6286
rect 6631 6252 6665 6286
rect 6699 6252 6733 6286
rect 6767 6252 6801 6286
rect 6835 6252 6869 6286
rect 6903 6252 6937 6286
rect 6971 6252 7005 6286
rect 7039 6252 7073 6286
rect 7107 6252 7141 6286
rect 7175 6252 7209 6286
rect 7243 6252 7277 6286
rect 7311 6252 7345 6286
rect 7379 6252 7413 6286
rect 7447 6252 7481 6286
rect 7515 6252 7549 6286
rect 7583 6252 7617 6286
rect 7651 6252 7685 6286
rect 7719 6252 7753 6286
rect 7787 6252 7821 6286
rect 7855 6252 7889 6286
rect 7923 6252 7957 6286
rect 7991 6252 8025 6286
rect 8059 6252 8093 6286
rect 8127 6252 8161 6286
rect 8195 6252 8229 6286
rect 8263 6252 8297 6286
rect 8331 6252 8365 6286
rect 8399 6252 8433 6286
rect 8467 6252 8501 6286
rect 8535 6252 8569 6286
rect 8603 6252 8637 6286
rect 8671 6252 8705 6286
rect 8739 6252 8773 6286
rect 8807 6252 8841 6286
rect 8875 6252 8909 6286
rect 8943 6252 8977 6286
rect 9011 6252 9045 6286
rect 9079 6252 9113 6286
rect 9147 6252 9181 6286
rect 9215 6252 9249 6286
rect 9283 6252 9317 6286
rect 9351 6252 9385 6286
rect 9419 6252 9453 6286
rect 9487 6252 9521 6286
rect 9555 6252 9589 6286
rect 9623 6252 9657 6286
rect 9691 6252 9725 6286
rect 9759 6252 9793 6286
rect 9827 6252 9861 6286
rect 9895 6252 9929 6286
rect 9963 6252 9997 6286
rect 10031 6252 10065 6286
rect 10099 6252 10133 6286
rect 10167 6252 10201 6286
rect 10235 6252 10269 6286
rect 10303 6252 10337 6286
rect 10371 6252 10405 6286
rect 10439 6252 10473 6286
rect 10507 6252 10541 6286
rect 10575 6252 10609 6286
rect 10643 6252 10677 6286
rect 10711 6252 10745 6286
rect 10779 6252 10813 6286
rect 10847 6252 10881 6286
rect 10915 6252 10949 6286
rect 10983 6252 11017 6286
rect 11051 6252 11085 6286
rect 11119 6252 11153 6286
rect 11187 6252 11221 6286
rect 11255 6252 11289 6286
rect 11323 6252 11357 6286
rect 11391 6252 11425 6286
rect 11459 6252 11493 6286
rect 11527 6252 11561 6286
rect 11595 6252 11629 6286
rect 11663 6252 11697 6286
rect 11731 6252 11765 6286
rect 11799 6252 11833 6286
rect 11867 6252 11901 6286
rect 11935 6252 11969 6286
rect 12003 6252 12037 6286
rect 12071 6252 12105 6286
rect 12139 6252 12173 6286
rect 12207 6252 12241 6286
rect 12275 6252 12309 6286
rect 12343 6252 12377 6286
rect 12411 6252 12445 6286
rect 12479 6252 12513 6286
rect 12547 6252 12581 6286
rect 12615 6252 12649 6286
rect 12683 6252 12717 6286
rect 12751 6252 12785 6286
rect 12819 6252 12853 6286
rect 12887 6252 12921 6286
rect 12955 6252 12989 6286
rect 13023 6252 13057 6286
rect 13091 6252 13125 6286
rect 13159 6252 13193 6286
rect 13227 6252 13261 6286
rect 13295 6252 13329 6286
rect 13363 6252 13397 6286
rect 13431 6252 13465 6286
rect 13499 6252 13533 6286
rect 13567 6252 13601 6286
rect 13635 6252 13669 6286
rect 13703 6252 13737 6286
rect 13771 6252 13805 6286
rect 13839 6252 13873 6286
rect 13907 6252 13941 6286
rect 13975 6252 14009 6286
rect 14043 6252 14077 6286
rect 14111 6252 14145 6286
rect 14179 6252 14213 6286
rect 14247 6252 14281 6286
rect 14315 6252 14349 6286
rect 14383 6252 14417 6286
rect 14451 6252 14485 6286
rect 14519 6252 14553 6286
rect 14587 6252 14621 6286
rect 14655 6252 14689 6286
rect 14723 6252 14757 6286
rect 14791 6252 14825 6286
rect 14859 6252 14893 6286
rect 14932 6251 14966 6285
rect 15000 6251 15034 6285
rect 15068 6251 15102 6285
rect 68 6178 102 6212
rect 137 6178 171 6212
rect 206 6178 240 6212
rect 275 6178 309 6212
rect 344 6178 378 6212
rect 413 6178 447 6212
rect 482 6178 516 6212
rect 551 6178 585 6212
rect 620 6178 654 6212
rect 689 6178 723 6212
rect 758 6178 792 6212
rect 827 6178 861 6212
rect 896 6178 930 6212
rect 965 6178 999 6212
rect 1034 6178 1068 6212
rect 1103 6178 1137 6212
rect 1172 6178 1206 6212
rect 1241 6178 1275 6212
rect 1310 6178 1344 6212
rect 1379 6178 1413 6212
rect 1448 6178 1482 6212
rect 1517 6178 1551 6212
rect 1586 6178 1620 6212
rect 1655 6178 1689 6212
rect 1724 6178 1758 6212
rect 1793 6178 1827 6212
rect 1862 6178 1896 6212
rect 1931 6178 1965 6212
rect 2000 6178 2034 6212
rect 2069 6178 2103 6212
rect 2138 6178 2172 6212
rect 2207 6178 2241 6212
rect 2276 6178 2310 6212
rect 2345 6178 2379 6212
rect 2414 6178 2448 6212
rect 2483 6178 2517 6212
rect 2551 6178 2585 6212
rect 2619 6178 2653 6212
rect 2687 6178 2721 6212
rect 2755 6178 2789 6212
rect 2823 6178 2857 6212
rect 2891 6178 2925 6212
rect 2959 6178 2993 6212
rect 3027 6178 3061 6212
rect 3095 6178 3129 6212
rect 3163 6178 3197 6212
rect 3231 6178 3265 6212
rect 3299 6178 3333 6212
rect 3367 6178 3401 6212
rect 3435 6178 3469 6212
rect 3503 6178 3537 6212
rect 3571 6178 3605 6212
rect 3639 6178 3673 6212
rect 3707 6178 3741 6212
rect 3775 6178 3809 6212
rect 3843 6178 3877 6212
rect 3911 6178 3945 6212
rect 3979 6178 4013 6212
rect 4047 6178 4081 6212
rect 4115 6178 4149 6212
rect 4183 6178 4217 6212
rect 4251 6178 4285 6212
rect 4319 6178 4353 6212
rect 4387 6178 4421 6212
rect 4455 6178 4489 6212
rect 4523 6178 4557 6212
rect 4591 6178 4625 6212
rect 4659 6178 4693 6212
rect 4727 6178 4761 6212
rect 4795 6178 4829 6212
rect 4863 6178 4897 6212
rect 4931 6178 4965 6212
rect 4999 6178 5033 6212
rect 5067 6178 5101 6212
rect 5135 6178 5169 6212
rect 5203 6178 5237 6212
rect 5271 6178 5305 6212
rect 5339 6178 5373 6212
rect 5407 6178 5441 6212
rect 5475 6178 5509 6212
rect 5543 6178 5577 6212
rect 5611 6178 5645 6212
rect 5679 6178 5713 6212
rect 5747 6178 5781 6212
rect 5815 6178 5849 6212
rect 5883 6178 5917 6212
rect 5951 6178 5985 6212
rect 6019 6178 6053 6212
rect 6087 6178 6121 6212
rect 6155 6178 6189 6212
rect 6223 6178 6257 6212
rect 6291 6178 6325 6212
rect 6359 6178 6393 6212
rect 6427 6178 6461 6212
rect 6495 6178 6529 6212
rect 6563 6178 6597 6212
rect 6631 6178 6665 6212
rect 6699 6178 6733 6212
rect 6767 6178 6801 6212
rect 6835 6178 6869 6212
rect 6903 6178 6937 6212
rect 6971 6178 7005 6212
rect 7039 6178 7073 6212
rect 7107 6178 7141 6212
rect 7175 6178 7209 6212
rect 7243 6178 7277 6212
rect 7311 6178 7345 6212
rect 7379 6178 7413 6212
rect 7447 6178 7481 6212
rect 7515 6178 7549 6212
rect 7583 6178 7617 6212
rect 7651 6178 7685 6212
rect 7719 6178 7753 6212
rect 7787 6178 7821 6212
rect 7855 6178 7889 6212
rect 7923 6178 7957 6212
rect 7991 6178 8025 6212
rect 8059 6178 8093 6212
rect 8127 6178 8161 6212
rect 8195 6178 8229 6212
rect 8263 6178 8297 6212
rect 8331 6178 8365 6212
rect 8399 6178 8433 6212
rect 8467 6178 8501 6212
rect 8535 6178 8569 6212
rect 8603 6178 8637 6212
rect 8671 6178 8705 6212
rect 8739 6178 8773 6212
rect 8807 6178 8841 6212
rect 8875 6178 8909 6212
rect 8943 6178 8977 6212
rect 9011 6178 9045 6212
rect 9079 6178 9113 6212
rect 9147 6178 9181 6212
rect 9215 6178 9249 6212
rect 9283 6178 9317 6212
rect 9351 6178 9385 6212
rect 9419 6178 9453 6212
rect 9487 6178 9521 6212
rect 9555 6178 9589 6212
rect 9623 6178 9657 6212
rect 9691 6178 9725 6212
rect 9759 6178 9793 6212
rect 9827 6178 9861 6212
rect 9895 6178 9929 6212
rect 9963 6178 9997 6212
rect 10031 6178 10065 6212
rect 10099 6178 10133 6212
rect 10167 6178 10201 6212
rect 10235 6178 10269 6212
rect 10303 6178 10337 6212
rect 10371 6178 10405 6212
rect 10439 6178 10473 6212
rect 10507 6178 10541 6212
rect 10575 6178 10609 6212
rect 10643 6178 10677 6212
rect 10711 6178 10745 6212
rect 10779 6178 10813 6212
rect 10847 6178 10881 6212
rect 10915 6178 10949 6212
rect 10983 6178 11017 6212
rect 11051 6178 11085 6212
rect 11119 6178 11153 6212
rect 11187 6178 11221 6212
rect 11255 6178 11289 6212
rect 11323 6178 11357 6212
rect 11391 6178 11425 6212
rect 11459 6178 11493 6212
rect 11527 6178 11561 6212
rect 11595 6178 11629 6212
rect 11663 6178 11697 6212
rect 11731 6178 11765 6212
rect 11799 6178 11833 6212
rect 11867 6178 11901 6212
rect 11935 6178 11969 6212
rect 12003 6178 12037 6212
rect 12071 6178 12105 6212
rect 12139 6178 12173 6212
rect 12207 6178 12241 6212
rect 12275 6178 12309 6212
rect 12343 6178 12377 6212
rect 12411 6178 12445 6212
rect 12479 6178 12513 6212
rect 12547 6178 12581 6212
rect 12615 6178 12649 6212
rect 12683 6178 12717 6212
rect 12751 6178 12785 6212
rect 12819 6178 12853 6212
rect 12887 6178 12921 6212
rect 12955 6178 12989 6212
rect 13023 6178 13057 6212
rect 13091 6178 13125 6212
rect 13159 6178 13193 6212
rect 13227 6178 13261 6212
rect 13295 6178 13329 6212
rect 13363 6178 13397 6212
rect 13431 6178 13465 6212
rect 13499 6178 13533 6212
rect 13567 6178 13601 6212
rect 13635 6178 13669 6212
rect 13703 6178 13737 6212
rect 13771 6178 13805 6212
rect 13839 6178 13873 6212
rect 13907 6178 13941 6212
rect 13975 6178 14009 6212
rect 14043 6178 14077 6212
rect 14111 6178 14145 6212
rect 14179 6178 14213 6212
rect 14247 6178 14281 6212
rect 14315 6178 14349 6212
rect 14383 6178 14417 6212
rect 14451 6178 14485 6212
rect 14519 6178 14553 6212
rect 14587 6178 14621 6212
rect 14655 6178 14689 6212
rect 14723 6178 14757 6212
rect 14791 6178 14825 6212
rect 14859 6178 14893 6212
rect 14932 6176 14966 6210
rect 15000 6176 15034 6210
rect 15068 6176 15102 6210
rect 68 6104 102 6138
rect 137 6104 171 6138
rect 206 6104 240 6138
rect 275 6104 309 6138
rect 344 6104 378 6138
rect 413 6104 447 6138
rect 482 6104 516 6138
rect 551 6104 585 6138
rect 620 6104 654 6138
rect 689 6104 723 6138
rect 758 6104 792 6138
rect 827 6104 861 6138
rect 896 6104 930 6138
rect 965 6104 999 6138
rect 1034 6104 1068 6138
rect 1103 6104 1137 6138
rect 1172 6104 1206 6138
rect 1241 6104 1275 6138
rect 1310 6104 1344 6138
rect 1379 6104 1413 6138
rect 1448 6104 1482 6138
rect 1517 6104 1551 6138
rect 1586 6104 1620 6138
rect 1655 6104 1689 6138
rect 1724 6104 1758 6138
rect 1793 6104 1827 6138
rect 1862 6104 1896 6138
rect 1931 6104 1965 6138
rect 2000 6104 2034 6138
rect 2069 6104 2103 6138
rect 2138 6104 2172 6138
rect 2207 6104 2241 6138
rect 2276 6104 2310 6138
rect 2345 6104 2379 6138
rect 2414 6104 2448 6138
rect 2483 6104 2517 6138
rect 2551 6104 2585 6138
rect 2619 6104 2653 6138
rect 2687 6104 2721 6138
rect 2755 6104 2789 6138
rect 2823 6104 2857 6138
rect 2891 6104 2925 6138
rect 2959 6104 2993 6138
rect 3027 6104 3061 6138
rect 3095 6104 3129 6138
rect 3163 6104 3197 6138
rect 3231 6104 3265 6138
rect 3299 6104 3333 6138
rect 3367 6104 3401 6138
rect 3435 6104 3469 6138
rect 3503 6104 3537 6138
rect 3571 6104 3605 6138
rect 3639 6104 3673 6138
rect 3707 6104 3741 6138
rect 3775 6104 3809 6138
rect 3843 6104 3877 6138
rect 3911 6104 3945 6138
rect 3979 6104 4013 6138
rect 4047 6104 4081 6138
rect 4115 6104 4149 6138
rect 4183 6104 4217 6138
rect 4251 6104 4285 6138
rect 4319 6104 4353 6138
rect 4387 6104 4421 6138
rect 4455 6104 4489 6138
rect 4523 6104 4557 6138
rect 4591 6104 4625 6138
rect 4659 6104 4693 6138
rect 4727 6104 4761 6138
rect 4795 6104 4829 6138
rect 4863 6104 4897 6138
rect 4931 6104 4965 6138
rect 4999 6104 5033 6138
rect 5067 6104 5101 6138
rect 5135 6104 5169 6138
rect 5203 6104 5237 6138
rect 5271 6104 5305 6138
rect 5339 6104 5373 6138
rect 5407 6104 5441 6138
rect 5475 6104 5509 6138
rect 5543 6104 5577 6138
rect 5611 6104 5645 6138
rect 5679 6104 5713 6138
rect 5747 6104 5781 6138
rect 5815 6104 5849 6138
rect 5883 6104 5917 6138
rect 5951 6104 5985 6138
rect 6019 6104 6053 6138
rect 6087 6104 6121 6138
rect 6155 6104 6189 6138
rect 6223 6104 6257 6138
rect 6291 6104 6325 6138
rect 6359 6104 6393 6138
rect 6427 6104 6461 6138
rect 6495 6104 6529 6138
rect 6563 6104 6597 6138
rect 6631 6104 6665 6138
rect 6699 6104 6733 6138
rect 6767 6104 6801 6138
rect 6835 6104 6869 6138
rect 6903 6104 6937 6138
rect 6971 6104 7005 6138
rect 7039 6104 7073 6138
rect 7107 6104 7141 6138
rect 7175 6104 7209 6138
rect 7243 6104 7277 6138
rect 7311 6104 7345 6138
rect 7379 6104 7413 6138
rect 7447 6104 7481 6138
rect 7515 6104 7549 6138
rect 7583 6104 7617 6138
rect 7651 6104 7685 6138
rect 7719 6104 7753 6138
rect 7787 6104 7821 6138
rect 7855 6104 7889 6138
rect 7923 6104 7957 6138
rect 7991 6104 8025 6138
rect 8059 6104 8093 6138
rect 8127 6104 8161 6138
rect 8195 6104 8229 6138
rect 8263 6104 8297 6138
rect 8331 6104 8365 6138
rect 8399 6104 8433 6138
rect 8467 6104 8501 6138
rect 8535 6104 8569 6138
rect 8603 6104 8637 6138
rect 8671 6104 8705 6138
rect 8739 6104 8773 6138
rect 8807 6104 8841 6138
rect 8875 6104 8909 6138
rect 8943 6104 8977 6138
rect 9011 6104 9045 6138
rect 9079 6104 9113 6138
rect 9147 6104 9181 6138
rect 9215 6104 9249 6138
rect 9283 6104 9317 6138
rect 9351 6104 9385 6138
rect 9419 6104 9453 6138
rect 9487 6104 9521 6138
rect 9555 6104 9589 6138
rect 9623 6104 9657 6138
rect 9691 6104 9725 6138
rect 9759 6104 9793 6138
rect 9827 6104 9861 6138
rect 9895 6104 9929 6138
rect 9963 6104 9997 6138
rect 10031 6104 10065 6138
rect 10099 6104 10133 6138
rect 10167 6104 10201 6138
rect 10235 6104 10269 6138
rect 10303 6104 10337 6138
rect 10371 6104 10405 6138
rect 10439 6104 10473 6138
rect 10507 6104 10541 6138
rect 10575 6104 10609 6138
rect 10643 6104 10677 6138
rect 10711 6104 10745 6138
rect 10779 6104 10813 6138
rect 10847 6104 10881 6138
rect 10915 6104 10949 6138
rect 10983 6104 11017 6138
rect 11051 6104 11085 6138
rect 11119 6104 11153 6138
rect 11187 6104 11221 6138
rect 11255 6104 11289 6138
rect 11323 6104 11357 6138
rect 11391 6104 11425 6138
rect 11459 6104 11493 6138
rect 11527 6104 11561 6138
rect 11595 6104 11629 6138
rect 11663 6104 11697 6138
rect 11731 6104 11765 6138
rect 11799 6104 11833 6138
rect 11867 6104 11901 6138
rect 11935 6104 11969 6138
rect 12003 6104 12037 6138
rect 12071 6104 12105 6138
rect 12139 6104 12173 6138
rect 12207 6104 12241 6138
rect 12275 6104 12309 6138
rect 12343 6104 12377 6138
rect 12411 6104 12445 6138
rect 12479 6104 12513 6138
rect 12547 6104 12581 6138
rect 12615 6104 12649 6138
rect 12683 6104 12717 6138
rect 12751 6104 12785 6138
rect 12819 6104 12853 6138
rect 12887 6104 12921 6138
rect 12955 6104 12989 6138
rect 13023 6104 13057 6138
rect 13091 6104 13125 6138
rect 13159 6104 13193 6138
rect 13227 6104 13261 6138
rect 13295 6104 13329 6138
rect 13363 6104 13397 6138
rect 13431 6104 13465 6138
rect 13499 6104 13533 6138
rect 13567 6104 13601 6138
rect 13635 6104 13669 6138
rect 13703 6104 13737 6138
rect 13771 6104 13805 6138
rect 13839 6104 13873 6138
rect 13907 6104 13941 6138
rect 13975 6104 14009 6138
rect 14043 6104 14077 6138
rect 14111 6104 14145 6138
rect 14179 6104 14213 6138
rect 14247 6104 14281 6138
rect 14315 6104 14349 6138
rect 14383 6104 14417 6138
rect 14451 6104 14485 6138
rect 14519 6104 14553 6138
rect 14587 6104 14621 6138
rect 14655 6104 14689 6138
rect 14723 6104 14757 6138
rect 14791 6104 14825 6138
rect 14859 6104 14893 6138
rect 14932 6101 14966 6135
rect 15000 6101 15034 6135
rect 15068 6101 15102 6135
rect 14932 6026 14966 6060
rect 15000 6026 15034 6060
rect 15068 6026 15102 6060
rect 15000 4628 15102 5954
rect 15000 4559 15034 4593
rect 15068 4559 15102 4593
rect 15000 4490 15034 4524
rect 15068 4490 15102 4524
rect 15000 4421 15034 4455
rect 15068 4421 15102 4455
rect 15000 4352 15034 4386
rect 15068 4352 15102 4386
rect 15000 4283 15034 4317
rect 15068 4283 15102 4317
rect 15000 4214 15034 4248
rect 15068 4214 15102 4248
rect 15000 4145 15034 4179
rect 15068 4145 15102 4179
rect 15000 4076 15034 4110
rect 15068 4076 15102 4110
rect 15000 4007 15034 4041
rect 15068 4007 15102 4041
rect 15000 3938 15034 3972
rect 15068 3938 15102 3972
rect 15000 3869 15034 3903
rect 15068 3869 15102 3903
rect 15000 3800 15034 3834
rect 15068 3800 15102 3834
rect 15000 3731 15034 3765
rect 15068 3731 15102 3765
rect 15000 3662 15034 3696
rect 15068 3662 15102 3696
rect 15000 3593 15034 3627
rect 15068 3593 15102 3627
rect 15000 3524 15034 3558
rect 15068 3524 15102 3558
rect 15000 3455 15034 3489
rect 15068 3455 15102 3489
rect 15000 3386 15034 3420
rect 15068 3386 15102 3420
rect 15000 3317 15034 3351
rect 15068 3317 15102 3351
rect 15000 3248 15034 3282
rect 15068 3248 15102 3282
rect 15000 3179 15034 3213
rect 15068 3179 15102 3213
rect 15000 3110 15034 3144
rect 15068 3110 15102 3144
rect 15000 3041 15034 3075
rect 15068 3041 15102 3075
rect 15000 2972 15034 3006
rect 15068 2972 15102 3006
rect 15000 2903 15034 2937
rect 15068 2903 15102 2937
rect 15000 2834 15034 2868
rect 15068 2834 15102 2868
rect 15000 2765 15034 2799
rect 15068 2765 15102 2799
rect 15000 2696 15034 2730
rect 15068 2696 15102 2730
rect 15000 2627 15034 2661
rect 15068 2627 15102 2661
rect 15000 2558 15034 2592
rect 15068 2558 15102 2592
rect 15000 2489 15034 2523
rect 15068 2489 15102 2523
rect 15000 2420 15034 2454
rect 15068 2420 15102 2454
rect 15000 2351 15034 2385
rect 15068 2351 15102 2385
rect 15000 2282 15034 2316
rect 15068 2282 15102 2316
rect 15000 2213 15034 2247
rect 15068 2213 15102 2247
rect 15000 2144 15034 2178
rect 15068 2144 15102 2178
rect 15000 2075 15034 2109
rect 15068 2075 15102 2109
rect 15000 2006 15034 2040
rect 15068 2006 15102 2040
rect 15000 1937 15034 1971
rect 15068 1937 15102 1971
rect 15000 1868 15034 1902
rect 15068 1868 15102 1902
rect 15000 1799 15034 1833
rect 15068 1799 15102 1833
rect 15000 1730 15034 1764
rect 15068 1730 15102 1764
rect 15000 1661 15034 1695
rect 15068 1661 15102 1695
rect 15000 1592 15034 1626
rect 15068 1592 15102 1626
rect 15000 1523 15034 1557
rect 15068 1523 15102 1557
rect 15000 1454 15034 1488
rect 15068 1454 15102 1488
rect 15000 1385 15034 1419
rect 15068 1385 15102 1419
rect 15000 1316 15034 1350
rect 15068 1316 15102 1350
rect 3577 1217 3611 1251
rect 3645 1217 3679 1251
rect 3713 1217 3747 1251
rect 3781 1217 3815 1251
rect 3849 1217 3883 1251
rect 3917 1217 3951 1251
rect 3985 1217 4019 1251
rect 4053 1217 4087 1251
rect 4121 1217 4155 1251
rect 4189 1217 4223 1251
rect 4257 1217 4291 1251
rect 4325 1217 4359 1251
rect 4393 1217 4427 1251
rect 4461 1217 4495 1251
rect 4529 1217 4563 1251
rect 4597 1217 4631 1251
rect 4665 1217 4699 1251
rect 4733 1217 4767 1251
rect 4801 1217 4835 1251
rect 4869 1217 4903 1251
rect 4937 1217 4971 1251
rect 5005 1217 5039 1251
rect 5073 1217 5107 1251
rect 5141 1217 5175 1251
rect 5209 1217 5243 1251
rect 5277 1217 5311 1251
rect 5345 1217 5379 1251
rect 5413 1217 5447 1251
rect 5481 1217 5515 1251
rect 5549 1217 5583 1251
rect 5617 1217 5651 1251
rect 5685 1217 5719 1251
rect 5753 1217 5787 1251
rect 5821 1217 5855 1251
rect 5889 1217 5923 1251
rect 5957 1217 5991 1251
rect 6025 1217 6059 1251
rect 6093 1217 6127 1251
rect 6161 1217 6195 1251
rect 6229 1217 6263 1251
rect 6297 1217 6331 1251
rect 6365 1217 6399 1251
rect 6433 1217 6467 1251
rect 6501 1217 6535 1251
rect 6569 1217 6603 1251
rect 6637 1217 6671 1251
rect 6705 1217 6739 1251
rect 6773 1217 6807 1251
rect 6841 1217 6875 1251
rect 6909 1217 6943 1251
rect 6988 1193 7022 1227
rect 7068 1223 7102 1257
rect 7137 1223 7171 1257
rect 7206 1223 7240 1257
rect 7275 1223 7309 1257
rect 7344 1223 7378 1257
rect 7413 1223 7447 1257
rect 7482 1223 7516 1257
rect 7551 1223 7585 1257
rect 7620 1223 7654 1257
rect 7689 1223 7723 1257
rect 7758 1223 7792 1257
rect 7827 1223 7861 1257
rect 7896 1223 7930 1257
rect 7965 1223 7999 1257
rect 8034 1223 8068 1257
rect 8103 1223 8137 1257
rect 8172 1223 8206 1257
rect 8241 1223 8275 1257
rect 8310 1223 8344 1257
rect 8379 1223 8413 1257
rect 8448 1223 8482 1257
rect 8517 1223 8551 1257
rect 8586 1223 8620 1257
rect 8655 1223 8689 1257
rect 8724 1223 8758 1257
rect 8793 1223 8827 1257
rect 8862 1223 8896 1257
rect 8931 1223 8965 1257
rect 9000 1223 9034 1257
rect 9069 1223 9103 1257
rect 9138 1223 9172 1257
rect 9207 1223 9241 1257
rect 9276 1223 9310 1257
rect 9345 1223 9379 1257
rect 9414 1223 9448 1257
rect 9483 1223 9517 1257
rect 9552 1223 9586 1257
rect 9621 1223 9655 1257
rect 9690 1223 9724 1257
rect 6988 1125 7022 1159
rect 7068 1155 7102 1189
rect 7137 1155 7171 1189
rect 7206 1155 7240 1189
rect 7275 1155 7309 1189
rect 7344 1155 7378 1189
rect 7413 1155 7447 1189
rect 7482 1155 7516 1189
rect 7551 1155 7585 1189
rect 7620 1155 7654 1189
rect 7689 1155 7723 1189
rect 7758 1155 7792 1189
rect 7827 1155 7861 1189
rect 7896 1155 7930 1189
rect 7965 1155 7999 1189
rect 8034 1155 8068 1189
rect 8103 1155 8137 1189
rect 8172 1155 8206 1189
rect 8241 1155 8275 1189
rect 8310 1155 8344 1189
rect 8379 1155 8413 1189
rect 8448 1155 8482 1189
rect 8517 1155 8551 1189
rect 8586 1155 8620 1189
rect 8655 1155 8689 1189
rect 8724 1155 8758 1189
rect 8793 1155 8827 1189
rect 8862 1155 8896 1189
rect 8931 1155 8965 1189
rect 9000 1155 9034 1189
rect 9069 1155 9103 1189
rect 9138 1155 9172 1189
rect 9207 1155 9241 1189
rect 9276 1155 9310 1189
rect 9345 1155 9379 1189
rect 9414 1155 9448 1189
rect 9483 1155 9517 1189
rect 9552 1155 9586 1189
rect 9621 1155 9655 1189
rect 9690 1155 9724 1189
rect 6988 1057 7022 1091
rect 7068 1087 7102 1121
rect 7137 1087 7171 1121
rect 7206 1087 7240 1121
rect 7275 1087 7309 1121
rect 7344 1087 7378 1121
rect 7413 1087 7447 1121
rect 7482 1087 7516 1121
rect 7551 1087 7585 1121
rect 7620 1087 7654 1121
rect 7689 1087 7723 1121
rect 7758 1087 7792 1121
rect 7827 1087 7861 1121
rect 7896 1087 7930 1121
rect 7965 1087 7999 1121
rect 8034 1087 8068 1121
rect 8103 1087 8137 1121
rect 8172 1087 8206 1121
rect 8241 1087 8275 1121
rect 8310 1087 8344 1121
rect 8379 1087 8413 1121
rect 8448 1087 8482 1121
rect 8517 1087 8551 1121
rect 8586 1087 8620 1121
rect 8655 1087 8689 1121
rect 8724 1087 8758 1121
rect 8793 1087 8827 1121
rect 8862 1087 8896 1121
rect 8931 1087 8965 1121
rect 9000 1087 9034 1121
rect 9069 1087 9103 1121
rect 9138 1087 9172 1121
rect 9207 1087 9241 1121
rect 9276 1087 9310 1121
rect 9345 1087 9379 1121
rect 9414 1087 9448 1121
rect 9483 1087 9517 1121
rect 9552 1087 9586 1121
rect 9621 1087 9655 1121
rect 9690 1087 9724 1121
rect 6988 989 7022 1023
rect 7068 1019 7102 1053
rect 7137 1019 7171 1053
rect 7206 1019 7240 1053
rect 7275 1019 7309 1053
rect 7344 1019 7378 1053
rect 7413 1019 7447 1053
rect 7482 1019 7516 1053
rect 7551 1019 7585 1053
rect 7620 1019 7654 1053
rect 7689 1019 7723 1053
rect 7758 1019 7792 1053
rect 7827 1019 7861 1053
rect 7896 1019 7930 1053
rect 7965 1019 7999 1053
rect 8034 1019 8068 1053
rect 8103 1019 8137 1053
rect 8172 1019 8206 1053
rect 8241 1019 8275 1053
rect 8310 1019 8344 1053
rect 8379 1019 8413 1053
rect 8448 1019 8482 1053
rect 8517 1019 8551 1053
rect 8586 1019 8620 1053
rect 8655 1019 8689 1053
rect 8724 1019 8758 1053
rect 8793 1019 8827 1053
rect 8862 1019 8896 1053
rect 8931 1019 8965 1053
rect 9000 1019 9034 1053
rect 9069 1019 9103 1053
rect 9138 1019 9172 1053
rect 9207 1019 9241 1053
rect 9276 1019 9310 1053
rect 9345 1019 9379 1053
rect 9414 1019 9448 1053
rect 9483 1019 9517 1053
rect 9552 1019 9586 1053
rect 9621 1019 9655 1053
rect 9690 1019 9724 1053
rect 9759 1019 14893 1257
rect 14932 1210 14966 1244
rect 15000 1210 15034 1244
rect 15068 1210 15102 1244
rect 14932 1138 14966 1172
rect 15000 1138 15034 1172
rect 15068 1138 15102 1172
rect 14932 1066 14966 1100
rect 15000 1066 15034 1100
rect 15068 1066 15102 1100
rect 14932 994 14966 1028
rect 15000 994 15034 1028
rect 15068 994 15102 1028
rect 6988 921 7022 955
rect 7067 913 7101 947
rect 7137 913 7171 947
rect 7207 913 7241 947
rect 7277 913 7311 947
rect 7347 913 7381 947
rect 7417 913 7451 947
rect 7487 913 7521 947
rect 7557 913 7591 947
rect 7627 913 7661 947
rect 7696 913 7730 947
rect 6988 853 7022 887
rect 7067 841 7101 875
rect 7137 841 7171 875
rect 7207 841 7241 875
rect 7277 841 7311 875
rect 7347 841 7381 875
rect 7417 841 7451 875
rect 7487 841 7521 875
rect 7557 841 7591 875
rect 7627 841 7661 875
rect 7696 841 7730 875
rect 6988 785 7022 819
rect 7067 769 7101 803
rect 7137 769 7171 803
rect 7207 769 7241 803
rect 7277 769 7311 803
rect 7347 769 7381 803
rect 7417 769 7451 803
rect 7487 769 7521 803
rect 7557 769 7591 803
rect 7627 769 7661 803
rect 7696 769 7730 803
rect 6988 717 7022 751
rect 7067 697 7101 731
rect 7137 697 7171 731
rect 7207 697 7241 731
rect 7277 697 7311 731
rect 7347 697 7381 731
rect 7417 697 7451 731
rect 7487 697 7521 731
rect 7557 697 7591 731
rect 7627 697 7661 731
rect 7696 697 7730 731
rect 6988 649 7022 683
rect 7067 625 7101 659
rect 7137 625 7171 659
rect 7207 625 7241 659
rect 7277 625 7311 659
rect 7347 625 7381 659
rect 7417 625 7451 659
rect 7487 625 7521 659
rect 7557 625 7591 659
rect 7627 625 7661 659
rect 7696 625 7730 659
rect 6988 581 7022 615
rect 7067 553 7101 587
rect 7137 553 7171 587
rect 7207 553 7241 587
rect 7277 553 7311 587
rect 7347 553 7381 587
rect 7417 553 7451 587
rect 7487 553 7521 587
rect 7557 553 7591 587
rect 7627 553 7661 587
rect 7696 553 7730 587
rect 6988 513 7022 547
rect 7067 481 7101 515
rect 7137 481 7171 515
rect 7207 481 7241 515
rect 7277 481 7311 515
rect 7347 481 7381 515
rect 7417 481 7451 515
rect 7487 481 7521 515
rect 7557 481 7591 515
rect 7627 481 7661 515
rect 7696 481 7730 515
rect 6988 445 7022 479
rect 6988 377 7022 411
rect 7067 409 7101 443
rect 7137 409 7171 443
rect 7207 409 7241 443
rect 7277 409 7311 443
rect 7347 409 7381 443
rect 7417 409 7451 443
rect 7487 409 7521 443
rect 7557 409 7591 443
rect 7627 409 7661 443
rect 7696 409 7730 443
rect 9711 913 9745 947
rect 9781 913 9815 947
rect 9851 913 9885 947
rect 9921 913 9955 947
rect 9991 913 10025 947
rect 10061 913 10095 947
rect 10131 913 10165 947
rect 10201 913 10235 947
rect 10271 913 10305 947
rect 10341 913 10375 947
rect 10411 913 10445 947
rect 10481 913 10515 947
rect 10551 913 10585 947
rect 10621 913 10655 947
rect 10691 913 10725 947
rect 10761 913 10795 947
rect 10831 913 10865 947
rect 10901 913 10935 947
rect 10971 913 11005 947
rect 11041 913 11075 947
rect 11111 913 11145 947
rect 11181 913 11215 947
rect 11251 913 11285 947
rect 11321 913 11355 947
rect 11391 913 11425 947
rect 11460 913 11494 947
rect 11529 913 11563 947
rect 11598 913 11632 947
rect 11680 921 11714 955
rect 11750 921 11784 955
rect 11820 921 11854 955
rect 11890 921 11924 955
rect 11960 921 11994 955
rect 12030 921 12064 955
rect 12099 921 12133 955
rect 12168 921 12202 955
rect 12237 921 12271 955
rect 12306 921 12340 955
rect 12375 921 12409 955
rect 12444 921 12478 955
rect 12513 921 12547 955
rect 12582 921 12616 955
rect 12651 921 12685 955
rect 12720 921 12754 955
rect 12789 921 12823 955
rect 12858 921 12892 955
rect 12927 921 12961 955
rect 12996 921 13030 955
rect 13065 921 13099 955
rect 13134 921 13168 955
rect 13203 921 13237 955
rect 13272 921 13306 955
rect 13341 921 13375 955
rect 13410 921 13444 955
rect 13479 921 13513 955
rect 13548 921 13582 955
rect 13617 921 13651 955
rect 13686 921 13720 955
rect 13755 921 13789 955
rect 13824 921 13858 955
rect 13893 921 13927 955
rect 13962 921 13996 955
rect 14031 921 14065 955
rect 14100 921 14134 955
rect 14169 921 14203 955
rect 14238 921 14272 955
rect 14307 921 14341 955
rect 14376 921 14410 955
rect 14445 921 14479 955
rect 14514 921 14548 955
rect 14583 921 14617 955
rect 14652 921 14686 955
rect 14721 921 14755 955
rect 14790 921 14824 955
rect 14859 921 14893 955
rect 14932 922 14966 956
rect 15000 922 15034 956
rect 15068 922 15102 956
rect 9711 841 9745 875
rect 9781 841 9815 875
rect 9851 841 9885 875
rect 9921 841 9955 875
rect 9991 841 10025 875
rect 10061 841 10095 875
rect 10131 841 10165 875
rect 10201 841 10235 875
rect 10271 841 10305 875
rect 10341 841 10375 875
rect 10411 841 10445 875
rect 10481 841 10515 875
rect 10551 841 10585 875
rect 10621 841 10655 875
rect 10691 841 10725 875
rect 10761 841 10795 875
rect 10831 841 10865 875
rect 10901 841 10935 875
rect 10971 841 11005 875
rect 11041 841 11075 875
rect 11111 841 11145 875
rect 11181 841 11215 875
rect 11251 841 11285 875
rect 11321 841 11355 875
rect 11391 841 11425 875
rect 11460 841 11494 875
rect 11529 841 11563 875
rect 11598 841 11632 875
rect 11680 841 11714 875
rect 11750 841 11784 875
rect 11820 841 11854 875
rect 11890 841 11924 875
rect 11960 841 11994 875
rect 12030 841 12064 875
rect 12099 841 12133 875
rect 12168 841 12202 875
rect 12237 841 12271 875
rect 12306 841 12340 875
rect 12375 841 12409 875
rect 12444 841 12478 875
rect 12513 841 12547 875
rect 12582 841 12616 875
rect 12651 841 12685 875
rect 12720 841 12754 875
rect 12789 841 12823 875
rect 12858 841 12892 875
rect 12927 841 12961 875
rect 12996 841 13030 875
rect 13065 841 13099 875
rect 13134 841 13168 875
rect 13203 841 13237 875
rect 13272 841 13306 875
rect 13341 841 13375 875
rect 13410 841 13444 875
rect 13479 841 13513 875
rect 13548 841 13582 875
rect 13617 841 13651 875
rect 13686 841 13720 875
rect 13755 841 13789 875
rect 13824 841 13858 875
rect 13893 841 13927 875
rect 13962 841 13996 875
rect 14031 841 14065 875
rect 14100 841 14134 875
rect 14169 841 14203 875
rect 14238 841 14272 875
rect 14307 841 14341 875
rect 14376 841 14410 875
rect 14445 841 14479 875
rect 14514 841 14548 875
rect 14583 841 14617 875
rect 14652 841 14686 875
rect 14721 841 14755 875
rect 14790 841 14824 875
rect 14859 841 14893 875
rect 14932 850 14966 884
rect 15000 850 15034 884
rect 15068 850 15102 884
rect 9711 769 9745 803
rect 9781 769 9815 803
rect 9851 769 9885 803
rect 9921 769 9955 803
rect 9991 769 10025 803
rect 10061 769 10095 803
rect 10131 769 10165 803
rect 10201 769 10235 803
rect 10271 769 10305 803
rect 10341 769 10375 803
rect 10411 769 10445 803
rect 10481 769 10515 803
rect 10551 769 10585 803
rect 10621 769 10655 803
rect 10691 769 10725 803
rect 10761 769 10795 803
rect 10831 769 10865 803
rect 10901 769 10935 803
rect 10971 769 11005 803
rect 11041 769 11075 803
rect 11111 769 11145 803
rect 11181 769 11215 803
rect 11251 769 11285 803
rect 11321 769 11355 803
rect 11391 769 11425 803
rect 11460 769 11494 803
rect 11529 769 11563 803
rect 11598 769 11632 803
rect 11680 761 11714 795
rect 11750 761 11784 795
rect 11820 761 11854 795
rect 11890 761 11924 795
rect 11960 761 11994 795
rect 12030 761 12064 795
rect 12099 761 12133 795
rect 12168 761 12202 795
rect 12237 761 12271 795
rect 12306 761 12340 795
rect 12375 761 12409 795
rect 12444 761 12478 795
rect 12513 761 12547 795
rect 12582 761 12616 795
rect 12651 761 12685 795
rect 12720 761 12754 795
rect 12789 761 12823 795
rect 12858 761 12892 795
rect 12927 761 12961 795
rect 12996 761 13030 795
rect 13065 761 13099 795
rect 13134 761 13168 795
rect 13203 761 13237 795
rect 13272 761 13306 795
rect 13341 761 13375 795
rect 13410 761 13444 795
rect 13479 761 13513 795
rect 13548 761 13582 795
rect 13617 761 13651 795
rect 13686 761 13720 795
rect 13755 761 13789 795
rect 13824 761 13858 795
rect 13893 761 13927 795
rect 13962 761 13996 795
rect 14031 761 14065 795
rect 14100 761 14134 795
rect 14169 761 14203 795
rect 14238 761 14272 795
rect 14307 761 14341 795
rect 14376 761 14410 795
rect 14445 761 14479 795
rect 14514 761 14548 795
rect 14583 761 14617 795
rect 14652 761 14686 795
rect 14721 761 14755 795
rect 14790 761 14824 795
rect 14859 761 14893 795
rect 14932 778 14966 812
rect 15000 778 15034 812
rect 15068 778 15102 812
rect 9711 697 9745 731
rect 9781 697 9815 731
rect 9851 697 9885 731
rect 9921 697 9955 731
rect 9991 697 10025 731
rect 10061 697 10095 731
rect 10131 697 10165 731
rect 10201 697 10235 731
rect 10271 697 10305 731
rect 10341 697 10375 731
rect 10411 697 10445 731
rect 10481 697 10515 731
rect 10551 697 10585 731
rect 10621 697 10655 731
rect 10691 697 10725 731
rect 10761 697 10795 731
rect 10831 697 10865 731
rect 10901 697 10935 731
rect 10971 697 11005 731
rect 11041 697 11075 731
rect 11111 697 11145 731
rect 11181 697 11215 731
rect 11251 697 11285 731
rect 11321 697 11355 731
rect 11391 697 11425 731
rect 11460 697 11494 731
rect 11529 697 11563 731
rect 11598 697 11632 731
rect 9711 625 9745 659
rect 9781 625 9815 659
rect 9851 625 9885 659
rect 9921 625 9955 659
rect 9991 625 10025 659
rect 10061 625 10095 659
rect 10131 625 10165 659
rect 10201 625 10235 659
rect 10271 625 10305 659
rect 10341 625 10375 659
rect 10411 625 10445 659
rect 10481 625 10515 659
rect 10551 625 10585 659
rect 10621 625 10655 659
rect 10691 625 10725 659
rect 10761 625 10795 659
rect 10831 625 10865 659
rect 10901 625 10935 659
rect 10971 625 11005 659
rect 11041 625 11075 659
rect 11111 625 11145 659
rect 11181 625 11215 659
rect 11251 625 11285 659
rect 11321 625 11355 659
rect 11391 625 11425 659
rect 11460 625 11494 659
rect 11529 625 11563 659
rect 11598 625 11632 659
rect 9711 553 9745 587
rect 9781 553 9815 587
rect 9851 553 9885 587
rect 9921 553 9955 587
rect 9991 553 10025 587
rect 10061 553 10095 587
rect 10131 553 10165 587
rect 10201 553 10235 587
rect 10271 553 10305 587
rect 10341 553 10375 587
rect 10411 553 10445 587
rect 10481 553 10515 587
rect 10551 553 10585 587
rect 10621 553 10655 587
rect 10691 553 10725 587
rect 10761 553 10795 587
rect 10831 553 10865 587
rect 10901 553 10935 587
rect 10971 553 11005 587
rect 11041 553 11075 587
rect 11111 553 11145 587
rect 11181 553 11215 587
rect 11251 553 11285 587
rect 11321 553 11355 587
rect 11391 553 11425 587
rect 11460 553 11494 587
rect 11529 553 11563 587
rect 11598 553 11632 587
rect 9711 481 9745 515
rect 9781 481 9815 515
rect 9851 481 9885 515
rect 9921 481 9955 515
rect 9991 481 10025 515
rect 10061 481 10095 515
rect 10131 481 10165 515
rect 10201 481 10235 515
rect 10271 481 10305 515
rect 10341 481 10375 515
rect 10411 481 10445 515
rect 10481 481 10515 515
rect 10551 481 10585 515
rect 10621 481 10655 515
rect 10691 481 10725 515
rect 10761 481 10795 515
rect 10831 481 10865 515
rect 10901 481 10935 515
rect 10971 481 11005 515
rect 11041 481 11075 515
rect 11111 481 11145 515
rect 11181 481 11215 515
rect 11251 481 11285 515
rect 11321 481 11355 515
rect 11391 481 11425 515
rect 11460 481 11494 515
rect 11529 481 11563 515
rect 11598 481 11632 515
rect 9711 409 9745 443
rect 9781 409 9815 443
rect 9851 409 9885 443
rect 9921 409 9955 443
rect 9991 409 10025 443
rect 10061 409 10095 443
rect 10131 409 10165 443
rect 10201 409 10235 443
rect 10271 409 10305 443
rect 10341 409 10375 443
rect 10411 409 10445 443
rect 10481 409 10515 443
rect 10551 409 10585 443
rect 10621 409 10655 443
rect 10691 409 10725 443
rect 10761 409 10795 443
rect 10831 409 10865 443
rect 10901 409 10935 443
rect 10971 409 11005 443
rect 11041 409 11075 443
rect 11111 409 11145 443
rect 11181 409 11215 443
rect 11251 409 11285 443
rect 11321 409 11355 443
rect 11391 409 11425 443
rect 11460 409 11494 443
rect 11529 409 11563 443
rect 11598 409 11632 443
rect 14932 706 14966 740
rect 15000 706 15034 740
rect 15068 706 15102 740
rect 14465 661 14499 695
rect 14543 661 14577 695
rect 14621 661 14655 695
rect 14698 661 14732 695
rect 14775 661 14809 695
rect 14852 661 14886 695
rect 14932 634 14966 668
rect 15000 634 15034 668
rect 15068 634 15102 668
rect 14465 575 14499 609
rect 14543 575 14577 609
rect 14621 575 14655 609
rect 14698 575 14732 609
rect 14775 575 14809 609
rect 14852 575 14886 609
rect 14932 562 14966 596
rect 15000 562 15034 596
rect 15068 562 15102 596
rect 14465 489 14499 523
rect 14543 489 14577 523
rect 14621 489 14655 523
rect 14698 489 14732 523
rect 14775 489 14809 523
rect 14852 489 14886 523
rect 14932 490 14966 524
rect 15000 490 15034 524
rect 15068 490 15102 524
rect 14465 403 14499 437
rect 14543 403 14577 437
rect 14621 403 14655 437
rect 14698 403 14732 437
rect 14775 403 14809 437
rect 14852 403 14886 437
rect 14932 418 14966 452
rect 15000 418 15034 452
rect 15068 418 15102 452
rect 6988 309 7022 343
rect 7056 333 7090 367
rect 7125 333 7159 367
rect 7194 333 7228 367
rect 7263 333 7297 367
rect 7332 333 7366 367
rect 7401 333 7435 367
rect 7470 333 7504 367
rect 7539 333 7573 367
rect 7608 333 7642 367
rect 7677 333 7711 367
rect 7746 333 7780 367
rect 7815 333 7849 367
rect 7884 333 7918 367
rect 7953 333 7987 367
rect 8022 333 8056 367
rect 8091 333 8125 367
rect 8160 333 8194 367
rect 8229 333 8263 367
rect 8298 333 8332 367
rect 8367 333 8401 367
rect 8436 333 8470 367
rect 8505 333 8539 367
rect 8574 333 8608 367
rect 8643 333 8677 367
rect 8712 333 8746 367
rect 8781 333 8815 367
rect 8850 333 8884 367
rect 8919 333 8953 367
rect 8988 333 9022 367
rect 9057 333 9091 367
rect 9126 333 9160 367
rect 9195 333 9229 367
rect 9264 333 9298 367
rect 9333 333 9367 367
rect 9402 333 9436 367
rect 9471 333 9505 367
rect 9540 333 9574 367
rect 9609 333 9643 367
rect 9678 333 9712 367
rect 9747 333 9781 367
rect 9816 333 9850 367
rect 9885 333 9919 367
rect 9954 333 9988 367
rect 10023 333 10057 367
rect 10092 333 10126 367
rect 10161 333 10195 367
rect 10230 333 10264 367
rect 10299 333 10333 367
rect 10368 333 10402 367
rect 10437 333 10471 367
rect 10506 333 10540 367
rect 10575 333 10609 367
rect 10643 333 10677 367
rect 10711 333 10745 367
rect 10779 333 10813 367
rect 10847 333 10881 367
rect 10915 333 10949 367
rect 10983 333 11017 367
rect 11051 333 11085 367
rect 11119 333 11153 367
rect 11187 333 11221 367
rect 11255 333 11289 367
rect 11323 333 11357 367
rect 11391 333 11425 367
rect 11459 333 11493 367
rect 11527 333 11561 367
rect 11595 333 11629 367
rect 11663 333 11697 367
rect 11731 333 11765 367
rect 11799 333 11833 367
rect 11867 333 11901 367
rect 11935 333 11969 367
rect 12003 333 12037 367
rect 12071 333 12105 367
rect 12139 333 12173 367
rect 12207 333 12241 367
rect 12275 333 12309 367
rect 12343 333 12377 367
rect 12411 333 12445 367
rect 12479 333 12513 367
rect 12547 333 12581 367
rect 12615 333 12649 367
rect 12683 333 12717 367
rect 12751 333 12785 367
rect 12819 333 12853 367
rect 12887 333 12921 367
rect 12955 333 12989 367
rect 13023 333 13057 367
rect 13091 333 13125 367
rect 13159 333 13193 367
rect 13227 333 13261 367
rect 13295 333 13329 367
rect 13363 333 13397 367
rect 13431 333 13465 367
rect 13499 333 13533 367
rect 13567 333 13601 367
rect 13635 333 13669 367
rect 13703 333 13737 367
rect 13771 333 13805 367
rect 13839 333 13873 367
rect 13907 333 13941 367
rect 13975 333 14009 367
rect 14043 333 14077 367
rect 14111 333 14145 367
rect 14179 333 14213 367
rect 14247 333 14281 367
rect 14315 333 14349 367
rect 14383 333 14417 367
rect 14451 333 14485 367
rect 14519 333 14553 367
rect 14587 333 14621 367
rect 14655 333 14689 367
rect 14723 333 14757 367
rect 14791 333 14825 367
rect 14859 333 14893 367
rect 14932 346 14966 380
rect 15000 346 15034 380
rect 15068 346 15102 380
rect 6988 241 7022 275
rect 7056 255 7090 289
rect 7125 255 7159 289
rect 7194 255 7228 289
rect 7263 255 7297 289
rect 7332 255 7366 289
rect 7401 255 7435 289
rect 7470 255 7504 289
rect 7539 255 7573 289
rect 7608 255 7642 289
rect 7677 255 7711 289
rect 7746 255 7780 289
rect 7815 255 7849 289
rect 7884 255 7918 289
rect 7953 255 7987 289
rect 8022 255 8056 289
rect 8091 255 8125 289
rect 8160 255 8194 289
rect 8229 255 8263 289
rect 8298 255 8332 289
rect 8367 255 8401 289
rect 8436 255 8470 289
rect 8505 255 8539 289
rect 8574 255 8608 289
rect 8643 255 8677 289
rect 8712 255 8746 289
rect 8781 255 8815 289
rect 8850 255 8884 289
rect 8919 255 8953 289
rect 8988 255 9022 289
rect 9057 255 9091 289
rect 9126 255 9160 289
rect 9195 255 9229 289
rect 9264 255 9298 289
rect 9333 255 9367 289
rect 9402 255 9436 289
rect 9471 255 9505 289
rect 9540 255 9574 289
rect 9609 255 9643 289
rect 9678 255 9712 289
rect 9747 255 9781 289
rect 9816 255 9850 289
rect 9885 255 9919 289
rect 9954 255 9988 289
rect 10023 255 10057 289
rect 10092 255 10126 289
rect 10161 255 10195 289
rect 10230 255 10264 289
rect 10299 255 10333 289
rect 10368 255 10402 289
rect 10437 255 10471 289
rect 10506 255 10540 289
rect 10575 255 10609 289
rect 10643 255 10677 289
rect 10711 255 10745 289
rect 10779 255 10813 289
rect 10847 255 10881 289
rect 10915 255 10949 289
rect 10983 255 11017 289
rect 11051 255 11085 289
rect 11119 255 11153 289
rect 11187 255 11221 289
rect 11255 255 11289 289
rect 11323 255 11357 289
rect 11391 255 11425 289
rect 11459 255 11493 289
rect 11527 255 11561 289
rect 11595 255 11629 289
rect 11663 255 11697 289
rect 11731 255 11765 289
rect 11799 255 11833 289
rect 11867 255 11901 289
rect 11935 255 11969 289
rect 12003 255 12037 289
rect 12071 255 12105 289
rect 12139 255 12173 289
rect 12207 255 12241 289
rect 12275 255 12309 289
rect 12343 255 12377 289
rect 12411 255 12445 289
rect 12479 255 12513 289
rect 12547 255 12581 289
rect 12615 255 12649 289
rect 12683 255 12717 289
rect 12751 255 12785 289
rect 12819 255 12853 289
rect 12887 255 12921 289
rect 12955 255 12989 289
rect 13023 255 13057 289
rect 13091 255 13125 289
rect 13159 255 13193 289
rect 13227 255 13261 289
rect 13295 255 13329 289
rect 13363 255 13397 289
rect 13431 255 13465 289
rect 13499 255 13533 289
rect 13567 255 13601 289
rect 13635 255 13669 289
rect 13703 255 13737 289
rect 13771 255 13805 289
rect 13839 255 13873 289
rect 13907 255 13941 289
rect 13975 255 14009 289
rect 14043 255 14077 289
rect 14111 255 14145 289
rect 14179 255 14213 289
rect 14247 255 14281 289
rect 14315 255 14349 289
rect 14383 255 14417 289
rect 14451 255 14485 289
rect 14519 255 14553 289
rect 14587 255 14621 289
rect 14655 255 14689 289
rect 14723 255 14757 289
rect 14791 255 14825 289
rect 14859 255 14893 289
rect 14932 274 14966 308
rect 15000 274 15034 308
rect 15068 274 15102 308
rect 6988 173 7022 207
rect 7056 177 7090 211
rect 7125 177 7159 211
rect 7194 177 7228 211
rect 7263 177 7297 211
rect 7332 177 7366 211
rect 7401 177 7435 211
rect 7470 177 7504 211
rect 7539 177 7573 211
rect 7608 177 7642 211
rect 7677 177 7711 211
rect 7746 177 7780 211
rect 7815 177 7849 211
rect 7884 177 7918 211
rect 7953 177 7987 211
rect 8022 177 8056 211
rect 8091 177 8125 211
rect 8160 177 8194 211
rect 8229 177 8263 211
rect 8298 177 8332 211
rect 8367 177 8401 211
rect 8436 177 8470 211
rect 8505 177 8539 211
rect 8574 177 8608 211
rect 8643 177 8677 211
rect 8712 177 8746 211
rect 8781 177 8815 211
rect 8850 177 8884 211
rect 8919 177 8953 211
rect 8988 177 9022 211
rect 9057 177 9091 211
rect 9126 177 9160 211
rect 9195 177 9229 211
rect 9264 177 9298 211
rect 9333 177 9367 211
rect 9402 177 9436 211
rect 9471 177 9505 211
rect 9540 177 9574 211
rect 9609 177 9643 211
rect 9678 177 9712 211
rect 9747 177 9781 211
rect 9816 177 9850 211
rect 9885 177 9919 211
rect 9954 177 9988 211
rect 10023 177 10057 211
rect 10092 177 10126 211
rect 10161 177 10195 211
rect 10230 177 10264 211
rect 10299 177 10333 211
rect 10368 177 10402 211
rect 10437 177 10471 211
rect 10506 177 10540 211
rect 10575 177 10609 211
rect 10643 177 10677 211
rect 10711 177 10745 211
rect 10779 177 10813 211
rect 10847 177 10881 211
rect 10915 177 10949 211
rect 10983 177 11017 211
rect 11051 177 11085 211
rect 11119 177 11153 211
rect 11187 177 11221 211
rect 11255 177 11289 211
rect 11323 177 11357 211
rect 11391 177 11425 211
rect 11459 177 11493 211
rect 11527 177 11561 211
rect 11595 177 11629 211
rect 11663 177 11697 211
rect 11731 177 11765 211
rect 11799 177 11833 211
rect 11867 177 11901 211
rect 11935 177 11969 211
rect 12003 177 12037 211
rect 12071 177 12105 211
rect 12139 177 12173 211
rect 12207 177 12241 211
rect 12275 177 12309 211
rect 12343 177 12377 211
rect 12411 177 12445 211
rect 12479 177 12513 211
rect 12547 177 12581 211
rect 12615 177 12649 211
rect 12683 177 12717 211
rect 12751 177 12785 211
rect 12819 177 12853 211
rect 12887 177 12921 211
rect 12955 177 12989 211
rect 13023 177 13057 211
rect 13091 177 13125 211
rect 13159 177 13193 211
rect 13227 177 13261 211
rect 13295 177 13329 211
rect 13363 177 13397 211
rect 13431 177 13465 211
rect 13499 177 13533 211
rect 13567 177 13601 211
rect 13635 177 13669 211
rect 13703 177 13737 211
rect 13771 177 13805 211
rect 13839 177 13873 211
rect 13907 177 13941 211
rect 13975 177 14009 211
rect 14043 177 14077 211
rect 14111 177 14145 211
rect 14179 177 14213 211
rect 14247 177 14281 211
rect 14315 177 14349 211
rect 14383 177 14417 211
rect 14451 177 14485 211
rect 14519 177 14553 211
rect 14587 177 14621 211
rect 14655 177 14689 211
rect 14723 177 14757 211
rect 14791 177 14825 211
rect 14859 177 14893 211
rect 14932 202 14966 236
rect 15000 202 15034 236
rect 15068 202 15102 236
rect 6988 105 7022 139
rect 7056 99 7090 133
rect 7125 99 7159 133
rect 7194 99 7228 133
rect 7263 99 7297 133
rect 7332 99 7366 133
rect 7401 99 7435 133
rect 7470 99 7504 133
rect 7539 99 7573 133
rect 7608 99 7642 133
rect 7677 99 7711 133
rect 7746 99 7780 133
rect 7815 99 7849 133
rect 7884 99 7918 133
rect 7953 99 7987 133
rect 8022 99 8056 133
rect 8091 99 8125 133
rect 8160 99 8194 133
rect 8229 99 8263 133
rect 8298 99 8332 133
rect 8367 99 8401 133
rect 8436 99 8470 133
rect 8505 99 8539 133
rect 8574 99 8608 133
rect 8643 99 8677 133
rect 8712 99 8746 133
rect 8781 99 8815 133
rect 8850 99 8884 133
rect 8919 99 8953 133
rect 8988 99 9022 133
rect 9057 99 9091 133
rect 9126 99 9160 133
rect 9195 99 9229 133
rect 9264 99 9298 133
rect 9333 99 9367 133
rect 9402 99 9436 133
rect 9471 99 9505 133
rect 9540 99 9574 133
rect 9609 99 9643 133
rect 9678 99 9712 133
rect 9747 99 9781 133
rect 9816 99 9850 133
rect 9885 99 9919 133
rect 9954 99 9988 133
rect 10023 99 10057 133
rect 10092 99 10126 133
rect 10161 99 10195 133
rect 10230 99 10264 133
rect 10299 99 10333 133
rect 10368 99 10402 133
rect 10437 99 10471 133
rect 10506 99 10540 133
rect 10575 99 10609 133
rect 10643 99 10677 133
rect 10711 99 10745 133
rect 10779 99 10813 133
rect 10847 99 10881 133
rect 10915 99 10949 133
rect 10983 99 11017 133
rect 11051 99 11085 133
rect 11119 99 11153 133
rect 11187 99 11221 133
rect 11255 99 11289 133
rect 11323 99 11357 133
rect 11391 99 11425 133
rect 11459 99 11493 133
rect 11527 99 11561 133
rect 11595 99 11629 133
rect 11663 99 11697 133
rect 11731 99 11765 133
rect 11799 99 11833 133
rect 11867 99 11901 133
rect 11935 99 11969 133
rect 12003 99 12037 133
rect 12071 99 12105 133
rect 12139 99 12173 133
rect 12207 99 12241 133
rect 12275 99 12309 133
rect 12343 99 12377 133
rect 12411 99 12445 133
rect 12479 99 12513 133
rect 12547 99 12581 133
rect 12615 99 12649 133
rect 12683 99 12717 133
rect 12751 99 12785 133
rect 12819 99 12853 133
rect 12887 99 12921 133
rect 12955 99 12989 133
rect 13023 99 13057 133
rect 13091 99 13125 133
rect 13159 99 13193 133
rect 13227 99 13261 133
rect 13295 99 13329 133
rect 13363 99 13397 133
rect 13431 99 13465 133
rect 13499 99 13533 133
rect 13567 99 13601 133
rect 13635 99 13669 133
rect 13703 99 13737 133
rect 13771 99 13805 133
rect 13839 99 13873 133
rect 13907 99 13941 133
rect 13975 99 14009 133
rect 14043 99 14077 133
rect 14111 99 14145 133
rect 14179 99 14213 133
rect 14247 99 14281 133
rect 14315 99 14349 133
rect 14383 99 14417 133
rect 14451 99 14485 133
rect 14519 99 14553 133
rect 14587 99 14621 133
rect 14655 99 14689 133
rect 14723 99 14757 133
rect 14791 99 14825 133
rect 14859 99 14893 133
rect 14932 130 14966 164
rect 15000 130 15034 164
rect 15068 130 15102 164
rect 14932 57 14966 91
rect 15000 57 15034 91
rect 15068 57 15102 91
rect 3632 -11 3666 23
rect 3700 -11 3734 23
rect 3768 -11 3802 23
rect 3836 -11 3870 23
rect 3904 -11 3938 23
rect 3972 -11 4006 23
rect 4040 -11 4074 23
rect 4108 -11 4142 23
rect 4176 -11 4210 23
rect 4244 -11 4278 23
rect 4312 -11 4346 23
rect 4380 -11 4414 23
rect 4448 -11 4482 23
rect 4516 -11 4550 23
rect 4584 -11 4618 23
rect 4652 -11 4686 23
rect 4720 -11 4754 23
rect 4788 -11 4822 23
rect 4856 -11 4890 23
rect 4924 -11 4958 23
rect 4992 -11 5026 23
rect 5060 -11 5094 23
rect 5128 -11 5162 23
rect 5196 -11 5230 23
rect 5264 -11 5298 23
rect 5332 -11 5366 23
rect 5400 -11 5434 23
rect 5468 -11 5502 23
rect 5536 -11 5570 23
rect 5604 -11 5638 23
rect 5672 -11 5706 23
rect 5740 -11 5774 23
rect 5808 -11 5842 23
rect 5876 -11 5910 23
rect 5944 -11 5978 23
rect 6012 -11 6046 23
rect 6080 -11 6114 23
rect 6148 -11 6182 23
rect 6216 -11 6250 23
rect 6284 -11 6318 23
rect 6352 -11 6386 23
rect 6420 -11 6454 23
rect 6488 -11 6522 23
rect 6556 -11 6590 23
rect 6624 -11 6658 23
rect 6692 -11 6726 23
rect 6760 -11 6794 23
rect 6828 -11 6862 23
rect 6896 -11 6930 23
rect 6964 -11 6998 23
rect 7056 21 7090 55
rect 7125 21 7159 55
rect 7194 21 7228 55
rect 7263 21 7297 55
rect 7332 21 7366 55
rect 7401 21 7435 55
rect 7470 21 7504 55
rect 7539 21 7573 55
rect 7608 21 7642 55
rect 7677 21 7711 55
rect 7746 21 7780 55
rect 7815 21 7849 55
rect 7884 21 7918 55
rect 7953 21 7987 55
rect 8022 21 8056 55
rect 8091 21 8125 55
rect 8160 21 8194 55
rect 8229 21 8263 55
rect 8298 21 8332 55
rect 8367 21 8401 55
rect 8436 21 8470 55
rect 8505 21 8539 55
rect 8574 21 8608 55
rect 8643 21 8677 55
rect 8712 21 8746 55
rect 8781 21 8815 55
rect 8850 21 8884 55
rect 8919 21 8953 55
rect 8988 21 9022 55
rect 9057 21 9091 55
rect 9126 21 9160 55
rect 9195 21 9229 55
rect 9264 21 9298 55
rect 9333 21 9367 55
rect 9402 21 9436 55
rect 9471 21 9505 55
rect 9540 21 9574 55
rect 9609 21 9643 55
rect 9678 21 9712 55
rect 9747 21 9781 55
rect 9816 21 9850 55
rect 9885 21 9919 55
rect 9954 21 9988 55
rect 10023 21 10057 55
rect 10092 21 10126 55
rect 10161 21 10195 55
rect 10230 21 10264 55
rect 10299 21 10333 55
rect 10368 21 10402 55
rect 10437 21 10471 55
rect 10506 21 10540 55
rect 10575 21 10609 55
rect 10643 21 10677 55
rect 10711 21 10745 55
rect 10779 21 10813 55
rect 10847 21 10881 55
rect 10915 21 10949 55
rect 10983 21 11017 55
rect 11051 21 11085 55
rect 11119 21 11153 55
rect 11187 21 11221 55
rect 11255 21 11289 55
rect 11323 21 11357 55
rect 11391 21 11425 55
rect 11459 21 11493 55
rect 11527 21 11561 55
rect 11595 21 11629 55
rect 11663 21 11697 55
rect 11731 21 11765 55
rect 11799 21 11833 55
rect 11867 21 11901 55
rect 11935 21 11969 55
rect 12003 21 12037 55
rect 12071 21 12105 55
rect 12139 21 12173 55
rect 12207 21 12241 55
rect 12275 21 12309 55
rect 12343 21 12377 55
rect 12411 21 12445 55
rect 12479 21 12513 55
rect 12547 21 12581 55
rect 12615 21 12649 55
rect 12683 21 12717 55
rect 12751 21 12785 55
rect 12819 21 12853 55
rect 12887 21 12921 55
rect 12955 21 12989 55
rect 13023 21 13057 55
rect 13091 21 13125 55
rect 13159 21 13193 55
rect 13227 21 13261 55
rect 13295 21 13329 55
rect 13363 21 13397 55
rect 13431 21 13465 55
rect 13499 21 13533 55
rect 13567 21 13601 55
rect 13635 21 13669 55
rect 13703 21 13737 55
rect 13771 21 13805 55
rect 13839 21 13873 55
rect 13907 21 13941 55
rect 13975 21 14009 55
rect 14043 21 14077 55
rect 14111 21 14145 55
rect 14179 21 14213 55
rect 14247 21 14281 55
rect 14315 21 14349 55
rect 14383 21 14417 55
rect 14451 21 14485 55
rect 14519 21 14553 55
rect 14587 21 14621 55
rect 14655 21 14689 55
rect 14723 21 14757 55
rect 14791 21 14825 55
rect 14859 21 14893 55
<< mvnsubdiffcont >>
rect 68 16459 102 16493
rect 139 16459 173 16493
rect 210 16459 244 16493
rect 281 16459 315 16493
rect 352 16459 386 16493
rect 444 16459 478 16493
rect 513 16459 547 16493
rect 582 16459 616 16493
rect 651 16459 685 16493
rect 720 16459 754 16493
rect 789 16459 823 16493
rect 858 16459 892 16493
rect 927 16459 961 16493
rect 996 16459 1030 16493
rect 1065 16459 1099 16493
rect 1134 16459 1168 16493
rect 1203 16459 1237 16493
rect 1272 16459 1306 16493
rect 1341 16459 1375 16493
rect 1410 16459 1444 16493
rect 1479 16459 1513 16493
rect 1548 16459 1582 16493
rect 1617 16459 1651 16493
rect 1686 16459 1720 16493
rect 1755 16459 1789 16493
rect 1824 16459 1858 16493
rect 1893 16459 1927 16493
rect 1962 16459 1996 16493
rect 2031 16459 2065 16493
rect 2100 16459 2134 16493
rect 2169 16459 2203 16493
rect 2238 16459 2272 16493
rect 2307 16459 2341 16493
rect 2376 16459 2410 16493
rect 2445 16459 2479 16493
rect 2514 16459 2548 16493
rect 2583 16459 2617 16493
rect 2652 16459 2686 16493
rect 2721 16459 2755 16493
rect 2790 16459 2824 16493
rect 2859 16459 2893 16493
rect 2928 16459 2962 16493
rect 2996 16459 3030 16493
rect 3064 16459 3098 16493
rect 3132 16459 3166 16493
rect 3200 16459 3234 16493
rect 3268 16459 3302 16493
rect 3336 16459 3370 16493
rect 3404 16459 3438 16493
rect 3472 16459 3506 16493
rect 3540 16459 3574 16493
rect 3608 16459 3642 16493
rect 3676 16459 3710 16493
rect 3744 16459 3778 16493
rect 3812 16459 3846 16493
rect 3880 16459 3914 16493
rect 3948 16459 3982 16493
rect 4016 16459 4050 16493
rect 4084 16459 4118 16493
rect 4152 16459 4186 16493
rect 4220 16459 4254 16493
rect 4288 16459 4322 16493
rect 4356 16459 4390 16493
rect 4424 16459 4458 16493
rect 4492 16459 4526 16493
rect 4560 16459 4594 16493
rect 4628 16459 4662 16493
rect 4696 16459 4730 16493
rect 4764 16459 4798 16493
rect 4832 16459 4866 16493
rect 4900 16459 4934 16493
rect 4968 16459 5002 16493
rect 5036 16459 5070 16493
rect 5104 16459 5138 16493
rect 5172 16459 5206 16493
rect 5240 16459 5274 16493
rect 5308 16459 5342 16493
rect 5376 16459 5410 16493
rect 5444 16459 5478 16493
rect 5512 16459 5546 16493
rect 5580 16459 5614 16493
rect 5648 16459 5682 16493
rect 5716 16459 5750 16493
rect 5784 16459 5818 16493
rect 5852 16459 5886 16493
rect 5920 16459 5954 16493
rect 5988 16459 6022 16493
rect 6056 16459 6090 16493
rect 6124 16459 6158 16493
rect 6192 16459 6226 16493
rect 6260 16459 6294 16493
rect 6328 16459 6362 16493
rect 6396 16459 6430 16493
rect 6464 16459 6498 16493
rect 6532 16459 6566 16493
rect 6600 16459 6634 16493
rect 6668 16459 6702 16493
rect 6736 16459 6770 16493
rect 6804 16459 6838 16493
rect 6872 16459 6906 16493
rect 6940 16459 6974 16493
rect 7008 16459 7042 16493
rect 7076 16459 7110 16493
rect 7144 16459 7178 16493
rect 7212 16459 7246 16493
rect 7280 16459 7314 16493
rect 7348 16459 7382 16493
rect 7416 16459 7450 16493
rect 7484 16459 7518 16493
rect 7552 16459 7586 16493
rect 7620 16459 7654 16493
rect 7688 16459 7722 16493
rect 7756 16459 7790 16493
rect 7824 16459 7858 16493
rect 7892 16459 7926 16493
rect 7960 16459 7994 16493
rect 8028 16459 8062 16493
rect 8096 16459 8130 16493
rect 8164 16459 8198 16493
rect 8232 16459 8266 16493
rect 8300 16459 8334 16493
rect 8368 16459 8402 16493
rect 8436 16459 8470 16493
rect 8504 16459 8538 16493
rect 8572 16459 8606 16493
rect 8640 16459 8674 16493
rect 8708 16459 8742 16493
rect 8776 16459 8810 16493
rect 8844 16459 8878 16493
rect 8912 16459 8946 16493
rect 8980 16459 9014 16493
rect 9048 16459 9082 16493
rect 9116 16459 9150 16493
rect 9184 16459 9218 16493
rect 9252 16459 9286 16493
rect 9320 16459 9354 16493
rect 9388 16459 9422 16493
rect 9456 16459 9490 16493
rect 9524 16459 9558 16493
rect 9592 16459 9626 16493
rect 9660 16459 9694 16493
rect 9728 16459 9762 16493
rect 9796 16459 9830 16493
rect 9864 16459 9898 16493
rect 9932 16459 9966 16493
rect 10000 16459 10034 16493
rect 10068 16459 10102 16493
rect 10136 16459 10170 16493
rect 10204 16459 10238 16493
rect 10272 16459 10306 16493
rect 10340 16459 10374 16493
rect 10408 16459 10442 16493
rect 10476 16459 10510 16493
rect 10544 16459 10578 16493
rect 10612 16459 10646 16493
rect 10680 16459 10714 16493
rect 10748 16459 10782 16493
rect 10816 16459 10850 16493
rect 10884 16459 10918 16493
rect 10952 16459 10986 16493
rect 11020 16459 11054 16493
rect 11088 16459 11122 16493
rect 11156 16459 11190 16493
rect 11224 16459 11258 16493
rect 11292 16459 11326 16493
rect 11360 16459 11394 16493
rect 11428 16459 11462 16493
rect 11496 16459 11530 16493
rect 11564 16459 11598 16493
rect 11632 16459 11666 16493
rect 11700 16459 11734 16493
rect 11768 16459 11802 16493
rect 11836 16459 11870 16493
rect 11904 16459 11938 16493
rect 11972 16459 12006 16493
rect 12040 16459 12074 16493
rect 12108 16459 12142 16493
rect 12176 16459 12210 16493
rect 12244 16459 12278 16493
rect 12312 16459 12346 16493
rect 12380 16459 12414 16493
rect 12448 16459 12482 16493
rect 12516 16459 12550 16493
rect 12584 16459 12618 16493
rect 12652 16459 12686 16493
rect 12720 16459 12754 16493
rect 12788 16459 12822 16493
rect 12856 16459 12890 16493
rect 12924 16459 12958 16493
rect 12992 16459 13026 16493
rect 13060 16459 13094 16493
rect 13128 16459 13162 16493
rect 13196 16459 13230 16493
rect 13264 16459 13298 16493
rect 13332 16459 13366 16493
rect 13400 16459 13434 16493
rect 13468 16459 13502 16493
rect 13536 16459 13570 16493
rect 13604 16459 13638 16493
rect 13672 16459 13706 16493
rect 13740 16459 13774 16493
rect 13808 16459 13842 16493
rect 13876 16459 13910 16493
rect 13944 16459 13978 16493
rect 14012 16459 14046 16493
rect 14080 16459 14114 16493
rect 14148 16459 14182 16493
rect 14216 16459 14250 16493
rect 14284 16459 14318 16493
rect 14352 16459 14386 16493
rect 14420 16469 14454 16503
rect 14492 16469 14526 16503
rect 14564 16469 14598 16503
rect 14636 16469 14670 16503
rect 14708 16469 14742 16503
rect 14780 16469 14814 16503
rect 14852 16469 14886 16503
rect 14924 16469 14958 16503
rect 14996 16469 15030 16503
rect 15068 16469 15102 16503
rect 68 16391 102 16425
rect 139 16391 173 16425
rect 210 16391 244 16425
rect 281 16391 315 16425
rect 352 16391 386 16425
rect 444 16389 478 16423
rect 513 16389 547 16423
rect 582 16389 616 16423
rect 651 16389 685 16423
rect 720 16389 754 16423
rect 789 16389 823 16423
rect 858 16389 892 16423
rect 927 16389 961 16423
rect 996 16389 1030 16423
rect 1065 16389 1099 16423
rect 1134 16389 1168 16423
rect 1203 16389 1237 16423
rect 1272 16389 1306 16423
rect 1341 16389 1375 16423
rect 1410 16389 1444 16423
rect 1479 16389 1513 16423
rect 1548 16389 1582 16423
rect 1617 16389 1651 16423
rect 1686 16389 1720 16423
rect 1755 16389 1789 16423
rect 1824 16389 1858 16423
rect 1893 16389 1927 16423
rect 1962 16389 1996 16423
rect 2031 16389 2065 16423
rect 2100 16389 2134 16423
rect 2169 16389 2203 16423
rect 2238 16389 2272 16423
rect 2307 16389 2341 16423
rect 2376 16389 2410 16423
rect 2445 16389 2479 16423
rect 2514 16389 2548 16423
rect 2583 16389 2617 16423
rect 2652 16389 2686 16423
rect 2721 16389 2755 16423
rect 2790 16389 2824 16423
rect 2859 16389 2893 16423
rect 2928 16389 2962 16423
rect 2996 16389 3030 16423
rect 3064 16389 3098 16423
rect 3132 16389 3166 16423
rect 3200 16389 3234 16423
rect 3268 16389 3302 16423
rect 3336 16389 3370 16423
rect 3404 16389 3438 16423
rect 3472 16389 3506 16423
rect 3540 16389 3574 16423
rect 3608 16389 3642 16423
rect 3676 16389 3710 16423
rect 3744 16389 3778 16423
rect 3812 16389 3846 16423
rect 3880 16389 3914 16423
rect 3948 16389 3982 16423
rect 4016 16389 4050 16423
rect 4084 16389 4118 16423
rect 4152 16389 4186 16423
rect 4220 16389 4254 16423
rect 4288 16389 4322 16423
rect 4356 16389 4390 16423
rect 4424 16389 4458 16423
rect 4492 16389 4526 16423
rect 4560 16389 4594 16423
rect 4628 16389 4662 16423
rect 4696 16389 4730 16423
rect 4764 16389 4798 16423
rect 4832 16389 4866 16423
rect 4900 16389 4934 16423
rect 4968 16389 5002 16423
rect 5036 16389 5070 16423
rect 5104 16389 5138 16423
rect 5172 16389 5206 16423
rect 5240 16389 5274 16423
rect 5308 16389 5342 16423
rect 5376 16389 5410 16423
rect 5444 16389 5478 16423
rect 5512 16389 5546 16423
rect 5580 16389 5614 16423
rect 5648 16389 5682 16423
rect 5716 16389 5750 16423
rect 5784 16389 5818 16423
rect 5852 16389 5886 16423
rect 5920 16389 5954 16423
rect 5988 16389 6022 16423
rect 6056 16389 6090 16423
rect 6124 16389 6158 16423
rect 6192 16389 6226 16423
rect 6260 16389 6294 16423
rect 6328 16389 6362 16423
rect 6396 16389 6430 16423
rect 6464 16389 6498 16423
rect 6532 16389 6566 16423
rect 6600 16389 6634 16423
rect 6668 16389 6702 16423
rect 6736 16389 6770 16423
rect 6804 16389 6838 16423
rect 6872 16389 6906 16423
rect 6940 16389 6974 16423
rect 7008 16389 7042 16423
rect 7076 16389 7110 16423
rect 7144 16389 7178 16423
rect 7212 16389 7246 16423
rect 7280 16389 7314 16423
rect 7348 16389 7382 16423
rect 7416 16389 7450 16423
rect 7484 16389 7518 16423
rect 7552 16389 7586 16423
rect 7620 16389 7654 16423
rect 7688 16389 7722 16423
rect 7756 16389 7790 16423
rect 7824 16389 7858 16423
rect 7892 16389 7926 16423
rect 7960 16389 7994 16423
rect 8028 16389 8062 16423
rect 8096 16389 8130 16423
rect 8164 16389 8198 16423
rect 8232 16389 8266 16423
rect 8300 16389 8334 16423
rect 8368 16389 8402 16423
rect 8436 16389 8470 16423
rect 8504 16389 8538 16423
rect 8572 16389 8606 16423
rect 8640 16389 8674 16423
rect 8708 16389 8742 16423
rect 8776 16389 8810 16423
rect 8844 16389 8878 16423
rect 8912 16389 8946 16423
rect 8980 16389 9014 16423
rect 9048 16389 9082 16423
rect 9116 16389 9150 16423
rect 9184 16389 9218 16423
rect 9252 16389 9286 16423
rect 9320 16389 9354 16423
rect 9388 16389 9422 16423
rect 9456 16389 9490 16423
rect 9524 16389 9558 16423
rect 9592 16389 9626 16423
rect 9660 16389 9694 16423
rect 9728 16389 9762 16423
rect 9796 16389 9830 16423
rect 9864 16389 9898 16423
rect 9932 16389 9966 16423
rect 10000 16389 10034 16423
rect 10068 16389 10102 16423
rect 10136 16389 10170 16423
rect 10204 16389 10238 16423
rect 10272 16389 10306 16423
rect 10340 16389 10374 16423
rect 10408 16389 10442 16423
rect 10476 16389 10510 16423
rect 10544 16389 10578 16423
rect 10612 16389 10646 16423
rect 10680 16389 10714 16423
rect 10748 16389 10782 16423
rect 10816 16389 10850 16423
rect 10884 16389 10918 16423
rect 10952 16389 10986 16423
rect 11020 16389 11054 16423
rect 11088 16389 11122 16423
rect 11156 16389 11190 16423
rect 11224 16389 11258 16423
rect 11292 16389 11326 16423
rect 11360 16389 11394 16423
rect 11428 16389 11462 16423
rect 11496 16389 11530 16423
rect 11564 16389 11598 16423
rect 11632 16389 11666 16423
rect 11700 16389 11734 16423
rect 11768 16389 11802 16423
rect 11836 16389 11870 16423
rect 11904 16389 11938 16423
rect 11972 16389 12006 16423
rect 12040 16389 12074 16423
rect 12108 16389 12142 16423
rect 12176 16389 12210 16423
rect 12244 16389 12278 16423
rect 12312 16389 12346 16423
rect 12380 16389 12414 16423
rect 12448 16389 12482 16423
rect 12516 16389 12550 16423
rect 12584 16389 12618 16423
rect 12652 16389 12686 16423
rect 12720 16389 12754 16423
rect 12788 16389 12822 16423
rect 12856 16389 12890 16423
rect 12924 16389 12958 16423
rect 12992 16389 13026 16423
rect 13060 16389 13094 16423
rect 13128 16389 13162 16423
rect 13196 16389 13230 16423
rect 13264 16389 13298 16423
rect 13332 16389 13366 16423
rect 13400 16389 13434 16423
rect 13468 16389 13502 16423
rect 13536 16389 13570 16423
rect 13604 16389 13638 16423
rect 13672 16389 13706 16423
rect 13740 16389 13774 16423
rect 13808 16389 13842 16423
rect 13876 16389 13910 16423
rect 13944 16389 13978 16423
rect 14012 16389 14046 16423
rect 14080 16389 14114 16423
rect 14148 16389 14182 16423
rect 14216 16389 14250 16423
rect 14284 16389 14318 16423
rect 14352 16389 14386 16423
rect 14420 16400 14454 16434
rect 14492 16400 14526 16434
rect 14564 16400 14598 16434
rect 14636 16400 14670 16434
rect 14708 16400 14742 16434
rect 14780 16400 14814 16434
rect 14852 16400 14886 16434
rect 14924 16400 14958 16434
rect 14996 16400 15030 16434
rect 15068 16400 15102 16434
rect 68 16323 102 16357
rect 139 16323 173 16357
rect 210 16323 244 16357
rect 281 16323 315 16357
rect 352 16323 386 16357
rect 444 16319 478 16353
rect 513 16319 547 16353
rect 582 16319 616 16353
rect 651 16319 685 16353
rect 720 16319 754 16353
rect 789 16319 823 16353
rect 858 16319 892 16353
rect 927 16319 961 16353
rect 996 16319 1030 16353
rect 1065 16319 1099 16353
rect 1134 16319 1168 16353
rect 1203 16319 1237 16353
rect 1272 16319 1306 16353
rect 1341 16319 1375 16353
rect 1410 16319 1444 16353
rect 1479 16319 1513 16353
rect 1548 16319 1582 16353
rect 1617 16319 1651 16353
rect 1686 16319 1720 16353
rect 1755 16319 1789 16353
rect 1824 16319 1858 16353
rect 1893 16319 1927 16353
rect 1962 16319 1996 16353
rect 2031 16319 2065 16353
rect 2100 16319 2134 16353
rect 2169 16319 2203 16353
rect 2238 16319 2272 16353
rect 2307 16319 2341 16353
rect 2376 16319 2410 16353
rect 2445 16319 2479 16353
rect 2514 16319 2548 16353
rect 2583 16319 2617 16353
rect 2652 16319 2686 16353
rect 2721 16319 2755 16353
rect 2790 16319 2824 16353
rect 2859 16319 2893 16353
rect 2928 16319 2962 16353
rect 2996 16319 3030 16353
rect 3064 16319 3098 16353
rect 3132 16319 3166 16353
rect 3200 16319 3234 16353
rect 3268 16319 3302 16353
rect 3336 16319 3370 16353
rect 3404 16319 3438 16353
rect 3472 16319 3506 16353
rect 3540 16319 3574 16353
rect 3608 16319 3642 16353
rect 3676 16319 3710 16353
rect 3744 16319 3778 16353
rect 3812 16319 3846 16353
rect 3880 16319 3914 16353
rect 3948 16319 3982 16353
rect 4016 16319 4050 16353
rect 4084 16319 4118 16353
rect 4152 16319 4186 16353
rect 4220 16319 4254 16353
rect 4288 16319 4322 16353
rect 4356 16319 4390 16353
rect 4424 16319 4458 16353
rect 4492 16319 4526 16353
rect 4560 16319 4594 16353
rect 4628 16319 4662 16353
rect 4696 16319 4730 16353
rect 4764 16319 4798 16353
rect 4832 16319 4866 16353
rect 4900 16319 4934 16353
rect 4968 16319 5002 16353
rect 5036 16319 5070 16353
rect 5104 16319 5138 16353
rect 5172 16319 5206 16353
rect 5240 16319 5274 16353
rect 5308 16319 5342 16353
rect 5376 16319 5410 16353
rect 5444 16319 5478 16353
rect 5512 16319 5546 16353
rect 5580 16319 5614 16353
rect 5648 16319 5682 16353
rect 5716 16319 5750 16353
rect 5784 16319 5818 16353
rect 5852 16319 5886 16353
rect 5920 16319 5954 16353
rect 5988 16319 6022 16353
rect 6056 16319 6090 16353
rect 6124 16319 6158 16353
rect 6192 16319 6226 16353
rect 6260 16319 6294 16353
rect 6328 16319 6362 16353
rect 6396 16319 6430 16353
rect 6464 16319 6498 16353
rect 6532 16319 6566 16353
rect 6600 16319 6634 16353
rect 6668 16319 6702 16353
rect 6736 16319 6770 16353
rect 6804 16319 6838 16353
rect 6872 16319 6906 16353
rect 6940 16319 6974 16353
rect 7008 16319 7042 16353
rect 7076 16319 7110 16353
rect 7144 16319 7178 16353
rect 7212 16319 7246 16353
rect 7280 16319 7314 16353
rect 7348 16319 7382 16353
rect 7416 16319 7450 16353
rect 7484 16319 7518 16353
rect 7552 16319 7586 16353
rect 7620 16319 7654 16353
rect 7688 16319 7722 16353
rect 7756 16319 7790 16353
rect 7824 16319 7858 16353
rect 7892 16319 7926 16353
rect 7960 16319 7994 16353
rect 8028 16319 8062 16353
rect 8096 16319 8130 16353
rect 8164 16319 8198 16353
rect 8232 16319 8266 16353
rect 8300 16319 8334 16353
rect 8368 16319 8402 16353
rect 8436 16319 8470 16353
rect 8504 16319 8538 16353
rect 8572 16319 8606 16353
rect 8640 16319 8674 16353
rect 8708 16319 8742 16353
rect 8776 16319 8810 16353
rect 8844 16319 8878 16353
rect 8912 16319 8946 16353
rect 8980 16319 9014 16353
rect 9048 16319 9082 16353
rect 9116 16319 9150 16353
rect 9184 16319 9218 16353
rect 9252 16319 9286 16353
rect 9320 16319 9354 16353
rect 9388 16319 9422 16353
rect 9456 16319 9490 16353
rect 9524 16319 9558 16353
rect 9592 16319 9626 16353
rect 9660 16319 9694 16353
rect 9728 16319 9762 16353
rect 9796 16319 9830 16353
rect 9864 16319 9898 16353
rect 9932 16319 9966 16353
rect 10000 16319 10034 16353
rect 10068 16319 10102 16353
rect 10136 16319 10170 16353
rect 10204 16319 10238 16353
rect 10272 16319 10306 16353
rect 10340 16319 10374 16353
rect 10408 16319 10442 16353
rect 10476 16319 10510 16353
rect 10544 16319 10578 16353
rect 10612 16319 10646 16353
rect 10680 16319 10714 16353
rect 10748 16319 10782 16353
rect 10816 16319 10850 16353
rect 10884 16319 10918 16353
rect 10952 16319 10986 16353
rect 11020 16319 11054 16353
rect 11088 16319 11122 16353
rect 11156 16319 11190 16353
rect 11224 16319 11258 16353
rect 11292 16319 11326 16353
rect 11360 16319 11394 16353
rect 11428 16319 11462 16353
rect 11496 16319 11530 16353
rect 11564 16319 11598 16353
rect 11632 16319 11666 16353
rect 11700 16319 11734 16353
rect 11768 16319 11802 16353
rect 11836 16319 11870 16353
rect 11904 16319 11938 16353
rect 11972 16319 12006 16353
rect 12040 16319 12074 16353
rect 12108 16319 12142 16353
rect 12176 16319 12210 16353
rect 12244 16319 12278 16353
rect 12312 16319 12346 16353
rect 12380 16319 12414 16353
rect 12448 16319 12482 16353
rect 12516 16319 12550 16353
rect 12584 16319 12618 16353
rect 12652 16319 12686 16353
rect 12720 16319 12754 16353
rect 12788 16319 12822 16353
rect 12856 16319 12890 16353
rect 12924 16319 12958 16353
rect 12992 16319 13026 16353
rect 13060 16319 13094 16353
rect 13128 16319 13162 16353
rect 13196 16319 13230 16353
rect 13264 16319 13298 16353
rect 13332 16319 13366 16353
rect 13400 16319 13434 16353
rect 13468 16319 13502 16353
rect 13536 16319 13570 16353
rect 13604 16319 13638 16353
rect 13672 16319 13706 16353
rect 13740 16319 13774 16353
rect 13808 16319 13842 16353
rect 13876 16319 13910 16353
rect 13944 16319 13978 16353
rect 14012 16319 14046 16353
rect 14080 16319 14114 16353
rect 14148 16319 14182 16353
rect 14216 16319 14250 16353
rect 14284 16319 14318 16353
rect 14352 16319 14386 16353
rect 14420 16331 14454 16365
rect 14492 16331 14526 16365
rect 14564 16331 14598 16365
rect 14636 16331 14670 16365
rect 14708 16331 14742 16365
rect 14780 16331 14814 16365
rect 14852 16331 14886 16365
rect 14924 16331 14958 16365
rect 14996 16331 15030 16365
rect 15068 16331 15102 16365
rect 68 16255 102 16289
rect 139 16255 173 16289
rect 210 16255 244 16289
rect 281 16255 315 16289
rect 352 16255 386 16289
rect 444 16249 478 16283
rect 513 16249 547 16283
rect 582 16249 616 16283
rect 651 16249 685 16283
rect 720 16249 754 16283
rect 789 16249 823 16283
rect 858 16249 892 16283
rect 927 16249 961 16283
rect 996 16249 1030 16283
rect 1065 16249 1099 16283
rect 1134 16249 1168 16283
rect 1203 16249 1237 16283
rect 1272 16249 1306 16283
rect 1341 16249 1375 16283
rect 1410 16249 1444 16283
rect 1479 16249 1513 16283
rect 1548 16249 1582 16283
rect 1617 16249 1651 16283
rect 1686 16249 1720 16283
rect 1755 16249 1789 16283
rect 1824 16249 1858 16283
rect 1893 16249 1927 16283
rect 1962 16249 1996 16283
rect 2031 16249 2065 16283
rect 2100 16249 2134 16283
rect 2169 16249 2203 16283
rect 2238 16249 2272 16283
rect 2307 16249 2341 16283
rect 2376 16249 2410 16283
rect 2445 16249 2479 16283
rect 2514 16249 2548 16283
rect 2583 16249 2617 16283
rect 2652 16249 2686 16283
rect 2721 16249 2755 16283
rect 2790 16249 2824 16283
rect 2859 16249 2893 16283
rect 2928 16249 2962 16283
rect 2996 16249 3030 16283
rect 3064 16249 3098 16283
rect 3132 16249 3166 16283
rect 3200 16249 3234 16283
rect 3268 16249 3302 16283
rect 3336 16249 3370 16283
rect 3404 16249 3438 16283
rect 3472 16249 3506 16283
rect 3540 16249 3574 16283
rect 3608 16249 3642 16283
rect 3676 16249 3710 16283
rect 3744 16249 3778 16283
rect 3812 16249 3846 16283
rect 3880 16249 3914 16283
rect 3948 16249 3982 16283
rect 4016 16249 4050 16283
rect 4084 16249 4118 16283
rect 4152 16249 4186 16283
rect 4220 16249 4254 16283
rect 4288 16249 4322 16283
rect 4356 16249 4390 16283
rect 4424 16249 4458 16283
rect 4492 16249 4526 16283
rect 4560 16249 4594 16283
rect 4628 16249 4662 16283
rect 4696 16249 4730 16283
rect 4764 16249 4798 16283
rect 4832 16249 4866 16283
rect 4900 16249 4934 16283
rect 4968 16249 5002 16283
rect 5036 16249 5070 16283
rect 5104 16249 5138 16283
rect 5172 16249 5206 16283
rect 5240 16249 5274 16283
rect 5308 16249 5342 16283
rect 5376 16249 5410 16283
rect 5444 16249 5478 16283
rect 5512 16249 5546 16283
rect 5580 16249 5614 16283
rect 5648 16249 5682 16283
rect 5716 16249 5750 16283
rect 5784 16249 5818 16283
rect 5852 16249 5886 16283
rect 5920 16249 5954 16283
rect 5988 16249 6022 16283
rect 6056 16249 6090 16283
rect 6124 16249 6158 16283
rect 6192 16249 6226 16283
rect 6260 16249 6294 16283
rect 6328 16249 6362 16283
rect 6396 16249 6430 16283
rect 6464 16249 6498 16283
rect 6532 16249 6566 16283
rect 6600 16249 6634 16283
rect 6668 16249 6702 16283
rect 6736 16249 6770 16283
rect 6804 16249 6838 16283
rect 6872 16249 6906 16283
rect 6940 16249 6974 16283
rect 7008 16249 7042 16283
rect 7076 16249 7110 16283
rect 7144 16249 7178 16283
rect 7212 16249 7246 16283
rect 7280 16249 7314 16283
rect 7348 16249 7382 16283
rect 7416 16249 7450 16283
rect 7484 16249 7518 16283
rect 7552 16249 7586 16283
rect 7620 16249 7654 16283
rect 7688 16249 7722 16283
rect 7756 16249 7790 16283
rect 7824 16249 7858 16283
rect 7892 16249 7926 16283
rect 7960 16249 7994 16283
rect 8028 16249 8062 16283
rect 8096 16249 8130 16283
rect 8164 16249 8198 16283
rect 8232 16249 8266 16283
rect 8300 16249 8334 16283
rect 8368 16249 8402 16283
rect 8436 16249 8470 16283
rect 8504 16249 8538 16283
rect 8572 16249 8606 16283
rect 8640 16249 8674 16283
rect 8708 16249 8742 16283
rect 8776 16249 8810 16283
rect 8844 16249 8878 16283
rect 8912 16249 8946 16283
rect 8980 16249 9014 16283
rect 9048 16249 9082 16283
rect 9116 16249 9150 16283
rect 9184 16249 9218 16283
rect 9252 16249 9286 16283
rect 9320 16249 9354 16283
rect 9388 16249 9422 16283
rect 9456 16249 9490 16283
rect 9524 16249 9558 16283
rect 9592 16249 9626 16283
rect 9660 16249 9694 16283
rect 9728 16249 9762 16283
rect 9796 16249 9830 16283
rect 9864 16249 9898 16283
rect 9932 16249 9966 16283
rect 10000 16249 10034 16283
rect 10068 16249 10102 16283
rect 10136 16249 10170 16283
rect 10204 16249 10238 16283
rect 10272 16249 10306 16283
rect 10340 16249 10374 16283
rect 10408 16249 10442 16283
rect 10476 16249 10510 16283
rect 10544 16249 10578 16283
rect 10612 16249 10646 16283
rect 10680 16249 10714 16283
rect 10748 16249 10782 16283
rect 10816 16249 10850 16283
rect 10884 16249 10918 16283
rect 10952 16249 10986 16283
rect 11020 16249 11054 16283
rect 11088 16249 11122 16283
rect 11156 16249 11190 16283
rect 11224 16249 11258 16283
rect 11292 16249 11326 16283
rect 11360 16249 11394 16283
rect 11428 16249 11462 16283
rect 11496 16249 11530 16283
rect 11564 16249 11598 16283
rect 11632 16249 11666 16283
rect 11700 16249 11734 16283
rect 11768 16249 11802 16283
rect 11836 16249 11870 16283
rect 11904 16249 11938 16283
rect 11972 16249 12006 16283
rect 12040 16249 12074 16283
rect 12108 16249 12142 16283
rect 12176 16249 12210 16283
rect 12244 16249 12278 16283
rect 12312 16249 12346 16283
rect 12380 16249 12414 16283
rect 12448 16249 12482 16283
rect 12516 16249 12550 16283
rect 12584 16249 12618 16283
rect 12652 16249 12686 16283
rect 12720 16249 12754 16283
rect 12788 16249 12822 16283
rect 12856 16249 12890 16283
rect 12924 16249 12958 16283
rect 12992 16249 13026 16283
rect 13060 16249 13094 16283
rect 13128 16249 13162 16283
rect 13196 16249 13230 16283
rect 13264 16249 13298 16283
rect 13332 16249 13366 16283
rect 13400 16249 13434 16283
rect 13468 16249 13502 16283
rect 13536 16249 13570 16283
rect 13604 16249 13638 16283
rect 13672 16249 13706 16283
rect 13740 16249 13774 16283
rect 13808 16249 13842 16283
rect 13876 16249 13910 16283
rect 13944 16249 13978 16283
rect 14012 16249 14046 16283
rect 14080 16249 14114 16283
rect 14148 16249 14182 16283
rect 14216 16249 14250 16283
rect 14284 16249 14318 16283
rect 14352 16249 14386 16283
rect 14420 16262 14454 16296
rect 14492 16262 14526 16296
rect 14564 16262 14598 16296
rect 14636 16262 14670 16296
rect 14708 16262 14742 16296
rect 14780 16262 14814 16296
rect 14852 16262 14886 16296
rect 14924 16262 14958 16296
rect 14996 16262 15030 16296
rect 15068 16262 15102 16296
rect 68 16187 102 16221
rect 139 16187 173 16221
rect 210 16187 244 16221
rect 281 16187 315 16221
rect 352 16187 386 16221
rect 444 16179 478 16213
rect 513 16179 547 16213
rect 582 16179 616 16213
rect 651 16179 685 16213
rect 720 16179 754 16213
rect 789 16179 823 16213
rect 858 16179 892 16213
rect 927 16179 961 16213
rect 996 16179 1030 16213
rect 1065 16179 1099 16213
rect 1134 16179 1168 16213
rect 1203 16179 1237 16213
rect 1272 16179 1306 16213
rect 1341 16179 1375 16213
rect 1410 16179 1444 16213
rect 1479 16179 1513 16213
rect 1548 16179 1582 16213
rect 1617 16179 1651 16213
rect 1686 16179 1720 16213
rect 1755 16179 1789 16213
rect 1824 16179 1858 16213
rect 1893 16179 1927 16213
rect 1962 16179 1996 16213
rect 2031 16179 2065 16213
rect 2100 16179 2134 16213
rect 2169 16179 2203 16213
rect 2238 16179 2272 16213
rect 2307 16179 2341 16213
rect 2376 16179 2410 16213
rect 2445 16179 2479 16213
rect 2514 16179 2548 16213
rect 2583 16179 2617 16213
rect 2652 16179 2686 16213
rect 2721 16179 2755 16213
rect 2790 16179 2824 16213
rect 2859 16179 2893 16213
rect 2928 16179 2962 16213
rect 2996 16179 3030 16213
rect 3064 16179 3098 16213
rect 3132 16179 3166 16213
rect 3200 16179 3234 16213
rect 3268 16179 3302 16213
rect 3336 16179 3370 16213
rect 3404 16179 3438 16213
rect 3472 16179 3506 16213
rect 3540 16179 3574 16213
rect 3608 16179 3642 16213
rect 3676 16179 3710 16213
rect 3744 16179 3778 16213
rect 3812 16179 3846 16213
rect 3880 16179 3914 16213
rect 3948 16179 3982 16213
rect 4016 16179 4050 16213
rect 4084 16179 4118 16213
rect 4152 16179 4186 16213
rect 4220 16179 4254 16213
rect 4288 16179 4322 16213
rect 4356 16179 4390 16213
rect 4424 16179 4458 16213
rect 4492 16179 4526 16213
rect 4560 16179 4594 16213
rect 4628 16179 4662 16213
rect 4696 16179 4730 16213
rect 4764 16179 4798 16213
rect 4832 16179 4866 16213
rect 4900 16179 4934 16213
rect 4968 16179 5002 16213
rect 5036 16179 5070 16213
rect 5104 16179 5138 16213
rect 5172 16179 5206 16213
rect 5240 16179 5274 16213
rect 5308 16179 5342 16213
rect 5376 16179 5410 16213
rect 5444 16179 5478 16213
rect 5512 16179 5546 16213
rect 5580 16179 5614 16213
rect 5648 16179 5682 16213
rect 5716 16179 5750 16213
rect 5784 16179 5818 16213
rect 5852 16179 5886 16213
rect 5920 16179 5954 16213
rect 5988 16179 6022 16213
rect 6056 16179 6090 16213
rect 6124 16179 6158 16213
rect 6192 16179 6226 16213
rect 6260 16179 6294 16213
rect 6328 16179 6362 16213
rect 6396 16179 6430 16213
rect 6464 16179 6498 16213
rect 6532 16179 6566 16213
rect 6600 16179 6634 16213
rect 6668 16179 6702 16213
rect 6736 16179 6770 16213
rect 6804 16179 6838 16213
rect 6872 16179 6906 16213
rect 6940 16179 6974 16213
rect 7008 16179 7042 16213
rect 7076 16179 7110 16213
rect 7144 16179 7178 16213
rect 7212 16179 7246 16213
rect 7280 16179 7314 16213
rect 7348 16179 7382 16213
rect 7416 16179 7450 16213
rect 7484 16179 7518 16213
rect 7552 16179 7586 16213
rect 7620 16179 7654 16213
rect 7688 16179 7722 16213
rect 7756 16179 7790 16213
rect 7824 16179 7858 16213
rect 7892 16179 7926 16213
rect 7960 16179 7994 16213
rect 8028 16179 8062 16213
rect 8096 16179 8130 16213
rect 8164 16179 8198 16213
rect 8232 16179 8266 16213
rect 8300 16179 8334 16213
rect 8368 16179 8402 16213
rect 8436 16179 8470 16213
rect 8504 16179 8538 16213
rect 8572 16179 8606 16213
rect 8640 16179 8674 16213
rect 8708 16179 8742 16213
rect 8776 16179 8810 16213
rect 8844 16179 8878 16213
rect 8912 16179 8946 16213
rect 8980 16179 9014 16213
rect 9048 16179 9082 16213
rect 9116 16179 9150 16213
rect 9184 16179 9218 16213
rect 9252 16179 9286 16213
rect 9320 16179 9354 16213
rect 9388 16179 9422 16213
rect 9456 16179 9490 16213
rect 9524 16179 9558 16213
rect 9592 16179 9626 16213
rect 9660 16179 9694 16213
rect 9728 16179 9762 16213
rect 9796 16179 9830 16213
rect 9864 16179 9898 16213
rect 9932 16179 9966 16213
rect 10000 16179 10034 16213
rect 10068 16179 10102 16213
rect 10136 16179 10170 16213
rect 10204 16179 10238 16213
rect 10272 16179 10306 16213
rect 10340 16179 10374 16213
rect 10408 16179 10442 16213
rect 10476 16179 10510 16213
rect 10544 16179 10578 16213
rect 10612 16179 10646 16213
rect 10680 16179 10714 16213
rect 10748 16179 10782 16213
rect 10816 16179 10850 16213
rect 10884 16179 10918 16213
rect 10952 16179 10986 16213
rect 11020 16179 11054 16213
rect 11088 16179 11122 16213
rect 11156 16179 11190 16213
rect 11224 16179 11258 16213
rect 11292 16179 11326 16213
rect 11360 16179 11394 16213
rect 11428 16179 11462 16213
rect 11496 16179 11530 16213
rect 11564 16179 11598 16213
rect 11632 16179 11666 16213
rect 11700 16179 11734 16213
rect 11768 16179 11802 16213
rect 11836 16179 11870 16213
rect 11904 16179 11938 16213
rect 11972 16179 12006 16213
rect 12040 16179 12074 16213
rect 12108 16179 12142 16213
rect 12176 16179 12210 16213
rect 12244 16179 12278 16213
rect 12312 16179 12346 16213
rect 12380 16179 12414 16213
rect 12448 16179 12482 16213
rect 12516 16179 12550 16213
rect 12584 16179 12618 16213
rect 12652 16179 12686 16213
rect 12720 16179 12754 16213
rect 12788 16179 12822 16213
rect 12856 16179 12890 16213
rect 12924 16179 12958 16213
rect 12992 16179 13026 16213
rect 13060 16179 13094 16213
rect 13128 16179 13162 16213
rect 13196 16179 13230 16213
rect 13264 16179 13298 16213
rect 13332 16179 13366 16213
rect 13400 16179 13434 16213
rect 13468 16179 13502 16213
rect 13536 16179 13570 16213
rect 13604 16179 13638 16213
rect 13672 16179 13706 16213
rect 13740 16179 13774 16213
rect 13808 16179 13842 16213
rect 13876 16179 13910 16213
rect 13944 16179 13978 16213
rect 14012 16179 14046 16213
rect 14080 16179 14114 16213
rect 14148 16179 14182 16213
rect 14216 16179 14250 16213
rect 14284 16179 14318 16213
rect 14352 16179 14386 16213
rect 14420 16193 14454 16227
rect 14492 16193 14526 16227
rect 14564 16193 14598 16227
rect 14636 16193 14670 16227
rect 14708 16193 14742 16227
rect 14780 16193 14814 16227
rect 14852 16193 14886 16227
rect 14924 16193 14958 16227
rect 14996 16193 15030 16227
rect 15068 16193 15102 16227
rect 68 16119 102 16153
rect 139 16119 173 16153
rect 210 16119 244 16153
rect 281 16119 315 16153
rect 352 16119 386 16153
rect 444 16109 478 16143
rect 513 16109 547 16143
rect 582 16109 616 16143
rect 651 16109 685 16143
rect 720 16109 754 16143
rect 789 16109 823 16143
rect 858 16109 892 16143
rect 927 16109 961 16143
rect 996 16109 1030 16143
rect 1065 16109 1099 16143
rect 1134 16109 1168 16143
rect 1203 16109 1237 16143
rect 1272 16109 1306 16143
rect 1341 16109 1375 16143
rect 1410 16109 1444 16143
rect 1479 16109 1513 16143
rect 1548 16109 1582 16143
rect 1617 16109 1651 16143
rect 1686 16109 1720 16143
rect 1755 16109 1789 16143
rect 1824 16109 1858 16143
rect 1893 16109 1927 16143
rect 1962 16109 1996 16143
rect 2031 16109 2065 16143
rect 2100 16109 2134 16143
rect 2169 16109 2203 16143
rect 2238 16109 2272 16143
rect 2307 16109 2341 16143
rect 2376 16109 2410 16143
rect 2445 16109 2479 16143
rect 2514 16109 2548 16143
rect 2583 16109 2617 16143
rect 2652 16109 2686 16143
rect 2721 16109 2755 16143
rect 2790 16109 2824 16143
rect 2859 16109 2893 16143
rect 2928 16109 2962 16143
rect 2996 16109 3030 16143
rect 3064 16109 3098 16143
rect 3132 16109 3166 16143
rect 3200 16109 3234 16143
rect 3268 16109 3302 16143
rect 3336 16109 3370 16143
rect 3404 16109 3438 16143
rect 3472 16109 3506 16143
rect 3540 16109 3574 16143
rect 3608 16109 3642 16143
rect 3676 16109 3710 16143
rect 3744 16109 3778 16143
rect 3812 16109 3846 16143
rect 3880 16109 3914 16143
rect 3948 16109 3982 16143
rect 4016 16109 4050 16143
rect 4084 16109 4118 16143
rect 4152 16109 4186 16143
rect 4220 16109 4254 16143
rect 4288 16109 4322 16143
rect 4356 16109 4390 16143
rect 4424 16109 4458 16143
rect 4492 16109 4526 16143
rect 4560 16109 4594 16143
rect 4628 16109 4662 16143
rect 4696 16109 4730 16143
rect 4764 16109 4798 16143
rect 4832 16109 4866 16143
rect 4900 16109 4934 16143
rect 4968 16109 5002 16143
rect 5036 16109 5070 16143
rect 5104 16109 5138 16143
rect 5172 16109 5206 16143
rect 5240 16109 5274 16143
rect 5308 16109 5342 16143
rect 5376 16109 5410 16143
rect 5444 16109 5478 16143
rect 5512 16109 5546 16143
rect 5580 16109 5614 16143
rect 5648 16109 5682 16143
rect 5716 16109 5750 16143
rect 5784 16109 5818 16143
rect 5852 16109 5886 16143
rect 5920 16109 5954 16143
rect 5988 16109 6022 16143
rect 6056 16109 6090 16143
rect 6124 16109 6158 16143
rect 6192 16109 6226 16143
rect 6260 16109 6294 16143
rect 6328 16109 6362 16143
rect 6396 16109 6430 16143
rect 6464 16109 6498 16143
rect 6532 16109 6566 16143
rect 6600 16109 6634 16143
rect 6668 16109 6702 16143
rect 6736 16109 6770 16143
rect 6804 16109 6838 16143
rect 6872 16109 6906 16143
rect 6940 16109 6974 16143
rect 7008 16109 7042 16143
rect 7076 16109 7110 16143
rect 7144 16109 7178 16143
rect 7212 16109 7246 16143
rect 7280 16109 7314 16143
rect 7348 16109 7382 16143
rect 7416 16109 7450 16143
rect 7484 16109 7518 16143
rect 7552 16109 7586 16143
rect 7620 16109 7654 16143
rect 7688 16109 7722 16143
rect 7756 16109 7790 16143
rect 7824 16109 7858 16143
rect 7892 16109 7926 16143
rect 7960 16109 7994 16143
rect 8028 16109 8062 16143
rect 8096 16109 8130 16143
rect 8164 16109 8198 16143
rect 8232 16109 8266 16143
rect 8300 16109 8334 16143
rect 8368 16109 8402 16143
rect 8436 16109 8470 16143
rect 8504 16109 8538 16143
rect 8572 16109 8606 16143
rect 8640 16109 8674 16143
rect 8708 16109 8742 16143
rect 8776 16109 8810 16143
rect 8844 16109 8878 16143
rect 8912 16109 8946 16143
rect 8980 16109 9014 16143
rect 9048 16109 9082 16143
rect 9116 16109 9150 16143
rect 9184 16109 9218 16143
rect 9252 16109 9286 16143
rect 9320 16109 9354 16143
rect 9388 16109 9422 16143
rect 9456 16109 9490 16143
rect 9524 16109 9558 16143
rect 9592 16109 9626 16143
rect 9660 16109 9694 16143
rect 9728 16109 9762 16143
rect 9796 16109 9830 16143
rect 9864 16109 9898 16143
rect 9932 16109 9966 16143
rect 10000 16109 10034 16143
rect 10068 16109 10102 16143
rect 10136 16109 10170 16143
rect 10204 16109 10238 16143
rect 10272 16109 10306 16143
rect 10340 16109 10374 16143
rect 10408 16109 10442 16143
rect 10476 16109 10510 16143
rect 10544 16109 10578 16143
rect 10612 16109 10646 16143
rect 10680 16109 10714 16143
rect 10748 16109 10782 16143
rect 10816 16109 10850 16143
rect 10884 16109 10918 16143
rect 10952 16109 10986 16143
rect 11020 16109 11054 16143
rect 11088 16109 11122 16143
rect 11156 16109 11190 16143
rect 11224 16109 11258 16143
rect 11292 16109 11326 16143
rect 11360 16109 11394 16143
rect 11428 16109 11462 16143
rect 11496 16109 11530 16143
rect 11564 16109 11598 16143
rect 11632 16109 11666 16143
rect 11700 16109 11734 16143
rect 11768 16109 11802 16143
rect 11836 16109 11870 16143
rect 11904 16109 11938 16143
rect 11972 16109 12006 16143
rect 12040 16109 12074 16143
rect 12108 16109 12142 16143
rect 12176 16109 12210 16143
rect 12244 16109 12278 16143
rect 12312 16109 12346 16143
rect 12380 16109 12414 16143
rect 12448 16109 12482 16143
rect 12516 16109 12550 16143
rect 12584 16109 12618 16143
rect 12652 16109 12686 16143
rect 12720 16109 12754 16143
rect 12788 16109 12822 16143
rect 12856 16109 12890 16143
rect 12924 16109 12958 16143
rect 12992 16109 13026 16143
rect 13060 16109 13094 16143
rect 13128 16109 13162 16143
rect 13196 16109 13230 16143
rect 13264 16109 13298 16143
rect 13332 16109 13366 16143
rect 13400 16109 13434 16143
rect 13468 16109 13502 16143
rect 13536 16109 13570 16143
rect 13604 16109 13638 16143
rect 13672 16109 13706 16143
rect 13740 16109 13774 16143
rect 13808 16109 13842 16143
rect 13876 16109 13910 16143
rect 13944 16109 13978 16143
rect 14012 16109 14046 16143
rect 14080 16109 14114 16143
rect 14148 16109 14182 16143
rect 14216 16109 14250 16143
rect 14284 16109 14318 16143
rect 14352 16109 14386 16143
rect 14420 16124 14454 16158
rect 14492 16124 14526 16158
rect 14564 16124 14598 16158
rect 14636 16124 14670 16158
rect 14708 16124 14742 16158
rect 14780 16124 14814 16158
rect 14852 16124 14886 16158
rect 14924 16124 14958 16158
rect 14996 16124 15030 16158
rect 15068 16124 15102 16158
rect 68 16051 102 16085
rect 139 16051 173 16085
rect 210 16051 244 16085
rect 281 16051 315 16085
rect 352 16051 386 16085
rect 444 16039 478 16073
rect 513 16039 547 16073
rect 582 16039 616 16073
rect 651 16039 685 16073
rect 720 16039 754 16073
rect 789 16039 823 16073
rect 858 16039 892 16073
rect 927 16039 961 16073
rect 996 16039 1030 16073
rect 1065 16039 1099 16073
rect 1134 16039 1168 16073
rect 1203 16039 1237 16073
rect 1272 16039 1306 16073
rect 1341 16039 1375 16073
rect 1410 16039 1444 16073
rect 1479 16039 1513 16073
rect 1548 16039 1582 16073
rect 1617 16039 1651 16073
rect 1686 16039 1720 16073
rect 1755 16039 1789 16073
rect 1824 16039 1858 16073
rect 1893 16039 1927 16073
rect 1962 16039 1996 16073
rect 2031 16039 2065 16073
rect 2100 16039 2134 16073
rect 2169 16039 2203 16073
rect 2238 16039 2272 16073
rect 2307 16039 2341 16073
rect 2376 16039 2410 16073
rect 2445 16039 2479 16073
rect 2514 16039 2548 16073
rect 2583 16039 2617 16073
rect 2652 16039 2686 16073
rect 2721 16039 2755 16073
rect 2790 16039 2824 16073
rect 2859 16039 2893 16073
rect 2928 16039 2962 16073
rect 2996 16039 3030 16073
rect 3064 16039 3098 16073
rect 3132 16039 3166 16073
rect 3200 16039 3234 16073
rect 3268 16039 3302 16073
rect 3336 16039 3370 16073
rect 3404 16039 3438 16073
rect 3472 16039 3506 16073
rect 3540 16039 3574 16073
rect 3608 16039 3642 16073
rect 3676 16039 3710 16073
rect 3744 16039 3778 16073
rect 3812 16039 3846 16073
rect 3880 16039 3914 16073
rect 3948 16039 3982 16073
rect 4016 16039 4050 16073
rect 4084 16039 4118 16073
rect 4152 16039 4186 16073
rect 4220 16039 4254 16073
rect 4288 16039 4322 16073
rect 4356 16039 4390 16073
rect 4424 16039 4458 16073
rect 4492 16039 4526 16073
rect 4560 16039 4594 16073
rect 4628 16039 4662 16073
rect 4696 16039 4730 16073
rect 4764 16039 4798 16073
rect 4832 16039 4866 16073
rect 4900 16039 4934 16073
rect 4968 16039 5002 16073
rect 5036 16039 5070 16073
rect 5104 16039 5138 16073
rect 5172 16039 5206 16073
rect 5240 16039 5274 16073
rect 5308 16039 5342 16073
rect 5376 16039 5410 16073
rect 5444 16039 5478 16073
rect 5512 16039 5546 16073
rect 5580 16039 5614 16073
rect 5648 16039 5682 16073
rect 5716 16039 5750 16073
rect 5784 16039 5818 16073
rect 5852 16039 5886 16073
rect 5920 16039 5954 16073
rect 5988 16039 6022 16073
rect 6056 16039 6090 16073
rect 6124 16039 6158 16073
rect 6192 16039 6226 16073
rect 6260 16039 6294 16073
rect 6328 16039 6362 16073
rect 6396 16039 6430 16073
rect 6464 16039 6498 16073
rect 6532 16039 6566 16073
rect 6600 16039 6634 16073
rect 6668 16039 6702 16073
rect 6736 16039 6770 16073
rect 6804 16039 6838 16073
rect 6872 16039 6906 16073
rect 6940 16039 6974 16073
rect 7008 16039 7042 16073
rect 7076 16039 7110 16073
rect 7144 16039 7178 16073
rect 7212 16039 7246 16073
rect 7280 16039 7314 16073
rect 7348 16039 7382 16073
rect 7416 16039 7450 16073
rect 7484 16039 7518 16073
rect 7552 16039 7586 16073
rect 7620 16039 7654 16073
rect 7688 16039 7722 16073
rect 7756 16039 7790 16073
rect 7824 16039 7858 16073
rect 7892 16039 7926 16073
rect 7960 16039 7994 16073
rect 8028 16039 8062 16073
rect 8096 16039 8130 16073
rect 8164 16039 8198 16073
rect 8232 16039 8266 16073
rect 8300 16039 8334 16073
rect 8368 16039 8402 16073
rect 8436 16039 8470 16073
rect 8504 16039 8538 16073
rect 8572 16039 8606 16073
rect 8640 16039 8674 16073
rect 8708 16039 8742 16073
rect 8776 16039 8810 16073
rect 8844 16039 8878 16073
rect 8912 16039 8946 16073
rect 8980 16039 9014 16073
rect 9048 16039 9082 16073
rect 9116 16039 9150 16073
rect 9184 16039 9218 16073
rect 9252 16039 9286 16073
rect 9320 16039 9354 16073
rect 9388 16039 9422 16073
rect 9456 16039 9490 16073
rect 9524 16039 9558 16073
rect 9592 16039 9626 16073
rect 9660 16039 9694 16073
rect 9728 16039 9762 16073
rect 9796 16039 9830 16073
rect 9864 16039 9898 16073
rect 9932 16039 9966 16073
rect 10000 16039 10034 16073
rect 10068 16039 10102 16073
rect 10136 16039 10170 16073
rect 10204 16039 10238 16073
rect 10272 16039 10306 16073
rect 10340 16039 10374 16073
rect 10408 16039 10442 16073
rect 10476 16039 10510 16073
rect 10544 16039 10578 16073
rect 10612 16039 10646 16073
rect 10680 16039 10714 16073
rect 10748 16039 10782 16073
rect 10816 16039 10850 16073
rect 10884 16039 10918 16073
rect 10952 16039 10986 16073
rect 11020 16039 11054 16073
rect 11088 16039 11122 16073
rect 11156 16039 11190 16073
rect 11224 16039 11258 16073
rect 11292 16039 11326 16073
rect 11360 16039 11394 16073
rect 11428 16039 11462 16073
rect 11496 16039 11530 16073
rect 11564 16039 11598 16073
rect 11632 16039 11666 16073
rect 11700 16039 11734 16073
rect 11768 16039 11802 16073
rect 11836 16039 11870 16073
rect 11904 16039 11938 16073
rect 11972 16039 12006 16073
rect 12040 16039 12074 16073
rect 12108 16039 12142 16073
rect 12176 16039 12210 16073
rect 12244 16039 12278 16073
rect 12312 16039 12346 16073
rect 12380 16039 12414 16073
rect 12448 16039 12482 16073
rect 12516 16039 12550 16073
rect 12584 16039 12618 16073
rect 12652 16039 12686 16073
rect 12720 16039 12754 16073
rect 12788 16039 12822 16073
rect 12856 16039 12890 16073
rect 12924 16039 12958 16073
rect 12992 16039 13026 16073
rect 13060 16039 13094 16073
rect 13128 16039 13162 16073
rect 13196 16039 13230 16073
rect 13264 16039 13298 16073
rect 13332 16039 13366 16073
rect 13400 16039 13434 16073
rect 13468 16039 13502 16073
rect 13536 16039 13570 16073
rect 13604 16039 13638 16073
rect 13672 16039 13706 16073
rect 13740 16039 13774 16073
rect 13808 16039 13842 16073
rect 13876 16039 13910 16073
rect 13944 16039 13978 16073
rect 14012 16039 14046 16073
rect 14080 16039 14114 16073
rect 14148 16039 14182 16073
rect 14216 16039 14250 16073
rect 14284 16039 14318 16073
rect 14352 16039 14386 16073
rect 14420 16055 14454 16089
rect 14492 16055 14526 16089
rect 14564 16055 14598 16089
rect 14636 16055 14670 16089
rect 14708 16055 14742 16089
rect 14780 16055 14814 16089
rect 14852 16055 14886 16089
rect 14924 16055 14958 16089
rect 14996 16055 15030 16089
rect 15068 16055 15102 16089
rect 68 15983 102 16017
rect 139 15983 173 16017
rect 210 15983 244 16017
rect 281 15983 315 16017
rect 352 15983 386 16017
rect 444 15969 478 16003
rect 513 15969 547 16003
rect 582 15969 616 16003
rect 651 15969 685 16003
rect 720 15969 754 16003
rect 789 15969 823 16003
rect 858 15969 892 16003
rect 927 15969 961 16003
rect 996 15969 1030 16003
rect 1065 15969 1099 16003
rect 1134 15969 1168 16003
rect 1203 15969 1237 16003
rect 1272 15969 1306 16003
rect 1341 15969 1375 16003
rect 1410 15969 1444 16003
rect 1479 15969 1513 16003
rect 1548 15969 1582 16003
rect 1617 15969 1651 16003
rect 1686 15969 1720 16003
rect 1755 15969 1789 16003
rect 1824 15969 1858 16003
rect 1893 15969 1927 16003
rect 1962 15969 1996 16003
rect 2031 15969 2065 16003
rect 2100 15969 2134 16003
rect 2169 15969 2203 16003
rect 2238 15969 2272 16003
rect 2307 15969 2341 16003
rect 2376 15969 2410 16003
rect 2445 15969 2479 16003
rect 2514 15969 2548 16003
rect 2583 15969 2617 16003
rect 2652 15969 2686 16003
rect 2721 15969 2755 16003
rect 2790 15969 2824 16003
rect 2859 15969 2893 16003
rect 2928 15969 2962 16003
rect 2996 15969 3030 16003
rect 3064 15969 3098 16003
rect 3132 15969 3166 16003
rect 3200 15969 3234 16003
rect 3268 15969 3302 16003
rect 3336 15969 3370 16003
rect 3404 15969 3438 16003
rect 3472 15969 3506 16003
rect 3540 15969 3574 16003
rect 3608 15969 3642 16003
rect 3676 15969 3710 16003
rect 3744 15969 3778 16003
rect 3812 15969 3846 16003
rect 3880 15969 3914 16003
rect 3948 15969 3982 16003
rect 4016 15969 4050 16003
rect 4084 15969 4118 16003
rect 4152 15969 4186 16003
rect 4220 15969 4254 16003
rect 4288 15969 4322 16003
rect 4356 15969 4390 16003
rect 4424 15969 4458 16003
rect 4492 15969 4526 16003
rect 4560 15969 4594 16003
rect 4628 15969 4662 16003
rect 4696 15969 4730 16003
rect 4764 15969 4798 16003
rect 4832 15969 4866 16003
rect 4900 15969 4934 16003
rect 4968 15969 5002 16003
rect 5036 15969 5070 16003
rect 5104 15969 5138 16003
rect 5172 15969 5206 16003
rect 5240 15969 5274 16003
rect 5308 15969 5342 16003
rect 5376 15969 5410 16003
rect 5444 15969 5478 16003
rect 5512 15969 5546 16003
rect 5580 15969 5614 16003
rect 5648 15969 5682 16003
rect 5716 15969 5750 16003
rect 5784 15969 5818 16003
rect 5852 15969 5886 16003
rect 5920 15969 5954 16003
rect 5988 15969 6022 16003
rect 6056 15969 6090 16003
rect 6124 15969 6158 16003
rect 6192 15969 6226 16003
rect 6260 15969 6294 16003
rect 6328 15969 6362 16003
rect 6396 15969 6430 16003
rect 6464 15969 6498 16003
rect 6532 15969 6566 16003
rect 6600 15969 6634 16003
rect 6668 15969 6702 16003
rect 6736 15969 6770 16003
rect 6804 15969 6838 16003
rect 6872 15969 6906 16003
rect 6940 15969 6974 16003
rect 7008 15969 7042 16003
rect 7076 15969 7110 16003
rect 7144 15969 7178 16003
rect 7212 15969 7246 16003
rect 7280 15969 7314 16003
rect 7348 15969 7382 16003
rect 7416 15969 7450 16003
rect 7484 15969 7518 16003
rect 7552 15969 7586 16003
rect 7620 15969 7654 16003
rect 7688 15969 7722 16003
rect 7756 15969 7790 16003
rect 7824 15969 7858 16003
rect 7892 15969 7926 16003
rect 7960 15969 7994 16003
rect 8028 15969 8062 16003
rect 8096 15969 8130 16003
rect 8164 15969 8198 16003
rect 8232 15969 8266 16003
rect 8300 15969 8334 16003
rect 8368 15969 8402 16003
rect 8436 15969 8470 16003
rect 8504 15969 8538 16003
rect 8572 15969 8606 16003
rect 8640 15969 8674 16003
rect 8708 15969 8742 16003
rect 8776 15969 8810 16003
rect 8844 15969 8878 16003
rect 8912 15969 8946 16003
rect 8980 15969 9014 16003
rect 9048 15969 9082 16003
rect 9116 15969 9150 16003
rect 9184 15969 9218 16003
rect 9252 15969 9286 16003
rect 9320 15969 9354 16003
rect 9388 15969 9422 16003
rect 9456 15969 9490 16003
rect 9524 15969 9558 16003
rect 9592 15969 9626 16003
rect 9660 15969 9694 16003
rect 9728 15969 9762 16003
rect 9796 15969 9830 16003
rect 9864 15969 9898 16003
rect 9932 15969 9966 16003
rect 10000 15969 10034 16003
rect 10068 15969 10102 16003
rect 10136 15969 10170 16003
rect 10204 15969 10238 16003
rect 10272 15969 10306 16003
rect 10340 15969 10374 16003
rect 10408 15969 10442 16003
rect 10476 15969 10510 16003
rect 10544 15969 10578 16003
rect 10612 15969 10646 16003
rect 10680 15969 10714 16003
rect 10748 15969 10782 16003
rect 10816 15969 10850 16003
rect 10884 15969 10918 16003
rect 10952 15969 10986 16003
rect 11020 15969 11054 16003
rect 11088 15969 11122 16003
rect 11156 15969 11190 16003
rect 11224 15969 11258 16003
rect 11292 15969 11326 16003
rect 11360 15969 11394 16003
rect 11428 15969 11462 16003
rect 11496 15969 11530 16003
rect 11564 15969 11598 16003
rect 11632 15969 11666 16003
rect 11700 15969 11734 16003
rect 11768 15969 11802 16003
rect 11836 15969 11870 16003
rect 11904 15969 11938 16003
rect 11972 15969 12006 16003
rect 12040 15969 12074 16003
rect 12108 15969 12142 16003
rect 12176 15969 12210 16003
rect 12244 15969 12278 16003
rect 12312 15969 12346 16003
rect 12380 15969 12414 16003
rect 12448 15969 12482 16003
rect 12516 15969 12550 16003
rect 12584 15969 12618 16003
rect 12652 15969 12686 16003
rect 12720 15969 12754 16003
rect 12788 15969 12822 16003
rect 12856 15969 12890 16003
rect 12924 15969 12958 16003
rect 12992 15969 13026 16003
rect 13060 15969 13094 16003
rect 13128 15969 13162 16003
rect 13196 15969 13230 16003
rect 13264 15969 13298 16003
rect 13332 15969 13366 16003
rect 13400 15969 13434 16003
rect 13468 15969 13502 16003
rect 13536 15969 13570 16003
rect 13604 15969 13638 16003
rect 13672 15969 13706 16003
rect 13740 15969 13774 16003
rect 13808 15969 13842 16003
rect 13876 15969 13910 16003
rect 13944 15969 13978 16003
rect 14012 15969 14046 16003
rect 14080 15969 14114 16003
rect 14148 15969 14182 16003
rect 14216 15969 14250 16003
rect 14284 15969 14318 16003
rect 14352 15969 14386 16003
rect 14420 15986 14454 16020
rect 14492 15986 14526 16020
rect 14564 15986 14598 16020
rect 14636 15986 14670 16020
rect 14708 15986 14742 16020
rect 14780 15986 14814 16020
rect 14852 15986 14886 16020
rect 14924 15986 14958 16020
rect 14996 15986 15030 16020
rect 15068 15986 15102 16020
rect 68 15915 102 15949
rect 139 15915 173 15949
rect 210 15915 244 15949
rect 281 15915 315 15949
rect 352 15915 386 15949
rect 444 15899 478 15933
rect 513 15899 547 15933
rect 582 15899 616 15933
rect 651 15899 685 15933
rect 720 15899 754 15933
rect 789 15899 823 15933
rect 858 15899 892 15933
rect 927 15899 961 15933
rect 996 15899 1030 15933
rect 1065 15899 1099 15933
rect 1134 15899 1168 15933
rect 1203 15899 1237 15933
rect 1272 15899 1306 15933
rect 1341 15899 1375 15933
rect 1410 15899 1444 15933
rect 1479 15899 1513 15933
rect 1548 15899 1582 15933
rect 1617 15899 1651 15933
rect 1686 15899 1720 15933
rect 1755 15899 1789 15933
rect 1824 15899 1858 15933
rect 1893 15899 1927 15933
rect 1962 15899 1996 15933
rect 2031 15899 2065 15933
rect 2100 15899 2134 15933
rect 2169 15899 2203 15933
rect 2238 15899 2272 15933
rect 2307 15899 2341 15933
rect 2376 15899 2410 15933
rect 2445 15899 2479 15933
rect 2514 15899 2548 15933
rect 2583 15899 2617 15933
rect 2652 15899 2686 15933
rect 2721 15899 2755 15933
rect 2790 15899 2824 15933
rect 2859 15899 2893 15933
rect 2928 15899 2962 15933
rect 2996 15899 3030 15933
rect 3064 15899 3098 15933
rect 3132 15899 3166 15933
rect 3200 15899 3234 15933
rect 3268 15899 3302 15933
rect 3336 15899 3370 15933
rect 3404 15899 3438 15933
rect 3472 15899 3506 15933
rect 3540 15899 3574 15933
rect 3608 15899 3642 15933
rect 3676 15899 3710 15933
rect 3744 15899 3778 15933
rect 3812 15899 3846 15933
rect 3880 15899 3914 15933
rect 3948 15899 3982 15933
rect 4016 15899 4050 15933
rect 4084 15899 4118 15933
rect 4152 15899 4186 15933
rect 4220 15899 4254 15933
rect 4288 15899 4322 15933
rect 4356 15899 4390 15933
rect 4424 15899 4458 15933
rect 4492 15899 4526 15933
rect 4560 15899 4594 15933
rect 4628 15899 4662 15933
rect 4696 15899 4730 15933
rect 4764 15899 4798 15933
rect 4832 15899 4866 15933
rect 4900 15899 4934 15933
rect 4968 15899 5002 15933
rect 5036 15899 5070 15933
rect 5104 15899 5138 15933
rect 5172 15899 5206 15933
rect 5240 15899 5274 15933
rect 5308 15899 5342 15933
rect 5376 15899 5410 15933
rect 5444 15899 5478 15933
rect 5512 15899 5546 15933
rect 5580 15899 5614 15933
rect 5648 15899 5682 15933
rect 5716 15899 5750 15933
rect 5784 15899 5818 15933
rect 5852 15899 5886 15933
rect 5920 15899 5954 15933
rect 5988 15899 6022 15933
rect 6056 15899 6090 15933
rect 6124 15899 6158 15933
rect 6192 15899 6226 15933
rect 6260 15899 6294 15933
rect 6328 15899 6362 15933
rect 6396 15899 6430 15933
rect 6464 15899 6498 15933
rect 6532 15899 6566 15933
rect 6600 15899 6634 15933
rect 6668 15899 6702 15933
rect 6736 15899 6770 15933
rect 6804 15899 6838 15933
rect 6872 15899 6906 15933
rect 6940 15899 6974 15933
rect 7008 15899 7042 15933
rect 7076 15899 7110 15933
rect 7144 15899 7178 15933
rect 7212 15899 7246 15933
rect 7280 15899 7314 15933
rect 7348 15899 7382 15933
rect 7416 15899 7450 15933
rect 7484 15899 7518 15933
rect 7552 15899 7586 15933
rect 7620 15899 7654 15933
rect 7688 15899 7722 15933
rect 7756 15899 7790 15933
rect 7824 15899 7858 15933
rect 7892 15899 7926 15933
rect 7960 15899 7994 15933
rect 8028 15899 8062 15933
rect 8096 15899 8130 15933
rect 8164 15899 8198 15933
rect 8232 15899 8266 15933
rect 8300 15899 8334 15933
rect 8368 15899 8402 15933
rect 8436 15899 8470 15933
rect 8504 15899 8538 15933
rect 8572 15899 8606 15933
rect 8640 15899 8674 15933
rect 8708 15899 8742 15933
rect 8776 15899 8810 15933
rect 8844 15899 8878 15933
rect 8912 15899 8946 15933
rect 8980 15899 9014 15933
rect 9048 15899 9082 15933
rect 9116 15899 9150 15933
rect 9184 15899 9218 15933
rect 9252 15899 9286 15933
rect 9320 15899 9354 15933
rect 9388 15899 9422 15933
rect 9456 15899 9490 15933
rect 9524 15899 9558 15933
rect 9592 15899 9626 15933
rect 9660 15899 9694 15933
rect 9728 15899 9762 15933
rect 9796 15899 9830 15933
rect 9864 15899 9898 15933
rect 9932 15899 9966 15933
rect 10000 15899 10034 15933
rect 10068 15899 10102 15933
rect 10136 15899 10170 15933
rect 10204 15899 10238 15933
rect 10272 15899 10306 15933
rect 10340 15899 10374 15933
rect 10408 15899 10442 15933
rect 10476 15899 10510 15933
rect 10544 15899 10578 15933
rect 10612 15899 10646 15933
rect 10680 15899 10714 15933
rect 10748 15899 10782 15933
rect 10816 15899 10850 15933
rect 10884 15899 10918 15933
rect 10952 15899 10986 15933
rect 11020 15899 11054 15933
rect 11088 15899 11122 15933
rect 11156 15899 11190 15933
rect 11224 15899 11258 15933
rect 11292 15899 11326 15933
rect 11360 15899 11394 15933
rect 11428 15899 11462 15933
rect 11496 15899 11530 15933
rect 11564 15899 11598 15933
rect 11632 15899 11666 15933
rect 11700 15899 11734 15933
rect 11768 15899 11802 15933
rect 11836 15899 11870 15933
rect 11904 15899 11938 15933
rect 11972 15899 12006 15933
rect 12040 15899 12074 15933
rect 12108 15899 12142 15933
rect 12176 15899 12210 15933
rect 12244 15899 12278 15933
rect 12312 15899 12346 15933
rect 12380 15899 12414 15933
rect 12448 15899 12482 15933
rect 12516 15899 12550 15933
rect 12584 15899 12618 15933
rect 12652 15899 12686 15933
rect 12720 15899 12754 15933
rect 12788 15899 12822 15933
rect 12856 15899 12890 15933
rect 12924 15899 12958 15933
rect 12992 15899 13026 15933
rect 13060 15899 13094 15933
rect 13128 15899 13162 15933
rect 13196 15899 13230 15933
rect 13264 15899 13298 15933
rect 13332 15899 13366 15933
rect 13400 15899 13434 15933
rect 13468 15899 13502 15933
rect 13536 15899 13570 15933
rect 13604 15899 13638 15933
rect 13672 15899 13706 15933
rect 13740 15899 13774 15933
rect 13808 15899 13842 15933
rect 13876 15899 13910 15933
rect 13944 15899 13978 15933
rect 14012 15899 14046 15933
rect 14080 15899 14114 15933
rect 14148 15899 14182 15933
rect 14216 15899 14250 15933
rect 14284 15899 14318 15933
rect 14352 15899 14386 15933
rect 14420 15917 14454 15951
rect 14492 15917 14526 15951
rect 14564 15917 14598 15951
rect 14636 15917 14670 15951
rect 14708 15917 14742 15951
rect 14780 15917 14814 15951
rect 14852 15917 14886 15951
rect 14924 15917 14958 15951
rect 14996 15917 15030 15951
rect 15068 15917 15102 15951
rect 68 15846 102 15880
rect 139 15846 173 15880
rect 210 15846 244 15880
rect 281 15846 315 15880
rect 352 15846 386 15880
rect 444 15829 478 15863
rect 513 15829 547 15863
rect 582 15829 616 15863
rect 651 15829 685 15863
rect 720 15829 754 15863
rect 789 15829 823 15863
rect 858 15829 892 15863
rect 927 15829 961 15863
rect 996 15829 1030 15863
rect 1065 15829 1099 15863
rect 1134 15829 1168 15863
rect 1203 15829 1237 15863
rect 1272 15829 1306 15863
rect 1341 15829 1375 15863
rect 1410 15829 1444 15863
rect 1479 15829 1513 15863
rect 1548 15829 1582 15863
rect 1617 15829 1651 15863
rect 1686 15829 1720 15863
rect 1755 15829 1789 15863
rect 1824 15829 1858 15863
rect 1893 15829 1927 15863
rect 1962 15829 1996 15863
rect 2031 15829 2065 15863
rect 2100 15829 2134 15863
rect 2169 15829 2203 15863
rect 2238 15829 2272 15863
rect 2307 15829 2341 15863
rect 2376 15829 2410 15863
rect 2445 15829 2479 15863
rect 2514 15829 2548 15863
rect 2583 15829 2617 15863
rect 2652 15829 2686 15863
rect 2721 15829 2755 15863
rect 2790 15829 2824 15863
rect 2859 15829 2893 15863
rect 2928 15829 2962 15863
rect 2996 15829 3030 15863
rect 3064 15829 3098 15863
rect 3132 15829 3166 15863
rect 3200 15829 3234 15863
rect 3268 15829 3302 15863
rect 3336 15829 3370 15863
rect 3404 15829 3438 15863
rect 3472 15829 3506 15863
rect 3540 15829 3574 15863
rect 3608 15829 3642 15863
rect 3676 15829 3710 15863
rect 3744 15829 3778 15863
rect 3812 15829 3846 15863
rect 3880 15829 3914 15863
rect 3948 15829 3982 15863
rect 4016 15829 4050 15863
rect 4084 15829 4118 15863
rect 4152 15829 4186 15863
rect 4220 15829 4254 15863
rect 4288 15829 4322 15863
rect 4356 15829 4390 15863
rect 4424 15829 4458 15863
rect 4492 15829 4526 15863
rect 4560 15829 4594 15863
rect 4628 15829 4662 15863
rect 4696 15829 4730 15863
rect 4764 15829 4798 15863
rect 4832 15829 4866 15863
rect 4900 15829 4934 15863
rect 4968 15829 5002 15863
rect 5036 15829 5070 15863
rect 5104 15829 5138 15863
rect 5172 15829 5206 15863
rect 5240 15829 5274 15863
rect 5308 15829 5342 15863
rect 5376 15829 5410 15863
rect 5444 15829 5478 15863
rect 5512 15829 5546 15863
rect 5580 15829 5614 15863
rect 5648 15829 5682 15863
rect 5716 15829 5750 15863
rect 5784 15829 5818 15863
rect 5852 15829 5886 15863
rect 5920 15829 5954 15863
rect 5988 15829 6022 15863
rect 6056 15829 6090 15863
rect 6124 15829 6158 15863
rect 6192 15829 6226 15863
rect 6260 15829 6294 15863
rect 6328 15829 6362 15863
rect 6396 15829 6430 15863
rect 6464 15829 6498 15863
rect 6532 15829 6566 15863
rect 6600 15829 6634 15863
rect 6668 15829 6702 15863
rect 6736 15829 6770 15863
rect 6804 15829 6838 15863
rect 6872 15829 6906 15863
rect 6940 15829 6974 15863
rect 7008 15829 7042 15863
rect 7076 15829 7110 15863
rect 7144 15829 7178 15863
rect 7212 15829 7246 15863
rect 7280 15829 7314 15863
rect 7348 15829 7382 15863
rect 7416 15829 7450 15863
rect 7484 15829 7518 15863
rect 7552 15829 7586 15863
rect 7620 15829 7654 15863
rect 7688 15829 7722 15863
rect 7756 15829 7790 15863
rect 7824 15829 7858 15863
rect 7892 15829 7926 15863
rect 7960 15829 7994 15863
rect 8028 15829 8062 15863
rect 8096 15829 8130 15863
rect 8164 15829 8198 15863
rect 8232 15829 8266 15863
rect 8300 15829 8334 15863
rect 8368 15829 8402 15863
rect 8436 15829 8470 15863
rect 8504 15829 8538 15863
rect 8572 15829 8606 15863
rect 8640 15829 8674 15863
rect 8708 15829 8742 15863
rect 8776 15829 8810 15863
rect 8844 15829 8878 15863
rect 8912 15829 8946 15863
rect 8980 15829 9014 15863
rect 9048 15829 9082 15863
rect 9116 15829 9150 15863
rect 9184 15829 9218 15863
rect 9252 15829 9286 15863
rect 9320 15829 9354 15863
rect 9388 15829 9422 15863
rect 9456 15829 9490 15863
rect 9524 15829 9558 15863
rect 9592 15829 9626 15863
rect 9660 15829 9694 15863
rect 9728 15829 9762 15863
rect 9796 15829 9830 15863
rect 9864 15829 9898 15863
rect 9932 15829 9966 15863
rect 10000 15829 10034 15863
rect 10068 15829 10102 15863
rect 10136 15829 10170 15863
rect 10204 15829 10238 15863
rect 10272 15829 10306 15863
rect 10340 15829 10374 15863
rect 10408 15829 10442 15863
rect 10476 15829 10510 15863
rect 10544 15829 10578 15863
rect 10612 15829 10646 15863
rect 10680 15829 10714 15863
rect 10748 15829 10782 15863
rect 10816 15829 10850 15863
rect 10884 15829 10918 15863
rect 10952 15829 10986 15863
rect 11020 15829 11054 15863
rect 11088 15829 11122 15863
rect 11156 15829 11190 15863
rect 11224 15829 11258 15863
rect 11292 15829 11326 15863
rect 11360 15829 11394 15863
rect 11428 15829 11462 15863
rect 11496 15829 11530 15863
rect 11564 15829 11598 15863
rect 11632 15829 11666 15863
rect 11700 15829 11734 15863
rect 11768 15829 11802 15863
rect 11836 15829 11870 15863
rect 11904 15829 11938 15863
rect 11972 15829 12006 15863
rect 12040 15829 12074 15863
rect 12108 15829 12142 15863
rect 12176 15829 12210 15863
rect 12244 15829 12278 15863
rect 12312 15829 12346 15863
rect 12380 15829 12414 15863
rect 12448 15829 12482 15863
rect 12516 15829 12550 15863
rect 12584 15829 12618 15863
rect 12652 15829 12686 15863
rect 12720 15829 12754 15863
rect 12788 15829 12822 15863
rect 12856 15829 12890 15863
rect 12924 15829 12958 15863
rect 12992 15829 13026 15863
rect 13060 15829 13094 15863
rect 13128 15829 13162 15863
rect 13196 15829 13230 15863
rect 13264 15829 13298 15863
rect 13332 15829 13366 15863
rect 13400 15829 13434 15863
rect 13468 15829 13502 15863
rect 13536 15829 13570 15863
rect 13604 15829 13638 15863
rect 13672 15829 13706 15863
rect 13740 15829 13774 15863
rect 13808 15829 13842 15863
rect 13876 15829 13910 15863
rect 13944 15829 13978 15863
rect 14012 15829 14046 15863
rect 14080 15829 14114 15863
rect 14148 15829 14182 15863
rect 14216 15829 14250 15863
rect 14284 15829 14318 15863
rect 14352 15829 14386 15863
rect 14420 15848 14454 15882
rect 14492 15848 14526 15882
rect 14564 15848 14598 15882
rect 14636 15848 14670 15882
rect 14708 15848 14742 15882
rect 14780 15848 14814 15882
rect 14852 15848 14886 15882
rect 14924 15848 14958 15882
rect 14996 15848 15030 15882
rect 15068 15848 15102 15882
rect 68 15777 102 15811
rect 139 15777 173 15811
rect 210 15777 244 15811
rect 281 15777 315 15811
rect 352 15777 386 15811
rect 444 15759 478 15793
rect 513 15759 547 15793
rect 582 15759 616 15793
rect 651 15759 685 15793
rect 720 15759 754 15793
rect 789 15759 823 15793
rect 858 15759 892 15793
rect 927 15759 961 15793
rect 996 15759 1030 15793
rect 1065 15759 1099 15793
rect 1134 15759 1168 15793
rect 1203 15759 1237 15793
rect 1272 15759 1306 15793
rect 1341 15759 1375 15793
rect 1410 15759 1444 15793
rect 1479 15759 1513 15793
rect 1548 15759 1582 15793
rect 1617 15759 1651 15793
rect 1686 15759 1720 15793
rect 1755 15759 1789 15793
rect 1824 15759 1858 15793
rect 1893 15759 1927 15793
rect 1962 15759 1996 15793
rect 2031 15759 2065 15793
rect 2100 15759 2134 15793
rect 2169 15759 2203 15793
rect 2238 15759 2272 15793
rect 2307 15759 2341 15793
rect 2376 15759 2410 15793
rect 2445 15759 2479 15793
rect 2514 15759 2548 15793
rect 2583 15759 2617 15793
rect 2652 15759 2686 15793
rect 2721 15759 2755 15793
rect 2790 15759 2824 15793
rect 2859 15759 2893 15793
rect 2928 15759 2962 15793
rect 2996 15759 3030 15793
rect 3064 15759 3098 15793
rect 3132 15759 3166 15793
rect 3200 15759 3234 15793
rect 3268 15759 3302 15793
rect 3336 15759 3370 15793
rect 3404 15759 3438 15793
rect 3472 15759 3506 15793
rect 3540 15759 3574 15793
rect 3608 15759 3642 15793
rect 3676 15759 3710 15793
rect 3744 15759 3778 15793
rect 3812 15759 3846 15793
rect 3880 15759 3914 15793
rect 3948 15759 3982 15793
rect 4016 15759 4050 15793
rect 4084 15759 4118 15793
rect 4152 15759 4186 15793
rect 4220 15759 4254 15793
rect 4288 15759 4322 15793
rect 4356 15759 4390 15793
rect 4424 15759 4458 15793
rect 4492 15759 4526 15793
rect 4560 15759 4594 15793
rect 4628 15759 4662 15793
rect 4696 15759 4730 15793
rect 4764 15759 4798 15793
rect 4832 15759 4866 15793
rect 4900 15759 4934 15793
rect 4968 15759 5002 15793
rect 5036 15759 5070 15793
rect 5104 15759 5138 15793
rect 5172 15759 5206 15793
rect 5240 15759 5274 15793
rect 5308 15759 5342 15793
rect 5376 15759 5410 15793
rect 5444 15759 5478 15793
rect 5512 15759 5546 15793
rect 5580 15759 5614 15793
rect 5648 15759 5682 15793
rect 5716 15759 5750 15793
rect 5784 15759 5818 15793
rect 5852 15759 5886 15793
rect 5920 15759 5954 15793
rect 5988 15759 6022 15793
rect 6056 15759 6090 15793
rect 6124 15759 6158 15793
rect 6192 15759 6226 15793
rect 6260 15759 6294 15793
rect 6328 15759 6362 15793
rect 6396 15759 6430 15793
rect 6464 15759 6498 15793
rect 6532 15759 6566 15793
rect 6600 15759 6634 15793
rect 6668 15759 6702 15793
rect 6736 15759 6770 15793
rect 6804 15759 6838 15793
rect 6872 15759 6906 15793
rect 6940 15759 6974 15793
rect 7008 15759 7042 15793
rect 7076 15759 7110 15793
rect 7144 15759 7178 15793
rect 7212 15759 7246 15793
rect 7280 15759 7314 15793
rect 7348 15759 7382 15793
rect 7416 15759 7450 15793
rect 7484 15759 7518 15793
rect 7552 15759 7586 15793
rect 7620 15759 7654 15793
rect 7688 15759 7722 15793
rect 7756 15759 7790 15793
rect 7824 15759 7858 15793
rect 7892 15759 7926 15793
rect 7960 15759 7994 15793
rect 8028 15759 8062 15793
rect 8096 15759 8130 15793
rect 8164 15759 8198 15793
rect 8232 15759 8266 15793
rect 8300 15759 8334 15793
rect 8368 15759 8402 15793
rect 8436 15759 8470 15793
rect 8504 15759 8538 15793
rect 8572 15759 8606 15793
rect 8640 15759 8674 15793
rect 8708 15759 8742 15793
rect 8776 15759 8810 15793
rect 8844 15759 8878 15793
rect 8912 15759 8946 15793
rect 8980 15759 9014 15793
rect 9048 15759 9082 15793
rect 9116 15759 9150 15793
rect 9184 15759 9218 15793
rect 9252 15759 9286 15793
rect 9320 15759 9354 15793
rect 9388 15759 9422 15793
rect 9456 15759 9490 15793
rect 9524 15759 9558 15793
rect 9592 15759 9626 15793
rect 9660 15759 9694 15793
rect 9728 15759 9762 15793
rect 9796 15759 9830 15793
rect 9864 15759 9898 15793
rect 9932 15759 9966 15793
rect 10000 15759 10034 15793
rect 10068 15759 10102 15793
rect 10136 15759 10170 15793
rect 10204 15759 10238 15793
rect 10272 15759 10306 15793
rect 10340 15759 10374 15793
rect 10408 15759 10442 15793
rect 10476 15759 10510 15793
rect 10544 15759 10578 15793
rect 10612 15759 10646 15793
rect 10680 15759 10714 15793
rect 10748 15759 10782 15793
rect 10816 15759 10850 15793
rect 10884 15759 10918 15793
rect 10952 15759 10986 15793
rect 11020 15759 11054 15793
rect 11088 15759 11122 15793
rect 11156 15759 11190 15793
rect 11224 15759 11258 15793
rect 11292 15759 11326 15793
rect 11360 15759 11394 15793
rect 11428 15759 11462 15793
rect 11496 15759 11530 15793
rect 11564 15759 11598 15793
rect 11632 15759 11666 15793
rect 11700 15759 11734 15793
rect 11768 15759 11802 15793
rect 11836 15759 11870 15793
rect 11904 15759 11938 15793
rect 11972 15759 12006 15793
rect 12040 15759 12074 15793
rect 12108 15759 12142 15793
rect 12176 15759 12210 15793
rect 12244 15759 12278 15793
rect 12312 15759 12346 15793
rect 12380 15759 12414 15793
rect 12448 15759 12482 15793
rect 12516 15759 12550 15793
rect 12584 15759 12618 15793
rect 12652 15759 12686 15793
rect 12720 15759 12754 15793
rect 12788 15759 12822 15793
rect 12856 15759 12890 15793
rect 12924 15759 12958 15793
rect 12992 15759 13026 15793
rect 13060 15759 13094 15793
rect 13128 15759 13162 15793
rect 13196 15759 13230 15793
rect 13264 15759 13298 15793
rect 13332 15759 13366 15793
rect 13400 15759 13434 15793
rect 13468 15759 13502 15793
rect 13536 15759 13570 15793
rect 13604 15759 13638 15793
rect 13672 15759 13706 15793
rect 13740 15759 13774 15793
rect 13808 15759 13842 15793
rect 13876 15759 13910 15793
rect 13944 15759 13978 15793
rect 14012 15759 14046 15793
rect 14080 15759 14114 15793
rect 14148 15759 14182 15793
rect 14216 15759 14250 15793
rect 14284 15759 14318 15793
rect 14352 15759 14386 15793
rect 14420 15779 14454 15813
rect 14492 15779 14526 15813
rect 14564 15779 14598 15813
rect 14636 15779 14670 15813
rect 14708 15779 14742 15813
rect 14780 15779 14814 15813
rect 14852 15779 14886 15813
rect 14924 15779 14958 15813
rect 14996 15779 15030 15813
rect 15068 15779 15102 15813
rect 68 15708 102 15742
rect 139 15708 173 15742
rect 210 15708 244 15742
rect 281 15708 315 15742
rect 352 15708 386 15742
rect 444 15689 478 15723
rect 513 15689 547 15723
rect 582 15689 616 15723
rect 651 15689 685 15723
rect 720 15689 754 15723
rect 789 15689 823 15723
rect 858 15689 892 15723
rect 927 15689 961 15723
rect 996 15689 1030 15723
rect 1065 15689 1099 15723
rect 1134 15689 1168 15723
rect 1203 15689 1237 15723
rect 1272 15689 1306 15723
rect 1341 15689 1375 15723
rect 1410 15689 1444 15723
rect 1479 15689 1513 15723
rect 1548 15689 1582 15723
rect 1617 15689 1651 15723
rect 1686 15689 1720 15723
rect 1755 15689 1789 15723
rect 1824 15689 1858 15723
rect 1893 15689 1927 15723
rect 1962 15689 1996 15723
rect 2031 15689 2065 15723
rect 2100 15689 2134 15723
rect 2169 15689 2203 15723
rect 2238 15689 2272 15723
rect 2307 15689 2341 15723
rect 2376 15689 2410 15723
rect 2445 15689 2479 15723
rect 2514 15689 2548 15723
rect 2583 15689 2617 15723
rect 2652 15689 2686 15723
rect 2721 15689 2755 15723
rect 2790 15689 2824 15723
rect 2859 15689 2893 15723
rect 2928 15689 2962 15723
rect 2996 15689 3030 15723
rect 3064 15689 3098 15723
rect 3132 15689 3166 15723
rect 3200 15689 3234 15723
rect 3268 15689 3302 15723
rect 3336 15689 3370 15723
rect 3404 15689 3438 15723
rect 3472 15689 3506 15723
rect 3540 15689 3574 15723
rect 3608 15689 3642 15723
rect 3676 15689 3710 15723
rect 3744 15689 3778 15723
rect 3812 15689 3846 15723
rect 3880 15689 3914 15723
rect 3948 15689 3982 15723
rect 4016 15689 4050 15723
rect 4084 15689 4118 15723
rect 4152 15689 4186 15723
rect 4220 15689 4254 15723
rect 4288 15689 4322 15723
rect 4356 15689 4390 15723
rect 4424 15689 4458 15723
rect 4492 15689 4526 15723
rect 4560 15689 4594 15723
rect 4628 15689 4662 15723
rect 4696 15689 4730 15723
rect 4764 15689 4798 15723
rect 4832 15689 4866 15723
rect 4900 15689 4934 15723
rect 4968 15689 5002 15723
rect 5036 15689 5070 15723
rect 5104 15689 5138 15723
rect 5172 15689 5206 15723
rect 5240 15689 5274 15723
rect 5308 15689 5342 15723
rect 5376 15689 5410 15723
rect 5444 15689 5478 15723
rect 5512 15689 5546 15723
rect 5580 15689 5614 15723
rect 5648 15689 5682 15723
rect 5716 15689 5750 15723
rect 5784 15689 5818 15723
rect 5852 15689 5886 15723
rect 5920 15689 5954 15723
rect 5988 15689 6022 15723
rect 6056 15689 6090 15723
rect 6124 15689 6158 15723
rect 6192 15689 6226 15723
rect 6260 15689 6294 15723
rect 6328 15689 6362 15723
rect 6396 15689 6430 15723
rect 6464 15689 6498 15723
rect 6532 15689 6566 15723
rect 6600 15689 6634 15723
rect 6668 15689 6702 15723
rect 6736 15689 6770 15723
rect 6804 15689 6838 15723
rect 6872 15689 6906 15723
rect 6940 15689 6974 15723
rect 7008 15689 7042 15723
rect 7076 15689 7110 15723
rect 7144 15689 7178 15723
rect 7212 15689 7246 15723
rect 7280 15689 7314 15723
rect 7348 15689 7382 15723
rect 7416 15689 7450 15723
rect 7484 15689 7518 15723
rect 7552 15689 7586 15723
rect 7620 15689 7654 15723
rect 7688 15689 7722 15723
rect 7756 15689 7790 15723
rect 7824 15689 7858 15723
rect 7892 15689 7926 15723
rect 7960 15689 7994 15723
rect 8028 15689 8062 15723
rect 8096 15689 8130 15723
rect 8164 15689 8198 15723
rect 8232 15689 8266 15723
rect 8300 15689 8334 15723
rect 8368 15689 8402 15723
rect 8436 15689 8470 15723
rect 8504 15689 8538 15723
rect 8572 15689 8606 15723
rect 8640 15689 8674 15723
rect 8708 15689 8742 15723
rect 8776 15689 8810 15723
rect 8844 15689 8878 15723
rect 8912 15689 8946 15723
rect 8980 15689 9014 15723
rect 9048 15689 9082 15723
rect 9116 15689 9150 15723
rect 9184 15689 9218 15723
rect 9252 15689 9286 15723
rect 9320 15689 9354 15723
rect 9388 15689 9422 15723
rect 9456 15689 9490 15723
rect 9524 15689 9558 15723
rect 9592 15689 9626 15723
rect 9660 15689 9694 15723
rect 9728 15689 9762 15723
rect 9796 15689 9830 15723
rect 9864 15689 9898 15723
rect 9932 15689 9966 15723
rect 10000 15689 10034 15723
rect 10068 15689 10102 15723
rect 10136 15689 10170 15723
rect 10204 15689 10238 15723
rect 10272 15689 10306 15723
rect 10340 15689 10374 15723
rect 10408 15689 10442 15723
rect 10476 15689 10510 15723
rect 10544 15689 10578 15723
rect 10612 15689 10646 15723
rect 10680 15689 10714 15723
rect 10748 15689 10782 15723
rect 10816 15689 10850 15723
rect 10884 15689 10918 15723
rect 10952 15689 10986 15723
rect 11020 15689 11054 15723
rect 11088 15689 11122 15723
rect 11156 15689 11190 15723
rect 11224 15689 11258 15723
rect 11292 15689 11326 15723
rect 11360 15689 11394 15723
rect 11428 15689 11462 15723
rect 11496 15689 11530 15723
rect 11564 15689 11598 15723
rect 11632 15689 11666 15723
rect 11700 15689 11734 15723
rect 11768 15689 11802 15723
rect 11836 15689 11870 15723
rect 11904 15689 11938 15723
rect 11972 15689 12006 15723
rect 12040 15689 12074 15723
rect 12108 15689 12142 15723
rect 12176 15689 12210 15723
rect 12244 15689 12278 15723
rect 12312 15689 12346 15723
rect 12380 15689 12414 15723
rect 12448 15689 12482 15723
rect 12516 15689 12550 15723
rect 12584 15689 12618 15723
rect 12652 15689 12686 15723
rect 12720 15689 12754 15723
rect 12788 15689 12822 15723
rect 12856 15689 12890 15723
rect 12924 15689 12958 15723
rect 12992 15689 13026 15723
rect 13060 15689 13094 15723
rect 13128 15689 13162 15723
rect 13196 15689 13230 15723
rect 13264 15689 13298 15723
rect 13332 15689 13366 15723
rect 13400 15689 13434 15723
rect 13468 15689 13502 15723
rect 13536 15689 13570 15723
rect 13604 15689 13638 15723
rect 13672 15689 13706 15723
rect 13740 15689 13774 15723
rect 13808 15689 13842 15723
rect 13876 15689 13910 15723
rect 13944 15689 13978 15723
rect 14012 15689 14046 15723
rect 14080 15689 14114 15723
rect 14148 15689 14182 15723
rect 14216 15689 14250 15723
rect 14284 15689 14318 15723
rect 14352 15689 14386 15723
rect 14420 15710 14454 15744
rect 14492 15710 14526 15744
rect 14564 15710 14598 15744
rect 14636 15710 14670 15744
rect 14708 15710 14742 15744
rect 14780 15710 14814 15744
rect 14852 15710 14886 15744
rect 14924 15710 14958 15744
rect 14996 15710 15030 15744
rect 15068 15710 15102 15744
rect 68 15639 102 15673
rect 139 15639 173 15673
rect 210 15639 244 15673
rect 281 15639 315 15673
rect 352 15639 386 15673
rect 12660 15617 12694 15651
rect 12730 15617 12764 15651
rect 12800 15617 12834 15651
rect 12869 15617 12903 15651
rect 12938 15617 12972 15651
rect 13007 15617 13041 15651
rect 13076 15617 13110 15651
rect 13145 15617 13179 15651
rect 13214 15617 13248 15651
rect 13283 15617 13317 15651
rect 13352 15617 13386 15651
rect 13421 15617 13455 15651
rect 13490 15617 13524 15651
rect 13559 15617 13593 15651
rect 13628 15617 13662 15651
rect 13697 15617 13731 15651
rect 13766 15617 13800 15651
rect 13835 15617 13869 15651
rect 13904 15617 13938 15651
rect 13973 15617 14007 15651
rect 14042 15617 14076 15651
rect 14111 15617 14145 15651
rect 14180 15617 14214 15651
rect 14249 15617 14283 15651
rect 14318 15617 14352 15651
rect 14420 15641 14454 15675
rect 14492 15641 14526 15675
rect 14564 15641 14598 15675
rect 14636 15641 14670 15675
rect 14708 15641 14742 15675
rect 14780 15641 14814 15675
rect 14852 15641 14886 15675
rect 14924 15641 14958 15675
rect 14996 15641 15030 15675
rect 15068 15641 15102 15675
rect 68 15570 102 15604
rect 139 15570 173 15604
rect 210 15570 244 15604
rect 281 15570 315 15604
rect 352 15570 386 15604
rect 420 15549 454 15583
rect 488 15549 522 15583
rect 594 15573 628 15607
rect 663 15573 697 15607
rect 732 15573 766 15607
rect 801 15573 835 15607
rect 870 15573 904 15607
rect 939 15573 973 15607
rect 1008 15573 1042 15607
rect 1077 15573 1111 15607
rect 1146 15573 1180 15607
rect 1215 15573 1249 15607
rect 1284 15573 1318 15607
rect 1353 15573 1387 15607
rect 1422 15573 1456 15607
rect 1491 15573 1525 15607
rect 1560 15573 1594 15607
rect 1629 15573 1663 15607
rect 1698 15573 1732 15607
rect 1767 15573 1801 15607
rect 1836 15573 1870 15607
rect 1904 15573 1938 15607
rect 1972 15573 2006 15607
rect 2040 15573 2074 15607
rect 2108 15573 2142 15607
rect 2176 15573 2210 15607
rect 2244 15573 2278 15607
rect 2312 15573 2346 15607
rect 2380 15573 2414 15607
rect 2448 15573 2482 15607
rect 2516 15573 2550 15607
rect 2584 15573 2618 15607
rect 2652 15573 2686 15607
rect 2720 15573 2754 15607
rect 2788 15573 2822 15607
rect 2856 15573 2890 15607
rect 2924 15573 2958 15607
rect 2992 15573 3026 15607
rect 3060 15573 3094 15607
rect 3128 15573 3162 15607
rect 3196 15573 3230 15607
rect 3264 15573 3298 15607
rect 3332 15573 3366 15607
rect 3400 15573 3434 15607
rect 3468 15573 3502 15607
rect 3536 15573 3570 15607
rect 3604 15573 3638 15607
rect 3672 15573 3706 15607
rect 3740 15573 3774 15607
rect 3808 15573 3842 15607
rect 3876 15573 3910 15607
rect 3944 15573 3978 15607
rect 4012 15573 4046 15607
rect 4080 15573 4114 15607
rect 4148 15573 4182 15607
rect 4216 15573 4250 15607
rect 4284 15573 4318 15607
rect 4352 15573 4386 15607
rect 4420 15573 4454 15607
rect 4488 15573 4522 15607
rect 4556 15573 4590 15607
rect 4624 15573 4658 15607
rect 4692 15573 4726 15607
rect 4760 15573 4794 15607
rect 4828 15573 4862 15607
rect 4896 15573 4930 15607
rect 4964 15573 4998 15607
rect 5032 15573 5066 15607
rect 5100 15573 5134 15607
rect 5168 15573 5202 15607
rect 5236 15573 5270 15607
rect 5304 15573 5338 15607
rect 5372 15573 5406 15607
rect 68 15501 102 15535
rect 139 15501 173 15535
rect 210 15501 244 15535
rect 281 15501 315 15535
rect 352 15501 386 15535
rect 420 15480 454 15514
rect 488 15480 522 15514
rect 68 15432 102 15466
rect 139 15432 173 15466
rect 210 15432 244 15466
rect 281 15432 315 15466
rect 352 15432 386 15466
rect 420 15411 454 15445
rect 488 15411 522 15445
rect 68 15363 102 15397
rect 139 15363 173 15397
rect 210 15363 244 15397
rect 281 15363 315 15397
rect 352 15363 386 15397
rect 420 15341 454 15375
rect 488 15341 522 15375
rect 68 15294 102 15328
rect 139 15294 173 15328
rect 210 15294 244 15328
rect 281 15294 315 15328
rect 352 15294 386 15328
rect 420 15271 454 15305
rect 488 15271 522 15305
rect 68 15225 102 15259
rect 139 15225 173 15259
rect 210 15225 244 15259
rect 281 15225 315 15259
rect 352 15225 386 15259
rect 420 15201 454 15235
rect 488 15201 522 15235
rect 68 15156 102 15190
rect 139 15156 173 15190
rect 210 15156 244 15190
rect 281 15156 315 15190
rect 352 15156 386 15190
rect 420 15131 454 15165
rect 488 15131 522 15165
rect 68 15087 102 15121
rect 139 15087 173 15121
rect 210 15087 244 15121
rect 281 15087 315 15121
rect 352 15087 386 15121
rect 420 15061 454 15095
rect 488 15061 522 15095
rect 68 15018 102 15052
rect 139 15018 173 15052
rect 210 15018 244 15052
rect 281 15018 315 15052
rect 352 15018 386 15052
rect 420 14991 454 15025
rect 488 14991 522 15025
rect 68 14949 102 14983
rect 139 14949 173 14983
rect 210 14949 244 14983
rect 281 14949 315 14983
rect 352 14949 386 14983
rect 420 14921 454 14955
rect 488 14921 522 14955
rect 68 14880 102 14914
rect 139 14880 173 14914
rect 210 14880 244 14914
rect 281 14880 315 14914
rect 352 14880 386 14914
rect 420 14851 454 14885
rect 488 14851 522 14885
rect 68 14811 102 14845
rect 139 14811 173 14845
rect 210 14811 244 14845
rect 281 14811 315 14845
rect 352 14811 386 14845
rect 12660 15547 12694 15581
rect 12730 15547 12764 15581
rect 12800 15547 12834 15581
rect 12869 15547 12903 15581
rect 12938 15547 12972 15581
rect 13007 15547 13041 15581
rect 13076 15547 13110 15581
rect 13145 15547 13179 15581
rect 13214 15547 13248 15581
rect 13283 15547 13317 15581
rect 13352 15547 13386 15581
rect 13421 15547 13455 15581
rect 13490 15547 13524 15581
rect 13559 15547 13593 15581
rect 13628 15547 13662 15581
rect 13697 15547 13731 15581
rect 13766 15547 13800 15581
rect 13835 15547 13869 15581
rect 13904 15547 13938 15581
rect 13973 15547 14007 15581
rect 14042 15547 14076 15581
rect 14111 15547 14145 15581
rect 14180 15547 14214 15581
rect 14249 15547 14283 15581
rect 14318 15547 14352 15581
rect 14420 15572 14454 15606
rect 14492 15572 14526 15606
rect 14564 15572 14598 15606
rect 14636 15572 14670 15606
rect 14708 15572 14742 15606
rect 14780 15572 14814 15606
rect 14852 15572 14886 15606
rect 14924 15572 14958 15606
rect 14996 15572 15030 15606
rect 15068 15572 15102 15606
rect 12660 15477 12694 15511
rect 12730 15477 12764 15511
rect 12800 15477 12834 15511
rect 12869 15477 12903 15511
rect 12938 15477 12972 15511
rect 13007 15477 13041 15511
rect 13076 15477 13110 15511
rect 13145 15477 13179 15511
rect 13214 15477 13248 15511
rect 13283 15477 13317 15511
rect 13352 15477 13386 15511
rect 13421 15477 13455 15511
rect 13490 15477 13524 15511
rect 13559 15477 13593 15511
rect 13628 15477 13662 15511
rect 13697 15477 13731 15511
rect 13766 15477 13800 15511
rect 13835 15477 13869 15511
rect 13904 15477 13938 15511
rect 13973 15477 14007 15511
rect 14042 15477 14076 15511
rect 14111 15477 14145 15511
rect 14180 15477 14214 15511
rect 14249 15477 14283 15511
rect 14318 15477 14352 15511
rect 14420 15503 14454 15537
rect 14492 15503 14526 15537
rect 14564 15503 14598 15537
rect 14636 15503 14670 15537
rect 14708 15503 14742 15537
rect 14780 15503 14814 15537
rect 14852 15503 14886 15537
rect 14924 15503 14958 15537
rect 14996 15503 15030 15537
rect 15068 15503 15102 15537
rect 12660 15407 12694 15441
rect 12730 15407 12764 15441
rect 12800 15407 12834 15441
rect 12869 15407 12903 15441
rect 12938 15407 12972 15441
rect 13007 15407 13041 15441
rect 13076 15407 13110 15441
rect 13145 15407 13179 15441
rect 13214 15407 13248 15441
rect 13283 15407 13317 15441
rect 13352 15407 13386 15441
rect 13421 15407 13455 15441
rect 13490 15407 13524 15441
rect 13559 15407 13593 15441
rect 13628 15407 13662 15441
rect 13697 15407 13731 15441
rect 13766 15407 13800 15441
rect 13835 15407 13869 15441
rect 13904 15407 13938 15441
rect 13973 15407 14007 15441
rect 14042 15407 14076 15441
rect 14111 15407 14145 15441
rect 14180 15407 14214 15441
rect 14249 15407 14283 15441
rect 14318 15407 14352 15441
rect 14420 15434 14454 15468
rect 14492 15434 14526 15468
rect 14564 15434 14598 15468
rect 14636 15434 14670 15468
rect 14708 15434 14742 15468
rect 14780 15434 14814 15468
rect 14852 15434 14886 15468
rect 14924 15434 14958 15468
rect 14996 15434 15030 15468
rect 15068 15434 15102 15468
rect 12660 15337 12694 15371
rect 12730 15337 12764 15371
rect 12800 15337 12834 15371
rect 12869 15337 12903 15371
rect 12938 15337 12972 15371
rect 13007 15337 13041 15371
rect 13076 15337 13110 15371
rect 13145 15337 13179 15371
rect 13214 15337 13248 15371
rect 13283 15337 13317 15371
rect 13352 15337 13386 15371
rect 13421 15337 13455 15371
rect 13490 15337 13524 15371
rect 13559 15337 13593 15371
rect 13628 15337 13662 15371
rect 13697 15337 13731 15371
rect 13766 15337 13800 15371
rect 13835 15337 13869 15371
rect 13904 15337 13938 15371
rect 13973 15337 14007 15371
rect 14042 15337 14076 15371
rect 14111 15337 14145 15371
rect 14180 15337 14214 15371
rect 14249 15337 14283 15371
rect 14318 15337 14352 15371
rect 14420 15365 14454 15399
rect 14492 15365 14526 15399
rect 14564 15365 14598 15399
rect 14636 15365 14670 15399
rect 14708 15365 14742 15399
rect 14780 15365 14814 15399
rect 14852 15365 14886 15399
rect 14924 15365 14958 15399
rect 14996 15365 15030 15399
rect 15068 15365 15102 15399
rect 12660 15267 12694 15301
rect 12730 15267 12764 15301
rect 12800 15267 12834 15301
rect 12869 15267 12903 15301
rect 12938 15267 12972 15301
rect 13007 15267 13041 15301
rect 13076 15267 13110 15301
rect 13145 15267 13179 15301
rect 13214 15267 13248 15301
rect 13283 15267 13317 15301
rect 13352 15267 13386 15301
rect 13421 15267 13455 15301
rect 13490 15267 13524 15301
rect 13559 15267 13593 15301
rect 13628 15267 13662 15301
rect 13697 15267 13731 15301
rect 13766 15267 13800 15301
rect 13835 15267 13869 15301
rect 13904 15267 13938 15301
rect 13973 15267 14007 15301
rect 14042 15267 14076 15301
rect 14111 15267 14145 15301
rect 14180 15267 14214 15301
rect 14249 15267 14283 15301
rect 14318 15267 14352 15301
rect 14420 15296 14454 15330
rect 14492 15296 14526 15330
rect 14564 15296 14598 15330
rect 14636 15296 14670 15330
rect 14708 15296 14742 15330
rect 14780 15296 14814 15330
rect 14852 15296 14886 15330
rect 14924 15296 14958 15330
rect 14996 15296 15030 15330
rect 15068 15296 15102 15330
rect 12660 15197 12694 15231
rect 12730 15197 12764 15231
rect 12800 15197 12834 15231
rect 12869 15197 12903 15231
rect 12938 15197 12972 15231
rect 13007 15197 13041 15231
rect 13076 15197 13110 15231
rect 13145 15197 13179 15231
rect 13214 15197 13248 15231
rect 13283 15197 13317 15231
rect 13352 15197 13386 15231
rect 13421 15197 13455 15231
rect 13490 15197 13524 15231
rect 13559 15197 13593 15231
rect 13628 15197 13662 15231
rect 13697 15197 13731 15231
rect 13766 15197 13800 15231
rect 13835 15197 13869 15231
rect 13904 15197 13938 15231
rect 13973 15197 14007 15231
rect 14042 15197 14076 15231
rect 14111 15197 14145 15231
rect 14180 15197 14214 15231
rect 14249 15197 14283 15231
rect 14318 15197 14352 15231
rect 14420 15227 14454 15261
rect 14492 15227 14526 15261
rect 14564 15227 14598 15261
rect 14636 15227 14670 15261
rect 14708 15227 14742 15261
rect 14780 15227 14814 15261
rect 14852 15227 14886 15261
rect 14924 15227 14958 15261
rect 14996 15227 15030 15261
rect 15068 15227 15102 15261
rect 12660 15127 12694 15161
rect 12730 15127 12764 15161
rect 12800 15127 12834 15161
rect 12869 15127 12903 15161
rect 12938 15127 12972 15161
rect 13007 15127 13041 15161
rect 13076 15127 13110 15161
rect 13145 15127 13179 15161
rect 13214 15127 13248 15161
rect 13283 15127 13317 15161
rect 13352 15127 13386 15161
rect 13421 15127 13455 15161
rect 13490 15127 13524 15161
rect 13559 15127 13593 15161
rect 13628 15127 13662 15161
rect 13697 15127 13731 15161
rect 13766 15127 13800 15161
rect 13835 15127 13869 15161
rect 13904 15127 13938 15161
rect 13973 15127 14007 15161
rect 14042 15127 14076 15161
rect 14111 15127 14145 15161
rect 14180 15127 14214 15161
rect 14249 15127 14283 15161
rect 14318 15127 14352 15161
rect 14420 15158 14454 15192
rect 14492 15158 14526 15192
rect 14564 15158 14598 15192
rect 14636 15158 14670 15192
rect 14708 15158 14742 15192
rect 14780 15158 14814 15192
rect 14852 15158 14886 15192
rect 14924 15158 14958 15192
rect 14996 15158 15030 15192
rect 15068 15158 15102 15192
rect 12660 15057 12694 15091
rect 12730 15057 12764 15091
rect 12800 15057 12834 15091
rect 12869 15057 12903 15091
rect 12938 15057 12972 15091
rect 13007 15057 13041 15091
rect 13076 15057 13110 15091
rect 13145 15057 13179 15091
rect 13214 15057 13248 15091
rect 13283 15057 13317 15091
rect 13352 15057 13386 15091
rect 13421 15057 13455 15091
rect 13490 15057 13524 15091
rect 13559 15057 13593 15091
rect 13628 15057 13662 15091
rect 13697 15057 13731 15091
rect 13766 15057 13800 15091
rect 13835 15057 13869 15091
rect 13904 15057 13938 15091
rect 13973 15057 14007 15091
rect 14042 15057 14076 15091
rect 14111 15057 14145 15091
rect 14180 15057 14214 15091
rect 14249 15057 14283 15091
rect 14318 15057 14352 15091
rect 14420 15089 14454 15123
rect 14492 15089 14526 15123
rect 14564 15089 14598 15123
rect 14636 15089 14670 15123
rect 14708 15089 14742 15123
rect 14780 15089 14814 15123
rect 14852 15089 14886 15123
rect 14924 15089 14958 15123
rect 14996 15089 15030 15123
rect 15068 15089 15102 15123
rect 12660 14987 12694 15021
rect 12730 14987 12764 15021
rect 12800 14987 12834 15021
rect 12869 14987 12903 15021
rect 12938 14987 12972 15021
rect 13007 14987 13041 15021
rect 13076 14987 13110 15021
rect 13145 14987 13179 15021
rect 13214 14987 13248 15021
rect 13283 14987 13317 15021
rect 13352 14987 13386 15021
rect 13421 14987 13455 15021
rect 13490 14987 13524 15021
rect 13559 14987 13593 15021
rect 13628 14987 13662 15021
rect 13697 14987 13731 15021
rect 13766 14987 13800 15021
rect 13835 14987 13869 15021
rect 13904 14987 13938 15021
rect 13973 14987 14007 15021
rect 14042 14987 14076 15021
rect 14111 14987 14145 15021
rect 14180 14987 14214 15021
rect 14249 14987 14283 15021
rect 14318 14987 14352 15021
rect 14420 15020 14454 15054
rect 14492 15020 14526 15054
rect 14564 15020 14598 15054
rect 14636 15020 14670 15054
rect 14708 15020 14742 15054
rect 14780 15020 14814 15054
rect 14852 15020 14886 15054
rect 14924 15020 14958 15054
rect 14996 15020 15030 15054
rect 15068 15020 15102 15054
rect 14420 14951 14454 14985
rect 14492 14951 14526 14985
rect 14564 14951 14598 14985
rect 14636 14951 14670 14985
rect 14708 14951 14742 14985
rect 14780 14951 14814 14985
rect 14852 14951 14886 14985
rect 14924 14951 14958 14985
rect 14996 14951 15030 14985
rect 15068 14951 15102 14985
rect 12660 14917 12694 14951
rect 12730 14917 12764 14951
rect 12800 14917 12834 14951
rect 12869 14917 12903 14951
rect 12938 14917 12972 14951
rect 13007 14917 13041 14951
rect 13076 14917 13110 14951
rect 13145 14917 13179 14951
rect 13214 14917 13248 14951
rect 13283 14917 13317 14951
rect 13352 14917 13386 14951
rect 13421 14917 13455 14951
rect 13490 14917 13524 14951
rect 13559 14917 13593 14951
rect 13628 14917 13662 14951
rect 13697 14917 13731 14951
rect 13766 14917 13800 14951
rect 13835 14917 13869 14951
rect 13904 14917 13938 14951
rect 13973 14917 14007 14951
rect 14042 14917 14076 14951
rect 14111 14917 14145 14951
rect 14180 14917 14214 14951
rect 14249 14917 14283 14951
rect 14318 14917 14352 14951
rect 14420 14882 14454 14916
rect 14492 14882 14526 14916
rect 14564 14882 14598 14916
rect 14636 14882 14670 14916
rect 14708 14882 14742 14916
rect 14780 14882 14814 14916
rect 14852 14882 14886 14916
rect 14924 14882 14958 14916
rect 14996 14882 15030 14916
rect 15068 14882 15102 14916
rect 12660 14847 12694 14881
rect 12730 14847 12764 14881
rect 12800 14847 12834 14881
rect 12869 14847 12903 14881
rect 12938 14847 12972 14881
rect 13007 14847 13041 14881
rect 13076 14847 13110 14881
rect 13145 14847 13179 14881
rect 13214 14847 13248 14881
rect 13283 14847 13317 14881
rect 13352 14847 13386 14881
rect 13421 14847 13455 14881
rect 13490 14847 13524 14881
rect 13559 14847 13593 14881
rect 13628 14847 13662 14881
rect 13697 14847 13731 14881
rect 13766 14847 13800 14881
rect 13835 14847 13869 14881
rect 13904 14847 13938 14881
rect 13973 14847 14007 14881
rect 14042 14847 14076 14881
rect 14111 14847 14145 14881
rect 14180 14847 14214 14881
rect 14249 14847 14283 14881
rect 14318 14847 14352 14881
rect 14420 14813 14454 14847
rect 14492 14813 14526 14847
rect 14564 14813 14598 14847
rect 14636 14813 14670 14847
rect 14708 14813 14742 14847
rect 14780 14813 14814 14847
rect 14852 14813 14886 14847
rect 14924 14813 14958 14847
rect 14996 14813 15030 14847
rect 15068 14813 15102 14847
rect 68 8740 102 8774
rect 138 8740 172 8774
rect 208 8740 242 8774
rect 278 8740 312 8774
rect 348 8740 382 8774
rect 418 8740 452 8774
rect 488 8740 522 8774
rect 558 8740 592 8774
rect 628 8740 662 8774
rect 698 8740 732 8774
rect 768 8740 802 8774
rect 838 8740 872 8774
rect 908 8740 942 8774
rect 978 8740 1012 8774
rect 1048 8740 1082 8774
rect 1118 8740 1152 8774
rect 1188 8740 1222 8774
rect 1258 8740 1292 8774
rect 1328 8740 1362 8774
rect 1398 8740 1432 8774
rect 1467 8740 1501 8774
rect 1536 8740 1570 8774
rect 1605 8740 1639 8774
rect 1674 8740 1708 8774
rect 1743 8740 1777 8774
rect 1812 8740 1846 8774
rect 1881 8740 1915 8774
rect 1950 8740 1984 8774
rect 2019 8740 2053 8774
rect 2088 8740 2122 8774
rect 2157 8740 2191 8774
rect 2226 8740 2260 8774
rect 2295 8740 2329 8774
rect 2364 8740 2398 8774
rect 2433 8740 2467 8774
rect 2502 8740 2536 8774
rect 2571 8740 2605 8774
rect 2640 8740 2674 8774
rect 2709 8740 2743 8774
rect 2778 8740 2812 8774
rect 2847 8740 2881 8774
rect 2933 8736 2967 8770
rect 3002 8736 3036 8770
rect 3071 8736 3105 8770
rect 3139 8736 3173 8770
rect 3207 8736 3241 8770
rect 3275 8736 3309 8770
rect 3343 8736 3377 8770
rect 3411 8736 3445 8770
rect 3479 8736 3513 8770
rect 3547 8736 3581 8770
rect 3615 8736 3649 8770
rect 3683 8736 3717 8770
rect 3751 8736 3785 8770
rect 3819 8736 3853 8770
rect 3887 8736 3921 8770
rect 3955 8736 3989 8770
rect 4023 8736 4057 8770
rect 4091 8736 4125 8770
rect 4159 8736 4193 8770
rect 4227 8736 4261 8770
rect 4295 8736 4329 8770
rect 4363 8736 4397 8770
rect 4431 8736 4465 8770
rect 4499 8736 4533 8770
rect 4567 8736 4601 8770
rect 4635 8736 4669 8770
rect 4703 8736 4737 8770
rect 4771 8736 4805 8770
rect 4839 8736 4873 8770
rect 4907 8736 4941 8770
rect 4975 8736 5009 8770
rect 5043 8736 5077 8770
rect 5111 8736 5145 8770
rect 5179 8736 5213 8770
rect 5247 8736 5281 8770
rect 5315 8736 5349 8770
rect 5383 8736 5417 8770
rect 5451 8736 5485 8770
rect 5519 8736 5553 8770
rect 5587 8736 5621 8770
rect 5655 8736 5689 8770
rect 5723 8736 5757 8770
rect 5791 8736 5825 8770
rect 5859 8736 5893 8770
rect 5927 8736 5961 8770
rect 5995 8736 6029 8770
rect 6063 8736 6097 8770
rect 6131 8736 6165 8770
rect 6199 8736 6233 8770
rect 6267 8736 6301 8770
rect 6335 8736 6369 8770
rect 6403 8736 6437 8770
rect 6471 8736 6505 8770
rect 6539 8736 6573 8770
rect 6607 8736 6641 8770
rect 6675 8736 6709 8770
rect 6743 8736 6777 8770
rect 6811 8736 6845 8770
rect 6879 8736 6913 8770
rect 6947 8736 6981 8770
rect 7015 8736 7049 8770
rect 7083 8736 7117 8770
rect 7151 8736 7185 8770
rect 7219 8736 7253 8770
rect 7287 8736 7321 8770
rect 7355 8736 7389 8770
rect 7423 8736 7457 8770
rect 7491 8736 7525 8770
rect 7559 8736 7593 8770
rect 7627 8736 7661 8770
rect 7695 8736 7729 8770
rect 7763 8736 7797 8770
rect 7831 8736 7865 8770
rect 7899 8736 7933 8770
rect 7967 8736 8001 8770
rect 8035 8736 8069 8770
rect 8103 8736 8137 8770
rect 8171 8736 8205 8770
rect 8239 8736 8273 8770
rect 8307 8736 8341 8770
rect 8393 8739 8427 8773
rect 8462 8739 8496 8773
rect 8531 8739 8565 8773
rect 8600 8739 8634 8773
rect 8669 8739 8703 8773
rect 8738 8739 8772 8773
rect 8807 8739 8841 8773
rect 8876 8739 8910 8773
rect 8945 8739 8979 8773
rect 9014 8739 9048 8773
rect 9083 8739 9117 8773
rect 9152 8739 9186 8773
rect 9220 8739 9254 8773
rect 9288 8739 9322 8773
rect 9356 8739 9390 8773
rect 9424 8739 9458 8773
rect 9492 8739 9526 8773
rect 9560 8739 9594 8773
rect 9628 8739 9662 8773
rect 9696 8739 9730 8773
rect 9764 8739 9798 8773
rect 9832 8739 9866 8773
rect 9900 8739 9934 8773
rect 9968 8739 10002 8773
rect 10036 8739 10070 8773
rect 10104 8739 10138 8773
rect 10172 8739 10206 8773
rect 10240 8739 10274 8773
rect 10308 8739 10342 8773
rect 10376 8739 10410 8773
rect 10444 8739 10478 8773
rect 10512 8739 10546 8773
rect 10580 8739 10614 8773
rect 10648 8739 10682 8773
rect 10716 8739 10750 8773
rect 10784 8739 10818 8773
rect 10852 8739 10886 8773
rect 10920 8739 10954 8773
rect 10988 8739 11022 8773
rect 11056 8739 11090 8773
rect 11124 8739 11158 8773
rect 11192 8739 11226 8773
rect 11260 8739 11294 8773
rect 11328 8739 11362 8773
rect 11396 8739 11430 8773
rect 11464 8739 11498 8773
rect 11532 8739 11566 8773
rect 11600 8739 11634 8773
rect 11668 8739 11702 8773
rect 11736 8739 11770 8773
rect 11804 8739 11838 8773
rect 11872 8739 11906 8773
rect 11940 8739 11974 8773
rect 12008 8739 12042 8773
rect 12076 8739 12110 8773
rect 12144 8739 12178 8773
rect 12212 8739 12246 8773
rect 12280 8739 12314 8773
rect 12348 8739 12382 8773
rect 12416 8739 12450 8773
rect 12484 8739 12518 8773
rect 12552 8739 12586 8773
rect 12620 8739 12654 8773
rect 12688 8739 12722 8773
rect 12756 8739 12790 8773
rect 12824 8739 12858 8773
rect 12892 8739 12926 8773
rect 12960 8739 12994 8773
rect 13028 8739 13062 8773
rect 13096 8739 13130 8773
rect 13164 8739 13198 8773
rect 13232 8739 13266 8773
rect 13300 8739 13334 8773
rect 13368 8739 13402 8773
rect 13436 8739 13470 8773
rect 13504 8739 13538 8773
rect 13572 8739 13606 8773
rect 13640 8739 13674 8773
rect 13708 8739 13742 8773
rect 13776 8739 13810 8773
rect 13844 8739 13878 8773
rect 13912 8739 13946 8773
rect 13980 8739 14014 8773
rect 14048 8739 14082 8773
rect 14116 8739 14150 8773
rect 14184 8739 14218 8773
rect 14252 8739 14286 8773
rect 14320 8739 14354 8773
rect 14388 8739 14422 8773
rect 14456 8739 14490 8773
rect 14524 8739 14558 8773
rect 14592 8739 14626 8773
rect 14660 8739 14694 8773
rect 14728 8739 14762 8773
rect 14796 8739 14830 8773
rect 14864 8739 14898 8773
rect 68 8666 102 8700
rect 138 8666 172 8700
rect 208 8666 242 8700
rect 278 8666 312 8700
rect 348 8666 382 8700
rect 418 8666 452 8700
rect 488 8666 522 8700
rect 558 8666 592 8700
rect 628 8666 662 8700
rect 698 8666 732 8700
rect 768 8666 802 8700
rect 838 8666 872 8700
rect 908 8666 942 8700
rect 978 8666 1012 8700
rect 1048 8666 1082 8700
rect 1118 8666 1152 8700
rect 1188 8666 1222 8700
rect 1258 8666 1292 8700
rect 1328 8666 1362 8700
rect 1398 8666 1432 8700
rect 1467 8666 1501 8700
rect 1536 8666 1570 8700
rect 1605 8666 1639 8700
rect 1674 8666 1708 8700
rect 1743 8666 1777 8700
rect 1812 8666 1846 8700
rect 1881 8666 1915 8700
rect 1950 8666 1984 8700
rect 2019 8666 2053 8700
rect 2088 8666 2122 8700
rect 2157 8666 2191 8700
rect 2226 8666 2260 8700
rect 2295 8666 2329 8700
rect 2364 8666 2398 8700
rect 2433 8666 2467 8700
rect 2502 8666 2536 8700
rect 2571 8666 2605 8700
rect 2640 8666 2674 8700
rect 2709 8666 2743 8700
rect 2778 8666 2812 8700
rect 2847 8666 2881 8700
rect 2933 8666 2967 8700
rect 3002 8666 3036 8700
rect 3071 8666 3105 8700
rect 3139 8666 3173 8700
rect 3207 8666 3241 8700
rect 3275 8666 3309 8700
rect 3343 8666 3377 8700
rect 3411 8666 3445 8700
rect 3479 8666 3513 8700
rect 3547 8666 3581 8700
rect 3615 8666 3649 8700
rect 3683 8666 3717 8700
rect 3751 8666 3785 8700
rect 3819 8666 3853 8700
rect 3887 8666 3921 8700
rect 3955 8666 3989 8700
rect 4023 8666 4057 8700
rect 4091 8666 4125 8700
rect 4159 8666 4193 8700
rect 4227 8666 4261 8700
rect 4295 8666 4329 8700
rect 4363 8666 4397 8700
rect 4431 8666 4465 8700
rect 4499 8666 4533 8700
rect 4567 8666 4601 8700
rect 4635 8666 4669 8700
rect 4703 8666 4737 8700
rect 4771 8666 4805 8700
rect 4839 8666 4873 8700
rect 4907 8666 4941 8700
rect 4975 8666 5009 8700
rect 5043 8666 5077 8700
rect 5111 8666 5145 8700
rect 5179 8666 5213 8700
rect 5247 8666 5281 8700
rect 5315 8666 5349 8700
rect 5383 8666 5417 8700
rect 5451 8666 5485 8700
rect 5519 8666 5553 8700
rect 5587 8666 5621 8700
rect 5655 8666 5689 8700
rect 5723 8666 5757 8700
rect 5791 8666 5825 8700
rect 5859 8666 5893 8700
rect 5927 8666 5961 8700
rect 5995 8666 6029 8700
rect 6063 8666 6097 8700
rect 6131 8666 6165 8700
rect 6199 8666 6233 8700
rect 6267 8666 6301 8700
rect 6335 8666 6369 8700
rect 6403 8666 6437 8700
rect 6471 8666 6505 8700
rect 6539 8666 6573 8700
rect 6607 8666 6641 8700
rect 6675 8666 6709 8700
rect 6743 8666 6777 8700
rect 6811 8666 6845 8700
rect 6879 8666 6913 8700
rect 6947 8666 6981 8700
rect 7015 8666 7049 8700
rect 7083 8666 7117 8700
rect 7151 8666 7185 8700
rect 7219 8666 7253 8700
rect 7287 8666 7321 8700
rect 7355 8666 7389 8700
rect 7423 8666 7457 8700
rect 7491 8666 7525 8700
rect 7559 8666 7593 8700
rect 7627 8666 7661 8700
rect 7695 8666 7729 8700
rect 7763 8666 7797 8700
rect 7831 8666 7865 8700
rect 7899 8666 7933 8700
rect 7967 8666 8001 8700
rect 8035 8666 8069 8700
rect 8103 8666 8137 8700
rect 8171 8666 8205 8700
rect 8239 8666 8273 8700
rect 8307 8666 8341 8700
rect 8393 8659 8427 8693
rect 8462 8659 8496 8693
rect 8531 8659 8565 8693
rect 8600 8659 8634 8693
rect 8669 8659 8703 8693
rect 8738 8659 8772 8693
rect 8807 8659 8841 8693
rect 8876 8659 8910 8693
rect 8945 8659 8979 8693
rect 9014 8659 9048 8693
rect 9083 8659 9117 8693
rect 9152 8659 9186 8693
rect 9220 8659 9254 8693
rect 9288 8659 9322 8693
rect 9356 8659 9390 8693
rect 9424 8659 9458 8693
rect 9492 8659 9526 8693
rect 9560 8659 9594 8693
rect 9628 8659 9662 8693
rect 9696 8659 9730 8693
rect 9764 8659 9798 8693
rect 9832 8659 9866 8693
rect 9900 8659 9934 8693
rect 9968 8659 10002 8693
rect 10036 8659 10070 8693
rect 10104 8659 10138 8693
rect 10172 8659 10206 8693
rect 10240 8659 10274 8693
rect 10308 8659 10342 8693
rect 10376 8659 10410 8693
rect 10444 8659 10478 8693
rect 10512 8659 10546 8693
rect 10580 8659 10614 8693
rect 10648 8659 10682 8693
rect 10716 8659 10750 8693
rect 10784 8659 10818 8693
rect 10852 8659 10886 8693
rect 10920 8659 10954 8693
rect 10988 8659 11022 8693
rect 11056 8659 11090 8693
rect 11124 8659 11158 8693
rect 11192 8659 11226 8693
rect 11260 8659 11294 8693
rect 11328 8659 11362 8693
rect 11396 8659 11430 8693
rect 11464 8659 11498 8693
rect 11532 8659 11566 8693
rect 11600 8659 11634 8693
rect 11668 8659 11702 8693
rect 11736 8659 11770 8693
rect 11804 8659 11838 8693
rect 11872 8659 11906 8693
rect 11940 8659 11974 8693
rect 12008 8659 12042 8693
rect 12076 8659 12110 8693
rect 12144 8659 12178 8693
rect 12212 8659 12246 8693
rect 12280 8659 12314 8693
rect 12348 8659 12382 8693
rect 12416 8659 12450 8693
rect 12484 8659 12518 8693
rect 12552 8659 12586 8693
rect 12620 8659 12654 8693
rect 12688 8659 12722 8693
rect 12756 8659 12790 8693
rect 12824 8659 12858 8693
rect 12892 8659 12926 8693
rect 12960 8659 12994 8693
rect 13028 8659 13062 8693
rect 13096 8659 13130 8693
rect 13164 8659 13198 8693
rect 13232 8659 13266 8693
rect 13300 8659 13334 8693
rect 13368 8659 13402 8693
rect 13436 8659 13470 8693
rect 13504 8659 13538 8693
rect 13572 8659 13606 8693
rect 13640 8659 13674 8693
rect 13708 8659 13742 8693
rect 13776 8659 13810 8693
rect 13844 8659 13878 8693
rect 13912 8659 13946 8693
rect 13980 8659 14014 8693
rect 14048 8659 14082 8693
rect 14116 8659 14150 8693
rect 14184 8659 14218 8693
rect 14252 8659 14286 8693
rect 14320 8659 14354 8693
rect 14388 8659 14422 8693
rect 14456 8659 14490 8693
rect 14524 8659 14558 8693
rect 14592 8659 14626 8693
rect 14660 8659 14694 8693
rect 14728 8659 14762 8693
rect 14796 8659 14830 8693
rect 14864 8659 14898 8693
rect 14932 8687 14966 8721
rect 15000 8687 15034 8721
rect 15068 8687 15102 8721
rect 68 8592 102 8626
rect 138 8592 172 8626
rect 208 8592 242 8626
rect 278 8592 312 8626
rect 348 8592 382 8626
rect 418 8592 452 8626
rect 488 8592 522 8626
rect 558 8592 592 8626
rect 628 8592 662 8626
rect 698 8592 732 8626
rect 768 8592 802 8626
rect 838 8592 872 8626
rect 908 8592 942 8626
rect 978 8592 1012 8626
rect 1048 8592 1082 8626
rect 1118 8592 1152 8626
rect 1188 8592 1222 8626
rect 1258 8592 1292 8626
rect 1328 8592 1362 8626
rect 1398 8592 1432 8626
rect 1467 8592 1501 8626
rect 1536 8592 1570 8626
rect 1605 8592 1639 8626
rect 1674 8592 1708 8626
rect 1743 8592 1777 8626
rect 1812 8592 1846 8626
rect 1881 8592 1915 8626
rect 1950 8592 1984 8626
rect 2019 8592 2053 8626
rect 2088 8592 2122 8626
rect 2157 8592 2191 8626
rect 2226 8592 2260 8626
rect 2295 8592 2329 8626
rect 2364 8592 2398 8626
rect 2433 8592 2467 8626
rect 2502 8592 2536 8626
rect 2571 8592 2605 8626
rect 2640 8592 2674 8626
rect 2709 8592 2743 8626
rect 2778 8592 2812 8626
rect 2847 8592 2881 8626
rect 2933 8596 2967 8630
rect 3002 8596 3036 8630
rect 3071 8596 3105 8630
rect 3139 8596 3173 8630
rect 3207 8596 3241 8630
rect 3275 8596 3309 8630
rect 3343 8596 3377 8630
rect 3411 8596 3445 8630
rect 3479 8596 3513 8630
rect 3547 8596 3581 8630
rect 3615 8596 3649 8630
rect 3683 8596 3717 8630
rect 3751 8596 3785 8630
rect 3819 8596 3853 8630
rect 3887 8596 3921 8630
rect 3955 8596 3989 8630
rect 4023 8596 4057 8630
rect 4091 8596 4125 8630
rect 4159 8596 4193 8630
rect 4227 8596 4261 8630
rect 4295 8596 4329 8630
rect 4363 8596 4397 8630
rect 4431 8596 4465 8630
rect 4499 8596 4533 8630
rect 4567 8596 4601 8630
rect 4635 8596 4669 8630
rect 4703 8596 4737 8630
rect 4771 8596 4805 8630
rect 4839 8596 4873 8630
rect 4907 8596 4941 8630
rect 4975 8596 5009 8630
rect 5043 8596 5077 8630
rect 5111 8596 5145 8630
rect 5179 8596 5213 8630
rect 5247 8596 5281 8630
rect 5315 8596 5349 8630
rect 5383 8596 5417 8630
rect 5451 8596 5485 8630
rect 5519 8596 5553 8630
rect 5587 8596 5621 8630
rect 5655 8596 5689 8630
rect 5723 8596 5757 8630
rect 5791 8596 5825 8630
rect 5859 8596 5893 8630
rect 5927 8596 5961 8630
rect 5995 8596 6029 8630
rect 6063 8596 6097 8630
rect 6131 8596 6165 8630
rect 6199 8596 6233 8630
rect 6267 8596 6301 8630
rect 6335 8596 6369 8630
rect 6403 8596 6437 8630
rect 6471 8596 6505 8630
rect 6539 8596 6573 8630
rect 6607 8596 6641 8630
rect 6675 8596 6709 8630
rect 6743 8596 6777 8630
rect 6811 8596 6845 8630
rect 6879 8596 6913 8630
rect 6947 8596 6981 8630
rect 7015 8596 7049 8630
rect 7083 8596 7117 8630
rect 7151 8596 7185 8630
rect 7219 8596 7253 8630
rect 7287 8596 7321 8630
rect 7355 8596 7389 8630
rect 7423 8596 7457 8630
rect 7491 8596 7525 8630
rect 7559 8596 7593 8630
rect 7627 8596 7661 8630
rect 7695 8596 7729 8630
rect 7763 8596 7797 8630
rect 7831 8596 7865 8630
rect 7899 8596 7933 8630
rect 7967 8596 8001 8630
rect 8035 8596 8069 8630
rect 8103 8596 8137 8630
rect 8171 8596 8205 8630
rect 8239 8596 8273 8630
rect 8307 8596 8341 8630
rect 14932 8615 14966 8649
rect 15000 8615 15034 8649
rect 15068 8615 15102 8649
rect 8393 8579 8427 8613
rect 8462 8579 8496 8613
rect 8531 8579 8565 8613
rect 8600 8579 8634 8613
rect 8669 8579 8703 8613
rect 8738 8579 8772 8613
rect 8807 8579 8841 8613
rect 8876 8579 8910 8613
rect 8945 8579 8979 8613
rect 9014 8579 9048 8613
rect 9083 8579 9117 8613
rect 9152 8579 9186 8613
rect 9220 8579 9254 8613
rect 9288 8579 9322 8613
rect 9356 8579 9390 8613
rect 9424 8579 9458 8613
rect 9492 8579 9526 8613
rect 9560 8579 9594 8613
rect 9628 8579 9662 8613
rect 9696 8579 9730 8613
rect 9764 8579 9798 8613
rect 9832 8579 9866 8613
rect 9900 8579 9934 8613
rect 9968 8579 10002 8613
rect 10036 8579 10070 8613
rect 10104 8579 10138 8613
rect 10172 8579 10206 8613
rect 10240 8579 10274 8613
rect 10308 8579 10342 8613
rect 10376 8579 10410 8613
rect 10444 8579 10478 8613
rect 10512 8579 10546 8613
rect 10580 8579 10614 8613
rect 10648 8579 10682 8613
rect 10716 8579 10750 8613
rect 10784 8579 10818 8613
rect 10852 8579 10886 8613
rect 10920 8579 10954 8613
rect 10988 8579 11022 8613
rect 11056 8579 11090 8613
rect 11124 8579 11158 8613
rect 11192 8579 11226 8613
rect 11260 8579 11294 8613
rect 11328 8579 11362 8613
rect 11396 8579 11430 8613
rect 11464 8579 11498 8613
rect 11532 8579 11566 8613
rect 11600 8579 11634 8613
rect 11668 8579 11702 8613
rect 11736 8579 11770 8613
rect 11804 8579 11838 8613
rect 11872 8579 11906 8613
rect 11940 8579 11974 8613
rect 12008 8579 12042 8613
rect 12076 8579 12110 8613
rect 12144 8579 12178 8613
rect 12212 8579 12246 8613
rect 12280 8579 12314 8613
rect 12348 8579 12382 8613
rect 12416 8579 12450 8613
rect 12484 8579 12518 8613
rect 12552 8579 12586 8613
rect 12620 8579 12654 8613
rect 12688 8579 12722 8613
rect 12756 8579 12790 8613
rect 12824 8579 12858 8613
rect 12892 8579 12926 8613
rect 12960 8579 12994 8613
rect 13028 8579 13062 8613
rect 13096 8579 13130 8613
rect 13164 8579 13198 8613
rect 13232 8579 13266 8613
rect 13300 8579 13334 8613
rect 13368 8579 13402 8613
rect 13436 8579 13470 8613
rect 13504 8579 13538 8613
rect 13572 8579 13606 8613
rect 13640 8579 13674 8613
rect 13708 8579 13742 8613
rect 13776 8579 13810 8613
rect 13844 8579 13878 8613
rect 13912 8579 13946 8613
rect 13980 8579 14014 8613
rect 14048 8579 14082 8613
rect 14116 8579 14150 8613
rect 14184 8579 14218 8613
rect 14252 8579 14286 8613
rect 14320 8579 14354 8613
rect 14388 8579 14422 8613
rect 14456 8579 14490 8613
rect 14524 8579 14558 8613
rect 14592 8579 14626 8613
rect 14660 8579 14694 8613
rect 14728 8579 14762 8613
rect 14796 8579 14830 8613
rect 14864 8579 14898 8613
rect 68 8518 102 8552
rect 138 8518 172 8552
rect 208 8518 242 8552
rect 278 8518 312 8552
rect 348 8518 382 8552
rect 418 8518 452 8552
rect 488 8518 522 8552
rect 558 8518 592 8552
rect 628 8518 662 8552
rect 698 8518 732 8552
rect 768 8518 802 8552
rect 838 8518 872 8552
rect 908 8518 942 8552
rect 978 8518 1012 8552
rect 1048 8518 1082 8552
rect 1118 8518 1152 8552
rect 1188 8518 1222 8552
rect 1258 8518 1292 8552
rect 1328 8518 1362 8552
rect 1398 8518 1432 8552
rect 1467 8518 1501 8552
rect 1536 8518 1570 8552
rect 1605 8518 1639 8552
rect 1674 8518 1708 8552
rect 1743 8518 1777 8552
rect 1812 8518 1846 8552
rect 1881 8518 1915 8552
rect 1950 8518 1984 8552
rect 2019 8518 2053 8552
rect 2088 8518 2122 8552
rect 2157 8518 2191 8552
rect 2226 8518 2260 8552
rect 2295 8518 2329 8552
rect 2364 8518 2398 8552
rect 2433 8518 2467 8552
rect 2502 8518 2536 8552
rect 2571 8518 2605 8552
rect 2640 8518 2674 8552
rect 2709 8518 2743 8552
rect 2778 8518 2812 8552
rect 2847 8518 2881 8552
rect 2933 8526 2967 8560
rect 3002 8526 3036 8560
rect 3071 8526 3105 8560
rect 3139 8526 3173 8560
rect 3207 8526 3241 8560
rect 3275 8526 3309 8560
rect 3343 8526 3377 8560
rect 3411 8526 3445 8560
rect 3479 8526 3513 8560
rect 3547 8526 3581 8560
rect 3615 8526 3649 8560
rect 3683 8526 3717 8560
rect 3751 8526 3785 8560
rect 3819 8526 3853 8560
rect 3887 8526 3921 8560
rect 3955 8526 3989 8560
rect 4023 8526 4057 8560
rect 4091 8526 4125 8560
rect 4159 8526 4193 8560
rect 4227 8526 4261 8560
rect 4295 8526 4329 8560
rect 4363 8526 4397 8560
rect 4431 8526 4465 8560
rect 4499 8526 4533 8560
rect 4567 8526 4601 8560
rect 4635 8526 4669 8560
rect 4703 8526 4737 8560
rect 4771 8526 4805 8560
rect 4839 8526 4873 8560
rect 4907 8526 4941 8560
rect 4975 8526 5009 8560
rect 5043 8526 5077 8560
rect 5111 8526 5145 8560
rect 5179 8526 5213 8560
rect 5247 8526 5281 8560
rect 5315 8526 5349 8560
rect 5383 8526 5417 8560
rect 5451 8526 5485 8560
rect 5519 8526 5553 8560
rect 5587 8526 5621 8560
rect 5655 8526 5689 8560
rect 5723 8526 5757 8560
rect 5791 8526 5825 8560
rect 5859 8526 5893 8560
rect 5927 8526 5961 8560
rect 5995 8526 6029 8560
rect 6063 8526 6097 8560
rect 6131 8526 6165 8560
rect 6199 8526 6233 8560
rect 6267 8526 6301 8560
rect 6335 8526 6369 8560
rect 6403 8526 6437 8560
rect 6471 8526 6505 8560
rect 6539 8526 6573 8560
rect 6607 8526 6641 8560
rect 6675 8526 6709 8560
rect 6743 8526 6777 8560
rect 6811 8526 6845 8560
rect 6879 8526 6913 8560
rect 6947 8526 6981 8560
rect 7015 8526 7049 8560
rect 7083 8526 7117 8560
rect 7151 8526 7185 8560
rect 7219 8526 7253 8560
rect 7287 8526 7321 8560
rect 7355 8526 7389 8560
rect 7423 8526 7457 8560
rect 7491 8526 7525 8560
rect 7559 8526 7593 8560
rect 7627 8526 7661 8560
rect 7695 8526 7729 8560
rect 7763 8526 7797 8560
rect 7831 8526 7865 8560
rect 7899 8526 7933 8560
rect 7967 8526 8001 8560
rect 8035 8526 8069 8560
rect 8103 8526 8137 8560
rect 8171 8526 8205 8560
rect 8239 8526 8273 8560
rect 8307 8526 8341 8560
rect 14932 8543 14966 8577
rect 15000 8543 15034 8577
rect 15068 8543 15102 8577
rect 8393 8499 8427 8533
rect 8462 8499 8496 8533
rect 8531 8499 8565 8533
rect 8600 8499 8634 8533
rect 8669 8499 8703 8533
rect 8738 8499 8772 8533
rect 8807 8499 8841 8533
rect 8876 8499 8910 8533
rect 8945 8499 8979 8533
rect 9014 8499 9048 8533
rect 9083 8499 9117 8533
rect 9152 8499 9186 8533
rect 9220 8499 9254 8533
rect 9288 8499 9322 8533
rect 9356 8499 9390 8533
rect 9424 8499 9458 8533
rect 9492 8499 9526 8533
rect 9560 8499 9594 8533
rect 9628 8499 9662 8533
rect 9696 8499 9730 8533
rect 9764 8499 9798 8533
rect 9832 8499 9866 8533
rect 9900 8499 9934 8533
rect 9968 8499 10002 8533
rect 10036 8499 10070 8533
rect 10104 8499 10138 8533
rect 10172 8499 10206 8533
rect 10240 8499 10274 8533
rect 10308 8499 10342 8533
rect 10376 8499 10410 8533
rect 10444 8499 10478 8533
rect 10512 8499 10546 8533
rect 10580 8499 10614 8533
rect 10648 8499 10682 8533
rect 10716 8499 10750 8533
rect 10784 8499 10818 8533
rect 10852 8499 10886 8533
rect 10920 8499 10954 8533
rect 10988 8499 11022 8533
rect 11056 8499 11090 8533
rect 11124 8499 11158 8533
rect 11192 8499 11226 8533
rect 11260 8499 11294 8533
rect 11328 8499 11362 8533
rect 11396 8499 11430 8533
rect 11464 8499 11498 8533
rect 11532 8499 11566 8533
rect 11600 8499 11634 8533
rect 11668 8499 11702 8533
rect 11736 8499 11770 8533
rect 11804 8499 11838 8533
rect 11872 8499 11906 8533
rect 11940 8499 11974 8533
rect 12008 8499 12042 8533
rect 12076 8499 12110 8533
rect 12144 8499 12178 8533
rect 12212 8499 12246 8533
rect 12280 8499 12314 8533
rect 12348 8499 12382 8533
rect 12416 8499 12450 8533
rect 12484 8499 12518 8533
rect 12552 8499 12586 8533
rect 12620 8499 12654 8533
rect 12688 8499 12722 8533
rect 12756 8499 12790 8533
rect 12824 8499 12858 8533
rect 12892 8499 12926 8533
rect 12960 8499 12994 8533
rect 13028 8499 13062 8533
rect 13096 8499 13130 8533
rect 13164 8499 13198 8533
rect 13232 8499 13266 8533
rect 13300 8499 13334 8533
rect 13368 8499 13402 8533
rect 13436 8499 13470 8533
rect 13504 8499 13538 8533
rect 13572 8499 13606 8533
rect 13640 8499 13674 8533
rect 13708 8499 13742 8533
rect 13776 8499 13810 8533
rect 13844 8499 13878 8533
rect 13912 8499 13946 8533
rect 13980 8499 14014 8533
rect 14048 8499 14082 8533
rect 14116 8499 14150 8533
rect 14184 8499 14218 8533
rect 14252 8499 14286 8533
rect 14320 8499 14354 8533
rect 14388 8499 14422 8533
rect 14456 8499 14490 8533
rect 14524 8499 14558 8533
rect 14592 8499 14626 8533
rect 14660 8499 14694 8533
rect 14728 8499 14762 8533
rect 14796 8499 14830 8533
rect 14864 8499 14898 8533
rect 68 8426 102 8460
rect 68 8358 102 8392
rect 2933 8456 2967 8490
rect 3002 8456 3036 8490
rect 3071 8456 3105 8490
rect 3139 8456 3173 8490
rect 3207 8456 3241 8490
rect 3275 8456 3309 8490
rect 3343 8456 3377 8490
rect 3411 8456 3445 8490
rect 3479 8456 3513 8490
rect 3547 8456 3581 8490
rect 3615 8456 3649 8490
rect 3683 8456 3717 8490
rect 3751 8456 3785 8490
rect 3819 8456 3853 8490
rect 3887 8456 3921 8490
rect 3955 8456 3989 8490
rect 4023 8456 4057 8490
rect 4091 8456 4125 8490
rect 4159 8456 4193 8490
rect 4227 8456 4261 8490
rect 4295 8456 4329 8490
rect 4363 8456 4397 8490
rect 4431 8456 4465 8490
rect 4499 8456 4533 8490
rect 4567 8456 4601 8490
rect 4635 8456 4669 8490
rect 4703 8456 4737 8490
rect 4771 8456 4805 8490
rect 4839 8456 4873 8490
rect 4907 8456 4941 8490
rect 4975 8456 5009 8490
rect 5043 8456 5077 8490
rect 5111 8456 5145 8490
rect 5179 8456 5213 8490
rect 5247 8456 5281 8490
rect 5315 8456 5349 8490
rect 5383 8456 5417 8490
rect 5451 8456 5485 8490
rect 5519 8456 5553 8490
rect 5587 8456 5621 8490
rect 5655 8456 5689 8490
rect 5723 8456 5757 8490
rect 5791 8456 5825 8490
rect 5859 8456 5893 8490
rect 5927 8456 5961 8490
rect 5995 8456 6029 8490
rect 6063 8456 6097 8490
rect 6131 8456 6165 8490
rect 6199 8456 6233 8490
rect 6267 8456 6301 8490
rect 6335 8456 6369 8490
rect 6403 8456 6437 8490
rect 6471 8456 6505 8490
rect 6539 8456 6573 8490
rect 6607 8456 6641 8490
rect 6675 8456 6709 8490
rect 6743 8456 6777 8490
rect 6811 8456 6845 8490
rect 6879 8456 6913 8490
rect 6947 8456 6981 8490
rect 7015 8456 7049 8490
rect 7083 8456 7117 8490
rect 7151 8456 7185 8490
rect 7219 8456 7253 8490
rect 7287 8456 7321 8490
rect 7355 8456 7389 8490
rect 7423 8456 7457 8490
rect 7491 8456 7525 8490
rect 7559 8456 7593 8490
rect 7627 8456 7661 8490
rect 7695 8456 7729 8490
rect 7763 8456 7797 8490
rect 7831 8456 7865 8490
rect 7899 8456 7933 8490
rect 7967 8456 8001 8490
rect 8035 8456 8069 8490
rect 8103 8456 8137 8490
rect 8171 8456 8205 8490
rect 8239 8456 8273 8490
rect 8307 8456 8341 8490
rect 14932 8471 14966 8505
rect 15000 8471 15034 8505
rect 15068 8471 15102 8505
rect 68 8290 102 8324
rect 2933 8386 2967 8420
rect 3002 8386 3036 8420
rect 3071 8386 3105 8420
rect 3139 8386 3173 8420
rect 3207 8386 3241 8420
rect 3275 8386 3309 8420
rect 3343 8386 3377 8420
rect 3411 8386 3445 8420
rect 3479 8386 3513 8420
rect 3547 8386 3581 8420
rect 3615 8386 3649 8420
rect 3683 8386 3717 8420
rect 3751 8386 3785 8420
rect 3819 8386 3853 8420
rect 3887 8386 3921 8420
rect 3955 8386 3989 8420
rect 4023 8386 4057 8420
rect 4091 8386 4125 8420
rect 4159 8386 4193 8420
rect 4227 8386 4261 8420
rect 4295 8386 4329 8420
rect 4363 8386 4397 8420
rect 4431 8386 4465 8420
rect 4499 8386 4533 8420
rect 4567 8386 4601 8420
rect 4635 8386 4669 8420
rect 4703 8386 4737 8420
rect 4771 8386 4805 8420
rect 4839 8386 4873 8420
rect 4907 8386 4941 8420
rect 4975 8386 5009 8420
rect 5043 8386 5077 8420
rect 5111 8386 5145 8420
rect 5179 8386 5213 8420
rect 5247 8386 5281 8420
rect 5315 8386 5349 8420
rect 5383 8386 5417 8420
rect 5451 8386 5485 8420
rect 5519 8386 5553 8420
rect 5587 8386 5621 8420
rect 5655 8386 5689 8420
rect 5723 8386 5757 8420
rect 5791 8386 5825 8420
rect 5859 8386 5893 8420
rect 5927 8386 5961 8420
rect 5995 8386 6029 8420
rect 6063 8386 6097 8420
rect 6131 8386 6165 8420
rect 6199 8386 6233 8420
rect 6267 8386 6301 8420
rect 6335 8386 6369 8420
rect 6403 8386 6437 8420
rect 6471 8386 6505 8420
rect 6539 8386 6573 8420
rect 6607 8386 6641 8420
rect 6675 8386 6709 8420
rect 6743 8386 6777 8420
rect 6811 8386 6845 8420
rect 6879 8386 6913 8420
rect 6947 8386 6981 8420
rect 7015 8386 7049 8420
rect 7083 8386 7117 8420
rect 7151 8386 7185 8420
rect 7219 8386 7253 8420
rect 7287 8386 7321 8420
rect 7355 8386 7389 8420
rect 7423 8386 7457 8420
rect 7491 8386 7525 8420
rect 7559 8386 7593 8420
rect 7627 8386 7661 8420
rect 7695 8386 7729 8420
rect 7763 8386 7797 8420
rect 7831 8386 7865 8420
rect 7899 8386 7933 8420
rect 7967 8386 8001 8420
rect 8035 8386 8069 8420
rect 8103 8386 8137 8420
rect 8171 8386 8205 8420
rect 8239 8386 8273 8420
rect 8307 8386 8341 8420
rect 8393 8419 8427 8453
rect 8462 8419 8496 8453
rect 8531 8419 8565 8453
rect 8600 8419 8634 8453
rect 8669 8419 8703 8453
rect 8738 8419 8772 8453
rect 8807 8419 8841 8453
rect 8876 8419 8910 8453
rect 8945 8419 8979 8453
rect 9014 8419 9048 8453
rect 9083 8419 9117 8453
rect 9152 8419 9186 8453
rect 9220 8419 9254 8453
rect 9288 8419 9322 8453
rect 9356 8419 9390 8453
rect 9424 8419 9458 8453
rect 9492 8419 9526 8453
rect 9560 8419 9594 8453
rect 9628 8419 9662 8453
rect 9696 8419 9730 8453
rect 9764 8419 9798 8453
rect 9832 8419 9866 8453
rect 9900 8419 9934 8453
rect 9968 8419 10002 8453
rect 10036 8419 10070 8453
rect 10104 8419 10138 8453
rect 10172 8419 10206 8453
rect 10240 8419 10274 8453
rect 10308 8419 10342 8453
rect 10376 8419 10410 8453
rect 10444 8419 10478 8453
rect 10512 8419 10546 8453
rect 10580 8419 10614 8453
rect 10648 8419 10682 8453
rect 10716 8419 10750 8453
rect 10784 8419 10818 8453
rect 10852 8419 10886 8453
rect 10920 8419 10954 8453
rect 10988 8419 11022 8453
rect 11056 8419 11090 8453
rect 11124 8419 11158 8453
rect 11192 8419 11226 8453
rect 11260 8419 11294 8453
rect 11328 8419 11362 8453
rect 11396 8419 11430 8453
rect 11464 8419 11498 8453
rect 11532 8419 11566 8453
rect 11600 8419 11634 8453
rect 11668 8419 11702 8453
rect 11736 8419 11770 8453
rect 11804 8419 11838 8453
rect 11872 8419 11906 8453
rect 11940 8419 11974 8453
rect 12008 8419 12042 8453
rect 12076 8419 12110 8453
rect 12144 8419 12178 8453
rect 12212 8419 12246 8453
rect 12280 8419 12314 8453
rect 12348 8419 12382 8453
rect 12416 8419 12450 8453
rect 12484 8419 12518 8453
rect 12552 8419 12586 8453
rect 12620 8419 12654 8453
rect 12688 8419 12722 8453
rect 12756 8419 12790 8453
rect 12824 8419 12858 8453
rect 12892 8419 12926 8453
rect 12960 8419 12994 8453
rect 13028 8419 13062 8453
rect 13096 8419 13130 8453
rect 13164 8419 13198 8453
rect 13232 8419 13266 8453
rect 13300 8419 13334 8453
rect 13368 8419 13402 8453
rect 13436 8419 13470 8453
rect 13504 8419 13538 8453
rect 13572 8419 13606 8453
rect 13640 8419 13674 8453
rect 13708 8419 13742 8453
rect 13776 8419 13810 8453
rect 13844 8419 13878 8453
rect 13912 8419 13946 8453
rect 13980 8419 14014 8453
rect 14048 8419 14082 8453
rect 14116 8419 14150 8453
rect 14184 8419 14218 8453
rect 14252 8419 14286 8453
rect 14320 8419 14354 8453
rect 14388 8419 14422 8453
rect 14456 8419 14490 8453
rect 14524 8419 14558 8453
rect 14592 8419 14626 8453
rect 14660 8419 14694 8453
rect 14728 8419 14762 8453
rect 14796 8419 14830 8453
rect 14864 8419 14898 8453
rect 14932 8399 14966 8433
rect 15000 8399 15034 8433
rect 15068 8399 15102 8433
rect 2933 8316 2967 8350
rect 3002 8316 3036 8350
rect 3071 8316 3105 8350
rect 3139 8316 3173 8350
rect 3207 8316 3241 8350
rect 3275 8316 3309 8350
rect 3343 8316 3377 8350
rect 3411 8316 3445 8350
rect 3479 8316 3513 8350
rect 3547 8316 3581 8350
rect 3615 8316 3649 8350
rect 3683 8316 3717 8350
rect 3751 8316 3785 8350
rect 3819 8316 3853 8350
rect 3887 8316 3921 8350
rect 3955 8316 3989 8350
rect 4023 8316 4057 8350
rect 4091 8316 4125 8350
rect 4159 8316 4193 8350
rect 4227 8316 4261 8350
rect 4295 8316 4329 8350
rect 4363 8316 4397 8350
rect 4431 8316 4465 8350
rect 4499 8316 4533 8350
rect 4567 8316 4601 8350
rect 4635 8316 4669 8350
rect 4703 8316 4737 8350
rect 4771 8316 4805 8350
rect 4839 8316 4873 8350
rect 4907 8316 4941 8350
rect 4975 8316 5009 8350
rect 5043 8316 5077 8350
rect 5111 8316 5145 8350
rect 5179 8316 5213 8350
rect 5247 8316 5281 8350
rect 5315 8316 5349 8350
rect 5383 8316 5417 8350
rect 5451 8316 5485 8350
rect 5519 8316 5553 8350
rect 5587 8316 5621 8350
rect 5655 8316 5689 8350
rect 5723 8316 5757 8350
rect 5791 8316 5825 8350
rect 5859 8316 5893 8350
rect 5927 8316 5961 8350
rect 5995 8316 6029 8350
rect 6063 8316 6097 8350
rect 6131 8316 6165 8350
rect 6199 8316 6233 8350
rect 6267 8316 6301 8350
rect 6335 8316 6369 8350
rect 6403 8316 6437 8350
rect 6471 8316 6505 8350
rect 6539 8316 6573 8350
rect 6607 8316 6641 8350
rect 6675 8316 6709 8350
rect 6743 8316 6777 8350
rect 6811 8316 6845 8350
rect 6879 8316 6913 8350
rect 6947 8316 6981 8350
rect 7015 8316 7049 8350
rect 7083 8316 7117 8350
rect 7151 8316 7185 8350
rect 7219 8316 7253 8350
rect 7287 8316 7321 8350
rect 7355 8316 7389 8350
rect 7423 8316 7457 8350
rect 7491 8316 7525 8350
rect 7559 8316 7593 8350
rect 7627 8316 7661 8350
rect 7695 8316 7729 8350
rect 7763 8316 7797 8350
rect 7831 8316 7865 8350
rect 7899 8316 7933 8350
rect 7967 8316 8001 8350
rect 8035 8316 8069 8350
rect 8103 8316 8137 8350
rect 8171 8316 8205 8350
rect 8239 8316 8273 8350
rect 8307 8316 8341 8350
rect 68 8222 102 8256
rect 13532 8323 13566 8357
rect 13603 8323 13637 8357
rect 13674 8323 13708 8357
rect 13744 8323 13778 8357
rect 13814 8323 13848 8357
rect 13884 8323 13918 8357
rect 13954 8323 13988 8357
rect 14024 8323 14058 8357
rect 14094 8323 14128 8357
rect 14164 8323 14198 8357
rect 14234 8323 14268 8357
rect 14304 8323 14338 8357
rect 14374 8323 14408 8357
rect 14444 8323 14478 8357
rect 14514 8323 14548 8357
rect 14584 8323 14618 8357
rect 14654 8323 14688 8357
rect 14724 8323 14758 8357
rect 14794 8323 14828 8357
rect 14864 8323 14898 8357
rect 14932 8327 14966 8361
rect 15000 8327 15034 8361
rect 15068 8327 15102 8361
rect 2933 8246 2967 8280
rect 3002 8246 3036 8280
rect 3071 8246 3105 8280
rect 3139 8246 3173 8280
rect 3207 8246 3241 8280
rect 3275 8246 3309 8280
rect 3343 8246 3377 8280
rect 3411 8246 3445 8280
rect 3479 8246 3513 8280
rect 3547 8246 3581 8280
rect 3615 8246 3649 8280
rect 3683 8246 3717 8280
rect 3751 8246 3785 8280
rect 3819 8246 3853 8280
rect 3887 8246 3921 8280
rect 3955 8246 3989 8280
rect 4023 8246 4057 8280
rect 4091 8246 4125 8280
rect 4159 8246 4193 8280
rect 4227 8246 4261 8280
rect 4295 8246 4329 8280
rect 4363 8246 4397 8280
rect 4431 8246 4465 8280
rect 4499 8246 4533 8280
rect 4567 8246 4601 8280
rect 4635 8246 4669 8280
rect 4703 8246 4737 8280
rect 4771 8246 4805 8280
rect 4839 8246 4873 8280
rect 4907 8246 4941 8280
rect 4975 8246 5009 8280
rect 5043 8246 5077 8280
rect 5111 8246 5145 8280
rect 5179 8246 5213 8280
rect 5247 8246 5281 8280
rect 5315 8246 5349 8280
rect 5383 8246 5417 8280
rect 5451 8246 5485 8280
rect 5519 8246 5553 8280
rect 5587 8246 5621 8280
rect 5655 8246 5689 8280
rect 5723 8246 5757 8280
rect 5791 8246 5825 8280
rect 5859 8246 5893 8280
rect 5927 8246 5961 8280
rect 5995 8246 6029 8280
rect 6063 8246 6097 8280
rect 6131 8246 6165 8280
rect 6199 8246 6233 8280
rect 6267 8246 6301 8280
rect 6335 8246 6369 8280
rect 6403 8246 6437 8280
rect 6471 8246 6505 8280
rect 6539 8246 6573 8280
rect 6607 8246 6641 8280
rect 6675 8246 6709 8280
rect 6743 8246 6777 8280
rect 6811 8246 6845 8280
rect 6879 8246 6913 8280
rect 6947 8246 6981 8280
rect 7015 8246 7049 8280
rect 7083 8246 7117 8280
rect 7151 8246 7185 8280
rect 7219 8246 7253 8280
rect 7287 8246 7321 8280
rect 7355 8246 7389 8280
rect 7423 8246 7457 8280
rect 7491 8246 7525 8280
rect 7559 8246 7593 8280
rect 7627 8246 7661 8280
rect 7695 8246 7729 8280
rect 7763 8246 7797 8280
rect 7831 8246 7865 8280
rect 7899 8246 7933 8280
rect 7967 8246 8001 8280
rect 8035 8246 8069 8280
rect 8103 8246 8137 8280
rect 8171 8246 8205 8280
rect 8239 8246 8273 8280
rect 8307 8246 8341 8280
rect 2933 8176 2967 8210
rect 3002 8176 3036 8210
rect 3071 8176 3105 8210
rect 3139 8176 3173 8210
rect 3207 8176 3241 8210
rect 3275 8176 3309 8210
rect 3343 8176 3377 8210
rect 3411 8176 3445 8210
rect 3479 8176 3513 8210
rect 3547 8176 3581 8210
rect 3615 8176 3649 8210
rect 3683 8176 3717 8210
rect 3751 8176 3785 8210
rect 3819 8176 3853 8210
rect 3887 8176 3921 8210
rect 3955 8176 3989 8210
rect 4023 8176 4057 8210
rect 4091 8176 4125 8210
rect 4159 8176 4193 8210
rect 4227 8176 4261 8210
rect 4295 8176 4329 8210
rect 4363 8176 4397 8210
rect 4431 8176 4465 8210
rect 4499 8176 4533 8210
rect 4567 8176 4601 8210
rect 4635 8176 4669 8210
rect 4703 8176 4737 8210
rect 4771 8176 4805 8210
rect 4839 8176 4873 8210
rect 4907 8176 4941 8210
rect 4975 8176 5009 8210
rect 5043 8176 5077 8210
rect 5111 8176 5145 8210
rect 5179 8176 5213 8210
rect 5247 8176 5281 8210
rect 5315 8176 5349 8210
rect 5383 8176 5417 8210
rect 5451 8176 5485 8210
rect 5519 8176 5553 8210
rect 5587 8176 5621 8210
rect 5655 8176 5689 8210
rect 5723 8176 5757 8210
rect 5791 8176 5825 8210
rect 5859 8176 5893 8210
rect 5927 8176 5961 8210
rect 5995 8176 6029 8210
rect 6063 8176 6097 8210
rect 6131 8176 6165 8210
rect 6199 8176 6233 8210
rect 6267 8176 6301 8210
rect 6335 8176 6369 8210
rect 6403 8176 6437 8210
rect 6471 8176 6505 8210
rect 6539 8176 6573 8210
rect 6607 8176 6641 8210
rect 6675 8176 6709 8210
rect 6743 8176 6777 8210
rect 6811 8176 6845 8210
rect 6879 8176 6913 8210
rect 6947 8176 6981 8210
rect 7015 8176 7049 8210
rect 7083 8176 7117 8210
rect 7151 8176 7185 8210
rect 7219 8176 7253 8210
rect 7287 8176 7321 8210
rect 7355 8176 7389 8210
rect 7423 8176 7457 8210
rect 7491 8176 7525 8210
rect 7559 8176 7593 8210
rect 7627 8176 7661 8210
rect 7695 8176 7729 8210
rect 7763 8176 7797 8210
rect 7831 8176 7865 8210
rect 7899 8176 7933 8210
rect 7967 8176 8001 8210
rect 8035 8176 8069 8210
rect 8103 8176 8137 8210
rect 8171 8176 8205 8210
rect 8239 8176 8273 8210
rect 8307 8176 8341 8210
rect 68 8123 102 8157
rect 138 8123 172 8157
rect 208 8123 242 8157
rect 278 8123 312 8157
rect 348 8123 382 8157
rect 418 8123 452 8157
rect 488 8123 522 8157
rect 558 8123 592 8157
rect 628 8123 662 8157
rect 698 8123 732 8157
rect 768 8123 802 8157
rect 838 8123 872 8157
rect 908 8123 942 8157
rect 978 8123 1012 8157
rect 1048 8123 1082 8157
rect 1118 8123 1152 8157
rect 1188 8123 1222 8157
rect 1258 8123 1292 8157
rect 1328 8123 1362 8157
rect 1398 8123 1432 8157
rect 1467 8123 1501 8157
rect 1536 8123 1570 8157
rect 1605 8123 1639 8157
rect 1674 8123 1708 8157
rect 1743 8123 1777 8157
rect 1812 8123 1846 8157
rect 1881 8123 1915 8157
rect 1950 8123 1984 8157
rect 2019 8123 2053 8157
rect 2088 8123 2122 8157
rect 2157 8123 2191 8157
rect 2226 8123 2260 8157
rect 2295 8123 2329 8157
rect 2364 8123 2398 8157
rect 2433 8123 2467 8157
rect 2502 8123 2536 8157
rect 2571 8123 2605 8157
rect 2640 8123 2674 8157
rect 2709 8123 2743 8157
rect 2778 8123 2812 8157
rect 2847 8123 2881 8157
rect 2933 8106 2967 8140
rect 3002 8106 3036 8140
rect 3071 8106 3105 8140
rect 3139 8106 3173 8140
rect 3207 8106 3241 8140
rect 3275 8106 3309 8140
rect 3343 8106 3377 8140
rect 3411 8106 3445 8140
rect 3479 8106 3513 8140
rect 3547 8106 3581 8140
rect 3615 8106 3649 8140
rect 3683 8106 3717 8140
rect 3751 8106 3785 8140
rect 3819 8106 3853 8140
rect 3887 8106 3921 8140
rect 3955 8106 3989 8140
rect 4023 8106 4057 8140
rect 4091 8106 4125 8140
rect 4159 8106 4193 8140
rect 4227 8106 4261 8140
rect 4295 8106 4329 8140
rect 4363 8106 4397 8140
rect 4431 8106 4465 8140
rect 4499 8106 4533 8140
rect 4567 8106 4601 8140
rect 4635 8106 4669 8140
rect 4703 8106 4737 8140
rect 4771 8106 4805 8140
rect 4839 8106 4873 8140
rect 4907 8106 4941 8140
rect 4975 8106 5009 8140
rect 5043 8106 5077 8140
rect 5111 8106 5145 8140
rect 5179 8106 5213 8140
rect 5247 8106 5281 8140
rect 5315 8106 5349 8140
rect 5383 8106 5417 8140
rect 5451 8106 5485 8140
rect 5519 8106 5553 8140
rect 5587 8106 5621 8140
rect 5655 8106 5689 8140
rect 5723 8106 5757 8140
rect 5791 8106 5825 8140
rect 5859 8106 5893 8140
rect 5927 8106 5961 8140
rect 5995 8106 6029 8140
rect 6063 8106 6097 8140
rect 6131 8106 6165 8140
rect 6199 8106 6233 8140
rect 6267 8106 6301 8140
rect 6335 8106 6369 8140
rect 6403 8106 6437 8140
rect 6471 8106 6505 8140
rect 6539 8106 6573 8140
rect 6607 8106 6641 8140
rect 6675 8106 6709 8140
rect 6743 8106 6777 8140
rect 6811 8106 6845 8140
rect 6879 8106 6913 8140
rect 6947 8106 6981 8140
rect 7015 8106 7049 8140
rect 7083 8106 7117 8140
rect 7151 8106 7185 8140
rect 7219 8106 7253 8140
rect 7287 8106 7321 8140
rect 7355 8106 7389 8140
rect 7423 8106 7457 8140
rect 7491 8106 7525 8140
rect 7559 8106 7593 8140
rect 7627 8106 7661 8140
rect 7695 8106 7729 8140
rect 7763 8106 7797 8140
rect 7831 8106 7865 8140
rect 7899 8106 7933 8140
rect 7967 8106 8001 8140
rect 8035 8106 8069 8140
rect 8103 8106 8137 8140
rect 8171 8106 8205 8140
rect 8239 8106 8273 8140
rect 8307 8106 8341 8140
rect 68 8048 102 8082
rect 138 8048 172 8082
rect 208 8048 242 8082
rect 278 8048 312 8082
rect 348 8048 382 8082
rect 418 8048 452 8082
rect 488 8048 522 8082
rect 558 8048 592 8082
rect 628 8048 662 8082
rect 698 8048 732 8082
rect 768 8048 802 8082
rect 838 8048 872 8082
rect 908 8048 942 8082
rect 978 8048 1012 8082
rect 1048 8048 1082 8082
rect 1118 8048 1152 8082
rect 1188 8048 1222 8082
rect 1258 8048 1292 8082
rect 1328 8048 1362 8082
rect 1398 8048 1432 8082
rect 1467 8048 1501 8082
rect 1536 8048 1570 8082
rect 1605 8048 1639 8082
rect 1674 8048 1708 8082
rect 1743 8048 1777 8082
rect 1812 8048 1846 8082
rect 1881 8048 1915 8082
rect 1950 8048 1984 8082
rect 2019 8048 2053 8082
rect 2088 8048 2122 8082
rect 2157 8048 2191 8082
rect 2226 8048 2260 8082
rect 2295 8048 2329 8082
rect 2364 8048 2398 8082
rect 2433 8048 2467 8082
rect 2502 8048 2536 8082
rect 2571 8048 2605 8082
rect 2640 8048 2674 8082
rect 2709 8048 2743 8082
rect 2778 8048 2812 8082
rect 2847 8048 2881 8082
rect 2933 8036 2967 8070
rect 3002 8036 3036 8070
rect 3071 8036 3105 8070
rect 3139 8036 3173 8070
rect 3207 8036 3241 8070
rect 3275 8036 3309 8070
rect 3343 8036 3377 8070
rect 3411 8036 3445 8070
rect 3479 8036 3513 8070
rect 3547 8036 3581 8070
rect 3615 8036 3649 8070
rect 3683 8036 3717 8070
rect 3751 8036 3785 8070
rect 3819 8036 3853 8070
rect 3887 8036 3921 8070
rect 3955 8036 3989 8070
rect 4023 8036 4057 8070
rect 4091 8036 4125 8070
rect 4159 8036 4193 8070
rect 4227 8036 4261 8070
rect 4295 8036 4329 8070
rect 4363 8036 4397 8070
rect 4431 8036 4465 8070
rect 4499 8036 4533 8070
rect 4567 8036 4601 8070
rect 4635 8036 4669 8070
rect 4703 8036 4737 8070
rect 4771 8036 4805 8070
rect 4839 8036 4873 8070
rect 4907 8036 4941 8070
rect 4975 8036 5009 8070
rect 5043 8036 5077 8070
rect 5111 8036 5145 8070
rect 5179 8036 5213 8070
rect 5247 8036 5281 8070
rect 5315 8036 5349 8070
rect 5383 8036 5417 8070
rect 5451 8036 5485 8070
rect 5519 8036 5553 8070
rect 5587 8036 5621 8070
rect 5655 8036 5689 8070
rect 5723 8036 5757 8070
rect 5791 8036 5825 8070
rect 5859 8036 5893 8070
rect 5927 8036 5961 8070
rect 5995 8036 6029 8070
rect 6063 8036 6097 8070
rect 6131 8036 6165 8070
rect 6199 8036 6233 8070
rect 6267 8036 6301 8070
rect 6335 8036 6369 8070
rect 6403 8036 6437 8070
rect 6471 8036 6505 8070
rect 6539 8036 6573 8070
rect 6607 8036 6641 8070
rect 6675 8036 6709 8070
rect 6743 8036 6777 8070
rect 6811 8036 6845 8070
rect 6879 8036 6913 8070
rect 6947 8036 6981 8070
rect 7015 8036 7049 8070
rect 7083 8036 7117 8070
rect 7151 8036 7185 8070
rect 7219 8036 7253 8070
rect 7287 8036 7321 8070
rect 7355 8036 7389 8070
rect 7423 8036 7457 8070
rect 7491 8036 7525 8070
rect 7559 8036 7593 8070
rect 7627 8036 7661 8070
rect 7695 8036 7729 8070
rect 7763 8036 7797 8070
rect 7831 8036 7865 8070
rect 7899 8036 7933 8070
rect 7967 8036 8001 8070
rect 8035 8036 8069 8070
rect 8103 8036 8137 8070
rect 8171 8036 8205 8070
rect 8239 8036 8273 8070
rect 8307 8036 8341 8070
rect 68 7973 102 8007
rect 138 7973 172 8007
rect 208 7973 242 8007
rect 278 7973 312 8007
rect 348 7973 382 8007
rect 418 7973 452 8007
rect 488 7973 522 8007
rect 558 7973 592 8007
rect 628 7973 662 8007
rect 698 7973 732 8007
rect 768 7973 802 8007
rect 838 7973 872 8007
rect 908 7973 942 8007
rect 978 7973 1012 8007
rect 1048 7973 1082 8007
rect 1118 7973 1152 8007
rect 1188 7973 1222 8007
rect 1258 7973 1292 8007
rect 1328 7973 1362 8007
rect 1398 7973 1432 8007
rect 1467 7973 1501 8007
rect 1536 7973 1570 8007
rect 1605 7973 1639 8007
rect 1674 7973 1708 8007
rect 1743 7973 1777 8007
rect 1812 7973 1846 8007
rect 1881 7973 1915 8007
rect 1950 7973 1984 8007
rect 2019 7973 2053 8007
rect 2088 7973 2122 8007
rect 2157 7973 2191 8007
rect 2226 7973 2260 8007
rect 2295 7973 2329 8007
rect 2364 7973 2398 8007
rect 2433 7973 2467 8007
rect 2502 7973 2536 8007
rect 2571 7973 2605 8007
rect 2640 7973 2674 8007
rect 2709 7973 2743 8007
rect 2778 7973 2812 8007
rect 2847 7973 2881 8007
rect 2933 7966 2967 8000
rect 3002 7966 3036 8000
rect 3071 7966 3105 8000
rect 3139 7966 3173 8000
rect 3207 7966 3241 8000
rect 3275 7966 3309 8000
rect 3343 7966 3377 8000
rect 3411 7966 3445 8000
rect 3479 7966 3513 8000
rect 3547 7966 3581 8000
rect 3615 7966 3649 8000
rect 3683 7966 3717 8000
rect 3751 7966 3785 8000
rect 3819 7966 3853 8000
rect 3887 7966 3921 8000
rect 3955 7966 3989 8000
rect 4023 7966 4057 8000
rect 4091 7966 4125 8000
rect 4159 7966 4193 8000
rect 4227 7966 4261 8000
rect 4295 7966 4329 8000
rect 4363 7966 4397 8000
rect 4431 7966 4465 8000
rect 4499 7966 4533 8000
rect 4567 7966 4601 8000
rect 4635 7966 4669 8000
rect 4703 7966 4737 8000
rect 4771 7966 4805 8000
rect 4839 7966 4873 8000
rect 4907 7966 4941 8000
rect 4975 7966 5009 8000
rect 5043 7966 5077 8000
rect 5111 7966 5145 8000
rect 5179 7966 5213 8000
rect 5247 7966 5281 8000
rect 5315 7966 5349 8000
rect 5383 7966 5417 8000
rect 5451 7966 5485 8000
rect 5519 7966 5553 8000
rect 5587 7966 5621 8000
rect 5655 7966 5689 8000
rect 5723 7966 5757 8000
rect 5791 7966 5825 8000
rect 5859 7966 5893 8000
rect 5927 7966 5961 8000
rect 5995 7966 6029 8000
rect 6063 7966 6097 8000
rect 6131 7966 6165 8000
rect 6199 7966 6233 8000
rect 6267 7966 6301 8000
rect 6335 7966 6369 8000
rect 6403 7966 6437 8000
rect 6471 7966 6505 8000
rect 6539 7966 6573 8000
rect 6607 7966 6641 8000
rect 6675 7966 6709 8000
rect 6743 7966 6777 8000
rect 6811 7966 6845 8000
rect 6879 7966 6913 8000
rect 6947 7966 6981 8000
rect 7015 7966 7049 8000
rect 7083 7966 7117 8000
rect 7151 7966 7185 8000
rect 7219 7966 7253 8000
rect 7287 7966 7321 8000
rect 7355 7966 7389 8000
rect 7423 7966 7457 8000
rect 7491 7966 7525 8000
rect 7559 7966 7593 8000
rect 7627 7966 7661 8000
rect 7695 7966 7729 8000
rect 7763 7966 7797 8000
rect 7831 7966 7865 8000
rect 7899 7966 7933 8000
rect 7967 7966 8001 8000
rect 8035 7966 8069 8000
rect 8103 7966 8137 8000
rect 8171 7966 8205 8000
rect 8239 7966 8273 8000
rect 8307 7966 8341 8000
rect 68 7898 102 7932
rect 138 7898 172 7932
rect 208 7898 242 7932
rect 278 7898 312 7932
rect 348 7898 382 7932
rect 418 7898 452 7932
rect 488 7898 522 7932
rect 558 7898 592 7932
rect 628 7898 662 7932
rect 698 7898 732 7932
rect 768 7898 802 7932
rect 838 7898 872 7932
rect 908 7898 942 7932
rect 978 7898 1012 7932
rect 1048 7898 1082 7932
rect 1118 7898 1152 7932
rect 1188 7898 1222 7932
rect 1258 7898 1292 7932
rect 1328 7898 1362 7932
rect 1398 7898 1432 7932
rect 1467 7898 1501 7932
rect 1536 7898 1570 7932
rect 1605 7898 1639 7932
rect 1674 7898 1708 7932
rect 1743 7898 1777 7932
rect 1812 7898 1846 7932
rect 1881 7898 1915 7932
rect 1950 7898 1984 7932
rect 2019 7898 2053 7932
rect 2088 7898 2122 7932
rect 2157 7898 2191 7932
rect 2226 7898 2260 7932
rect 2295 7898 2329 7932
rect 2364 7898 2398 7932
rect 2433 7898 2467 7932
rect 2502 7898 2536 7932
rect 2571 7898 2605 7932
rect 2640 7898 2674 7932
rect 2709 7898 2743 7932
rect 2778 7898 2812 7932
rect 2847 7898 2881 7932
rect 2933 7896 2967 7930
rect 3002 7896 3036 7930
rect 3071 7896 3105 7930
rect 3139 7896 3173 7930
rect 3207 7896 3241 7930
rect 3275 7896 3309 7930
rect 3343 7896 3377 7930
rect 3411 7896 3445 7930
rect 3479 7896 3513 7930
rect 3547 7896 3581 7930
rect 3615 7896 3649 7930
rect 3683 7896 3717 7930
rect 3751 7896 3785 7930
rect 3819 7896 3853 7930
rect 3887 7896 3921 7930
rect 3955 7896 3989 7930
rect 4023 7896 4057 7930
rect 4091 7896 4125 7930
rect 4159 7896 4193 7930
rect 4227 7896 4261 7930
rect 4295 7896 4329 7930
rect 4363 7896 4397 7930
rect 4431 7896 4465 7930
rect 4499 7896 4533 7930
rect 4567 7896 4601 7930
rect 4635 7896 4669 7930
rect 4703 7896 4737 7930
rect 4771 7896 4805 7930
rect 4839 7896 4873 7930
rect 4907 7896 4941 7930
rect 4975 7896 5009 7930
rect 5043 7896 5077 7930
rect 5111 7896 5145 7930
rect 5179 7896 5213 7930
rect 5247 7896 5281 7930
rect 5315 7896 5349 7930
rect 5383 7896 5417 7930
rect 5451 7896 5485 7930
rect 5519 7896 5553 7930
rect 5587 7896 5621 7930
rect 5655 7896 5689 7930
rect 5723 7896 5757 7930
rect 5791 7896 5825 7930
rect 5859 7896 5893 7930
rect 5927 7896 5961 7930
rect 5995 7896 6029 7930
rect 6063 7896 6097 7930
rect 6131 7896 6165 7930
rect 6199 7896 6233 7930
rect 6267 7896 6301 7930
rect 6335 7896 6369 7930
rect 6403 7896 6437 7930
rect 6471 7896 6505 7930
rect 6539 7896 6573 7930
rect 6607 7896 6641 7930
rect 6675 7896 6709 7930
rect 6743 7896 6777 7930
rect 6811 7896 6845 7930
rect 6879 7896 6913 7930
rect 6947 7896 6981 7930
rect 7015 7896 7049 7930
rect 7083 7896 7117 7930
rect 7151 7896 7185 7930
rect 7219 7896 7253 7930
rect 7287 7896 7321 7930
rect 7355 7896 7389 7930
rect 7423 7896 7457 7930
rect 7491 7896 7525 7930
rect 7559 7896 7593 7930
rect 7627 7896 7661 7930
rect 7695 7896 7729 7930
rect 7763 7896 7797 7930
rect 7831 7896 7865 7930
rect 7899 7896 7933 7930
rect 7967 7896 8001 7930
rect 8035 7896 8069 7930
rect 8103 7896 8137 7930
rect 8171 7896 8205 7930
rect 8239 7896 8273 7930
rect 8307 7896 8341 7930
rect 13532 8249 13566 8283
rect 13603 8249 13637 8283
rect 13674 8249 13708 8283
rect 13744 8249 13778 8283
rect 13814 8249 13848 8283
rect 13884 8249 13918 8283
rect 13954 8249 13988 8283
rect 14024 8249 14058 8283
rect 14094 8249 14128 8283
rect 14164 8249 14198 8283
rect 14234 8249 14268 8283
rect 14304 8249 14338 8283
rect 14374 8249 14408 8283
rect 14444 8249 14478 8283
rect 14514 8249 14548 8283
rect 14584 8249 14618 8283
rect 14654 8249 14688 8283
rect 14724 8249 14758 8283
rect 14794 8249 14828 8283
rect 14864 8249 14898 8283
rect 14932 8255 14966 8289
rect 15000 8255 15034 8289
rect 15068 8255 15102 8289
rect 13532 8175 13566 8209
rect 13603 8175 13637 8209
rect 13674 8175 13708 8209
rect 13744 8175 13778 8209
rect 13814 8175 13848 8209
rect 13884 8175 13918 8209
rect 13954 8175 13988 8209
rect 14024 8175 14058 8209
rect 14094 8175 14128 8209
rect 14164 8175 14198 8209
rect 14234 8175 14268 8209
rect 14304 8175 14338 8209
rect 14374 8175 14408 8209
rect 14444 8175 14478 8209
rect 14514 8175 14548 8209
rect 14584 8175 14618 8209
rect 14654 8175 14688 8209
rect 14724 8175 14758 8209
rect 14794 8175 14828 8209
rect 14864 8175 14898 8209
rect 14932 8183 14966 8217
rect 15000 8183 15034 8217
rect 15068 8183 15102 8217
rect 13532 8101 13566 8135
rect 13603 8101 13637 8135
rect 13674 8101 13708 8135
rect 13744 8101 13778 8135
rect 13814 8101 13848 8135
rect 13884 8101 13918 8135
rect 13954 8101 13988 8135
rect 14024 8101 14058 8135
rect 14094 8101 14128 8135
rect 14164 8101 14198 8135
rect 14234 8101 14268 8135
rect 14304 8101 14338 8135
rect 14374 8101 14408 8135
rect 14444 8101 14478 8135
rect 14514 8101 14548 8135
rect 14584 8101 14618 8135
rect 14654 8101 14688 8135
rect 14724 8101 14758 8135
rect 14794 8101 14828 8135
rect 14864 8101 14898 8135
rect 14932 8111 14966 8145
rect 15000 8111 15034 8145
rect 15068 8111 15102 8145
rect 13532 8027 13566 8061
rect 13603 8027 13637 8061
rect 13674 8027 13708 8061
rect 13744 8027 13778 8061
rect 13814 8027 13848 8061
rect 13884 8027 13918 8061
rect 13954 8027 13988 8061
rect 14024 8027 14058 8061
rect 14094 8027 14128 8061
rect 14164 8027 14198 8061
rect 14234 8027 14268 8061
rect 14304 8027 14338 8061
rect 14374 8027 14408 8061
rect 14444 8027 14478 8061
rect 14514 8027 14548 8061
rect 14584 8027 14618 8061
rect 14654 8027 14688 8061
rect 14724 8027 14758 8061
rect 14794 8027 14828 8061
rect 14864 8027 14898 8061
rect 14932 8039 14966 8073
rect 15000 8039 15034 8073
rect 15068 8039 15102 8073
rect 13532 7953 13566 7987
rect 13603 7953 13637 7987
rect 13674 7953 13708 7987
rect 13744 7953 13778 7987
rect 13814 7953 13848 7987
rect 13884 7953 13918 7987
rect 13954 7953 13988 7987
rect 14024 7953 14058 7987
rect 14094 7953 14128 7987
rect 14164 7953 14198 7987
rect 14234 7953 14268 7987
rect 14304 7953 14338 7987
rect 14374 7953 14408 7987
rect 14444 7953 14478 7987
rect 14514 7953 14548 7987
rect 14584 7953 14618 7987
rect 14654 7953 14688 7987
rect 14724 7953 14758 7987
rect 14794 7953 14828 7987
rect 14864 7953 14898 7987
rect 14932 7967 14966 8001
rect 15000 7967 15034 8001
rect 15068 7967 15102 8001
rect 68 7823 102 7857
rect 138 7823 172 7857
rect 208 7823 242 7857
rect 278 7823 312 7857
rect 348 7823 382 7857
rect 418 7823 452 7857
rect 488 7823 522 7857
rect 558 7823 592 7857
rect 628 7823 662 7857
rect 698 7823 732 7857
rect 768 7823 802 7857
rect 838 7823 872 7857
rect 908 7823 942 7857
rect 978 7823 1012 7857
rect 1048 7823 1082 7857
rect 1118 7823 1152 7857
rect 1188 7823 1222 7857
rect 1258 7823 1292 7857
rect 1328 7823 1362 7857
rect 1398 7823 1432 7857
rect 1467 7823 1501 7857
rect 1536 7823 1570 7857
rect 1605 7823 1639 7857
rect 1674 7823 1708 7857
rect 1743 7823 1777 7857
rect 1812 7823 1846 7857
rect 1881 7823 1915 7857
rect 1950 7823 1984 7857
rect 2019 7823 2053 7857
rect 2088 7823 2122 7857
rect 2157 7823 2191 7857
rect 2226 7823 2260 7857
rect 2295 7823 2329 7857
rect 2364 7823 2398 7857
rect 2433 7823 2467 7857
rect 2502 7823 2536 7857
rect 2571 7823 2605 7857
rect 2640 7823 2674 7857
rect 2709 7823 2743 7857
rect 2778 7823 2812 7857
rect 2847 7823 2881 7857
rect 2933 7826 2967 7860
rect 3002 7826 3036 7860
rect 3071 7826 3105 7860
rect 3139 7826 3173 7860
rect 3207 7826 3241 7860
rect 3275 7826 3309 7860
rect 3343 7826 3377 7860
rect 3411 7826 3445 7860
rect 3479 7826 3513 7860
rect 3547 7826 3581 7860
rect 3615 7826 3649 7860
rect 3683 7826 3717 7860
rect 3751 7826 3785 7860
rect 3819 7826 3853 7860
rect 3887 7826 3921 7860
rect 3955 7826 3989 7860
rect 4023 7826 4057 7860
rect 4091 7826 4125 7860
rect 4159 7826 4193 7860
rect 4227 7826 4261 7860
rect 4295 7826 4329 7860
rect 4363 7826 4397 7860
rect 4431 7826 4465 7860
rect 4499 7826 4533 7860
rect 4567 7826 4601 7860
rect 4635 7826 4669 7860
rect 4703 7826 4737 7860
rect 4771 7826 4805 7860
rect 4839 7826 4873 7860
rect 4907 7826 4941 7860
rect 4975 7826 5009 7860
rect 5043 7826 5077 7860
rect 5111 7826 5145 7860
rect 5179 7826 5213 7860
rect 5247 7826 5281 7860
rect 5315 7826 5349 7860
rect 5383 7826 5417 7860
rect 5451 7826 5485 7860
rect 5519 7826 5553 7860
rect 5587 7826 5621 7860
rect 5655 7826 5689 7860
rect 5723 7826 5757 7860
rect 5791 7826 5825 7860
rect 5859 7826 5893 7860
rect 5927 7826 5961 7860
rect 5995 7826 6029 7860
rect 6063 7826 6097 7860
rect 6131 7826 6165 7860
rect 6199 7826 6233 7860
rect 6267 7826 6301 7860
rect 6335 7826 6369 7860
rect 6403 7826 6437 7860
rect 6471 7826 6505 7860
rect 6539 7826 6573 7860
rect 6607 7826 6641 7860
rect 6675 7826 6709 7860
rect 6743 7826 6777 7860
rect 6811 7826 6845 7860
rect 6879 7826 6913 7860
rect 6947 7826 6981 7860
rect 7015 7826 7049 7860
rect 7083 7826 7117 7860
rect 7151 7826 7185 7860
rect 7219 7826 7253 7860
rect 7287 7826 7321 7860
rect 7355 7826 7389 7860
rect 7423 7826 7457 7860
rect 7491 7826 7525 7860
rect 7559 7826 7593 7860
rect 7627 7826 7661 7860
rect 7695 7826 7729 7860
rect 7763 7826 7797 7860
rect 7831 7826 7865 7860
rect 7899 7826 7933 7860
rect 7967 7826 8001 7860
rect 8035 7826 8069 7860
rect 8103 7826 8137 7860
rect 8171 7826 8205 7860
rect 8239 7826 8273 7860
rect 8307 7826 8341 7860
rect 13532 7879 13566 7913
rect 13603 7879 13637 7913
rect 13674 7879 13708 7913
rect 13744 7879 13778 7913
rect 13814 7879 13848 7913
rect 13884 7879 13918 7913
rect 13954 7879 13988 7913
rect 14024 7879 14058 7913
rect 14094 7879 14128 7913
rect 14164 7879 14198 7913
rect 14234 7879 14268 7913
rect 14304 7879 14338 7913
rect 14374 7879 14408 7913
rect 14444 7879 14478 7913
rect 14514 7879 14548 7913
rect 14584 7879 14618 7913
rect 14654 7879 14688 7913
rect 14724 7879 14758 7913
rect 14794 7879 14828 7913
rect 14864 7879 14898 7913
rect 14932 7895 14966 7929
rect 15000 7895 15034 7929
rect 15068 7895 15102 7929
rect 13532 7805 13566 7839
rect 13603 7805 13637 7839
rect 13674 7805 13708 7839
rect 13744 7805 13778 7839
rect 13814 7805 13848 7839
rect 13884 7805 13918 7839
rect 13954 7805 13988 7839
rect 14024 7805 14058 7839
rect 14094 7805 14128 7839
rect 14164 7805 14198 7839
rect 14234 7805 14268 7839
rect 14304 7805 14338 7839
rect 14374 7805 14408 7839
rect 14444 7805 14478 7839
rect 14514 7805 14548 7839
rect 14584 7805 14618 7839
rect 14654 7805 14688 7839
rect 14724 7805 14758 7839
rect 14794 7805 14828 7839
rect 14864 7805 14898 7839
rect 14932 7823 14966 7857
rect 15000 7823 15034 7857
rect 15068 7823 15102 7857
rect 14932 7751 14966 7785
rect 15000 7751 15034 7785
rect 15068 7751 15102 7785
rect 68 7715 102 7749
rect 137 7715 171 7749
rect 206 7715 240 7749
rect 275 7715 309 7749
rect 344 7715 378 7749
rect 413 7715 447 7749
rect 482 7715 516 7749
rect 551 7715 585 7749
rect 620 7715 654 7749
rect 689 7715 723 7749
rect 758 7715 792 7749
rect 827 7715 861 7749
rect 896 7715 930 7749
rect 965 7715 999 7749
rect 1034 7715 1068 7749
rect 1103 7715 1137 7749
rect 1172 7715 1206 7749
rect 1241 7715 1275 7749
rect 1310 7715 1344 7749
rect 1379 7715 1413 7749
rect 1448 7715 1482 7749
rect 1517 7715 1551 7749
rect 1586 7715 1620 7749
rect 1655 7715 1689 7749
rect 1724 7715 1758 7749
rect 1793 7715 1827 7749
rect 1862 7715 1896 7749
rect 1931 7715 1965 7749
rect 2000 7715 2034 7749
rect 2069 7715 2103 7749
rect 2138 7715 2172 7749
rect 2207 7715 2241 7749
rect 2276 7715 2310 7749
rect 2345 7715 2379 7749
rect 2414 7715 2448 7749
rect 2483 7715 2517 7749
rect 2552 7715 2586 7749
rect 2621 7715 2655 7749
rect 2690 7715 2724 7749
rect 2759 7715 2793 7749
rect 2828 7715 2862 7749
rect 2896 7715 2930 7749
rect 2964 7715 2998 7749
rect 3032 7715 3066 7749
rect 3100 7715 3134 7749
rect 3168 7715 3202 7749
rect 3236 7715 3270 7749
rect 3304 7715 3338 7749
rect 3372 7715 3406 7749
rect 3440 7715 3474 7749
rect 3508 7715 3542 7749
rect 3576 7715 3610 7749
rect 3644 7715 3678 7749
rect 3712 7715 3746 7749
rect 3780 7715 3814 7749
rect 3848 7715 3882 7749
rect 3916 7715 3950 7749
rect 3984 7715 4018 7749
rect 4052 7715 4086 7749
rect 4120 7715 4154 7749
rect 4188 7715 4222 7749
rect 4256 7715 4290 7749
rect 4324 7715 4358 7749
rect 4392 7715 4426 7749
rect 4460 7715 4494 7749
rect 4528 7715 4562 7749
rect 4596 7715 4630 7749
rect 4664 7715 4698 7749
rect 4732 7715 4766 7749
rect 4800 7715 4834 7749
rect 4868 7715 4902 7749
rect 4936 7715 4970 7749
rect 5004 7715 5038 7749
rect 5072 7715 5106 7749
rect 5140 7715 5174 7749
rect 5208 7715 5242 7749
rect 5276 7715 5310 7749
rect 5344 7715 5378 7749
rect 5412 7715 5446 7749
rect 5480 7715 5514 7749
rect 5548 7715 5582 7749
rect 5616 7715 5650 7749
rect 5684 7715 5718 7749
rect 5752 7715 5786 7749
rect 5820 7715 5854 7749
rect 5888 7715 5922 7749
rect 5956 7715 5990 7749
rect 6024 7715 6058 7749
rect 6092 7715 6126 7749
rect 6160 7715 6194 7749
rect 6228 7715 6262 7749
rect 6296 7715 6330 7749
rect 6364 7715 6398 7749
rect 6432 7715 6466 7749
rect 6500 7715 6534 7749
rect 6568 7715 6602 7749
rect 6636 7715 6670 7749
rect 6704 7715 6738 7749
rect 6772 7715 6806 7749
rect 6840 7715 6874 7749
rect 6908 7715 6942 7749
rect 6976 7715 7010 7749
rect 7044 7715 7078 7749
rect 7112 7715 7146 7749
rect 7180 7715 7214 7749
rect 7248 7715 7282 7749
rect 7316 7715 7350 7749
rect 7384 7715 7418 7749
rect 7452 7715 7486 7749
rect 7520 7715 7554 7749
rect 7588 7715 7622 7749
rect 7656 7715 7690 7749
rect 7724 7715 7758 7749
rect 7792 7715 7826 7749
rect 7860 7715 7894 7749
rect 7928 7715 7962 7749
rect 7996 7715 8030 7749
rect 8064 7715 8098 7749
rect 8132 7715 8166 7749
rect 8200 7715 8234 7749
rect 8268 7715 8302 7749
rect 8336 7715 8370 7749
rect 8404 7715 8438 7749
rect 8472 7715 8506 7749
rect 8540 7715 8574 7749
rect 8608 7715 8642 7749
rect 8676 7715 8710 7749
rect 8744 7715 8778 7749
rect 8812 7715 8846 7749
rect 8880 7715 8914 7749
rect 8948 7715 8982 7749
rect 9016 7715 9050 7749
rect 9084 7715 9118 7749
rect 9152 7715 9186 7749
rect 9220 7715 9254 7749
rect 9288 7715 9322 7749
rect 9356 7715 9390 7749
rect 9424 7715 9458 7749
rect 9492 7715 9526 7749
rect 9560 7715 9594 7749
rect 9628 7715 9662 7749
rect 9696 7715 9730 7749
rect 9764 7715 9798 7749
rect 9832 7715 9866 7749
rect 9900 7715 9934 7749
rect 9968 7715 10002 7749
rect 10036 7715 10070 7749
rect 10104 7715 10138 7749
rect 10172 7715 10206 7749
rect 10240 7715 10274 7749
rect 10308 7715 10342 7749
rect 10376 7715 10410 7749
rect 10444 7715 10478 7749
rect 10512 7715 10546 7749
rect 10580 7715 10614 7749
rect 10648 7715 10682 7749
rect 10716 7715 10750 7749
rect 10784 7715 10818 7749
rect 10852 7715 10886 7749
rect 10920 7715 10954 7749
rect 10988 7715 11022 7749
rect 11056 7715 11090 7749
rect 11124 7715 11158 7749
rect 11192 7715 11226 7749
rect 11260 7715 11294 7749
rect 11328 7715 11362 7749
rect 11396 7715 11430 7749
rect 11464 7715 11498 7749
rect 11532 7715 11566 7749
rect 11600 7715 11634 7749
rect 11668 7715 11702 7749
rect 11736 7715 11770 7749
rect 11804 7715 11838 7749
rect 11872 7715 11906 7749
rect 11940 7715 11974 7749
rect 12008 7715 12042 7749
rect 12076 7715 12110 7749
rect 12144 7715 12178 7749
rect 12212 7715 12246 7749
rect 12280 7715 12314 7749
rect 12348 7715 12382 7749
rect 12416 7715 12450 7749
rect 12484 7715 12518 7749
rect 12552 7715 12586 7749
rect 12620 7715 12654 7749
rect 12688 7715 12722 7749
rect 12756 7715 12790 7749
rect 12824 7715 12858 7749
rect 12892 7715 12926 7749
rect 12960 7715 12994 7749
rect 13028 7715 13062 7749
rect 13096 7715 13130 7749
rect 13164 7715 13198 7749
rect 13232 7715 13266 7749
rect 13300 7715 13334 7749
rect 13368 7715 13402 7749
rect 13436 7715 13470 7749
rect 13504 7715 13538 7749
rect 13572 7715 13606 7749
rect 13640 7715 13674 7749
rect 13708 7715 13742 7749
rect 13776 7715 13810 7749
rect 13844 7715 13878 7749
rect 13912 7715 13946 7749
rect 13980 7715 14014 7749
rect 14048 7715 14082 7749
rect 14116 7715 14150 7749
rect 14184 7715 14218 7749
rect 14252 7715 14286 7749
rect 14320 7715 14354 7749
rect 14388 7715 14422 7749
rect 14456 7715 14490 7749
rect 14524 7715 14558 7749
rect 14592 7715 14626 7749
rect 14660 7715 14694 7749
rect 14728 7715 14762 7749
rect 14796 7715 14830 7749
rect 14864 7715 14898 7749
rect 14932 7679 14966 7713
rect 15000 7679 15034 7713
rect 15068 7679 15102 7713
rect 68 7608 102 7642
rect 137 7608 171 7642
rect 206 7608 240 7642
rect 275 7608 309 7642
rect 344 7608 378 7642
rect 413 7608 447 7642
rect 482 7608 516 7642
rect 551 7608 585 7642
rect 620 7608 654 7642
rect 689 7608 723 7642
rect 758 7608 792 7642
rect 827 7608 861 7642
rect 896 7608 930 7642
rect 965 7608 999 7642
rect 1033 7608 1067 7642
rect 1101 7608 1135 7642
rect 1169 7608 1203 7642
rect 1237 7608 1271 7642
rect 1305 7608 1339 7642
rect 1373 7608 1407 7642
rect 1441 7608 1475 7642
rect 1509 7608 1543 7642
rect 1577 7608 1611 7642
rect 1645 7608 1679 7642
rect 1713 7608 1747 7642
rect 1781 7608 1815 7642
rect 1849 7608 1883 7642
rect 1917 7608 1951 7642
rect 1985 7608 2019 7642
rect 2053 7608 2087 7642
rect 2121 7608 2155 7642
rect 2189 7608 2223 7642
rect 2257 7608 2291 7642
rect 2325 7608 2359 7642
rect 2393 7608 2427 7642
rect 2461 7608 2495 7642
rect 2529 7608 2563 7642
rect 2597 7608 2631 7642
rect 2665 7608 2699 7642
rect 68 7536 102 7570
rect 137 7536 171 7570
rect 206 7536 240 7570
rect 275 7536 309 7570
rect 344 7536 378 7570
rect 413 7536 447 7570
rect 482 7536 516 7570
rect 551 7536 585 7570
rect 620 7536 654 7570
rect 689 7536 723 7570
rect 758 7536 792 7570
rect 827 7536 861 7570
rect 896 7536 930 7570
rect 965 7536 999 7570
rect 1033 7536 1067 7570
rect 1101 7536 1135 7570
rect 1169 7536 1203 7570
rect 1237 7536 1271 7570
rect 1305 7536 1339 7570
rect 1373 7536 1407 7570
rect 1441 7536 1475 7570
rect 1509 7536 1543 7570
rect 1577 7536 1611 7570
rect 1645 7536 1679 7570
rect 1713 7536 1747 7570
rect 1781 7536 1815 7570
rect 1849 7536 1883 7570
rect 1917 7536 1951 7570
rect 1985 7536 2019 7570
rect 2053 7536 2087 7570
rect 2121 7536 2155 7570
rect 2189 7536 2223 7570
rect 2257 7536 2291 7570
rect 2325 7536 2359 7570
rect 2393 7536 2427 7570
rect 2461 7536 2495 7570
rect 2529 7536 2563 7570
rect 2597 7536 2631 7570
rect 2665 7536 2699 7570
rect 68 7464 102 7498
rect 137 7464 171 7498
rect 206 7464 240 7498
rect 275 7464 309 7498
rect 344 7464 378 7498
rect 413 7464 447 7498
rect 482 7464 516 7498
rect 551 7464 585 7498
rect 620 7464 654 7498
rect 689 7464 723 7498
rect 758 7464 792 7498
rect 827 7464 861 7498
rect 896 7464 930 7498
rect 965 7464 999 7498
rect 1033 7464 1067 7498
rect 1101 7464 1135 7498
rect 1169 7464 1203 7498
rect 1237 7464 1271 7498
rect 1305 7464 1339 7498
rect 1373 7464 1407 7498
rect 1441 7464 1475 7498
rect 1509 7464 1543 7498
rect 1577 7464 1611 7498
rect 1645 7464 1679 7498
rect 1713 7464 1747 7498
rect 1781 7464 1815 7498
rect 1849 7464 1883 7498
rect 1917 7464 1951 7498
rect 1985 7464 2019 7498
rect 2053 7464 2087 7498
rect 2121 7464 2155 7498
rect 2189 7464 2223 7498
rect 2257 7464 2291 7498
rect 2325 7464 2359 7498
rect 2393 7464 2427 7498
rect 2461 7464 2495 7498
rect 2529 7464 2563 7498
rect 2597 7464 2631 7498
rect 2665 7464 2699 7498
rect 68 7392 102 7426
rect 137 7392 171 7426
rect 206 7392 240 7426
rect 275 7392 309 7426
rect 344 7392 378 7426
rect 413 7392 447 7426
rect 482 7392 516 7426
rect 551 7392 585 7426
rect 620 7392 654 7426
rect 689 7392 723 7426
rect 758 7392 792 7426
rect 827 7392 861 7426
rect 896 7392 930 7426
rect 965 7392 999 7426
rect 1033 7392 1067 7426
rect 1101 7392 1135 7426
rect 1169 7392 1203 7426
rect 1237 7392 1271 7426
rect 1305 7392 1339 7426
rect 1373 7392 1407 7426
rect 1441 7392 1475 7426
rect 1509 7392 1543 7426
rect 1577 7392 1611 7426
rect 1645 7392 1679 7426
rect 1713 7392 1747 7426
rect 1781 7392 1815 7426
rect 1849 7392 1883 7426
rect 1917 7392 1951 7426
rect 1985 7392 2019 7426
rect 2053 7392 2087 7426
rect 2121 7392 2155 7426
rect 2189 7392 2223 7426
rect 2257 7392 2291 7426
rect 2325 7392 2359 7426
rect 2393 7392 2427 7426
rect 2461 7392 2495 7426
rect 2529 7392 2563 7426
rect 2597 7392 2631 7426
rect 2665 7392 2699 7426
rect 68 7320 102 7354
rect 137 7320 171 7354
rect 206 7320 240 7354
rect 275 7320 309 7354
rect 344 7320 378 7354
rect 413 7320 447 7354
rect 482 7320 516 7354
rect 551 7320 585 7354
rect 620 7320 654 7354
rect 689 7320 723 7354
rect 758 7320 792 7354
rect 827 7320 861 7354
rect 896 7320 930 7354
rect 965 7320 999 7354
rect 1033 7320 1067 7354
rect 1101 7320 1135 7354
rect 1169 7320 1203 7354
rect 1237 7320 1271 7354
rect 1305 7320 1339 7354
rect 1373 7320 1407 7354
rect 1441 7320 1475 7354
rect 1509 7320 1543 7354
rect 1577 7320 1611 7354
rect 1645 7320 1679 7354
rect 1713 7320 1747 7354
rect 1781 7320 1815 7354
rect 1849 7320 1883 7354
rect 1917 7320 1951 7354
rect 1985 7320 2019 7354
rect 2053 7320 2087 7354
rect 2121 7320 2155 7354
rect 2189 7320 2223 7354
rect 2257 7320 2291 7354
rect 2325 7320 2359 7354
rect 2393 7320 2427 7354
rect 2461 7320 2495 7354
rect 2529 7320 2563 7354
rect 2597 7320 2631 7354
rect 2665 7320 2699 7354
rect 12524 7606 12558 7640
rect 12593 7606 12627 7640
rect 12662 7606 12696 7640
rect 12731 7606 12765 7640
rect 12800 7606 12834 7640
rect 12869 7606 12903 7640
rect 12938 7606 12972 7640
rect 13007 7606 13041 7640
rect 13076 7606 13110 7640
rect 13145 7606 13179 7640
rect 13214 7606 13248 7640
rect 13283 7606 13317 7640
rect 13352 7606 13386 7640
rect 13421 7606 13455 7640
rect 13490 7606 13524 7640
rect 13559 7606 13593 7640
rect 13628 7606 13662 7640
rect 13697 7606 13731 7640
rect 13766 7606 13800 7640
rect 13835 7606 13869 7640
rect 13904 7606 13938 7640
rect 13973 7606 14007 7640
rect 14042 7606 14076 7640
rect 14111 7606 14145 7640
rect 14180 7606 14214 7640
rect 14249 7606 14283 7640
rect 14318 7606 14352 7640
rect 14387 7606 14421 7640
rect 14456 7606 14490 7640
rect 14524 7606 14558 7640
rect 14592 7606 14626 7640
rect 14660 7606 14694 7640
rect 14728 7606 14762 7640
rect 14796 7606 14830 7640
rect 14864 7606 14898 7640
rect 14932 7607 14966 7641
rect 15000 7607 15034 7641
rect 15068 7607 15102 7641
rect 12524 7522 12558 7556
rect 12593 7522 12627 7556
rect 12662 7522 12696 7556
rect 12731 7522 12765 7556
rect 12800 7522 12834 7556
rect 12869 7522 12903 7556
rect 12938 7522 12972 7556
rect 13007 7522 13041 7556
rect 13076 7522 13110 7556
rect 13145 7522 13179 7556
rect 13214 7522 13248 7556
rect 13283 7522 13317 7556
rect 13352 7522 13386 7556
rect 13421 7522 13455 7556
rect 13490 7522 13524 7556
rect 13559 7522 13593 7556
rect 13628 7522 13662 7556
rect 13697 7522 13731 7556
rect 13766 7522 13800 7556
rect 13835 7522 13869 7556
rect 13904 7522 13938 7556
rect 13973 7522 14007 7556
rect 14042 7522 14076 7556
rect 14111 7522 14145 7556
rect 14180 7522 14214 7556
rect 14249 7522 14283 7556
rect 14318 7522 14352 7556
rect 14387 7522 14421 7556
rect 14456 7522 14490 7556
rect 14524 7522 14558 7556
rect 14592 7522 14626 7556
rect 14660 7522 14694 7556
rect 14728 7522 14762 7556
rect 14796 7522 14830 7556
rect 14864 7522 14898 7556
rect 14932 7535 14966 7569
rect 15000 7535 15034 7569
rect 15068 7535 15102 7569
rect 12524 7438 12558 7472
rect 12593 7438 12627 7472
rect 12662 7438 12696 7472
rect 12731 7438 12765 7472
rect 12800 7438 12834 7472
rect 12869 7438 12903 7472
rect 12938 7438 12972 7472
rect 13007 7438 13041 7472
rect 13076 7438 13110 7472
rect 13145 7438 13179 7472
rect 13214 7438 13248 7472
rect 13283 7438 13317 7472
rect 13352 7438 13386 7472
rect 13421 7438 13455 7472
rect 13490 7438 13524 7472
rect 13559 7438 13593 7472
rect 13628 7438 13662 7472
rect 13697 7438 13731 7472
rect 13766 7438 13800 7472
rect 13835 7438 13869 7472
rect 13904 7438 13938 7472
rect 13973 7438 14007 7472
rect 14042 7438 14076 7472
rect 14111 7438 14145 7472
rect 14180 7438 14214 7472
rect 14249 7438 14283 7472
rect 14318 7438 14352 7472
rect 14387 7438 14421 7472
rect 14456 7438 14490 7472
rect 14524 7438 14558 7472
rect 14592 7438 14626 7472
rect 14660 7438 14694 7472
rect 14728 7438 14762 7472
rect 14796 7438 14830 7472
rect 14864 7438 14898 7472
rect 14932 7463 14966 7497
rect 15000 7463 15034 7497
rect 15068 7463 15102 7497
rect 14932 7391 14966 7425
rect 15000 7391 15034 7425
rect 15068 7391 15102 7425
rect 12524 7354 12558 7388
rect 12593 7354 12627 7388
rect 12662 7354 12696 7388
rect 12731 7354 12765 7388
rect 12800 7354 12834 7388
rect 12869 7354 12903 7388
rect 12938 7354 12972 7388
rect 13007 7354 13041 7388
rect 13076 7354 13110 7388
rect 13145 7354 13179 7388
rect 13214 7354 13248 7388
rect 13283 7354 13317 7388
rect 13352 7354 13386 7388
rect 13421 7354 13455 7388
rect 13490 7354 13524 7388
rect 13559 7354 13593 7388
rect 13628 7354 13662 7388
rect 13697 7354 13731 7388
rect 13766 7354 13800 7388
rect 13835 7354 13869 7388
rect 13904 7354 13938 7388
rect 13973 7354 14007 7388
rect 14042 7354 14076 7388
rect 14111 7354 14145 7388
rect 14180 7354 14214 7388
rect 14249 7354 14283 7388
rect 14318 7354 14352 7388
rect 14387 7354 14421 7388
rect 14456 7354 14490 7388
rect 14524 7354 14558 7388
rect 14592 7354 14626 7388
rect 14660 7354 14694 7388
rect 14728 7354 14762 7388
rect 14796 7354 14830 7388
rect 14864 7354 14898 7388
rect 14932 7319 14966 7353
rect 15000 7319 15034 7353
rect 15068 7319 15102 7353
rect 68 7248 102 7282
rect 137 7248 171 7282
rect 206 7248 240 7282
rect 275 7248 309 7282
rect 344 7248 378 7282
rect 413 7248 447 7282
rect 482 7248 516 7282
rect 551 7248 585 7282
rect 620 7248 654 7282
rect 689 7248 723 7282
rect 758 7248 792 7282
rect 827 7248 861 7282
rect 896 7248 930 7282
rect 965 7248 999 7282
rect 1033 7248 1067 7282
rect 1101 7248 1135 7282
rect 1169 7248 1203 7282
rect 1237 7248 1271 7282
rect 1305 7248 1339 7282
rect 1373 7248 1407 7282
rect 1441 7248 1475 7282
rect 1509 7248 1543 7282
rect 1577 7248 1611 7282
rect 1645 7248 1679 7282
rect 1713 7248 1747 7282
rect 1781 7248 1815 7282
rect 1849 7248 1883 7282
rect 1917 7248 1951 7282
rect 1985 7248 2019 7282
rect 2053 7248 2087 7282
rect 2121 7248 2155 7282
rect 2189 7248 2223 7282
rect 2257 7248 2291 7282
rect 2325 7248 2359 7282
rect 2393 7248 2427 7282
rect 2461 7248 2495 7282
rect 2529 7248 2563 7282
rect 2597 7248 2631 7282
rect 2665 7248 2699 7282
rect 68 7176 102 7210
rect 137 7176 171 7210
rect 206 7176 240 7210
rect 275 7176 309 7210
rect 344 7176 378 7210
rect 413 7176 447 7210
rect 482 7176 516 7210
rect 551 7176 585 7210
rect 620 7176 654 7210
rect 689 7176 723 7210
rect 758 7176 792 7210
rect 827 7176 861 7210
rect 896 7176 930 7210
rect 965 7176 999 7210
rect 1033 7176 1067 7210
rect 1101 7176 1135 7210
rect 1169 7176 1203 7210
rect 1237 7176 1271 7210
rect 1305 7176 1339 7210
rect 1373 7176 1407 7210
rect 1441 7176 1475 7210
rect 1509 7176 1543 7210
rect 1577 7176 1611 7210
rect 1645 7176 1679 7210
rect 1713 7176 1747 7210
rect 1781 7176 1815 7210
rect 1849 7176 1883 7210
rect 1917 7176 1951 7210
rect 1985 7176 2019 7210
rect 2053 7176 2087 7210
rect 2121 7176 2155 7210
rect 2189 7176 2223 7210
rect 2257 7176 2291 7210
rect 2325 7176 2359 7210
rect 2393 7176 2427 7210
rect 2461 7176 2495 7210
rect 2529 7176 2563 7210
rect 2597 7176 2631 7210
rect 2665 7176 2699 7210
rect 68 7104 102 7138
rect 137 7104 171 7138
rect 206 7104 240 7138
rect 275 7104 309 7138
rect 344 7104 378 7138
rect 413 7104 447 7138
rect 482 7104 516 7138
rect 551 7104 585 7138
rect 620 7104 654 7138
rect 689 7104 723 7138
rect 758 7104 792 7138
rect 827 7104 861 7138
rect 896 7104 930 7138
rect 965 7104 999 7138
rect 1033 7104 1067 7138
rect 1101 7104 1135 7138
rect 1169 7104 1203 7138
rect 1237 7104 1271 7138
rect 1305 7104 1339 7138
rect 1373 7104 1407 7138
rect 1441 7104 1475 7138
rect 1509 7104 1543 7138
rect 1577 7104 1611 7138
rect 1645 7104 1679 7138
rect 1713 7104 1747 7138
rect 1781 7104 1815 7138
rect 1849 7104 1883 7138
rect 1917 7104 1951 7138
rect 1985 7104 2019 7138
rect 2053 7104 2087 7138
rect 2121 7104 2155 7138
rect 2189 7104 2223 7138
rect 2257 7104 2291 7138
rect 2325 7104 2359 7138
rect 2393 7104 2427 7138
rect 2461 7104 2495 7138
rect 2529 7104 2563 7138
rect 2597 7104 2631 7138
rect 2665 7104 2699 7138
rect 68 7032 102 7066
rect 137 7032 171 7066
rect 206 7032 240 7066
rect 275 7032 309 7066
rect 344 7032 378 7066
rect 413 7032 447 7066
rect 482 7032 516 7066
rect 551 7032 585 7066
rect 620 7032 654 7066
rect 689 7032 723 7066
rect 758 7032 792 7066
rect 827 7032 861 7066
rect 896 7032 930 7066
rect 965 7032 999 7066
rect 1033 7032 1067 7066
rect 1101 7032 1135 7066
rect 1169 7032 1203 7066
rect 1237 7032 1271 7066
rect 1305 7032 1339 7066
rect 1373 7032 1407 7066
rect 1441 7032 1475 7066
rect 1509 7032 1543 7066
rect 1577 7032 1611 7066
rect 1645 7032 1679 7066
rect 1713 7032 1747 7066
rect 1781 7032 1815 7066
rect 1849 7032 1883 7066
rect 1917 7032 1951 7066
rect 1985 7032 2019 7066
rect 2053 7032 2087 7066
rect 2121 7032 2155 7066
rect 2189 7032 2223 7066
rect 2257 7032 2291 7066
rect 2325 7032 2359 7066
rect 2393 7032 2427 7066
rect 2461 7032 2495 7066
rect 2529 7032 2563 7066
rect 2597 7032 2631 7066
rect 2665 7032 2699 7066
rect 8210 7248 8244 7282
rect 8279 7248 8313 7282
rect 8348 7248 8382 7282
rect 8417 7248 8451 7282
rect 8486 7248 8520 7282
rect 8555 7248 8589 7282
rect 8624 7248 8658 7282
rect 8693 7248 8727 7282
rect 8762 7248 8796 7282
rect 8831 7248 8865 7282
rect 8900 7248 8934 7282
rect 8969 7248 9003 7282
rect 9038 7248 9072 7282
rect 9107 7248 9141 7282
rect 9176 7248 9210 7282
rect 9245 7248 9279 7282
rect 9314 7248 9348 7282
rect 9383 7248 9417 7282
rect 9452 7248 9486 7282
rect 9521 7248 9555 7282
rect 9590 7248 9624 7282
rect 9659 7248 9693 7282
rect 9728 7248 9762 7282
rect 9797 7248 9831 7282
rect 9866 7248 9900 7282
rect 9935 7248 9969 7282
rect 10004 7248 10038 7282
rect 10073 7248 10107 7282
rect 10142 7248 10176 7282
rect 10211 7248 10245 7282
rect 10280 7248 10314 7282
rect 10349 7248 10383 7282
rect 10418 7248 10452 7282
rect 10487 7248 10521 7282
rect 10556 7248 10590 7282
rect 10625 7248 10659 7282
rect 10694 7248 10728 7282
rect 10763 7248 10797 7282
rect 10832 7248 10866 7282
rect 10901 7248 10935 7282
rect 10970 7248 11004 7282
rect 11039 7248 11073 7282
rect 11108 7248 11142 7282
rect 11177 7248 11211 7282
rect 11246 7248 11280 7282
rect 11315 7248 11349 7282
rect 11384 7248 11418 7282
rect 11453 7248 11487 7282
rect 11522 7248 11556 7282
rect 11591 7248 11625 7282
rect 11660 7248 11694 7282
rect 11729 7248 11763 7282
rect 11798 7248 11832 7282
rect 11867 7248 11901 7282
rect 11936 7248 11970 7282
rect 12005 7248 12039 7282
rect 12074 7248 12108 7282
rect 12143 7248 12177 7282
rect 12212 7248 12246 7282
rect 12280 7248 12314 7282
rect 12348 7248 12382 7282
rect 12416 7248 12450 7282
rect 12484 7248 12518 7282
rect 12552 7248 12586 7282
rect 12620 7248 12654 7282
rect 12688 7248 12722 7282
rect 12756 7248 12790 7282
rect 12824 7248 12858 7282
rect 12892 7248 12926 7282
rect 12960 7248 12994 7282
rect 13028 7248 13062 7282
rect 13096 7248 13130 7282
rect 13164 7248 13198 7282
rect 13232 7248 13266 7282
rect 13300 7248 13334 7282
rect 13368 7248 13402 7282
rect 13436 7248 13470 7282
rect 13504 7248 13538 7282
rect 13572 7248 13606 7282
rect 13640 7248 13674 7282
rect 13708 7248 13742 7282
rect 13776 7248 13810 7282
rect 13844 7248 13878 7282
rect 13912 7248 13946 7282
rect 13980 7248 14014 7282
rect 14048 7248 14082 7282
rect 14116 7248 14150 7282
rect 14184 7248 14218 7282
rect 14252 7248 14286 7282
rect 14320 7248 14354 7282
rect 14388 7248 14422 7282
rect 14456 7248 14490 7282
rect 14524 7248 14558 7282
rect 14592 7248 14626 7282
rect 14660 7248 14694 7282
rect 14728 7248 14762 7282
rect 14796 7248 14830 7282
rect 14864 7248 14898 7282
rect 14932 7247 14966 7281
rect 15000 7247 15034 7281
rect 15068 7247 15102 7281
rect 8210 7176 8244 7210
rect 8279 7176 8313 7210
rect 8348 7176 8382 7210
rect 8417 7176 8451 7210
rect 8486 7176 8520 7210
rect 8555 7176 8589 7210
rect 8624 7176 8658 7210
rect 8693 7176 8727 7210
rect 8762 7176 8796 7210
rect 8831 7176 8865 7210
rect 8900 7176 8934 7210
rect 8969 7176 9003 7210
rect 9038 7176 9072 7210
rect 9107 7176 9141 7210
rect 9176 7176 9210 7210
rect 9245 7176 9279 7210
rect 9314 7176 9348 7210
rect 9383 7176 9417 7210
rect 9452 7176 9486 7210
rect 9521 7176 9555 7210
rect 9590 7176 9624 7210
rect 9659 7176 9693 7210
rect 9728 7176 9762 7210
rect 9797 7176 9831 7210
rect 9866 7176 9900 7210
rect 9935 7176 9969 7210
rect 10004 7176 10038 7210
rect 10073 7176 10107 7210
rect 10142 7176 10176 7210
rect 10211 7176 10245 7210
rect 10280 7176 10314 7210
rect 10349 7176 10383 7210
rect 10418 7176 10452 7210
rect 10487 7176 10521 7210
rect 10556 7176 10590 7210
rect 10625 7176 10659 7210
rect 10694 7176 10728 7210
rect 10763 7176 10797 7210
rect 10832 7176 10866 7210
rect 10901 7176 10935 7210
rect 10970 7176 11004 7210
rect 11039 7176 11073 7210
rect 11108 7176 11142 7210
rect 11177 7176 11211 7210
rect 11246 7176 11280 7210
rect 11315 7176 11349 7210
rect 11384 7176 11418 7210
rect 11453 7176 11487 7210
rect 11522 7176 11556 7210
rect 11591 7176 11625 7210
rect 11660 7176 11694 7210
rect 11729 7176 11763 7210
rect 11798 7176 11832 7210
rect 11867 7176 11901 7210
rect 11936 7176 11970 7210
rect 12005 7176 12039 7210
rect 12074 7176 12108 7210
rect 12143 7176 12177 7210
rect 12212 7176 12246 7210
rect 12280 7176 12314 7210
rect 12348 7176 12382 7210
rect 12416 7176 12450 7210
rect 12484 7176 12518 7210
rect 12552 7176 12586 7210
rect 12620 7176 12654 7210
rect 12688 7176 12722 7210
rect 12756 7176 12790 7210
rect 12824 7176 12858 7210
rect 12892 7176 12926 7210
rect 12960 7176 12994 7210
rect 13028 7176 13062 7210
rect 13096 7176 13130 7210
rect 13164 7176 13198 7210
rect 13232 7176 13266 7210
rect 13300 7176 13334 7210
rect 13368 7176 13402 7210
rect 13436 7176 13470 7210
rect 13504 7176 13538 7210
rect 13572 7176 13606 7210
rect 13640 7176 13674 7210
rect 13708 7176 13742 7210
rect 13776 7176 13810 7210
rect 13844 7176 13878 7210
rect 13912 7176 13946 7210
rect 13980 7176 14014 7210
rect 14048 7176 14082 7210
rect 14116 7176 14150 7210
rect 14184 7176 14218 7210
rect 14252 7176 14286 7210
rect 14320 7176 14354 7210
rect 14388 7176 14422 7210
rect 14456 7176 14490 7210
rect 14524 7176 14558 7210
rect 14592 7176 14626 7210
rect 14660 7176 14694 7210
rect 14728 7176 14762 7210
rect 14796 7176 14830 7210
rect 14864 7176 14898 7210
rect 14932 7175 14966 7209
rect 15000 7175 15034 7209
rect 15068 7175 15102 7209
rect 8210 7104 8244 7138
rect 8279 7104 8313 7138
rect 8348 7104 8382 7138
rect 8417 7104 8451 7138
rect 8486 7104 8520 7138
rect 8555 7104 8589 7138
rect 8624 7104 8658 7138
rect 8693 7104 8727 7138
rect 8762 7104 8796 7138
rect 8831 7104 8865 7138
rect 8900 7104 8934 7138
rect 8969 7104 9003 7138
rect 9038 7104 9072 7138
rect 9107 7104 9141 7138
rect 9176 7104 9210 7138
rect 9245 7104 9279 7138
rect 9314 7104 9348 7138
rect 9383 7104 9417 7138
rect 9452 7104 9486 7138
rect 9521 7104 9555 7138
rect 9590 7104 9624 7138
rect 9659 7104 9693 7138
rect 9728 7104 9762 7138
rect 9797 7104 9831 7138
rect 9866 7104 9900 7138
rect 9935 7104 9969 7138
rect 10004 7104 10038 7138
rect 10073 7104 10107 7138
rect 10142 7104 10176 7138
rect 10211 7104 10245 7138
rect 10280 7104 10314 7138
rect 10349 7104 10383 7138
rect 10418 7104 10452 7138
rect 10487 7104 10521 7138
rect 10556 7104 10590 7138
rect 10625 7104 10659 7138
rect 10694 7104 10728 7138
rect 10763 7104 10797 7138
rect 10832 7104 10866 7138
rect 10901 7104 10935 7138
rect 10970 7104 11004 7138
rect 11039 7104 11073 7138
rect 11108 7104 11142 7138
rect 11177 7104 11211 7138
rect 11246 7104 11280 7138
rect 11315 7104 11349 7138
rect 11384 7104 11418 7138
rect 11453 7104 11487 7138
rect 11522 7104 11556 7138
rect 11591 7104 11625 7138
rect 11660 7104 11694 7138
rect 11729 7104 11763 7138
rect 11798 7104 11832 7138
rect 11867 7104 11901 7138
rect 11936 7104 11970 7138
rect 12005 7104 12039 7138
rect 12074 7104 12108 7138
rect 12143 7104 12177 7138
rect 12212 7104 12246 7138
rect 12280 7104 12314 7138
rect 12348 7104 12382 7138
rect 12416 7104 12450 7138
rect 12484 7104 12518 7138
rect 12552 7104 12586 7138
rect 12620 7104 12654 7138
rect 12688 7104 12722 7138
rect 12756 7104 12790 7138
rect 12824 7104 12858 7138
rect 12892 7104 12926 7138
rect 12960 7104 12994 7138
rect 13028 7104 13062 7138
rect 13096 7104 13130 7138
rect 13164 7104 13198 7138
rect 13232 7104 13266 7138
rect 13300 7104 13334 7138
rect 13368 7104 13402 7138
rect 13436 7104 13470 7138
rect 13504 7104 13538 7138
rect 13572 7104 13606 7138
rect 13640 7104 13674 7138
rect 13708 7104 13742 7138
rect 13776 7104 13810 7138
rect 13844 7104 13878 7138
rect 13912 7104 13946 7138
rect 13980 7104 14014 7138
rect 14048 7104 14082 7138
rect 14116 7104 14150 7138
rect 14184 7104 14218 7138
rect 14252 7104 14286 7138
rect 14320 7104 14354 7138
rect 14388 7104 14422 7138
rect 14456 7104 14490 7138
rect 14524 7104 14558 7138
rect 14592 7104 14626 7138
rect 14660 7104 14694 7138
rect 14728 7104 14762 7138
rect 14796 7104 14830 7138
rect 14864 7104 14898 7138
rect 14932 7103 14966 7137
rect 15000 7103 15034 7137
rect 15068 7103 15102 7137
rect 2757 7013 2791 7047
rect 2825 7013 2859 7047
rect 2893 7013 2927 7047
rect 2961 7013 2995 7047
rect 3029 7013 3063 7047
rect 3097 7013 3131 7047
rect 3165 7013 3199 7047
rect 3233 7013 3267 7047
rect 3301 7013 3335 7047
rect 3369 7013 3403 7047
rect 3437 7013 3471 7047
rect 3505 7013 3539 7047
rect 3573 7013 3607 7047
rect 3641 7013 3675 7047
rect 3709 7013 3743 7047
rect 3777 7013 3811 7047
rect 3845 7013 3879 7047
rect 3913 7013 3947 7047
rect 3981 7013 4015 7047
rect 4049 7013 4083 7047
rect 4117 7013 4151 7047
rect 4185 7013 4219 7047
rect 4253 7013 4287 7047
rect 4321 7013 4355 7047
rect 4389 7013 4423 7047
rect 4457 7013 4491 7047
rect 4525 7013 4559 7047
rect 4593 7013 4627 7047
rect 4661 7013 4695 7047
rect 4729 7013 4763 7047
rect 4797 7013 4831 7047
rect 4865 7013 4899 7047
rect 4933 7013 4967 7047
rect 5001 7013 5035 7047
rect 5069 7013 5103 7047
rect 5137 7013 5171 7047
rect 5205 7013 5239 7047
rect 5273 7013 5307 7047
rect 5341 7013 5375 7047
rect 5409 7013 5443 7047
rect 5477 7013 5511 7047
rect 5545 7013 5579 7047
rect 5613 7013 5647 7047
rect 5681 7013 5715 7047
rect 5749 7013 5783 7047
rect 5817 7013 5851 7047
rect 5885 7013 5919 7047
rect 5953 7013 5987 7047
rect 6021 7013 6055 7047
rect 6089 7013 6123 7047
rect 6157 7013 6191 7047
rect 6225 7013 6259 7047
rect 6293 7013 6327 7047
rect 6361 7013 6395 7047
rect 6429 7013 6463 7047
rect 6497 7013 6531 7047
rect 6565 7013 6599 7047
rect 6633 7013 6667 7047
rect 6701 7013 6735 7047
rect 6769 7013 6803 7047
rect 6837 7013 6871 7047
rect 6905 7013 6939 7047
rect 6973 7013 7007 7047
rect 7041 7013 7075 7047
rect 7109 7013 7143 7047
rect 7177 7013 7211 7047
rect 7245 7013 7279 7047
rect 7313 7013 7347 7047
rect 7381 7013 7415 7047
rect 7449 7013 7483 7047
rect 7517 7013 7551 7047
rect 7585 7013 7619 7047
rect 7653 7013 7687 7047
rect 8210 7032 8244 7066
rect 8279 7032 8313 7066
rect 8348 7032 8382 7066
rect 8417 7032 8451 7066
rect 8486 7032 8520 7066
rect 8555 7032 8589 7066
rect 8624 7032 8658 7066
rect 8693 7032 8727 7066
rect 8762 7032 8796 7066
rect 8831 7032 8865 7066
rect 8900 7032 8934 7066
rect 8969 7032 9003 7066
rect 9038 7032 9072 7066
rect 9107 7032 9141 7066
rect 9176 7032 9210 7066
rect 9245 7032 9279 7066
rect 9314 7032 9348 7066
rect 9383 7032 9417 7066
rect 9452 7032 9486 7066
rect 9521 7032 9555 7066
rect 9590 7032 9624 7066
rect 9659 7032 9693 7066
rect 9728 7032 9762 7066
rect 9797 7032 9831 7066
rect 9866 7032 9900 7066
rect 9935 7032 9969 7066
rect 10004 7032 10038 7066
rect 10073 7032 10107 7066
rect 10142 7032 10176 7066
rect 10211 7032 10245 7066
rect 10280 7032 10314 7066
rect 10349 7032 10383 7066
rect 10418 7032 10452 7066
rect 10487 7032 10521 7066
rect 10556 7032 10590 7066
rect 10625 7032 10659 7066
rect 10694 7032 10728 7066
rect 10763 7032 10797 7066
rect 10832 7032 10866 7066
rect 10901 7032 10935 7066
rect 10970 7032 11004 7066
rect 11039 7032 11073 7066
rect 11108 7032 11142 7066
rect 11177 7032 11211 7066
rect 11246 7032 11280 7066
rect 11315 7032 11349 7066
rect 11384 7032 11418 7066
rect 11453 7032 11487 7066
rect 11522 7032 11556 7066
rect 11591 7032 11625 7066
rect 11660 7032 11694 7066
rect 11729 7032 11763 7066
rect 11798 7032 11832 7066
rect 11867 7032 11901 7066
rect 11936 7032 11970 7066
rect 12005 7032 12039 7066
rect 12074 7032 12108 7066
rect 12143 7032 12177 7066
rect 12212 7032 12246 7066
rect 12280 7032 12314 7066
rect 12348 7032 12382 7066
rect 12416 7032 12450 7066
rect 12484 7032 12518 7066
rect 12552 7032 12586 7066
rect 12620 7032 12654 7066
rect 12688 7032 12722 7066
rect 12756 7032 12790 7066
rect 12824 7032 12858 7066
rect 12892 7032 12926 7066
rect 12960 7032 12994 7066
rect 13028 7032 13062 7066
rect 13096 7032 13130 7066
rect 13164 7032 13198 7066
rect 13232 7032 13266 7066
rect 13300 7032 13334 7066
rect 13368 7032 13402 7066
rect 13436 7032 13470 7066
rect 13504 7032 13538 7066
rect 13572 7032 13606 7066
rect 13640 7032 13674 7066
rect 13708 7032 13742 7066
rect 13776 7032 13810 7066
rect 13844 7032 13878 7066
rect 13912 7032 13946 7066
rect 13980 7032 14014 7066
rect 14048 7032 14082 7066
rect 14116 7032 14150 7066
rect 14184 7032 14218 7066
rect 14252 7032 14286 7066
rect 14320 7032 14354 7066
rect 14388 7032 14422 7066
rect 14456 7032 14490 7066
rect 14524 7032 14558 7066
rect 14592 7032 14626 7066
rect 14660 7032 14694 7066
rect 14728 7032 14762 7066
rect 14796 7032 14830 7066
rect 14864 7032 14898 7066
rect 14932 7031 14966 7065
rect 15000 7031 15034 7065
rect 15068 7031 15102 7065
rect 3597 1031 3631 1065
rect 3666 1031 3700 1065
rect 3735 1031 3769 1065
rect 3804 1031 3838 1065
rect 3873 1031 3907 1065
rect 3942 1031 3976 1065
rect 4011 1031 4045 1065
rect 4080 1031 4114 1065
rect 4149 1031 4183 1065
rect 4218 1031 4252 1065
rect 4287 1031 4321 1065
rect 4356 1031 4390 1065
rect 4425 1031 4459 1065
rect 4494 1031 4528 1065
rect 4563 1031 4597 1065
rect 4632 1031 4666 1065
rect 4701 1031 4735 1065
rect 4770 1031 4804 1065
rect 4839 1031 4873 1065
rect 4908 1031 4942 1065
rect 4977 1031 5011 1065
rect 5046 1031 5080 1065
rect 5115 1031 5149 1065
rect 5184 1031 5218 1065
rect 5253 1031 5287 1065
rect 5322 1031 5356 1065
rect 5392 1031 5426 1065
rect 5462 1031 5496 1065
rect 5532 1031 5566 1065
rect 5602 1031 5636 1065
rect 5672 1031 5706 1065
rect 5742 1031 5776 1065
rect 5812 1031 5846 1065
rect 5882 1031 5916 1065
rect 5952 1031 5986 1065
rect 6022 1031 6056 1065
rect 6092 1031 6126 1065
rect 6162 1031 6196 1065
rect 6232 1031 6266 1065
rect 6302 1031 6336 1065
rect 6372 1031 6406 1065
rect 6442 1031 6476 1065
rect 6512 1031 6546 1065
rect 6582 1031 6616 1065
rect 6652 1031 6686 1065
rect 6722 1031 6756 1065
rect 6790 932 6824 966
rect 6790 811 6824 845
rect 6790 743 6824 777
rect 6790 675 6824 709
rect 6790 607 6824 641
rect 6790 539 6824 573
rect 6790 471 6824 505
rect 6790 403 6824 437
rect 6790 335 6824 369
rect 6790 267 6824 301
rect 3632 175 3666 209
rect 3700 175 3734 209
rect 3768 175 3802 209
rect 3836 175 3870 209
rect 3904 175 3938 209
rect 3972 175 4006 209
rect 4040 175 4074 209
rect 4108 175 4142 209
rect 4176 175 4210 209
rect 4244 175 4278 209
rect 4312 175 4346 209
rect 4380 175 4414 209
rect 4448 175 4482 209
rect 4516 175 4550 209
rect 4584 175 4618 209
rect 4652 175 4686 209
rect 4720 175 4754 209
rect 4788 175 4822 209
rect 4856 175 4890 209
rect 4924 175 4958 209
rect 4992 175 5026 209
rect 5060 175 5094 209
rect 5128 175 5162 209
rect 5196 175 5230 209
rect 5264 175 5298 209
rect 5332 175 5366 209
rect 5400 175 5434 209
rect 5468 175 5502 209
rect 5536 175 5570 209
rect 5604 175 5638 209
rect 5672 175 5706 209
rect 5740 175 5774 209
rect 5808 175 5842 209
rect 5876 175 5910 209
rect 5944 175 5978 209
rect 6012 175 6046 209
rect 6080 175 6114 209
rect 6148 175 6182 209
rect 6216 175 6250 209
rect 6284 175 6318 209
rect 6352 175 6386 209
rect 6420 175 6454 209
rect 6488 175 6522 209
rect 6556 175 6590 209
rect 6624 175 6658 209
rect 6692 175 6726 209
rect 6790 199 6824 233
<< poly >>
rect 756 15140 782 15260
rect 1782 15203 1892 15260
rect 1782 15169 1820 15203
rect 1854 15169 1892 15203
rect 1782 15140 1892 15169
rect 2892 15203 3013 15260
rect 2892 15169 2939 15203
rect 2973 15169 3013 15203
rect 2892 15140 3013 15169
rect 4013 15203 4134 15260
rect 4013 15169 4060 15203
rect 4094 15169 4134 15203
rect 4013 15140 4134 15169
rect 5134 15140 5160 15260
rect 234 8355 421 8388
rect 234 8321 251 8355
rect 285 8321 319 8355
rect 353 8321 387 8355
rect 234 8288 421 8321
rect 2461 8355 2648 8388
rect 2495 8321 2529 8355
rect 2563 8321 2597 8355
rect 2631 8321 2648 8355
rect 2461 8288 2648 8321
rect 8490 8239 8612 8286
rect 8490 7933 8510 8239
rect 8490 7886 8612 7933
rect 9612 8239 9714 8286
rect 9612 7886 9714 7933
rect 10314 8239 10416 8286
rect 10314 7886 10416 7933
rect 10816 8239 10934 8286
rect 10918 7933 10934 8239
rect 10816 7886 10934 7933
rect 3622 885 3726 904
rect 3622 851 3644 885
rect 3678 851 3726 885
rect 3622 813 3726 851
rect 3622 779 3644 813
rect 3678 804 3726 813
rect 5126 865 5256 904
rect 5126 831 5174 865
rect 5208 831 5256 865
rect 5126 804 5256 831
rect 6656 888 6760 904
rect 6656 854 6704 888
rect 6738 854 6760 888
rect 6656 816 6760 854
rect 6656 804 6704 816
rect 3678 779 3700 804
rect 3622 748 3700 779
rect 5152 796 5230 804
rect 5152 762 5174 796
rect 5208 762 5230 796
rect 5152 748 5230 762
rect 6682 782 6704 804
rect 6738 782 6760 816
rect 6682 748 6760 782
rect 3622 741 3726 748
rect 3622 707 3644 741
rect 3678 707 3726 741
rect 3622 670 3726 707
rect 3622 636 3644 670
rect 3678 648 3726 670
rect 5126 727 5256 748
rect 5126 693 5174 727
rect 5208 693 5256 727
rect 5126 658 5256 693
rect 5126 648 5174 658
rect 3678 636 3700 648
rect 3622 599 3700 636
rect 3622 565 3644 599
rect 3678 592 3700 599
rect 5152 624 5174 648
rect 5208 648 5256 658
rect 6656 744 6760 748
rect 6656 710 6704 744
rect 6738 710 6760 744
rect 6656 672 6760 710
rect 6656 648 6704 672
rect 5208 624 5230 648
rect 5152 592 5230 624
rect 6682 638 6704 648
rect 6738 638 6760 672
rect 6682 600 6760 638
rect 6682 592 6704 600
rect 3678 565 3726 592
rect 3622 528 3726 565
rect 3622 494 3644 528
rect 3678 494 3726 528
rect 3622 492 3726 494
rect 5126 590 5256 592
rect 5126 556 5174 590
rect 5208 556 5256 590
rect 5126 522 5256 556
rect 5126 492 5174 522
rect 3622 457 3700 492
rect 3622 423 3644 457
rect 3678 436 3700 457
rect 5152 488 5174 492
rect 5208 492 5256 522
rect 6656 566 6704 592
rect 6738 566 6760 600
rect 6656 528 6760 566
rect 6656 494 6704 528
rect 6738 494 6760 528
rect 6656 492 6760 494
rect 5208 488 5230 492
rect 5152 454 5230 488
rect 5152 436 5174 454
rect 3678 423 3726 436
rect 3622 386 3726 423
rect 3622 352 3644 386
rect 3678 352 3726 386
rect 3622 336 3726 352
rect 5126 420 5174 436
rect 5208 436 5230 454
rect 6682 457 6760 492
rect 6682 436 6704 457
rect 5208 420 5256 436
rect 5126 386 5256 420
rect 5126 352 5174 386
rect 5208 352 5256 386
rect 5126 336 5256 352
rect 6656 423 6704 436
rect 6738 423 6760 457
rect 6656 386 6760 423
rect 6656 352 6704 386
rect 6738 352 6760 386
rect 6656 336 6760 352
<< polycont >>
rect 1820 15169 1854 15203
rect 2939 15169 2973 15203
rect 4060 15169 4094 15203
rect 251 8321 285 8355
rect 319 8321 353 8355
rect 387 8321 421 8355
rect 2461 8321 2495 8355
rect 2529 8321 2563 8355
rect 2597 8321 2631 8355
rect 8510 7933 8612 8239
rect 9612 7933 9714 8239
rect 10314 7933 10416 8239
rect 10816 7933 10918 8239
rect 3644 851 3678 885
rect 3644 779 3678 813
rect 5174 831 5208 865
rect 6704 854 6738 888
rect 5174 762 5208 796
rect 6704 782 6738 816
rect 3644 707 3678 741
rect 3644 636 3678 670
rect 5174 693 5208 727
rect 3644 565 3678 599
rect 5174 624 5208 658
rect 6704 710 6738 744
rect 6704 638 6738 672
rect 3644 494 3678 528
rect 5174 556 5208 590
rect 3644 423 3678 457
rect 5174 488 5208 522
rect 6704 566 6738 600
rect 6704 494 6738 528
rect 3644 352 3678 386
rect 5174 420 5208 454
rect 5174 352 5208 386
rect 6704 423 6738 457
rect 6704 352 6738 386
<< npolyres >>
rect 421 8288 2461 8388
rect 8612 7886 9612 8286
rect 9714 7886 10314 8286
rect 10416 7886 10816 8286
<< locali >>
rect 67 16503 15106 16527
rect 67 16493 14420 16503
rect 14454 16493 14492 16503
rect 14526 16493 14564 16503
rect 14598 16493 14636 16503
rect 14670 16493 14708 16503
rect 14742 16493 14780 16503
rect 14814 16493 14852 16503
rect 14886 16493 14924 16503
rect 67 16459 68 16493
rect 102 16459 131 16493
rect 173 16459 204 16493
rect 244 16459 277 16493
rect 315 16459 350 16493
rect 386 16459 423 16493
rect 478 16459 496 16493
rect 547 16459 569 16493
rect 616 16459 642 16493
rect 685 16459 715 16493
rect 754 16459 788 16493
rect 823 16459 858 16493
rect 895 16459 927 16493
rect 968 16459 996 16493
rect 1041 16459 1065 16493
rect 1113 16459 1134 16493
rect 1185 16459 1203 16493
rect 1257 16459 1272 16493
rect 1329 16459 1341 16493
rect 1401 16459 1410 16493
rect 1473 16459 1479 16493
rect 1545 16459 1548 16493
rect 1582 16459 1583 16493
rect 1651 16459 1655 16493
rect 1720 16459 1727 16493
rect 1789 16459 1799 16493
rect 1858 16459 1871 16493
rect 1927 16459 1943 16493
rect 1996 16459 2015 16493
rect 2065 16459 2087 16493
rect 2134 16459 2159 16493
rect 2203 16459 2231 16493
rect 2272 16459 2303 16493
rect 2341 16459 2375 16493
rect 2410 16459 2445 16493
rect 2481 16459 2514 16493
rect 2553 16459 2583 16493
rect 2625 16459 2652 16493
rect 2697 16459 2721 16493
rect 2769 16459 2790 16493
rect 2841 16459 2859 16493
rect 2913 16459 2928 16493
rect 2985 16459 2996 16493
rect 3057 16459 3064 16493
rect 3129 16459 3132 16493
rect 3166 16459 3167 16493
rect 3234 16459 3239 16493
rect 3302 16459 3311 16493
rect 3370 16459 3383 16493
rect 3438 16459 3455 16493
rect 3506 16459 3527 16493
rect 3574 16459 3599 16493
rect 3642 16459 3671 16493
rect 3710 16459 3743 16493
rect 3778 16459 3812 16493
rect 3849 16459 3880 16493
rect 3921 16459 3948 16493
rect 3993 16459 4016 16493
rect 4065 16459 4084 16493
rect 4137 16459 4152 16493
rect 4209 16459 4220 16493
rect 4281 16459 4288 16493
rect 4353 16459 4356 16493
rect 4390 16459 4391 16493
rect 4458 16459 4463 16493
rect 4526 16459 4535 16493
rect 4594 16459 4607 16493
rect 4662 16459 4679 16493
rect 4730 16459 4751 16493
rect 4798 16459 4823 16493
rect 4866 16459 4895 16493
rect 4934 16459 4967 16493
rect 5002 16459 5036 16493
rect 5073 16459 5104 16493
rect 5145 16459 5172 16493
rect 5217 16459 5240 16493
rect 5289 16459 5308 16493
rect 5361 16459 5376 16493
rect 5433 16459 5444 16493
rect 5505 16459 5512 16493
rect 5577 16459 5580 16493
rect 5614 16459 5615 16493
rect 5682 16459 5687 16493
rect 5750 16459 5759 16493
rect 5818 16459 5831 16493
rect 5886 16459 5903 16493
rect 5954 16459 5975 16493
rect 6022 16459 6047 16493
rect 6090 16459 6119 16493
rect 6158 16459 6191 16493
rect 6226 16459 6260 16493
rect 6297 16459 6328 16493
rect 6369 16459 6396 16493
rect 6441 16459 6464 16493
rect 6513 16459 6532 16493
rect 6585 16459 6600 16493
rect 6657 16459 6668 16493
rect 6729 16459 6736 16493
rect 6801 16459 6804 16493
rect 6838 16459 6839 16493
rect 6906 16459 6911 16493
rect 6974 16459 6983 16493
rect 7042 16459 7055 16493
rect 7110 16459 7127 16493
rect 7178 16459 7199 16493
rect 7246 16459 7271 16493
rect 7314 16459 7343 16493
rect 7382 16459 7415 16493
rect 7450 16459 7484 16493
rect 7521 16459 7552 16493
rect 7593 16459 7620 16493
rect 7665 16459 7688 16493
rect 7737 16459 7756 16493
rect 7809 16459 7824 16493
rect 7881 16459 7892 16493
rect 7953 16459 7960 16493
rect 8025 16459 8028 16493
rect 8062 16459 8063 16493
rect 8130 16459 8135 16493
rect 8198 16459 8207 16493
rect 8266 16459 8279 16493
rect 8334 16459 8351 16493
rect 8402 16459 8423 16493
rect 8470 16459 8495 16493
rect 8538 16459 8567 16493
rect 8606 16459 8639 16493
rect 8674 16459 8708 16493
rect 8745 16459 8776 16493
rect 8817 16459 8844 16493
rect 8889 16459 8912 16493
rect 8961 16459 8980 16493
rect 9033 16459 9048 16493
rect 9105 16459 9116 16493
rect 9177 16459 9184 16493
rect 9249 16459 9252 16493
rect 9286 16459 9287 16493
rect 9354 16459 9359 16493
rect 9422 16459 9431 16493
rect 9490 16459 9503 16493
rect 9558 16459 9575 16493
rect 9626 16459 9647 16493
rect 9694 16459 9719 16493
rect 9762 16459 9791 16493
rect 9830 16459 9863 16493
rect 9898 16459 9932 16493
rect 9969 16459 10000 16493
rect 10041 16459 10068 16493
rect 10113 16459 10136 16493
rect 10185 16459 10204 16493
rect 10257 16459 10272 16493
rect 10329 16459 10340 16493
rect 10401 16459 10408 16493
rect 10473 16459 10476 16493
rect 10510 16459 10511 16493
rect 10578 16459 10583 16493
rect 10646 16459 10655 16493
rect 10714 16459 10727 16493
rect 10782 16459 10799 16493
rect 10850 16459 10871 16493
rect 10918 16459 10943 16493
rect 10986 16459 11015 16493
rect 11054 16459 11087 16493
rect 11122 16459 11156 16493
rect 11193 16459 11224 16493
rect 11265 16459 11292 16493
rect 11337 16459 11360 16493
rect 11409 16459 11428 16493
rect 11481 16459 11496 16493
rect 11553 16459 11564 16493
rect 11625 16459 11632 16493
rect 11697 16459 11700 16493
rect 11734 16459 11735 16493
rect 11802 16459 11807 16493
rect 11870 16459 11879 16493
rect 11938 16459 11951 16493
rect 12006 16459 12023 16493
rect 12074 16459 12095 16493
rect 12142 16459 12167 16493
rect 12210 16459 12239 16493
rect 12278 16459 12311 16493
rect 12346 16459 12380 16493
rect 12417 16459 12448 16493
rect 12489 16459 12516 16493
rect 12561 16459 12584 16493
rect 12633 16459 12652 16493
rect 12705 16459 12720 16493
rect 12777 16459 12788 16493
rect 12849 16459 12856 16493
rect 12921 16459 12924 16493
rect 12958 16459 12959 16493
rect 13026 16459 13031 16493
rect 13094 16459 13103 16493
rect 13162 16459 13175 16493
rect 13230 16459 13247 16493
rect 13298 16459 13319 16493
rect 13366 16459 13391 16493
rect 13434 16459 13463 16493
rect 13502 16459 13535 16493
rect 13570 16459 13604 16493
rect 13641 16459 13672 16493
rect 13713 16459 13740 16493
rect 13785 16459 13808 16493
rect 13857 16459 13876 16493
rect 13929 16459 13944 16493
rect 14001 16459 14012 16493
rect 14073 16459 14080 16493
rect 14145 16459 14148 16493
rect 14182 16459 14183 16493
rect 14250 16459 14255 16493
rect 14318 16459 14327 16493
rect 14386 16459 14399 16493
rect 14454 16469 14471 16493
rect 14526 16469 14543 16493
rect 14598 16469 14615 16493
rect 14670 16469 14687 16493
rect 14742 16469 14759 16493
rect 14814 16469 14831 16493
rect 14886 16469 14903 16493
rect 14958 16469 14996 16503
rect 15030 16469 15068 16503
rect 15102 16469 15106 16503
rect 14433 16459 14471 16469
rect 14505 16459 14543 16469
rect 14577 16459 14615 16469
rect 14649 16459 14687 16469
rect 14721 16459 14759 16469
rect 14793 16459 14831 16469
rect 14865 16459 14903 16469
rect 14937 16459 15106 16469
rect 67 16434 15106 16459
rect 67 16425 14420 16434
rect 67 16405 68 16425
rect 102 16405 139 16425
rect 102 16391 131 16405
rect 173 16391 210 16425
rect 244 16391 281 16425
rect 315 16391 352 16425
rect 386 16423 14420 16425
rect 386 16391 444 16423
rect 93 16371 131 16391
rect 165 16389 444 16391
rect 478 16389 513 16423
rect 547 16389 582 16423
rect 616 16389 651 16423
rect 685 16389 720 16423
rect 754 16389 789 16423
rect 823 16389 858 16423
rect 892 16389 927 16423
rect 961 16389 996 16423
rect 1030 16389 1065 16423
rect 1099 16389 1134 16423
rect 1168 16389 1203 16423
rect 1237 16389 1272 16423
rect 1306 16389 1341 16423
rect 1375 16389 1410 16423
rect 1444 16389 1479 16423
rect 1513 16389 1548 16423
rect 1582 16389 1617 16423
rect 1651 16389 1686 16423
rect 1720 16389 1755 16423
rect 1789 16389 1824 16423
rect 1858 16389 1893 16423
rect 1927 16389 1962 16423
rect 1996 16389 2031 16423
rect 2065 16389 2100 16423
rect 2134 16389 2169 16423
rect 2203 16389 2238 16423
rect 2272 16389 2307 16423
rect 2341 16389 2376 16423
rect 2410 16389 2445 16423
rect 2479 16389 2514 16423
rect 2548 16389 2583 16423
rect 2617 16389 2652 16423
rect 2686 16389 2721 16423
rect 2755 16389 2790 16423
rect 2824 16389 2859 16423
rect 2893 16389 2928 16423
rect 2962 16389 2996 16423
rect 3030 16389 3064 16423
rect 3098 16389 3132 16423
rect 3166 16389 3200 16423
rect 3234 16389 3268 16423
rect 3302 16389 3336 16423
rect 3370 16389 3404 16423
rect 3438 16389 3472 16423
rect 3506 16389 3540 16423
rect 3574 16389 3608 16423
rect 3642 16389 3676 16423
rect 3710 16389 3744 16423
rect 3778 16389 3812 16423
rect 3846 16389 3880 16423
rect 3914 16389 3948 16423
rect 3982 16389 4016 16423
rect 4050 16389 4084 16423
rect 4118 16389 4152 16423
rect 4186 16389 4220 16423
rect 4254 16389 4288 16423
rect 4322 16389 4356 16423
rect 4390 16389 4424 16423
rect 4458 16389 4492 16423
rect 4526 16389 4560 16423
rect 4594 16389 4628 16423
rect 4662 16389 4696 16423
rect 4730 16389 4764 16423
rect 4798 16389 4832 16423
rect 4866 16389 4900 16423
rect 4934 16389 4968 16423
rect 5002 16389 5036 16423
rect 5070 16389 5104 16423
rect 5138 16389 5172 16423
rect 5206 16389 5240 16423
rect 5274 16389 5308 16423
rect 5342 16389 5376 16423
rect 5410 16389 5444 16423
rect 5478 16389 5512 16423
rect 5546 16389 5580 16423
rect 5614 16389 5648 16423
rect 5682 16389 5716 16423
rect 5750 16389 5784 16423
rect 5818 16389 5852 16423
rect 5886 16389 5920 16423
rect 5954 16389 5988 16423
rect 6022 16389 6056 16423
rect 6090 16389 6124 16423
rect 6158 16389 6192 16423
rect 6226 16389 6260 16423
rect 6294 16389 6328 16423
rect 6362 16389 6396 16423
rect 6430 16389 6464 16423
rect 6498 16389 6532 16423
rect 6566 16389 6600 16423
rect 6634 16389 6668 16423
rect 6702 16389 6736 16423
rect 6770 16389 6804 16423
rect 6838 16389 6872 16423
rect 6906 16389 6940 16423
rect 6974 16389 7008 16423
rect 7042 16389 7076 16423
rect 7110 16389 7144 16423
rect 7178 16389 7212 16423
rect 7246 16389 7280 16423
rect 7314 16389 7348 16423
rect 7382 16389 7416 16423
rect 7450 16389 7484 16423
rect 7518 16389 7552 16423
rect 7586 16389 7620 16423
rect 7654 16389 7688 16423
rect 7722 16389 7756 16423
rect 7790 16389 7824 16423
rect 7858 16389 7892 16423
rect 7926 16389 7960 16423
rect 7994 16389 8028 16423
rect 8062 16389 8096 16423
rect 8130 16389 8164 16423
rect 8198 16389 8232 16423
rect 8266 16389 8300 16423
rect 8334 16389 8368 16423
rect 8402 16389 8436 16423
rect 8470 16389 8504 16423
rect 8538 16389 8572 16423
rect 8606 16389 8640 16423
rect 8674 16389 8708 16423
rect 8742 16389 8776 16423
rect 8810 16389 8844 16423
rect 8878 16389 8912 16423
rect 8946 16389 8980 16423
rect 9014 16389 9048 16423
rect 9082 16389 9116 16423
rect 9150 16389 9184 16423
rect 9218 16389 9252 16423
rect 9286 16389 9320 16423
rect 9354 16389 9388 16423
rect 9422 16389 9456 16423
rect 9490 16389 9524 16423
rect 9558 16389 9592 16423
rect 9626 16389 9660 16423
rect 9694 16389 9728 16423
rect 9762 16389 9796 16423
rect 9830 16389 9864 16423
rect 9898 16389 9932 16423
rect 9966 16389 10000 16423
rect 10034 16389 10068 16423
rect 10102 16389 10136 16423
rect 10170 16389 10204 16423
rect 10238 16389 10272 16423
rect 10306 16389 10340 16423
rect 10374 16389 10408 16423
rect 10442 16389 10476 16423
rect 10510 16389 10544 16423
rect 10578 16389 10612 16423
rect 10646 16389 10680 16423
rect 10714 16389 10748 16423
rect 10782 16389 10816 16423
rect 10850 16389 10884 16423
rect 10918 16389 10952 16423
rect 10986 16389 11020 16423
rect 11054 16389 11088 16423
rect 11122 16389 11156 16423
rect 11190 16389 11224 16423
rect 11258 16389 11292 16423
rect 11326 16389 11360 16423
rect 11394 16389 11428 16423
rect 11462 16389 11496 16423
rect 11530 16389 11564 16423
rect 11598 16389 11632 16423
rect 11666 16389 11700 16423
rect 11734 16389 11768 16423
rect 11802 16389 11836 16423
rect 11870 16389 11904 16423
rect 11938 16389 11972 16423
rect 12006 16389 12040 16423
rect 12074 16389 12108 16423
rect 12142 16389 12176 16423
rect 12210 16389 12244 16423
rect 12278 16389 12312 16423
rect 12346 16389 12380 16423
rect 12414 16389 12448 16423
rect 12482 16389 12516 16423
rect 12550 16389 12584 16423
rect 12618 16389 12652 16423
rect 12686 16389 12720 16423
rect 12754 16389 12788 16423
rect 12822 16389 12856 16423
rect 12890 16389 12924 16423
rect 12958 16389 12992 16423
rect 13026 16389 13060 16423
rect 13094 16389 13128 16423
rect 13162 16389 13196 16423
rect 13230 16389 13264 16423
rect 13298 16389 13332 16423
rect 13366 16389 13400 16423
rect 13434 16389 13468 16423
rect 13502 16389 13536 16423
rect 13570 16389 13604 16423
rect 13638 16389 13672 16423
rect 13706 16389 13740 16423
rect 13774 16389 13808 16423
rect 13842 16389 13876 16423
rect 13910 16389 13944 16423
rect 13978 16389 14012 16423
rect 14046 16389 14080 16423
rect 14114 16389 14148 16423
rect 14182 16389 14216 16423
rect 14250 16389 14284 16423
rect 14318 16389 14352 16423
rect 14386 16400 14420 16423
rect 14454 16400 14492 16434
rect 14526 16400 14564 16434
rect 14598 16400 14636 16434
rect 14670 16400 14708 16434
rect 14742 16400 14780 16434
rect 14814 16400 14852 16434
rect 14886 16400 14924 16434
rect 14958 16400 14996 16434
rect 15030 16400 15068 16434
rect 15102 16400 15106 16434
rect 14386 16389 15106 16400
rect 165 16371 15106 16389
rect 67 16365 15106 16371
rect 67 16357 14420 16365
rect 67 16323 68 16357
rect 102 16323 139 16357
rect 173 16323 210 16357
rect 244 16323 281 16357
rect 315 16323 352 16357
rect 386 16353 14420 16357
rect 386 16323 444 16353
rect 67 16319 444 16323
rect 478 16319 513 16353
rect 547 16319 582 16353
rect 616 16319 651 16353
rect 685 16319 720 16353
rect 754 16319 789 16353
rect 823 16319 858 16353
rect 892 16319 927 16353
rect 961 16319 996 16353
rect 1030 16319 1065 16353
rect 1099 16319 1134 16353
rect 1168 16319 1203 16353
rect 1237 16319 1272 16353
rect 1306 16319 1341 16353
rect 1375 16319 1410 16353
rect 1444 16319 1479 16353
rect 1513 16319 1548 16353
rect 1582 16319 1617 16353
rect 1651 16319 1686 16353
rect 1720 16319 1755 16353
rect 1789 16319 1824 16353
rect 1858 16319 1893 16353
rect 1927 16319 1962 16353
rect 1996 16319 2031 16353
rect 2065 16319 2100 16353
rect 2134 16319 2169 16353
rect 2203 16319 2238 16353
rect 2272 16319 2307 16353
rect 2341 16319 2376 16353
rect 2410 16319 2445 16353
rect 2479 16319 2514 16353
rect 2548 16319 2583 16353
rect 2617 16319 2652 16353
rect 2686 16319 2721 16353
rect 2755 16319 2790 16353
rect 2824 16319 2859 16353
rect 2893 16319 2928 16353
rect 2962 16319 2996 16353
rect 3030 16319 3064 16353
rect 3098 16319 3132 16353
rect 3166 16319 3200 16353
rect 3234 16319 3268 16353
rect 3302 16319 3336 16353
rect 3370 16319 3404 16353
rect 3438 16319 3472 16353
rect 3506 16319 3540 16353
rect 3574 16319 3608 16353
rect 3642 16319 3676 16353
rect 3710 16319 3744 16353
rect 3778 16319 3812 16353
rect 3846 16319 3880 16353
rect 3914 16319 3948 16353
rect 3982 16319 4016 16353
rect 4050 16319 4084 16353
rect 4118 16319 4152 16353
rect 4186 16319 4220 16353
rect 4254 16319 4288 16353
rect 4322 16319 4356 16353
rect 4390 16319 4424 16353
rect 4458 16319 4492 16353
rect 4526 16319 4560 16353
rect 4594 16319 4628 16353
rect 4662 16319 4696 16353
rect 4730 16319 4764 16353
rect 4798 16319 4832 16353
rect 4866 16319 4900 16353
rect 4934 16319 4968 16353
rect 5002 16319 5036 16353
rect 5070 16319 5104 16353
rect 5138 16319 5172 16353
rect 5206 16319 5240 16353
rect 5274 16319 5308 16353
rect 5342 16319 5376 16353
rect 5410 16319 5444 16353
rect 5478 16319 5512 16353
rect 5546 16319 5580 16353
rect 5614 16319 5648 16353
rect 5682 16319 5716 16353
rect 5750 16319 5784 16353
rect 5818 16319 5852 16353
rect 5886 16319 5920 16353
rect 5954 16319 5988 16353
rect 6022 16319 6056 16353
rect 6090 16319 6124 16353
rect 6158 16319 6192 16353
rect 6226 16319 6260 16353
rect 6294 16319 6328 16353
rect 6362 16319 6396 16353
rect 6430 16319 6464 16353
rect 6498 16319 6532 16353
rect 6566 16319 6600 16353
rect 6634 16319 6668 16353
rect 6702 16319 6736 16353
rect 6770 16319 6804 16353
rect 6838 16319 6872 16353
rect 6906 16319 6940 16353
rect 6974 16319 7008 16353
rect 7042 16319 7076 16353
rect 7110 16319 7144 16353
rect 7178 16319 7212 16353
rect 7246 16319 7280 16353
rect 7314 16319 7348 16353
rect 7382 16319 7416 16353
rect 7450 16319 7484 16353
rect 7518 16319 7552 16353
rect 7586 16319 7620 16353
rect 7654 16319 7688 16353
rect 7722 16319 7756 16353
rect 7790 16319 7824 16353
rect 7858 16319 7892 16353
rect 7926 16319 7960 16353
rect 7994 16319 8028 16353
rect 8062 16319 8096 16353
rect 8130 16319 8164 16353
rect 8198 16319 8232 16353
rect 8266 16319 8300 16353
rect 8334 16319 8368 16353
rect 8402 16319 8436 16353
rect 8470 16319 8504 16353
rect 8538 16319 8572 16353
rect 8606 16319 8640 16353
rect 8674 16319 8708 16353
rect 8742 16319 8776 16353
rect 8810 16319 8844 16353
rect 8878 16319 8912 16353
rect 8946 16319 8980 16353
rect 9014 16319 9048 16353
rect 9082 16319 9116 16353
rect 9150 16319 9184 16353
rect 9218 16319 9252 16353
rect 9286 16319 9320 16353
rect 9354 16319 9388 16353
rect 9422 16319 9456 16353
rect 9490 16319 9524 16353
rect 9558 16319 9592 16353
rect 9626 16319 9660 16353
rect 9694 16319 9728 16353
rect 9762 16319 9796 16353
rect 9830 16319 9864 16353
rect 9898 16319 9932 16353
rect 9966 16319 10000 16353
rect 10034 16319 10068 16353
rect 10102 16319 10136 16353
rect 10170 16319 10204 16353
rect 10238 16319 10272 16353
rect 10306 16319 10340 16353
rect 10374 16319 10408 16353
rect 10442 16319 10476 16353
rect 10510 16319 10544 16353
rect 10578 16319 10612 16353
rect 10646 16319 10680 16353
rect 10714 16319 10748 16353
rect 10782 16319 10816 16353
rect 10850 16319 10884 16353
rect 10918 16319 10952 16353
rect 10986 16319 11020 16353
rect 11054 16319 11088 16353
rect 11122 16319 11156 16353
rect 11190 16319 11224 16353
rect 11258 16319 11292 16353
rect 11326 16319 11360 16353
rect 11394 16319 11428 16353
rect 11462 16319 11496 16353
rect 11530 16319 11564 16353
rect 11598 16319 11632 16353
rect 11666 16319 11700 16353
rect 11734 16319 11768 16353
rect 11802 16319 11836 16353
rect 11870 16319 11904 16353
rect 11938 16319 11972 16353
rect 12006 16319 12040 16353
rect 12074 16319 12108 16353
rect 12142 16319 12176 16353
rect 12210 16319 12244 16353
rect 12278 16319 12312 16353
rect 12346 16319 12380 16353
rect 12414 16319 12448 16353
rect 12482 16319 12516 16353
rect 12550 16319 12584 16353
rect 12618 16319 12652 16353
rect 12686 16319 12720 16353
rect 12754 16319 12788 16353
rect 12822 16319 12856 16353
rect 12890 16319 12924 16353
rect 12958 16319 12992 16353
rect 13026 16319 13060 16353
rect 13094 16319 13128 16353
rect 13162 16319 13196 16353
rect 13230 16319 13264 16353
rect 13298 16319 13332 16353
rect 13366 16319 13400 16353
rect 13434 16319 13468 16353
rect 13502 16319 13536 16353
rect 13570 16319 13604 16353
rect 13638 16319 13672 16353
rect 13706 16319 13740 16353
rect 13774 16319 13808 16353
rect 13842 16319 13876 16353
rect 13910 16319 13944 16353
rect 13978 16319 14012 16353
rect 14046 16319 14080 16353
rect 14114 16319 14148 16353
rect 14182 16319 14216 16353
rect 14250 16319 14284 16353
rect 14318 16319 14352 16353
rect 14386 16331 14420 16353
rect 14454 16331 14492 16365
rect 14526 16331 14564 16365
rect 14598 16331 14636 16365
rect 14670 16331 14708 16365
rect 14742 16331 14780 16365
rect 14814 16331 14852 16365
rect 14886 16331 14924 16365
rect 14958 16331 14996 16365
rect 15030 16331 15068 16365
rect 15102 16331 15106 16365
rect 14386 16319 15106 16331
rect 67 16296 15106 16319
rect 67 16289 14420 16296
rect 67 16255 68 16289
rect 102 16255 139 16289
rect 173 16255 210 16289
rect 244 16255 281 16289
rect 315 16255 352 16289
rect 386 16283 14420 16289
rect 386 16255 444 16283
rect 67 16249 444 16255
rect 478 16249 513 16283
rect 547 16249 582 16283
rect 616 16249 651 16283
rect 685 16249 720 16283
rect 754 16249 789 16283
rect 823 16249 858 16283
rect 892 16249 927 16283
rect 961 16249 996 16283
rect 1030 16249 1065 16283
rect 1099 16249 1134 16283
rect 1168 16249 1203 16283
rect 1237 16249 1272 16283
rect 1306 16249 1341 16283
rect 1375 16249 1410 16283
rect 1444 16249 1479 16283
rect 1513 16249 1548 16283
rect 1582 16249 1617 16283
rect 1651 16249 1686 16283
rect 1720 16249 1755 16283
rect 1789 16249 1824 16283
rect 1858 16249 1893 16283
rect 1927 16249 1962 16283
rect 1996 16249 2031 16283
rect 2065 16249 2100 16283
rect 2134 16249 2169 16283
rect 2203 16249 2238 16283
rect 2272 16249 2307 16283
rect 2341 16249 2376 16283
rect 2410 16249 2445 16283
rect 2479 16249 2514 16283
rect 2548 16249 2583 16283
rect 2617 16249 2652 16283
rect 2686 16249 2721 16283
rect 2755 16249 2790 16283
rect 2824 16249 2859 16283
rect 2893 16249 2928 16283
rect 2962 16249 2996 16283
rect 3030 16249 3064 16283
rect 3098 16249 3132 16283
rect 3166 16249 3200 16283
rect 3234 16249 3268 16283
rect 3302 16249 3336 16283
rect 3370 16249 3404 16283
rect 3438 16249 3472 16283
rect 3506 16249 3540 16283
rect 3574 16249 3608 16283
rect 3642 16249 3676 16283
rect 3710 16249 3744 16283
rect 3778 16249 3812 16283
rect 3846 16249 3880 16283
rect 3914 16249 3948 16283
rect 3982 16249 4016 16283
rect 4050 16249 4084 16283
rect 4118 16249 4152 16283
rect 4186 16249 4220 16283
rect 4254 16249 4288 16283
rect 4322 16249 4356 16283
rect 4390 16249 4424 16283
rect 4458 16249 4492 16283
rect 4526 16249 4560 16283
rect 4594 16249 4628 16283
rect 4662 16249 4696 16283
rect 4730 16249 4764 16283
rect 4798 16249 4832 16283
rect 4866 16249 4900 16283
rect 4934 16249 4968 16283
rect 5002 16249 5036 16283
rect 5070 16249 5104 16283
rect 5138 16249 5172 16283
rect 5206 16249 5240 16283
rect 5274 16249 5308 16283
rect 5342 16249 5376 16283
rect 5410 16249 5444 16283
rect 5478 16249 5512 16283
rect 5546 16249 5580 16283
rect 5614 16249 5648 16283
rect 5682 16249 5716 16283
rect 5750 16249 5784 16283
rect 5818 16249 5852 16283
rect 5886 16249 5920 16283
rect 5954 16249 5988 16283
rect 6022 16249 6056 16283
rect 6090 16249 6124 16283
rect 6158 16249 6192 16283
rect 6226 16249 6260 16283
rect 6294 16249 6328 16283
rect 6362 16249 6396 16283
rect 6430 16249 6464 16283
rect 6498 16249 6532 16283
rect 6566 16249 6600 16283
rect 6634 16249 6668 16283
rect 6702 16249 6736 16283
rect 6770 16249 6804 16283
rect 6838 16249 6872 16283
rect 6906 16249 6940 16283
rect 6974 16249 7008 16283
rect 7042 16249 7076 16283
rect 7110 16249 7144 16283
rect 7178 16249 7212 16283
rect 7246 16249 7280 16283
rect 7314 16249 7348 16283
rect 7382 16249 7416 16283
rect 7450 16249 7484 16283
rect 7518 16249 7552 16283
rect 7586 16249 7620 16283
rect 7654 16249 7688 16283
rect 7722 16249 7756 16283
rect 7790 16249 7824 16283
rect 7858 16249 7892 16283
rect 7926 16249 7960 16283
rect 7994 16249 8028 16283
rect 8062 16249 8096 16283
rect 8130 16249 8164 16283
rect 8198 16249 8232 16283
rect 8266 16249 8300 16283
rect 8334 16249 8368 16283
rect 8402 16249 8436 16283
rect 8470 16249 8504 16283
rect 8538 16249 8572 16283
rect 8606 16249 8640 16283
rect 8674 16249 8708 16283
rect 8742 16249 8776 16283
rect 8810 16249 8844 16283
rect 8878 16249 8912 16283
rect 8946 16249 8980 16283
rect 9014 16249 9048 16283
rect 9082 16249 9116 16283
rect 9150 16249 9184 16283
rect 9218 16249 9252 16283
rect 9286 16249 9320 16283
rect 9354 16249 9388 16283
rect 9422 16249 9456 16283
rect 9490 16249 9524 16283
rect 9558 16249 9592 16283
rect 9626 16249 9660 16283
rect 9694 16249 9728 16283
rect 9762 16249 9796 16283
rect 9830 16249 9864 16283
rect 9898 16249 9932 16283
rect 9966 16249 10000 16283
rect 10034 16249 10068 16283
rect 10102 16249 10136 16283
rect 10170 16249 10204 16283
rect 10238 16249 10272 16283
rect 10306 16249 10340 16283
rect 10374 16249 10408 16283
rect 10442 16249 10476 16283
rect 10510 16249 10544 16283
rect 10578 16249 10612 16283
rect 10646 16249 10680 16283
rect 10714 16249 10748 16283
rect 10782 16249 10816 16283
rect 10850 16249 10884 16283
rect 10918 16249 10952 16283
rect 10986 16249 11020 16283
rect 11054 16249 11088 16283
rect 11122 16249 11156 16283
rect 11190 16249 11224 16283
rect 11258 16249 11292 16283
rect 11326 16249 11360 16283
rect 11394 16249 11428 16283
rect 11462 16249 11496 16283
rect 11530 16249 11564 16283
rect 11598 16249 11632 16283
rect 11666 16249 11700 16283
rect 11734 16249 11768 16283
rect 11802 16249 11836 16283
rect 11870 16249 11904 16283
rect 11938 16249 11972 16283
rect 12006 16249 12040 16283
rect 12074 16249 12108 16283
rect 12142 16249 12176 16283
rect 12210 16249 12244 16283
rect 12278 16249 12312 16283
rect 12346 16249 12380 16283
rect 12414 16249 12448 16283
rect 12482 16249 12516 16283
rect 12550 16249 12584 16283
rect 12618 16249 12652 16283
rect 12686 16249 12720 16283
rect 12754 16249 12788 16283
rect 12822 16249 12856 16283
rect 12890 16249 12924 16283
rect 12958 16249 12992 16283
rect 13026 16249 13060 16283
rect 13094 16249 13128 16283
rect 13162 16249 13196 16283
rect 13230 16249 13264 16283
rect 13298 16249 13332 16283
rect 13366 16249 13400 16283
rect 13434 16249 13468 16283
rect 13502 16249 13536 16283
rect 13570 16249 13604 16283
rect 13638 16249 13672 16283
rect 13706 16249 13740 16283
rect 13774 16249 13808 16283
rect 13842 16249 13876 16283
rect 13910 16249 13944 16283
rect 13978 16249 14012 16283
rect 14046 16249 14080 16283
rect 14114 16249 14148 16283
rect 14182 16249 14216 16283
rect 14250 16249 14284 16283
rect 14318 16249 14352 16283
rect 14386 16262 14420 16283
rect 14454 16262 14492 16296
rect 14526 16262 14564 16296
rect 14598 16262 14636 16296
rect 14670 16262 14708 16296
rect 14742 16262 14780 16296
rect 14814 16262 14852 16296
rect 14886 16262 14924 16296
rect 14958 16262 14996 16296
rect 15030 16262 15068 16296
rect 15102 16262 15106 16296
rect 14386 16249 15106 16262
rect 67 16227 15106 16249
rect 67 16221 14420 16227
rect 67 16187 68 16221
rect 102 16187 139 16221
rect 173 16187 210 16221
rect 244 16187 281 16221
rect 315 16187 352 16221
rect 386 16213 14420 16221
rect 386 16187 444 16213
rect 67 16179 444 16187
rect 478 16179 513 16213
rect 547 16179 582 16213
rect 616 16179 651 16213
rect 685 16179 720 16213
rect 754 16179 789 16213
rect 823 16179 858 16213
rect 892 16179 927 16213
rect 961 16179 996 16213
rect 1030 16179 1065 16213
rect 1099 16179 1134 16213
rect 1168 16179 1203 16213
rect 1237 16179 1272 16213
rect 1306 16179 1341 16213
rect 1375 16179 1410 16213
rect 1444 16179 1479 16213
rect 1513 16179 1548 16213
rect 1582 16179 1617 16213
rect 1651 16179 1686 16213
rect 1720 16179 1755 16213
rect 1789 16179 1824 16213
rect 1858 16179 1893 16213
rect 1927 16179 1962 16213
rect 1996 16179 2031 16213
rect 2065 16179 2100 16213
rect 2134 16179 2169 16213
rect 2203 16179 2238 16213
rect 2272 16179 2307 16213
rect 2341 16179 2376 16213
rect 2410 16179 2445 16213
rect 2479 16179 2514 16213
rect 2548 16179 2583 16213
rect 2617 16179 2652 16213
rect 2686 16179 2721 16213
rect 2755 16179 2790 16213
rect 2824 16179 2859 16213
rect 2893 16179 2928 16213
rect 2962 16179 2996 16213
rect 3030 16179 3064 16213
rect 3098 16179 3132 16213
rect 3166 16179 3200 16213
rect 3234 16179 3268 16213
rect 3302 16179 3336 16213
rect 3370 16179 3404 16213
rect 3438 16179 3472 16213
rect 3506 16179 3540 16213
rect 3574 16179 3608 16213
rect 3642 16179 3676 16213
rect 3710 16179 3744 16213
rect 3778 16179 3812 16213
rect 3846 16179 3880 16213
rect 3914 16179 3948 16213
rect 3982 16179 4016 16213
rect 4050 16179 4084 16213
rect 4118 16179 4152 16213
rect 4186 16179 4220 16213
rect 4254 16179 4288 16213
rect 4322 16179 4356 16213
rect 4390 16179 4424 16213
rect 4458 16179 4492 16213
rect 4526 16179 4560 16213
rect 4594 16179 4628 16213
rect 4662 16179 4696 16213
rect 4730 16179 4764 16213
rect 4798 16179 4832 16213
rect 4866 16179 4900 16213
rect 4934 16179 4968 16213
rect 5002 16179 5036 16213
rect 5070 16179 5104 16213
rect 5138 16179 5172 16213
rect 5206 16179 5240 16213
rect 5274 16179 5308 16213
rect 5342 16179 5376 16213
rect 5410 16179 5444 16213
rect 5478 16179 5512 16213
rect 5546 16179 5580 16213
rect 5614 16179 5648 16213
rect 5682 16179 5716 16213
rect 5750 16179 5784 16213
rect 5818 16179 5852 16213
rect 5886 16179 5920 16213
rect 5954 16179 5988 16213
rect 6022 16179 6056 16213
rect 6090 16179 6124 16213
rect 6158 16179 6192 16213
rect 6226 16179 6260 16213
rect 6294 16179 6328 16213
rect 6362 16179 6396 16213
rect 6430 16179 6464 16213
rect 6498 16179 6532 16213
rect 6566 16179 6600 16213
rect 6634 16179 6668 16213
rect 6702 16179 6736 16213
rect 6770 16179 6804 16213
rect 6838 16179 6872 16213
rect 6906 16179 6940 16213
rect 6974 16179 7008 16213
rect 7042 16179 7076 16213
rect 7110 16179 7144 16213
rect 7178 16179 7212 16213
rect 7246 16179 7280 16213
rect 7314 16179 7348 16213
rect 7382 16179 7416 16213
rect 7450 16179 7484 16213
rect 7518 16179 7552 16213
rect 7586 16179 7620 16213
rect 7654 16179 7688 16213
rect 7722 16179 7756 16213
rect 7790 16179 7824 16213
rect 7858 16179 7892 16213
rect 7926 16179 7960 16213
rect 7994 16179 8028 16213
rect 8062 16179 8096 16213
rect 8130 16179 8164 16213
rect 8198 16179 8232 16213
rect 8266 16179 8300 16213
rect 8334 16179 8368 16213
rect 8402 16179 8436 16213
rect 8470 16179 8504 16213
rect 8538 16179 8572 16213
rect 8606 16179 8640 16213
rect 8674 16179 8708 16213
rect 8742 16179 8776 16213
rect 8810 16179 8844 16213
rect 8878 16179 8912 16213
rect 8946 16179 8980 16213
rect 9014 16179 9048 16213
rect 9082 16179 9116 16213
rect 9150 16179 9184 16213
rect 9218 16179 9252 16213
rect 9286 16179 9320 16213
rect 9354 16179 9388 16213
rect 9422 16179 9456 16213
rect 9490 16179 9524 16213
rect 9558 16179 9592 16213
rect 9626 16179 9660 16213
rect 9694 16179 9728 16213
rect 9762 16179 9796 16213
rect 9830 16179 9864 16213
rect 9898 16179 9932 16213
rect 9966 16179 10000 16213
rect 10034 16179 10068 16213
rect 10102 16179 10136 16213
rect 10170 16179 10204 16213
rect 10238 16179 10272 16213
rect 10306 16179 10340 16213
rect 10374 16179 10408 16213
rect 10442 16179 10476 16213
rect 10510 16179 10544 16213
rect 10578 16179 10612 16213
rect 10646 16179 10680 16213
rect 10714 16179 10748 16213
rect 10782 16179 10816 16213
rect 10850 16179 10884 16213
rect 10918 16179 10952 16213
rect 10986 16179 11020 16213
rect 11054 16179 11088 16213
rect 11122 16179 11156 16213
rect 11190 16179 11224 16213
rect 11258 16179 11292 16213
rect 11326 16179 11360 16213
rect 11394 16179 11428 16213
rect 11462 16179 11496 16213
rect 11530 16179 11564 16213
rect 11598 16179 11632 16213
rect 11666 16179 11700 16213
rect 11734 16179 11768 16213
rect 11802 16179 11836 16213
rect 11870 16179 11904 16213
rect 11938 16179 11972 16213
rect 12006 16179 12040 16213
rect 12074 16179 12108 16213
rect 12142 16179 12176 16213
rect 12210 16179 12244 16213
rect 12278 16179 12312 16213
rect 12346 16179 12380 16213
rect 12414 16179 12448 16213
rect 12482 16179 12516 16213
rect 12550 16179 12584 16213
rect 12618 16179 12652 16213
rect 12686 16179 12720 16213
rect 12754 16179 12788 16213
rect 12822 16179 12856 16213
rect 12890 16179 12924 16213
rect 12958 16179 12992 16213
rect 13026 16179 13060 16213
rect 13094 16179 13128 16213
rect 13162 16179 13196 16213
rect 13230 16179 13264 16213
rect 13298 16179 13332 16213
rect 13366 16179 13400 16213
rect 13434 16179 13468 16213
rect 13502 16179 13536 16213
rect 13570 16179 13604 16213
rect 13638 16179 13672 16213
rect 13706 16179 13740 16213
rect 13774 16179 13808 16213
rect 13842 16179 13876 16213
rect 13910 16179 13944 16213
rect 13978 16179 14012 16213
rect 14046 16179 14080 16213
rect 14114 16179 14148 16213
rect 14182 16179 14216 16213
rect 14250 16179 14284 16213
rect 14318 16179 14352 16213
rect 14386 16193 14420 16213
rect 14454 16193 14492 16227
rect 14526 16193 14564 16227
rect 14598 16193 14636 16227
rect 14670 16193 14708 16227
rect 14742 16193 14780 16227
rect 14814 16193 14852 16227
rect 14886 16193 14924 16227
rect 14958 16193 14996 16227
rect 15030 16193 15068 16227
rect 15102 16193 15106 16227
rect 14386 16179 15106 16193
rect 67 16158 15106 16179
rect 67 16153 14420 16158
rect 67 16119 68 16153
rect 102 16119 139 16153
rect 173 16119 210 16153
rect 244 16119 281 16153
rect 315 16119 352 16153
rect 386 16143 14420 16153
rect 386 16119 444 16143
rect 67 16109 444 16119
rect 478 16109 513 16143
rect 547 16109 582 16143
rect 616 16109 651 16143
rect 685 16109 720 16143
rect 754 16109 789 16143
rect 823 16109 858 16143
rect 892 16109 927 16143
rect 961 16109 996 16143
rect 1030 16109 1065 16143
rect 1099 16109 1134 16143
rect 1168 16109 1203 16143
rect 1237 16109 1272 16143
rect 1306 16109 1341 16143
rect 1375 16109 1410 16143
rect 1444 16109 1479 16143
rect 1513 16109 1548 16143
rect 1582 16109 1617 16143
rect 1651 16109 1686 16143
rect 1720 16109 1755 16143
rect 1789 16109 1824 16143
rect 1858 16109 1893 16143
rect 1927 16109 1962 16143
rect 1996 16109 2031 16143
rect 2065 16109 2100 16143
rect 2134 16109 2169 16143
rect 2203 16109 2238 16143
rect 2272 16109 2307 16143
rect 2341 16109 2376 16143
rect 2410 16109 2445 16143
rect 2479 16109 2514 16143
rect 2548 16109 2583 16143
rect 2617 16109 2652 16143
rect 2686 16109 2721 16143
rect 2755 16109 2790 16143
rect 2824 16109 2859 16143
rect 2893 16109 2928 16143
rect 2962 16109 2996 16143
rect 3030 16109 3064 16143
rect 3098 16109 3132 16143
rect 3166 16109 3200 16143
rect 3234 16109 3268 16143
rect 3302 16109 3336 16143
rect 3370 16109 3404 16143
rect 3438 16109 3472 16143
rect 3506 16109 3540 16143
rect 3574 16109 3608 16143
rect 3642 16109 3676 16143
rect 3710 16109 3744 16143
rect 3778 16109 3812 16143
rect 3846 16109 3880 16143
rect 3914 16109 3948 16143
rect 3982 16109 4016 16143
rect 4050 16109 4084 16143
rect 4118 16109 4152 16143
rect 4186 16109 4220 16143
rect 4254 16109 4288 16143
rect 4322 16109 4356 16143
rect 4390 16109 4424 16143
rect 4458 16109 4492 16143
rect 4526 16109 4560 16143
rect 4594 16109 4628 16143
rect 4662 16109 4696 16143
rect 4730 16109 4764 16143
rect 4798 16109 4832 16143
rect 4866 16109 4900 16143
rect 4934 16109 4968 16143
rect 5002 16109 5036 16143
rect 5070 16109 5104 16143
rect 5138 16109 5172 16143
rect 5206 16109 5240 16143
rect 5274 16109 5308 16143
rect 5342 16109 5376 16143
rect 5410 16109 5444 16143
rect 5478 16109 5512 16143
rect 5546 16109 5580 16143
rect 5614 16109 5648 16143
rect 5682 16109 5716 16143
rect 5750 16109 5784 16143
rect 5818 16109 5852 16143
rect 5886 16109 5920 16143
rect 5954 16109 5988 16143
rect 6022 16109 6056 16143
rect 6090 16109 6124 16143
rect 6158 16109 6192 16143
rect 6226 16109 6260 16143
rect 6294 16109 6328 16143
rect 6362 16109 6396 16143
rect 6430 16109 6464 16143
rect 6498 16109 6532 16143
rect 6566 16109 6600 16143
rect 6634 16109 6668 16143
rect 6702 16109 6736 16143
rect 6770 16109 6804 16143
rect 6838 16109 6872 16143
rect 6906 16109 6940 16143
rect 6974 16109 7008 16143
rect 7042 16109 7076 16143
rect 7110 16109 7144 16143
rect 7178 16109 7212 16143
rect 7246 16109 7280 16143
rect 7314 16109 7348 16143
rect 7382 16109 7416 16143
rect 7450 16109 7484 16143
rect 7518 16109 7552 16143
rect 7586 16109 7620 16143
rect 7654 16109 7688 16143
rect 7722 16109 7756 16143
rect 7790 16109 7824 16143
rect 7858 16109 7892 16143
rect 7926 16109 7960 16143
rect 7994 16109 8028 16143
rect 8062 16109 8096 16143
rect 8130 16109 8164 16143
rect 8198 16109 8232 16143
rect 8266 16109 8300 16143
rect 8334 16109 8368 16143
rect 8402 16109 8436 16143
rect 8470 16109 8504 16143
rect 8538 16109 8572 16143
rect 8606 16109 8640 16143
rect 8674 16109 8708 16143
rect 8742 16109 8776 16143
rect 8810 16109 8844 16143
rect 8878 16109 8912 16143
rect 8946 16109 8980 16143
rect 9014 16109 9048 16143
rect 9082 16109 9116 16143
rect 9150 16109 9184 16143
rect 9218 16109 9252 16143
rect 9286 16109 9320 16143
rect 9354 16109 9388 16143
rect 9422 16109 9456 16143
rect 9490 16109 9524 16143
rect 9558 16109 9592 16143
rect 9626 16109 9660 16143
rect 9694 16109 9728 16143
rect 9762 16109 9796 16143
rect 9830 16109 9864 16143
rect 9898 16109 9932 16143
rect 9966 16109 10000 16143
rect 10034 16109 10068 16143
rect 10102 16109 10136 16143
rect 10170 16109 10204 16143
rect 10238 16109 10272 16143
rect 10306 16109 10340 16143
rect 10374 16109 10408 16143
rect 10442 16109 10476 16143
rect 10510 16109 10544 16143
rect 10578 16109 10612 16143
rect 10646 16109 10680 16143
rect 10714 16109 10748 16143
rect 10782 16109 10816 16143
rect 10850 16109 10884 16143
rect 10918 16109 10952 16143
rect 10986 16109 11020 16143
rect 11054 16109 11088 16143
rect 11122 16109 11156 16143
rect 11190 16109 11224 16143
rect 11258 16109 11292 16143
rect 11326 16109 11360 16143
rect 11394 16109 11428 16143
rect 11462 16109 11496 16143
rect 11530 16109 11564 16143
rect 11598 16109 11632 16143
rect 11666 16109 11700 16143
rect 11734 16109 11768 16143
rect 11802 16109 11836 16143
rect 11870 16109 11904 16143
rect 11938 16109 11972 16143
rect 12006 16109 12040 16143
rect 12074 16109 12108 16143
rect 12142 16109 12176 16143
rect 12210 16109 12244 16143
rect 12278 16109 12312 16143
rect 12346 16109 12380 16143
rect 12414 16109 12448 16143
rect 12482 16109 12516 16143
rect 12550 16109 12584 16143
rect 12618 16109 12652 16143
rect 12686 16109 12720 16143
rect 12754 16109 12788 16143
rect 12822 16109 12856 16143
rect 12890 16109 12924 16143
rect 12958 16109 12992 16143
rect 13026 16109 13060 16143
rect 13094 16109 13128 16143
rect 13162 16109 13196 16143
rect 13230 16109 13264 16143
rect 13298 16109 13332 16143
rect 13366 16109 13400 16143
rect 13434 16109 13468 16143
rect 13502 16109 13536 16143
rect 13570 16109 13604 16143
rect 13638 16109 13672 16143
rect 13706 16109 13740 16143
rect 13774 16109 13808 16143
rect 13842 16109 13876 16143
rect 13910 16109 13944 16143
rect 13978 16109 14012 16143
rect 14046 16109 14080 16143
rect 14114 16109 14148 16143
rect 14182 16109 14216 16143
rect 14250 16109 14284 16143
rect 14318 16109 14352 16143
rect 14386 16124 14420 16143
rect 14454 16124 14492 16158
rect 14526 16124 14564 16158
rect 14598 16124 14636 16158
rect 14670 16124 14708 16158
rect 14742 16124 14780 16158
rect 14814 16124 14852 16158
rect 14886 16124 14924 16158
rect 14958 16124 14996 16158
rect 15030 16124 15068 16158
rect 15102 16124 15106 16158
rect 14386 16109 15106 16124
rect 67 16089 15106 16109
rect 67 16085 14420 16089
rect 67 16051 68 16085
rect 102 16051 139 16085
rect 173 16051 210 16085
rect 244 16051 281 16085
rect 315 16051 352 16085
rect 386 16073 14420 16085
rect 386 16051 444 16073
rect 67 16039 444 16051
rect 478 16039 513 16073
rect 547 16039 582 16073
rect 616 16039 651 16073
rect 685 16039 720 16073
rect 754 16039 789 16073
rect 823 16039 858 16073
rect 892 16039 927 16073
rect 961 16039 996 16073
rect 1030 16039 1065 16073
rect 1099 16039 1134 16073
rect 1168 16039 1203 16073
rect 1237 16039 1272 16073
rect 1306 16039 1341 16073
rect 1375 16039 1410 16073
rect 1444 16039 1479 16073
rect 1513 16039 1548 16073
rect 1582 16039 1617 16073
rect 1651 16039 1686 16073
rect 1720 16039 1755 16073
rect 1789 16039 1824 16073
rect 1858 16039 1893 16073
rect 1927 16039 1962 16073
rect 1996 16039 2031 16073
rect 2065 16039 2100 16073
rect 2134 16039 2169 16073
rect 2203 16039 2238 16073
rect 2272 16039 2307 16073
rect 2341 16039 2376 16073
rect 2410 16039 2445 16073
rect 2479 16039 2514 16073
rect 2548 16039 2583 16073
rect 2617 16039 2652 16073
rect 2686 16039 2721 16073
rect 2755 16039 2790 16073
rect 2824 16039 2859 16073
rect 2893 16039 2928 16073
rect 2962 16039 2996 16073
rect 3030 16039 3064 16073
rect 3098 16039 3132 16073
rect 3166 16039 3200 16073
rect 3234 16039 3268 16073
rect 3302 16039 3336 16073
rect 3370 16039 3404 16073
rect 3438 16039 3472 16073
rect 3506 16039 3540 16073
rect 3574 16039 3608 16073
rect 3642 16039 3676 16073
rect 3710 16039 3744 16073
rect 3778 16039 3812 16073
rect 3846 16039 3880 16073
rect 3914 16039 3948 16073
rect 3982 16039 4016 16073
rect 4050 16039 4084 16073
rect 4118 16039 4152 16073
rect 4186 16039 4220 16073
rect 4254 16039 4288 16073
rect 4322 16039 4356 16073
rect 4390 16039 4424 16073
rect 4458 16039 4492 16073
rect 4526 16039 4560 16073
rect 4594 16039 4628 16073
rect 4662 16039 4696 16073
rect 4730 16039 4764 16073
rect 4798 16039 4832 16073
rect 4866 16039 4900 16073
rect 4934 16039 4968 16073
rect 5002 16039 5036 16073
rect 5070 16039 5104 16073
rect 5138 16039 5172 16073
rect 5206 16039 5240 16073
rect 5274 16039 5308 16073
rect 5342 16039 5376 16073
rect 5410 16039 5444 16073
rect 5478 16039 5512 16073
rect 5546 16039 5580 16073
rect 5614 16039 5648 16073
rect 5682 16039 5716 16073
rect 5750 16039 5784 16073
rect 5818 16039 5852 16073
rect 5886 16039 5920 16073
rect 5954 16039 5988 16073
rect 6022 16039 6056 16073
rect 6090 16039 6124 16073
rect 6158 16039 6192 16073
rect 6226 16039 6260 16073
rect 6294 16039 6328 16073
rect 6362 16039 6396 16073
rect 6430 16039 6464 16073
rect 6498 16039 6532 16073
rect 6566 16039 6600 16073
rect 6634 16039 6668 16073
rect 6702 16039 6736 16073
rect 6770 16039 6804 16073
rect 6838 16039 6872 16073
rect 6906 16039 6940 16073
rect 6974 16039 7008 16073
rect 7042 16039 7076 16073
rect 7110 16039 7144 16073
rect 7178 16039 7212 16073
rect 7246 16039 7280 16073
rect 7314 16039 7348 16073
rect 7382 16039 7416 16073
rect 7450 16039 7484 16073
rect 7518 16039 7552 16073
rect 7586 16039 7620 16073
rect 7654 16039 7688 16073
rect 7722 16039 7756 16073
rect 7790 16039 7824 16073
rect 7858 16039 7892 16073
rect 7926 16039 7960 16073
rect 7994 16039 8028 16073
rect 8062 16039 8096 16073
rect 8130 16039 8164 16073
rect 8198 16039 8232 16073
rect 8266 16039 8300 16073
rect 8334 16039 8368 16073
rect 8402 16039 8436 16073
rect 8470 16039 8504 16073
rect 8538 16039 8572 16073
rect 8606 16039 8640 16073
rect 8674 16039 8708 16073
rect 8742 16039 8776 16073
rect 8810 16039 8844 16073
rect 8878 16039 8912 16073
rect 8946 16039 8980 16073
rect 9014 16039 9048 16073
rect 9082 16039 9116 16073
rect 9150 16039 9184 16073
rect 9218 16039 9252 16073
rect 9286 16039 9320 16073
rect 9354 16039 9388 16073
rect 9422 16039 9456 16073
rect 9490 16039 9524 16073
rect 9558 16039 9592 16073
rect 9626 16039 9660 16073
rect 9694 16039 9728 16073
rect 9762 16039 9796 16073
rect 9830 16039 9864 16073
rect 9898 16039 9932 16073
rect 9966 16039 10000 16073
rect 10034 16039 10068 16073
rect 10102 16039 10136 16073
rect 10170 16039 10204 16073
rect 10238 16039 10272 16073
rect 10306 16039 10340 16073
rect 10374 16039 10408 16073
rect 10442 16039 10476 16073
rect 10510 16039 10544 16073
rect 10578 16039 10612 16073
rect 10646 16039 10680 16073
rect 10714 16039 10748 16073
rect 10782 16039 10816 16073
rect 10850 16039 10884 16073
rect 10918 16039 10952 16073
rect 10986 16039 11020 16073
rect 11054 16039 11088 16073
rect 11122 16039 11156 16073
rect 11190 16039 11224 16073
rect 11258 16039 11292 16073
rect 11326 16039 11360 16073
rect 11394 16039 11428 16073
rect 11462 16039 11496 16073
rect 11530 16039 11564 16073
rect 11598 16039 11632 16073
rect 11666 16039 11700 16073
rect 11734 16039 11768 16073
rect 11802 16039 11836 16073
rect 11870 16039 11904 16073
rect 11938 16039 11972 16073
rect 12006 16039 12040 16073
rect 12074 16039 12108 16073
rect 12142 16039 12176 16073
rect 12210 16039 12244 16073
rect 12278 16039 12312 16073
rect 12346 16039 12380 16073
rect 12414 16039 12448 16073
rect 12482 16039 12516 16073
rect 12550 16039 12584 16073
rect 12618 16039 12652 16073
rect 12686 16039 12720 16073
rect 12754 16039 12788 16073
rect 12822 16039 12856 16073
rect 12890 16039 12924 16073
rect 12958 16039 12992 16073
rect 13026 16039 13060 16073
rect 13094 16039 13128 16073
rect 13162 16039 13196 16073
rect 13230 16039 13264 16073
rect 13298 16039 13332 16073
rect 13366 16039 13400 16073
rect 13434 16039 13468 16073
rect 13502 16039 13536 16073
rect 13570 16039 13604 16073
rect 13638 16039 13672 16073
rect 13706 16039 13740 16073
rect 13774 16039 13808 16073
rect 13842 16039 13876 16073
rect 13910 16039 13944 16073
rect 13978 16039 14012 16073
rect 14046 16039 14080 16073
rect 14114 16039 14148 16073
rect 14182 16039 14216 16073
rect 14250 16039 14284 16073
rect 14318 16039 14352 16073
rect 14386 16055 14420 16073
rect 14454 16055 14492 16089
rect 14526 16055 14564 16089
rect 14598 16055 14636 16089
rect 14670 16055 14708 16089
rect 14742 16055 14780 16089
rect 14814 16055 14852 16089
rect 14886 16055 14924 16089
rect 14958 16055 14996 16089
rect 15030 16055 15068 16089
rect 15102 16055 15106 16089
rect 14386 16039 15106 16055
rect 67 16020 15106 16039
rect 67 16017 14420 16020
rect 67 15983 68 16017
rect 102 15983 139 16017
rect 173 15983 210 16017
rect 244 15983 281 16017
rect 315 15983 352 16017
rect 386 16003 14420 16017
rect 386 15983 444 16003
rect 67 15969 444 15983
rect 478 15969 513 16003
rect 547 15969 582 16003
rect 616 15969 651 16003
rect 685 15969 720 16003
rect 754 15969 789 16003
rect 823 15969 858 16003
rect 892 15969 927 16003
rect 961 15969 996 16003
rect 1030 15969 1065 16003
rect 1099 15969 1134 16003
rect 1168 15969 1203 16003
rect 1237 15969 1272 16003
rect 1306 15969 1341 16003
rect 1375 15969 1410 16003
rect 1444 15969 1479 16003
rect 1513 15969 1548 16003
rect 1582 15969 1617 16003
rect 1651 15969 1686 16003
rect 1720 15969 1755 16003
rect 1789 15969 1824 16003
rect 1858 15969 1893 16003
rect 1927 15969 1962 16003
rect 1996 15969 2031 16003
rect 2065 15969 2100 16003
rect 2134 15969 2169 16003
rect 2203 15969 2238 16003
rect 2272 15969 2307 16003
rect 2341 15969 2376 16003
rect 2410 15969 2445 16003
rect 2479 15969 2514 16003
rect 2548 15969 2583 16003
rect 2617 15969 2652 16003
rect 2686 15969 2721 16003
rect 2755 15969 2790 16003
rect 2824 15969 2859 16003
rect 2893 15969 2928 16003
rect 2962 15969 2996 16003
rect 3030 15969 3064 16003
rect 3098 15969 3132 16003
rect 3166 15969 3200 16003
rect 3234 15969 3268 16003
rect 3302 15969 3336 16003
rect 3370 15969 3404 16003
rect 3438 15969 3472 16003
rect 3506 15969 3540 16003
rect 3574 15969 3608 16003
rect 3642 15969 3676 16003
rect 3710 15969 3744 16003
rect 3778 15969 3812 16003
rect 3846 15969 3880 16003
rect 3914 15980 3948 16003
rect 3982 15980 4016 16003
rect 4050 15980 4084 16003
rect 4118 15980 4152 16003
rect 4186 15980 4220 16003
rect 4254 15980 4288 16003
rect 4322 15980 4356 16003
rect 3916 15969 3948 15980
rect 3989 15969 4016 15980
rect 4062 15969 4084 15980
rect 4135 15969 4152 15980
rect 4208 15969 4220 15980
rect 4281 15969 4288 15980
rect 4354 15969 4356 15980
rect 4390 15980 4424 16003
rect 4458 15980 4492 16003
rect 4526 15980 4560 16003
rect 4594 15980 4628 16003
rect 4662 15980 4696 16003
rect 4730 15980 4764 16003
rect 4798 15980 4832 16003
rect 4390 15969 4393 15980
rect 4458 15969 4466 15980
rect 4526 15969 4539 15980
rect 4594 15969 4612 15980
rect 4662 15969 4685 15980
rect 4730 15969 4758 15980
rect 4798 15969 4831 15980
rect 4866 15969 4900 16003
rect 4934 15980 4968 16003
rect 5002 15980 5036 16003
rect 5070 15980 5104 16003
rect 5138 15980 5172 16003
rect 5206 15980 5240 16003
rect 5274 15980 5308 16003
rect 4938 15969 4968 15980
rect 5011 15969 5036 15980
rect 5084 15969 5104 15980
rect 5157 15969 5172 15980
rect 5230 15969 5240 15980
rect 5303 15969 5308 15980
rect 5342 15980 5376 16003
rect 67 15949 3882 15969
rect 67 15915 68 15949
rect 102 15915 139 15949
rect 173 15915 210 15949
rect 244 15915 281 15949
rect 315 15915 352 15949
rect 386 15946 3882 15949
rect 3916 15946 3955 15969
rect 3989 15946 4028 15969
rect 4062 15946 4101 15969
rect 4135 15946 4174 15969
rect 4208 15946 4247 15969
rect 4281 15946 4320 15969
rect 4354 15946 4393 15969
rect 4427 15946 4466 15969
rect 4500 15946 4539 15969
rect 4573 15946 4612 15969
rect 4646 15946 4685 15969
rect 4719 15946 4758 15969
rect 4792 15946 4831 15969
rect 4865 15946 4904 15969
rect 4938 15946 4977 15969
rect 5011 15946 5050 15969
rect 5084 15946 5123 15969
rect 5157 15946 5196 15969
rect 5230 15946 5269 15969
rect 5303 15946 5342 15969
rect 5410 15980 5444 16003
rect 5478 15980 5512 16003
rect 5546 15980 5580 16003
rect 5614 15980 5648 16003
rect 5682 15980 5716 16003
rect 5750 15980 5784 16003
rect 5410 15969 5415 15980
rect 5478 15969 5488 15980
rect 5546 15969 5561 15980
rect 5614 15969 5634 15980
rect 5682 15969 5707 15980
rect 5750 15969 5780 15980
rect 5818 15969 5852 16003
rect 5886 15980 5920 16003
rect 5954 15980 5988 16003
rect 6022 15980 6056 16003
rect 6090 15980 6124 16003
rect 6158 15980 6192 16003
rect 6226 15980 6260 16003
rect 6294 15980 6328 16003
rect 5887 15969 5920 15980
rect 5960 15969 5988 15980
rect 6033 15969 6056 15980
rect 6106 15969 6124 15980
rect 6179 15969 6192 15980
rect 6252 15969 6260 15980
rect 6325 15969 6328 15980
rect 6362 15980 6396 16003
rect 6430 15980 6464 16003
rect 6498 15980 6532 16003
rect 6566 15980 6600 16003
rect 6634 15980 6668 16003
rect 6702 15980 6736 16003
rect 6770 15980 6804 16003
rect 6362 15969 6364 15980
rect 6430 15969 6437 15980
rect 6498 15969 6510 15980
rect 6566 15969 6583 15980
rect 6634 15969 6656 15980
rect 6702 15969 6729 15980
rect 6770 15969 6802 15980
rect 6838 15969 6872 16003
rect 6906 15980 6940 16003
rect 6974 15980 7008 16003
rect 7042 15980 7076 16003
rect 7110 15980 7144 16003
rect 7178 15980 7212 16003
rect 7246 15980 7280 16003
rect 7314 15980 7348 16003
rect 6909 15969 6940 15980
rect 6982 15969 7008 15980
rect 7055 15969 7076 15980
rect 7128 15969 7144 15980
rect 7201 15969 7212 15980
rect 7274 15969 7280 15980
rect 7347 15969 7348 15980
rect 7382 15980 7416 16003
rect 7450 15980 7484 16003
rect 7518 15980 7552 16003
rect 7586 15980 7620 16003
rect 7654 15980 7688 16003
rect 7722 15980 7756 16003
rect 7382 15969 7386 15980
rect 7450 15969 7459 15980
rect 7518 15969 7532 15980
rect 7586 15969 7605 15980
rect 7654 15969 7678 15980
rect 7722 15969 7751 15980
rect 7790 15969 7824 16003
rect 7858 15969 7892 16003
rect 7926 15980 7960 16003
rect 7994 15980 8028 16003
rect 8062 15980 8096 16003
rect 8130 15980 8164 16003
rect 8198 15980 8232 16003
rect 8266 15980 8300 16003
rect 7931 15969 7960 15980
rect 8004 15969 8028 15980
rect 8077 15969 8096 15980
rect 8150 15969 8164 15980
rect 8223 15969 8232 15980
rect 8296 15969 8300 15980
rect 8334 15980 8368 16003
rect 8402 15980 8436 16003
rect 8470 15980 8504 16003
rect 8538 15980 8572 16003
rect 8606 15980 8640 16003
rect 8674 15980 8708 16003
rect 8742 15980 8776 16003
rect 8810 15980 8844 16003
rect 8334 15969 8335 15980
rect 8402 15969 8408 15980
rect 8470 15969 8481 15980
rect 8538 15969 8554 15980
rect 8606 15969 8627 15980
rect 8674 15969 8699 15980
rect 8742 15969 8771 15980
rect 8810 15969 8843 15980
rect 8878 15969 8912 16003
rect 8946 15980 8980 16003
rect 9014 15980 9048 16003
rect 9082 15980 9116 16003
rect 9150 15980 9184 16003
rect 9218 15980 9252 16003
rect 9286 15980 9320 16003
rect 9354 15980 9388 16003
rect 9422 15980 9456 16003
rect 8949 15969 8980 15980
rect 9021 15969 9048 15980
rect 9093 15969 9116 15980
rect 9165 15969 9184 15980
rect 9237 15969 9252 15980
rect 9309 15969 9320 15980
rect 9381 15969 9388 15980
rect 9453 15969 9456 15980
rect 9490 15980 9524 16003
rect 9558 15980 9592 16003
rect 9626 15980 9660 16003
rect 9694 15980 9728 16003
rect 9762 15980 9796 16003
rect 9830 15980 9864 16003
rect 9898 15980 9932 16003
rect 9966 15980 10000 16003
rect 10034 15980 10068 16003
rect 9490 15969 9491 15980
rect 9558 15969 9563 15980
rect 9626 15969 9635 15980
rect 9694 15969 9707 15980
rect 9762 15969 9779 15980
rect 9830 15969 9851 15980
rect 9898 15969 9923 15980
rect 9966 15969 9995 15980
rect 10034 15969 10067 15980
rect 10102 15969 10136 16003
rect 10170 15980 10204 16003
rect 10238 15980 10272 16003
rect 10306 15980 10340 16003
rect 10374 15980 10408 16003
rect 10442 15980 10476 16003
rect 10510 15980 10544 16003
rect 10578 15980 10612 16003
rect 10646 15980 10680 16003
rect 10173 15969 10204 15980
rect 10245 15969 10272 15980
rect 10317 15969 10340 15980
rect 10389 15969 10408 15980
rect 10461 15969 10476 15980
rect 10533 15969 10544 15980
rect 10605 15969 10612 15980
rect 10677 15969 10680 15980
rect 10714 15980 10748 16003
rect 10782 15980 10816 16003
rect 10850 15980 10884 16003
rect 10918 15980 10952 16003
rect 10986 15980 11020 16003
rect 11054 15980 11088 16003
rect 11122 15980 11156 16003
rect 11190 15980 11224 16003
rect 11258 15980 11292 16003
rect 10714 15969 10715 15980
rect 10782 15969 10787 15980
rect 10850 15969 10859 15980
rect 10918 15969 10931 15980
rect 10986 15969 11003 15980
rect 11054 15969 11075 15980
rect 11122 15969 11147 15980
rect 11190 15969 11219 15980
rect 11258 15969 11291 15980
rect 11326 15969 11360 16003
rect 11394 15980 11428 16003
rect 11462 15980 11496 16003
rect 11530 15980 11564 16003
rect 11598 15980 11632 16003
rect 11666 15980 11700 16003
rect 11734 15980 11768 16003
rect 11802 15980 11836 16003
rect 11870 15980 11904 16003
rect 11397 15969 11428 15980
rect 11469 15969 11496 15980
rect 11541 15969 11564 15980
rect 11613 15969 11632 15980
rect 11685 15969 11700 15980
rect 11757 15969 11768 15980
rect 11829 15969 11836 15980
rect 11901 15969 11904 15980
rect 11938 15980 11972 16003
rect 12006 15980 12040 16003
rect 12074 15980 12108 16003
rect 12142 15980 12176 16003
rect 12210 15980 12244 16003
rect 12278 15980 12312 16003
rect 12346 15980 12380 16003
rect 12414 15980 12448 16003
rect 12482 15980 12516 16003
rect 11938 15969 11939 15980
rect 12006 15969 12011 15980
rect 12074 15969 12083 15980
rect 12142 15969 12155 15980
rect 12210 15969 12227 15980
rect 12278 15969 12299 15980
rect 12346 15969 12371 15980
rect 12414 15969 12443 15980
rect 12482 15969 12515 15980
rect 12550 15969 12584 16003
rect 12618 15980 12652 16003
rect 12686 15980 12720 16003
rect 12754 15980 12788 16003
rect 12822 15980 12856 16003
rect 12890 15980 12924 16003
rect 12958 15980 12992 16003
rect 13026 15980 13060 16003
rect 13094 15980 13128 16003
rect 12621 15969 12652 15980
rect 12693 15969 12720 15980
rect 12765 15969 12788 15980
rect 12837 15969 12856 15980
rect 12909 15969 12924 15980
rect 12981 15969 12992 15980
rect 13053 15969 13060 15980
rect 13125 15969 13128 15980
rect 13162 15980 13196 16003
rect 13230 15980 13264 16003
rect 13298 15980 13332 16003
rect 13366 15980 13400 16003
rect 13434 15980 13468 16003
rect 13502 15980 13536 16003
rect 13570 15980 13604 16003
rect 13638 15980 13672 16003
rect 13706 15980 13740 16003
rect 13162 15969 13163 15980
rect 13230 15969 13235 15980
rect 13298 15969 13307 15980
rect 13366 15969 13379 15980
rect 13434 15969 13451 15980
rect 13502 15969 13523 15980
rect 13570 15969 13595 15980
rect 13638 15969 13667 15980
rect 13706 15969 13739 15980
rect 13774 15969 13808 16003
rect 13842 15980 13876 16003
rect 13910 15980 13944 16003
rect 13978 15980 14012 16003
rect 14046 15980 14080 16003
rect 14114 15980 14148 16003
rect 14182 15980 14216 16003
rect 14250 15980 14284 16003
rect 14318 15980 14352 16003
rect 13845 15969 13876 15980
rect 13917 15969 13944 15980
rect 13989 15969 14012 15980
rect 14061 15969 14080 15980
rect 14133 15969 14148 15980
rect 14205 15969 14216 15980
rect 14277 15969 14284 15980
rect 14349 15969 14352 15980
rect 14386 15986 14420 16003
rect 14454 15986 14492 16020
rect 14526 15986 14564 16020
rect 14598 15986 14636 16020
rect 14670 15986 14708 16020
rect 14742 15986 14780 16020
rect 14814 15986 14852 16020
rect 14886 15986 14924 16020
rect 14958 15986 14996 16020
rect 15030 15986 15068 16020
rect 15102 15986 15106 16020
rect 14386 15980 15106 15986
rect 14386 15969 14387 15980
rect 5376 15946 5415 15969
rect 5449 15946 5488 15969
rect 5522 15946 5561 15969
rect 5595 15946 5634 15969
rect 5668 15946 5707 15969
rect 5741 15946 5780 15969
rect 5814 15946 5853 15969
rect 5887 15946 5926 15969
rect 5960 15946 5999 15969
rect 6033 15946 6072 15969
rect 6106 15946 6145 15969
rect 6179 15946 6218 15969
rect 6252 15946 6291 15969
rect 6325 15946 6364 15969
rect 6398 15946 6437 15969
rect 6471 15946 6510 15969
rect 6544 15946 6583 15969
rect 6617 15946 6656 15969
rect 6690 15946 6729 15969
rect 6763 15946 6802 15969
rect 6836 15946 6875 15969
rect 6909 15946 6948 15969
rect 6982 15946 7021 15969
rect 7055 15946 7094 15969
rect 7128 15946 7167 15969
rect 7201 15946 7240 15969
rect 7274 15946 7313 15969
rect 7347 15946 7386 15969
rect 7420 15946 7459 15969
rect 7493 15946 7532 15969
rect 7566 15946 7605 15969
rect 7639 15946 7678 15969
rect 7712 15946 7751 15969
rect 7785 15946 7824 15969
rect 7858 15946 7897 15969
rect 7931 15946 7970 15969
rect 8004 15946 8043 15969
rect 8077 15946 8116 15969
rect 8150 15946 8189 15969
rect 8223 15946 8262 15969
rect 8296 15946 8335 15969
rect 8369 15946 8408 15969
rect 8442 15946 8481 15969
rect 8515 15946 8554 15969
rect 8588 15946 8627 15969
rect 8661 15946 8699 15969
rect 8733 15946 8771 15969
rect 8805 15946 8843 15969
rect 8877 15946 8915 15969
rect 8949 15946 8987 15969
rect 9021 15946 9059 15969
rect 9093 15946 9131 15969
rect 9165 15946 9203 15969
rect 9237 15946 9275 15969
rect 9309 15946 9347 15969
rect 9381 15946 9419 15969
rect 9453 15946 9491 15969
rect 9525 15946 9563 15969
rect 9597 15946 9635 15969
rect 9669 15946 9707 15969
rect 9741 15946 9779 15969
rect 9813 15946 9851 15969
rect 9885 15946 9923 15969
rect 9957 15946 9995 15969
rect 10029 15946 10067 15969
rect 10101 15946 10139 15969
rect 10173 15946 10211 15969
rect 10245 15946 10283 15969
rect 10317 15946 10355 15969
rect 10389 15946 10427 15969
rect 10461 15946 10499 15969
rect 10533 15946 10571 15969
rect 10605 15946 10643 15969
rect 10677 15946 10715 15969
rect 10749 15946 10787 15969
rect 10821 15946 10859 15969
rect 10893 15946 10931 15969
rect 10965 15946 11003 15969
rect 11037 15946 11075 15969
rect 11109 15946 11147 15969
rect 11181 15946 11219 15969
rect 11253 15946 11291 15969
rect 11325 15946 11363 15969
rect 11397 15946 11435 15969
rect 11469 15946 11507 15969
rect 11541 15946 11579 15969
rect 11613 15946 11651 15969
rect 11685 15946 11723 15969
rect 11757 15946 11795 15969
rect 11829 15946 11867 15969
rect 11901 15946 11939 15969
rect 11973 15946 12011 15969
rect 12045 15946 12083 15969
rect 12117 15946 12155 15969
rect 12189 15946 12227 15969
rect 12261 15946 12299 15969
rect 12333 15946 12371 15969
rect 12405 15946 12443 15969
rect 12477 15946 12515 15969
rect 12549 15946 12587 15969
rect 12621 15946 12659 15969
rect 12693 15946 12731 15969
rect 12765 15946 12803 15969
rect 12837 15946 12875 15969
rect 12909 15946 12947 15969
rect 12981 15946 13019 15969
rect 13053 15946 13091 15969
rect 13125 15946 13163 15969
rect 13197 15946 13235 15969
rect 13269 15946 13307 15969
rect 13341 15946 13379 15969
rect 13413 15946 13451 15969
rect 13485 15946 13523 15969
rect 13557 15946 13595 15969
rect 13629 15946 13667 15969
rect 13701 15946 13739 15969
rect 13773 15946 13811 15969
rect 13845 15946 13883 15969
rect 13917 15946 13955 15969
rect 13989 15946 14027 15969
rect 14061 15946 14099 15969
rect 14133 15946 14171 15969
rect 14205 15946 14243 15969
rect 14277 15946 14315 15969
rect 14349 15946 14387 15969
rect 14421 15951 14459 15980
rect 14493 15951 14531 15980
rect 14565 15951 14603 15980
rect 14637 15951 14675 15980
rect 14709 15951 14747 15980
rect 14781 15951 14819 15980
rect 14853 15951 14891 15980
rect 14925 15951 15106 15980
rect 14454 15946 14459 15951
rect 14526 15946 14531 15951
rect 14598 15946 14603 15951
rect 14670 15946 14675 15951
rect 14742 15946 14747 15951
rect 14814 15946 14819 15951
rect 14886 15946 14891 15951
rect 386 15933 14420 15946
rect 386 15915 444 15933
rect 67 15899 444 15915
rect 478 15899 513 15933
rect 547 15899 582 15933
rect 616 15899 651 15933
rect 685 15899 720 15933
rect 754 15899 789 15933
rect 823 15899 858 15933
rect 892 15899 927 15933
rect 961 15899 996 15933
rect 1030 15899 1065 15933
rect 1099 15899 1134 15933
rect 1168 15899 1203 15933
rect 1237 15899 1272 15933
rect 1306 15899 1341 15933
rect 1375 15899 1410 15933
rect 1444 15899 1479 15933
rect 1513 15899 1548 15933
rect 1582 15899 1617 15933
rect 1651 15899 1686 15933
rect 1720 15899 1755 15933
rect 1789 15899 1824 15933
rect 1858 15899 1893 15933
rect 1927 15899 1962 15933
rect 1996 15899 2031 15933
rect 2065 15899 2100 15933
rect 2134 15899 2169 15933
rect 2203 15899 2238 15933
rect 2272 15899 2307 15933
rect 2341 15899 2376 15933
rect 2410 15899 2445 15933
rect 2479 15899 2514 15933
rect 2548 15899 2583 15933
rect 2617 15899 2652 15933
rect 2686 15899 2721 15933
rect 2755 15899 2790 15933
rect 2824 15899 2859 15933
rect 2893 15899 2928 15933
rect 2962 15899 2996 15933
rect 3030 15899 3064 15933
rect 3098 15899 3132 15933
rect 3166 15899 3200 15933
rect 3234 15899 3268 15933
rect 3302 15899 3336 15933
rect 3370 15899 3404 15933
rect 3438 15899 3472 15933
rect 3506 15899 3540 15933
rect 3574 15899 3608 15933
rect 3642 15899 3676 15933
rect 3710 15899 3744 15933
rect 3778 15899 3812 15933
rect 3846 15899 3880 15933
rect 3914 15906 3948 15933
rect 3982 15906 4016 15933
rect 4050 15906 4084 15933
rect 4118 15906 4152 15933
rect 4186 15906 4220 15933
rect 4254 15906 4288 15933
rect 4322 15906 4356 15933
rect 3916 15899 3948 15906
rect 3989 15899 4016 15906
rect 4062 15899 4084 15906
rect 4135 15899 4152 15906
rect 4208 15899 4220 15906
rect 4281 15899 4288 15906
rect 4354 15899 4356 15906
rect 4390 15906 4424 15933
rect 4458 15906 4492 15933
rect 4526 15906 4560 15933
rect 4594 15906 4628 15933
rect 4662 15906 4696 15933
rect 4730 15906 4764 15933
rect 4798 15906 4832 15933
rect 4390 15899 4393 15906
rect 4458 15899 4466 15906
rect 4526 15899 4539 15906
rect 4594 15899 4612 15906
rect 4662 15899 4685 15906
rect 4730 15899 4758 15906
rect 4798 15899 4831 15906
rect 4866 15899 4900 15933
rect 4934 15906 4968 15933
rect 5002 15906 5036 15933
rect 5070 15906 5104 15933
rect 5138 15906 5172 15933
rect 5206 15906 5240 15933
rect 5274 15906 5308 15933
rect 4938 15899 4968 15906
rect 5011 15899 5036 15906
rect 5084 15899 5104 15906
rect 5157 15899 5172 15906
rect 5230 15899 5240 15906
rect 5303 15899 5308 15906
rect 5342 15906 5376 15933
rect 67 15880 3882 15899
rect 67 15846 68 15880
rect 102 15846 139 15880
rect 173 15846 210 15880
rect 244 15846 281 15880
rect 315 15846 352 15880
rect 386 15872 3882 15880
rect 3916 15872 3955 15899
rect 3989 15872 4028 15899
rect 4062 15872 4101 15899
rect 4135 15872 4174 15899
rect 4208 15872 4247 15899
rect 4281 15872 4320 15899
rect 4354 15872 4393 15899
rect 4427 15872 4466 15899
rect 4500 15872 4539 15899
rect 4573 15872 4612 15899
rect 4646 15872 4685 15899
rect 4719 15872 4758 15899
rect 4792 15872 4831 15899
rect 4865 15872 4904 15899
rect 4938 15872 4977 15899
rect 5011 15872 5050 15899
rect 5084 15872 5123 15899
rect 5157 15872 5196 15899
rect 5230 15872 5269 15899
rect 5303 15872 5342 15899
rect 5410 15906 5444 15933
rect 5478 15906 5512 15933
rect 5546 15906 5580 15933
rect 5614 15906 5648 15933
rect 5682 15906 5716 15933
rect 5750 15906 5784 15933
rect 5410 15899 5415 15906
rect 5478 15899 5488 15906
rect 5546 15899 5561 15906
rect 5614 15899 5634 15906
rect 5682 15899 5707 15906
rect 5750 15899 5780 15906
rect 5818 15899 5852 15933
rect 5886 15906 5920 15933
rect 5954 15906 5988 15933
rect 6022 15906 6056 15933
rect 6090 15906 6124 15933
rect 6158 15906 6192 15933
rect 6226 15906 6260 15933
rect 6294 15906 6328 15933
rect 5887 15899 5920 15906
rect 5960 15899 5988 15906
rect 6033 15899 6056 15906
rect 6106 15899 6124 15906
rect 6179 15899 6192 15906
rect 6252 15899 6260 15906
rect 6325 15899 6328 15906
rect 6362 15906 6396 15933
rect 6430 15906 6464 15933
rect 6498 15906 6532 15933
rect 6566 15906 6600 15933
rect 6634 15906 6668 15933
rect 6702 15906 6736 15933
rect 6770 15906 6804 15933
rect 6362 15899 6364 15906
rect 6430 15899 6437 15906
rect 6498 15899 6510 15906
rect 6566 15899 6583 15906
rect 6634 15899 6656 15906
rect 6702 15899 6729 15906
rect 6770 15899 6802 15906
rect 6838 15899 6872 15933
rect 6906 15906 6940 15933
rect 6974 15906 7008 15933
rect 7042 15906 7076 15933
rect 7110 15906 7144 15933
rect 7178 15906 7212 15933
rect 7246 15906 7280 15933
rect 7314 15906 7348 15933
rect 6909 15899 6940 15906
rect 6982 15899 7008 15906
rect 7055 15899 7076 15906
rect 7128 15899 7144 15906
rect 7201 15899 7212 15906
rect 7274 15899 7280 15906
rect 7347 15899 7348 15906
rect 7382 15906 7416 15933
rect 7450 15906 7484 15933
rect 7518 15906 7552 15933
rect 7586 15906 7620 15933
rect 7654 15906 7688 15933
rect 7722 15906 7756 15933
rect 7382 15899 7386 15906
rect 7450 15899 7459 15906
rect 7518 15899 7532 15906
rect 7586 15899 7605 15906
rect 7654 15899 7678 15906
rect 7722 15899 7751 15906
rect 7790 15899 7824 15933
rect 7858 15899 7892 15933
rect 7926 15906 7960 15933
rect 7994 15906 8028 15933
rect 8062 15906 8096 15933
rect 8130 15906 8164 15933
rect 8198 15906 8232 15933
rect 8266 15906 8300 15933
rect 7931 15899 7960 15906
rect 8004 15899 8028 15906
rect 8077 15899 8096 15906
rect 8150 15899 8164 15906
rect 8223 15899 8232 15906
rect 8296 15899 8300 15906
rect 8334 15906 8368 15933
rect 8402 15906 8436 15933
rect 8470 15906 8504 15933
rect 8538 15906 8572 15933
rect 8606 15906 8640 15933
rect 8674 15906 8708 15933
rect 8742 15906 8776 15933
rect 8810 15906 8844 15933
rect 8334 15899 8335 15906
rect 8402 15899 8408 15906
rect 8470 15899 8481 15906
rect 8538 15899 8554 15906
rect 8606 15899 8627 15906
rect 8674 15899 8699 15906
rect 8742 15899 8771 15906
rect 8810 15899 8843 15906
rect 8878 15899 8912 15933
rect 8946 15906 8980 15933
rect 9014 15906 9048 15933
rect 9082 15906 9116 15933
rect 9150 15906 9184 15933
rect 9218 15906 9252 15933
rect 9286 15906 9320 15933
rect 9354 15906 9388 15933
rect 9422 15906 9456 15933
rect 8949 15899 8980 15906
rect 9021 15899 9048 15906
rect 9093 15899 9116 15906
rect 9165 15899 9184 15906
rect 9237 15899 9252 15906
rect 9309 15899 9320 15906
rect 9381 15899 9388 15906
rect 9453 15899 9456 15906
rect 9490 15906 9524 15933
rect 9558 15906 9592 15933
rect 9626 15906 9660 15933
rect 9694 15906 9728 15933
rect 9762 15906 9796 15933
rect 9830 15906 9864 15933
rect 9898 15906 9932 15933
rect 9966 15906 10000 15933
rect 10034 15906 10068 15933
rect 9490 15899 9491 15906
rect 9558 15899 9563 15906
rect 9626 15899 9635 15906
rect 9694 15899 9707 15906
rect 9762 15899 9779 15906
rect 9830 15899 9851 15906
rect 9898 15899 9923 15906
rect 9966 15899 9995 15906
rect 10034 15899 10067 15906
rect 10102 15899 10136 15933
rect 10170 15906 10204 15933
rect 10238 15906 10272 15933
rect 10306 15906 10340 15933
rect 10374 15906 10408 15933
rect 10442 15906 10476 15933
rect 10510 15906 10544 15933
rect 10578 15906 10612 15933
rect 10646 15906 10680 15933
rect 10173 15899 10204 15906
rect 10245 15899 10272 15906
rect 10317 15899 10340 15906
rect 10389 15899 10408 15906
rect 10461 15899 10476 15906
rect 10533 15899 10544 15906
rect 10605 15899 10612 15906
rect 10677 15899 10680 15906
rect 10714 15906 10748 15933
rect 10782 15906 10816 15933
rect 10850 15906 10884 15933
rect 10918 15906 10952 15933
rect 10986 15906 11020 15933
rect 11054 15906 11088 15933
rect 11122 15906 11156 15933
rect 11190 15906 11224 15933
rect 11258 15906 11292 15933
rect 10714 15899 10715 15906
rect 10782 15899 10787 15906
rect 10850 15899 10859 15906
rect 10918 15899 10931 15906
rect 10986 15899 11003 15906
rect 11054 15899 11075 15906
rect 11122 15899 11147 15906
rect 11190 15899 11219 15906
rect 11258 15899 11291 15906
rect 11326 15899 11360 15933
rect 11394 15906 11428 15933
rect 11462 15906 11496 15933
rect 11530 15906 11564 15933
rect 11598 15906 11632 15933
rect 11666 15906 11700 15933
rect 11734 15906 11768 15933
rect 11802 15906 11836 15933
rect 11870 15906 11904 15933
rect 11397 15899 11428 15906
rect 11469 15899 11496 15906
rect 11541 15899 11564 15906
rect 11613 15899 11632 15906
rect 11685 15899 11700 15906
rect 11757 15899 11768 15906
rect 11829 15899 11836 15906
rect 11901 15899 11904 15906
rect 11938 15906 11972 15933
rect 12006 15906 12040 15933
rect 12074 15906 12108 15933
rect 12142 15906 12176 15933
rect 12210 15906 12244 15933
rect 12278 15906 12312 15933
rect 12346 15906 12380 15933
rect 12414 15906 12448 15933
rect 12482 15906 12516 15933
rect 11938 15899 11939 15906
rect 12006 15899 12011 15906
rect 12074 15899 12083 15906
rect 12142 15899 12155 15906
rect 12210 15899 12227 15906
rect 12278 15899 12299 15906
rect 12346 15899 12371 15906
rect 12414 15899 12443 15906
rect 12482 15899 12515 15906
rect 12550 15899 12584 15933
rect 12618 15906 12652 15933
rect 12686 15906 12720 15933
rect 12754 15906 12788 15933
rect 12822 15906 12856 15933
rect 12890 15906 12924 15933
rect 12958 15906 12992 15933
rect 13026 15906 13060 15933
rect 13094 15906 13128 15933
rect 12621 15899 12652 15906
rect 12693 15899 12720 15906
rect 12765 15899 12788 15906
rect 12837 15899 12856 15906
rect 12909 15899 12924 15906
rect 12981 15899 12992 15906
rect 13053 15899 13060 15906
rect 13125 15899 13128 15906
rect 13162 15906 13196 15933
rect 13230 15906 13264 15933
rect 13298 15906 13332 15933
rect 13366 15906 13400 15933
rect 13434 15906 13468 15933
rect 13502 15906 13536 15933
rect 13570 15906 13604 15933
rect 13638 15906 13672 15933
rect 13706 15906 13740 15933
rect 13162 15899 13163 15906
rect 13230 15899 13235 15906
rect 13298 15899 13307 15906
rect 13366 15899 13379 15906
rect 13434 15899 13451 15906
rect 13502 15899 13523 15906
rect 13570 15899 13595 15906
rect 13638 15899 13667 15906
rect 13706 15899 13739 15906
rect 13774 15899 13808 15933
rect 13842 15906 13876 15933
rect 13910 15906 13944 15933
rect 13978 15906 14012 15933
rect 14046 15906 14080 15933
rect 14114 15906 14148 15933
rect 14182 15906 14216 15933
rect 14250 15906 14284 15933
rect 14318 15906 14352 15933
rect 13845 15899 13876 15906
rect 13917 15899 13944 15906
rect 13989 15899 14012 15906
rect 14061 15899 14080 15906
rect 14133 15899 14148 15906
rect 14205 15899 14216 15906
rect 14277 15899 14284 15906
rect 14349 15899 14352 15906
rect 14386 15917 14420 15933
rect 14454 15917 14492 15946
rect 14526 15917 14564 15946
rect 14598 15917 14636 15946
rect 14670 15917 14708 15946
rect 14742 15917 14780 15946
rect 14814 15917 14852 15946
rect 14886 15917 14924 15946
rect 14958 15917 14996 15951
rect 15030 15917 15068 15951
rect 15102 15917 15106 15951
rect 14386 15906 15106 15917
rect 14386 15899 14387 15906
rect 5376 15872 5415 15899
rect 5449 15872 5488 15899
rect 5522 15872 5561 15899
rect 5595 15872 5634 15899
rect 5668 15872 5707 15899
rect 5741 15872 5780 15899
rect 5814 15872 5853 15899
rect 5887 15872 5926 15899
rect 5960 15872 5999 15899
rect 6033 15872 6072 15899
rect 6106 15872 6145 15899
rect 6179 15872 6218 15899
rect 6252 15872 6291 15899
rect 6325 15872 6364 15899
rect 6398 15872 6437 15899
rect 6471 15872 6510 15899
rect 6544 15872 6583 15899
rect 6617 15872 6656 15899
rect 6690 15872 6729 15899
rect 6763 15872 6802 15899
rect 6836 15872 6875 15899
rect 6909 15872 6948 15899
rect 6982 15872 7021 15899
rect 7055 15872 7094 15899
rect 7128 15872 7167 15899
rect 7201 15872 7240 15899
rect 7274 15872 7313 15899
rect 7347 15872 7386 15899
rect 7420 15872 7459 15899
rect 7493 15872 7532 15899
rect 7566 15872 7605 15899
rect 7639 15872 7678 15899
rect 7712 15872 7751 15899
rect 7785 15872 7824 15899
rect 7858 15872 7897 15899
rect 7931 15872 7970 15899
rect 8004 15872 8043 15899
rect 8077 15872 8116 15899
rect 8150 15872 8189 15899
rect 8223 15872 8262 15899
rect 8296 15872 8335 15899
rect 8369 15872 8408 15899
rect 8442 15872 8481 15899
rect 8515 15872 8554 15899
rect 8588 15872 8627 15899
rect 8661 15872 8699 15899
rect 8733 15872 8771 15899
rect 8805 15872 8843 15899
rect 8877 15872 8915 15899
rect 8949 15872 8987 15899
rect 9021 15872 9059 15899
rect 9093 15872 9131 15899
rect 9165 15872 9203 15899
rect 9237 15872 9275 15899
rect 9309 15872 9347 15899
rect 9381 15872 9419 15899
rect 9453 15872 9491 15899
rect 9525 15872 9563 15899
rect 9597 15872 9635 15899
rect 9669 15872 9707 15899
rect 9741 15872 9779 15899
rect 9813 15872 9851 15899
rect 9885 15872 9923 15899
rect 9957 15872 9995 15899
rect 10029 15872 10067 15899
rect 10101 15872 10139 15899
rect 10173 15872 10211 15899
rect 10245 15872 10283 15899
rect 10317 15872 10355 15899
rect 10389 15872 10427 15899
rect 10461 15872 10499 15899
rect 10533 15872 10571 15899
rect 10605 15872 10643 15899
rect 10677 15872 10715 15899
rect 10749 15872 10787 15899
rect 10821 15872 10859 15899
rect 10893 15872 10931 15899
rect 10965 15872 11003 15899
rect 11037 15872 11075 15899
rect 11109 15872 11147 15899
rect 11181 15872 11219 15899
rect 11253 15872 11291 15899
rect 11325 15872 11363 15899
rect 11397 15872 11435 15899
rect 11469 15872 11507 15899
rect 11541 15872 11579 15899
rect 11613 15872 11651 15899
rect 11685 15872 11723 15899
rect 11757 15872 11795 15899
rect 11829 15872 11867 15899
rect 11901 15872 11939 15899
rect 11973 15872 12011 15899
rect 12045 15872 12083 15899
rect 12117 15872 12155 15899
rect 12189 15872 12227 15899
rect 12261 15872 12299 15899
rect 12333 15872 12371 15899
rect 12405 15872 12443 15899
rect 12477 15872 12515 15899
rect 12549 15872 12587 15899
rect 12621 15872 12659 15899
rect 12693 15872 12731 15899
rect 12765 15872 12803 15899
rect 12837 15872 12875 15899
rect 12909 15872 12947 15899
rect 12981 15872 13019 15899
rect 13053 15872 13091 15899
rect 13125 15872 13163 15899
rect 13197 15872 13235 15899
rect 13269 15872 13307 15899
rect 13341 15872 13379 15899
rect 13413 15872 13451 15899
rect 13485 15872 13523 15899
rect 13557 15872 13595 15899
rect 13629 15872 13667 15899
rect 13701 15872 13739 15899
rect 13773 15872 13811 15899
rect 13845 15872 13883 15899
rect 13917 15872 13955 15899
rect 13989 15872 14027 15899
rect 14061 15872 14099 15899
rect 14133 15872 14171 15899
rect 14205 15872 14243 15899
rect 14277 15872 14315 15899
rect 14349 15872 14387 15899
rect 14421 15882 14459 15906
rect 14493 15882 14531 15906
rect 14565 15882 14603 15906
rect 14637 15882 14675 15906
rect 14709 15882 14747 15906
rect 14781 15882 14819 15906
rect 14853 15882 14891 15906
rect 14925 15882 15106 15906
rect 14454 15872 14459 15882
rect 14526 15872 14531 15882
rect 14598 15872 14603 15882
rect 14670 15872 14675 15882
rect 14742 15872 14747 15882
rect 14814 15872 14819 15882
rect 14886 15872 14891 15882
rect 386 15863 14420 15872
rect 386 15846 444 15863
rect 67 15829 444 15846
rect 478 15829 513 15863
rect 547 15829 582 15863
rect 616 15829 651 15863
rect 685 15829 720 15863
rect 754 15829 789 15863
rect 823 15829 858 15863
rect 892 15829 927 15863
rect 961 15829 996 15863
rect 1030 15829 1065 15863
rect 1099 15829 1134 15863
rect 1168 15829 1203 15863
rect 1237 15829 1272 15863
rect 1306 15829 1341 15863
rect 1375 15829 1410 15863
rect 1444 15829 1479 15863
rect 1513 15829 1548 15863
rect 1582 15829 1617 15863
rect 1651 15829 1686 15863
rect 1720 15829 1755 15863
rect 1789 15829 1824 15863
rect 1858 15829 1893 15863
rect 1927 15829 1962 15863
rect 1996 15829 2031 15863
rect 2065 15829 2100 15863
rect 2134 15829 2169 15863
rect 2203 15829 2238 15863
rect 2272 15829 2307 15863
rect 2341 15829 2376 15863
rect 2410 15829 2445 15863
rect 2479 15829 2514 15863
rect 2548 15829 2583 15863
rect 2617 15829 2652 15863
rect 2686 15829 2721 15863
rect 2755 15829 2790 15863
rect 2824 15829 2859 15863
rect 2893 15829 2928 15863
rect 2962 15829 2996 15863
rect 3030 15829 3064 15863
rect 3098 15829 3132 15863
rect 3166 15829 3200 15863
rect 3234 15829 3268 15863
rect 3302 15829 3336 15863
rect 3370 15829 3404 15863
rect 3438 15829 3472 15863
rect 3506 15829 3540 15863
rect 3574 15829 3608 15863
rect 3642 15829 3676 15863
rect 3710 15829 3744 15863
rect 3778 15829 3812 15863
rect 3846 15829 3880 15863
rect 3914 15832 3948 15863
rect 3982 15832 4016 15863
rect 4050 15832 4084 15863
rect 4118 15832 4152 15863
rect 4186 15832 4220 15863
rect 4254 15832 4288 15863
rect 4322 15832 4356 15863
rect 3916 15829 3948 15832
rect 3989 15829 4016 15832
rect 4062 15829 4084 15832
rect 4135 15829 4152 15832
rect 4208 15829 4220 15832
rect 4281 15829 4288 15832
rect 4354 15829 4356 15832
rect 4390 15832 4424 15863
rect 4458 15832 4492 15863
rect 4526 15832 4560 15863
rect 4594 15832 4628 15863
rect 4662 15832 4696 15863
rect 4730 15832 4764 15863
rect 4798 15832 4832 15863
rect 4390 15829 4393 15832
rect 4458 15829 4466 15832
rect 4526 15829 4539 15832
rect 4594 15829 4612 15832
rect 4662 15829 4685 15832
rect 4730 15829 4758 15832
rect 4798 15829 4831 15832
rect 4866 15829 4900 15863
rect 4934 15832 4968 15863
rect 5002 15832 5036 15863
rect 5070 15832 5104 15863
rect 5138 15832 5172 15863
rect 5206 15832 5240 15863
rect 5274 15832 5308 15863
rect 4938 15829 4968 15832
rect 5011 15829 5036 15832
rect 5084 15829 5104 15832
rect 5157 15829 5172 15832
rect 5230 15829 5240 15832
rect 5303 15829 5308 15832
rect 5342 15832 5376 15863
rect 67 15811 3882 15829
rect 67 15777 68 15811
rect 102 15789 139 15811
rect 133 15777 139 15789
rect 173 15777 210 15811
rect 244 15777 281 15811
rect 315 15777 352 15811
rect 386 15798 3882 15811
rect 3916 15798 3955 15829
rect 3989 15798 4028 15829
rect 4062 15798 4101 15829
rect 4135 15798 4174 15829
rect 4208 15798 4247 15829
rect 4281 15798 4320 15829
rect 4354 15798 4393 15829
rect 4427 15798 4466 15829
rect 4500 15798 4539 15829
rect 4573 15798 4612 15829
rect 4646 15798 4685 15829
rect 4719 15798 4758 15829
rect 4792 15798 4831 15829
rect 4865 15798 4904 15829
rect 4938 15798 4977 15829
rect 5011 15798 5050 15829
rect 5084 15798 5123 15829
rect 5157 15798 5196 15829
rect 5230 15798 5269 15829
rect 5303 15798 5342 15829
rect 5410 15832 5444 15863
rect 5478 15832 5512 15863
rect 5546 15832 5580 15863
rect 5614 15832 5648 15863
rect 5682 15832 5716 15863
rect 5750 15832 5784 15863
rect 5410 15829 5415 15832
rect 5478 15829 5488 15832
rect 5546 15829 5561 15832
rect 5614 15829 5634 15832
rect 5682 15829 5707 15832
rect 5750 15829 5780 15832
rect 5818 15829 5852 15863
rect 5886 15832 5920 15863
rect 5954 15832 5988 15863
rect 6022 15832 6056 15863
rect 6090 15832 6124 15863
rect 6158 15832 6192 15863
rect 6226 15832 6260 15863
rect 6294 15832 6328 15863
rect 5887 15829 5920 15832
rect 5960 15829 5988 15832
rect 6033 15829 6056 15832
rect 6106 15829 6124 15832
rect 6179 15829 6192 15832
rect 6252 15829 6260 15832
rect 6325 15829 6328 15832
rect 6362 15832 6396 15863
rect 6430 15832 6464 15863
rect 6498 15832 6532 15863
rect 6566 15832 6600 15863
rect 6634 15832 6668 15863
rect 6702 15832 6736 15863
rect 6770 15832 6804 15863
rect 6362 15829 6364 15832
rect 6430 15829 6437 15832
rect 6498 15829 6510 15832
rect 6566 15829 6583 15832
rect 6634 15829 6656 15832
rect 6702 15829 6729 15832
rect 6770 15829 6802 15832
rect 6838 15829 6872 15863
rect 6906 15832 6940 15863
rect 6974 15832 7008 15863
rect 7042 15832 7076 15863
rect 7110 15832 7144 15863
rect 7178 15832 7212 15863
rect 7246 15832 7280 15863
rect 7314 15832 7348 15863
rect 6909 15829 6940 15832
rect 6982 15829 7008 15832
rect 7055 15829 7076 15832
rect 7128 15829 7144 15832
rect 7201 15829 7212 15832
rect 7274 15829 7280 15832
rect 7347 15829 7348 15832
rect 7382 15832 7416 15863
rect 7450 15832 7484 15863
rect 7518 15832 7552 15863
rect 7586 15832 7620 15863
rect 7654 15832 7688 15863
rect 7722 15832 7756 15863
rect 7382 15829 7386 15832
rect 7450 15829 7459 15832
rect 7518 15829 7532 15832
rect 7586 15829 7605 15832
rect 7654 15829 7678 15832
rect 7722 15829 7751 15832
rect 7790 15829 7824 15863
rect 7858 15829 7892 15863
rect 7926 15832 7960 15863
rect 7994 15832 8028 15863
rect 8062 15832 8096 15863
rect 8130 15832 8164 15863
rect 8198 15832 8232 15863
rect 8266 15832 8300 15863
rect 7931 15829 7960 15832
rect 8004 15829 8028 15832
rect 8077 15829 8096 15832
rect 8150 15829 8164 15832
rect 8223 15829 8232 15832
rect 8296 15829 8300 15832
rect 8334 15832 8368 15863
rect 8402 15832 8436 15863
rect 8470 15832 8504 15863
rect 8538 15832 8572 15863
rect 8606 15832 8640 15863
rect 8674 15832 8708 15863
rect 8742 15832 8776 15863
rect 8810 15832 8844 15863
rect 8334 15829 8335 15832
rect 8402 15829 8408 15832
rect 8470 15829 8481 15832
rect 8538 15829 8554 15832
rect 8606 15829 8627 15832
rect 8674 15829 8699 15832
rect 8742 15829 8771 15832
rect 8810 15829 8843 15832
rect 8878 15829 8912 15863
rect 8946 15832 8980 15863
rect 9014 15832 9048 15863
rect 9082 15832 9116 15863
rect 9150 15832 9184 15863
rect 9218 15832 9252 15863
rect 9286 15832 9320 15863
rect 9354 15832 9388 15863
rect 9422 15832 9456 15863
rect 8949 15829 8980 15832
rect 9021 15829 9048 15832
rect 9093 15829 9116 15832
rect 9165 15829 9184 15832
rect 9237 15829 9252 15832
rect 9309 15829 9320 15832
rect 9381 15829 9388 15832
rect 9453 15829 9456 15832
rect 9490 15832 9524 15863
rect 9558 15832 9592 15863
rect 9626 15832 9660 15863
rect 9694 15832 9728 15863
rect 9762 15832 9796 15863
rect 9830 15832 9864 15863
rect 9898 15832 9932 15863
rect 9966 15832 10000 15863
rect 10034 15832 10068 15863
rect 9490 15829 9491 15832
rect 9558 15829 9563 15832
rect 9626 15829 9635 15832
rect 9694 15829 9707 15832
rect 9762 15829 9779 15832
rect 9830 15829 9851 15832
rect 9898 15829 9923 15832
rect 9966 15829 9995 15832
rect 10034 15829 10067 15832
rect 10102 15829 10136 15863
rect 10170 15832 10204 15863
rect 10238 15832 10272 15863
rect 10306 15832 10340 15863
rect 10374 15832 10408 15863
rect 10442 15832 10476 15863
rect 10510 15832 10544 15863
rect 10578 15832 10612 15863
rect 10646 15832 10680 15863
rect 10173 15829 10204 15832
rect 10245 15829 10272 15832
rect 10317 15829 10340 15832
rect 10389 15829 10408 15832
rect 10461 15829 10476 15832
rect 10533 15829 10544 15832
rect 10605 15829 10612 15832
rect 10677 15829 10680 15832
rect 10714 15832 10748 15863
rect 10782 15832 10816 15863
rect 10850 15832 10884 15863
rect 10918 15832 10952 15863
rect 10986 15832 11020 15863
rect 11054 15832 11088 15863
rect 11122 15832 11156 15863
rect 11190 15832 11224 15863
rect 11258 15832 11292 15863
rect 10714 15829 10715 15832
rect 10782 15829 10787 15832
rect 10850 15829 10859 15832
rect 10918 15829 10931 15832
rect 10986 15829 11003 15832
rect 11054 15829 11075 15832
rect 11122 15829 11147 15832
rect 11190 15829 11219 15832
rect 11258 15829 11291 15832
rect 11326 15829 11360 15863
rect 11394 15832 11428 15863
rect 11462 15832 11496 15863
rect 11530 15832 11564 15863
rect 11598 15832 11632 15863
rect 11666 15832 11700 15863
rect 11734 15832 11768 15863
rect 11802 15832 11836 15863
rect 11870 15832 11904 15863
rect 11397 15829 11428 15832
rect 11469 15829 11496 15832
rect 11541 15829 11564 15832
rect 11613 15829 11632 15832
rect 11685 15829 11700 15832
rect 11757 15829 11768 15832
rect 11829 15829 11836 15832
rect 11901 15829 11904 15832
rect 11938 15832 11972 15863
rect 12006 15832 12040 15863
rect 12074 15832 12108 15863
rect 12142 15832 12176 15863
rect 12210 15832 12244 15863
rect 12278 15832 12312 15863
rect 12346 15832 12380 15863
rect 12414 15832 12448 15863
rect 12482 15832 12516 15863
rect 11938 15829 11939 15832
rect 12006 15829 12011 15832
rect 12074 15829 12083 15832
rect 12142 15829 12155 15832
rect 12210 15829 12227 15832
rect 12278 15829 12299 15832
rect 12346 15829 12371 15832
rect 12414 15829 12443 15832
rect 12482 15829 12515 15832
rect 12550 15829 12584 15863
rect 12618 15832 12652 15863
rect 12686 15832 12720 15863
rect 12754 15832 12788 15863
rect 12822 15832 12856 15863
rect 12890 15832 12924 15863
rect 12958 15832 12992 15863
rect 13026 15832 13060 15863
rect 13094 15832 13128 15863
rect 12621 15829 12652 15832
rect 12693 15829 12720 15832
rect 12765 15829 12788 15832
rect 12837 15829 12856 15832
rect 12909 15829 12924 15832
rect 12981 15829 12992 15832
rect 13053 15829 13060 15832
rect 13125 15829 13128 15832
rect 13162 15832 13196 15863
rect 13230 15832 13264 15863
rect 13298 15832 13332 15863
rect 13366 15832 13400 15863
rect 13434 15832 13468 15863
rect 13502 15832 13536 15863
rect 13570 15832 13604 15863
rect 13638 15832 13672 15863
rect 13706 15832 13740 15863
rect 13162 15829 13163 15832
rect 13230 15829 13235 15832
rect 13298 15829 13307 15832
rect 13366 15829 13379 15832
rect 13434 15829 13451 15832
rect 13502 15829 13523 15832
rect 13570 15829 13595 15832
rect 13638 15829 13667 15832
rect 13706 15829 13739 15832
rect 13774 15829 13808 15863
rect 13842 15832 13876 15863
rect 13910 15832 13944 15863
rect 13978 15832 14012 15863
rect 14046 15832 14080 15863
rect 14114 15832 14148 15863
rect 14182 15832 14216 15863
rect 14250 15832 14284 15863
rect 14318 15832 14352 15863
rect 13845 15829 13876 15832
rect 13917 15829 13944 15832
rect 13989 15829 14012 15832
rect 14061 15829 14080 15832
rect 14133 15829 14148 15832
rect 14205 15829 14216 15832
rect 14277 15829 14284 15832
rect 14349 15829 14352 15832
rect 14386 15848 14420 15863
rect 14454 15848 14492 15872
rect 14526 15848 14564 15872
rect 14598 15848 14636 15872
rect 14670 15848 14708 15872
rect 14742 15848 14780 15872
rect 14814 15848 14852 15872
rect 14886 15848 14924 15872
rect 14958 15848 14996 15882
rect 15030 15848 15068 15882
rect 15102 15848 15106 15882
rect 14386 15832 15106 15848
rect 14386 15829 14387 15832
rect 5376 15798 5415 15829
rect 5449 15798 5488 15829
rect 5522 15798 5561 15829
rect 5595 15798 5634 15829
rect 5668 15798 5707 15829
rect 5741 15798 5780 15829
rect 5814 15798 5853 15829
rect 5887 15798 5926 15829
rect 5960 15798 5999 15829
rect 6033 15798 6072 15829
rect 6106 15798 6145 15829
rect 6179 15798 6218 15829
rect 6252 15798 6291 15829
rect 6325 15798 6364 15829
rect 6398 15798 6437 15829
rect 6471 15798 6510 15829
rect 6544 15798 6583 15829
rect 6617 15798 6656 15829
rect 6690 15798 6729 15829
rect 6763 15798 6802 15829
rect 6836 15798 6875 15829
rect 6909 15798 6948 15829
rect 6982 15798 7021 15829
rect 7055 15798 7094 15829
rect 7128 15798 7167 15829
rect 7201 15798 7240 15829
rect 7274 15798 7313 15829
rect 7347 15798 7386 15829
rect 7420 15798 7459 15829
rect 7493 15798 7532 15829
rect 7566 15798 7605 15829
rect 7639 15798 7678 15829
rect 7712 15798 7751 15829
rect 7785 15798 7824 15829
rect 7858 15798 7897 15829
rect 7931 15798 7970 15829
rect 8004 15798 8043 15829
rect 8077 15798 8116 15829
rect 8150 15798 8189 15829
rect 8223 15798 8262 15829
rect 8296 15798 8335 15829
rect 8369 15798 8408 15829
rect 8442 15798 8481 15829
rect 8515 15798 8554 15829
rect 8588 15798 8627 15829
rect 8661 15798 8699 15829
rect 8733 15798 8771 15829
rect 8805 15798 8843 15829
rect 8877 15798 8915 15829
rect 8949 15798 8987 15829
rect 9021 15798 9059 15829
rect 9093 15798 9131 15829
rect 9165 15798 9203 15829
rect 9237 15798 9275 15829
rect 9309 15798 9347 15829
rect 9381 15798 9419 15829
rect 9453 15798 9491 15829
rect 9525 15798 9563 15829
rect 9597 15798 9635 15829
rect 9669 15798 9707 15829
rect 9741 15798 9779 15829
rect 9813 15798 9851 15829
rect 9885 15798 9923 15829
rect 9957 15798 9995 15829
rect 10029 15798 10067 15829
rect 10101 15798 10139 15829
rect 10173 15798 10211 15829
rect 10245 15798 10283 15829
rect 10317 15798 10355 15829
rect 10389 15798 10427 15829
rect 10461 15798 10499 15829
rect 10533 15798 10571 15829
rect 10605 15798 10643 15829
rect 10677 15798 10715 15829
rect 10749 15798 10787 15829
rect 10821 15798 10859 15829
rect 10893 15798 10931 15829
rect 10965 15798 11003 15829
rect 11037 15798 11075 15829
rect 11109 15798 11147 15829
rect 11181 15798 11219 15829
rect 11253 15798 11291 15829
rect 11325 15798 11363 15829
rect 11397 15798 11435 15829
rect 11469 15798 11507 15829
rect 11541 15798 11579 15829
rect 11613 15798 11651 15829
rect 11685 15798 11723 15829
rect 11757 15798 11795 15829
rect 11829 15798 11867 15829
rect 11901 15798 11939 15829
rect 11973 15798 12011 15829
rect 12045 15798 12083 15829
rect 12117 15798 12155 15829
rect 12189 15798 12227 15829
rect 12261 15798 12299 15829
rect 12333 15798 12371 15829
rect 12405 15798 12443 15829
rect 12477 15798 12515 15829
rect 12549 15798 12587 15829
rect 12621 15798 12659 15829
rect 12693 15798 12731 15829
rect 12765 15798 12803 15829
rect 12837 15798 12875 15829
rect 12909 15798 12947 15829
rect 12981 15798 13019 15829
rect 13053 15798 13091 15829
rect 13125 15798 13163 15829
rect 13197 15798 13235 15829
rect 13269 15798 13307 15829
rect 13341 15798 13379 15829
rect 13413 15798 13451 15829
rect 13485 15798 13523 15829
rect 13557 15798 13595 15829
rect 13629 15798 13667 15829
rect 13701 15798 13739 15829
rect 13773 15798 13811 15829
rect 13845 15798 13883 15829
rect 13917 15798 13955 15829
rect 13989 15798 14027 15829
rect 14061 15798 14099 15829
rect 14133 15798 14171 15829
rect 14205 15798 14243 15829
rect 14277 15798 14315 15829
rect 14349 15798 14387 15829
rect 14421 15813 14459 15832
rect 14493 15813 14531 15832
rect 14565 15813 14603 15832
rect 14637 15813 14675 15832
rect 14709 15813 14747 15832
rect 14781 15813 14819 15832
rect 14853 15813 14891 15832
rect 14925 15813 15106 15832
rect 14454 15798 14459 15813
rect 14526 15798 14531 15813
rect 14598 15798 14603 15813
rect 14670 15798 14675 15813
rect 14742 15798 14747 15813
rect 14814 15798 14819 15813
rect 14886 15798 14891 15813
rect 386 15793 14420 15798
rect 386 15777 444 15793
rect 67 15755 99 15777
rect 133 15759 444 15777
rect 478 15759 513 15793
rect 547 15759 582 15793
rect 616 15759 651 15793
rect 685 15759 720 15793
rect 754 15759 789 15793
rect 823 15759 858 15793
rect 892 15759 927 15793
rect 961 15759 996 15793
rect 1030 15759 1065 15793
rect 1099 15759 1134 15793
rect 1168 15759 1203 15793
rect 1237 15759 1272 15793
rect 1306 15759 1341 15793
rect 1375 15759 1410 15793
rect 1444 15759 1479 15793
rect 1513 15759 1548 15793
rect 1582 15759 1617 15793
rect 1651 15759 1686 15793
rect 1720 15759 1755 15793
rect 1789 15759 1824 15793
rect 1858 15759 1893 15793
rect 1927 15759 1962 15793
rect 1996 15759 2031 15793
rect 2065 15759 2100 15793
rect 2134 15759 2169 15793
rect 2203 15759 2238 15793
rect 2272 15759 2307 15793
rect 2341 15759 2376 15793
rect 2410 15759 2445 15793
rect 2479 15759 2514 15793
rect 2548 15759 2583 15793
rect 2617 15759 2652 15793
rect 2686 15759 2721 15793
rect 2755 15759 2790 15793
rect 2824 15759 2859 15793
rect 2893 15759 2928 15793
rect 2962 15759 2996 15793
rect 3030 15759 3064 15793
rect 3098 15759 3132 15793
rect 3166 15759 3200 15793
rect 3234 15759 3268 15793
rect 3302 15759 3336 15793
rect 3370 15759 3404 15793
rect 3438 15759 3472 15793
rect 3506 15759 3540 15793
rect 3574 15759 3608 15793
rect 3642 15759 3676 15793
rect 3710 15759 3744 15793
rect 3778 15759 3812 15793
rect 3846 15759 3880 15793
rect 3914 15759 3948 15793
rect 3982 15759 4016 15793
rect 4050 15759 4084 15793
rect 4118 15759 4152 15793
rect 4186 15759 4220 15793
rect 4254 15759 4288 15793
rect 4322 15759 4356 15793
rect 4390 15759 4424 15793
rect 4458 15759 4492 15793
rect 4526 15759 4560 15793
rect 4594 15759 4628 15793
rect 4662 15759 4696 15793
rect 4730 15759 4764 15793
rect 4798 15759 4832 15793
rect 4866 15759 4900 15793
rect 4934 15759 4968 15793
rect 5002 15759 5036 15793
rect 5070 15759 5104 15793
rect 5138 15759 5172 15793
rect 5206 15759 5240 15793
rect 5274 15759 5308 15793
rect 5342 15759 5376 15793
rect 5410 15759 5444 15793
rect 5478 15759 5512 15793
rect 5546 15759 5580 15793
rect 5614 15759 5648 15793
rect 5682 15759 5716 15793
rect 5750 15759 5784 15793
rect 5818 15759 5852 15793
rect 5886 15759 5920 15793
rect 5954 15759 5988 15793
rect 6022 15759 6056 15793
rect 6090 15759 6124 15793
rect 6158 15759 6192 15793
rect 6226 15759 6260 15793
rect 6294 15759 6328 15793
rect 6362 15759 6396 15793
rect 6430 15759 6464 15793
rect 6498 15759 6532 15793
rect 6566 15759 6600 15793
rect 6634 15759 6668 15793
rect 6702 15759 6736 15793
rect 6770 15759 6804 15793
rect 6838 15759 6872 15793
rect 6906 15759 6940 15793
rect 6974 15759 7008 15793
rect 7042 15759 7076 15793
rect 7110 15759 7144 15793
rect 7178 15759 7212 15793
rect 7246 15759 7280 15793
rect 7314 15759 7348 15793
rect 7382 15759 7416 15793
rect 7450 15759 7484 15793
rect 7518 15759 7552 15793
rect 7586 15759 7620 15793
rect 7654 15759 7688 15793
rect 7722 15759 7756 15793
rect 7790 15759 7824 15793
rect 7858 15759 7892 15793
rect 7926 15759 7960 15793
rect 7994 15759 8028 15793
rect 8062 15759 8096 15793
rect 8130 15759 8164 15793
rect 8198 15759 8232 15793
rect 8266 15759 8300 15793
rect 8334 15759 8368 15793
rect 8402 15759 8436 15793
rect 8470 15759 8504 15793
rect 8538 15759 8572 15793
rect 8606 15759 8640 15793
rect 8674 15759 8708 15793
rect 8742 15759 8776 15793
rect 8810 15759 8844 15793
rect 8878 15759 8912 15793
rect 8946 15759 8980 15793
rect 9014 15759 9048 15793
rect 9082 15759 9116 15793
rect 9150 15759 9184 15793
rect 9218 15759 9252 15793
rect 9286 15759 9320 15793
rect 9354 15759 9388 15793
rect 9422 15759 9456 15793
rect 9490 15759 9524 15793
rect 9558 15759 9592 15793
rect 9626 15759 9660 15793
rect 9694 15759 9728 15793
rect 9762 15759 9796 15793
rect 9830 15759 9864 15793
rect 9898 15759 9932 15793
rect 9966 15759 10000 15793
rect 10034 15759 10068 15793
rect 10102 15759 10136 15793
rect 10170 15759 10204 15793
rect 10238 15759 10272 15793
rect 10306 15759 10340 15793
rect 10374 15759 10408 15793
rect 10442 15759 10476 15793
rect 10510 15759 10544 15793
rect 10578 15759 10612 15793
rect 10646 15759 10680 15793
rect 10714 15759 10748 15793
rect 10782 15759 10816 15793
rect 10850 15759 10884 15793
rect 10918 15759 10952 15793
rect 10986 15759 11020 15793
rect 11054 15759 11088 15793
rect 11122 15759 11156 15793
rect 11190 15759 11224 15793
rect 11258 15759 11292 15793
rect 11326 15759 11360 15793
rect 11394 15759 11428 15793
rect 11462 15759 11496 15793
rect 11530 15759 11564 15793
rect 11598 15759 11632 15793
rect 11666 15759 11700 15793
rect 11734 15759 11768 15793
rect 11802 15759 11836 15793
rect 11870 15759 11904 15793
rect 11938 15759 11972 15793
rect 12006 15759 12040 15793
rect 12074 15759 12108 15793
rect 12142 15759 12176 15793
rect 12210 15759 12244 15793
rect 12278 15759 12312 15793
rect 12346 15759 12380 15793
rect 12414 15759 12448 15793
rect 12482 15759 12516 15793
rect 12550 15759 12584 15793
rect 12618 15759 12652 15793
rect 12686 15759 12720 15793
rect 12754 15759 12788 15793
rect 12822 15759 12856 15793
rect 12890 15759 12924 15793
rect 12958 15759 12992 15793
rect 13026 15759 13060 15793
rect 13094 15759 13128 15793
rect 13162 15759 13196 15793
rect 13230 15759 13264 15793
rect 13298 15759 13332 15793
rect 13366 15759 13400 15793
rect 13434 15759 13468 15793
rect 13502 15759 13536 15793
rect 13570 15759 13604 15793
rect 13638 15759 13672 15793
rect 13706 15759 13740 15793
rect 13774 15759 13808 15793
rect 13842 15759 13876 15793
rect 13910 15759 13944 15793
rect 13978 15759 14012 15793
rect 14046 15759 14080 15793
rect 14114 15759 14148 15793
rect 14182 15759 14216 15793
rect 14250 15759 14284 15793
rect 14318 15759 14352 15793
rect 14386 15779 14420 15793
rect 14454 15779 14492 15798
rect 14526 15779 14564 15798
rect 14598 15779 14636 15798
rect 14670 15779 14708 15798
rect 14742 15779 14780 15798
rect 14814 15779 14852 15798
rect 14886 15779 14924 15798
rect 14958 15779 14996 15813
rect 15030 15779 15068 15813
rect 15102 15779 15106 15813
rect 14386 15759 15106 15779
rect 133 15755 15106 15759
rect 67 15744 15106 15755
rect 67 15742 14420 15744
rect 67 15708 68 15742
rect 102 15717 139 15742
rect 173 15717 210 15742
rect 133 15708 139 15717
rect 205 15708 210 15717
rect 244 15708 281 15742
rect 315 15708 352 15742
rect 386 15737 14420 15742
rect 386 15723 3620 15737
rect 3654 15723 3692 15737
rect 3726 15723 3764 15737
rect 3798 15723 3836 15737
rect 3870 15723 3908 15737
rect 3942 15723 3980 15737
rect 4014 15723 4052 15737
rect 4086 15723 4124 15737
rect 4158 15723 4196 15737
rect 4230 15723 4268 15737
rect 4302 15723 4340 15737
rect 4374 15723 4412 15737
rect 4446 15723 4484 15737
rect 4518 15723 4557 15737
rect 4591 15723 4630 15737
rect 4664 15723 4703 15737
rect 4737 15723 4776 15737
rect 4810 15723 4849 15737
rect 4883 15723 4922 15737
rect 4956 15723 4995 15737
rect 5029 15723 5068 15737
rect 5102 15723 5141 15737
rect 5175 15723 5214 15737
rect 5248 15723 5287 15737
rect 5321 15723 5360 15737
rect 5394 15723 14420 15737
rect 386 15719 444 15723
rect 478 15719 513 15723
rect 547 15719 582 15723
rect 616 15719 651 15723
rect 685 15719 720 15723
rect 386 15708 427 15719
rect 67 15683 99 15708
rect 133 15683 171 15708
rect 205 15685 427 15708
rect 478 15689 500 15719
rect 547 15689 573 15719
rect 616 15689 646 15719
rect 685 15689 719 15719
rect 754 15689 789 15723
rect 823 15719 858 15723
rect 892 15719 927 15723
rect 961 15719 996 15723
rect 1030 15719 1065 15723
rect 1099 15719 1134 15723
rect 1168 15719 1203 15723
rect 1237 15719 1272 15723
rect 1306 15719 1341 15723
rect 826 15689 858 15719
rect 899 15689 927 15719
rect 972 15689 996 15719
rect 1045 15689 1065 15719
rect 1118 15689 1134 15719
rect 1191 15689 1203 15719
rect 1264 15689 1272 15719
rect 1337 15689 1341 15719
rect 1375 15719 1410 15723
rect 1375 15689 1376 15719
rect 461 15685 500 15689
rect 534 15685 573 15689
rect 607 15685 646 15689
rect 680 15685 719 15689
rect 753 15685 792 15689
rect 826 15685 865 15689
rect 899 15685 938 15689
rect 972 15685 1011 15689
rect 1045 15685 1084 15689
rect 1118 15685 1157 15689
rect 1191 15685 1230 15689
rect 1264 15685 1303 15689
rect 1337 15685 1376 15689
rect 1444 15719 1479 15723
rect 1513 15719 1548 15723
rect 1582 15719 1617 15723
rect 1651 15719 1686 15723
rect 1720 15719 1755 15723
rect 1789 15719 1824 15723
rect 1858 15719 1893 15723
rect 1927 15719 1962 15723
rect 1996 15719 2031 15723
rect 2065 15719 2100 15723
rect 1444 15689 1449 15719
rect 1513 15689 1521 15719
rect 1582 15689 1593 15719
rect 1651 15689 1665 15719
rect 1720 15689 1737 15719
rect 1789 15689 1809 15719
rect 1858 15689 1881 15719
rect 1927 15689 1953 15719
rect 1996 15689 2025 15719
rect 2065 15689 2097 15719
rect 2134 15689 2169 15723
rect 2203 15689 2238 15723
rect 2272 15719 2307 15723
rect 2341 15719 2376 15723
rect 2410 15719 2445 15723
rect 2479 15719 2514 15723
rect 2548 15719 2583 15723
rect 2617 15719 2652 15723
rect 2686 15719 2721 15723
rect 2755 15719 2790 15723
rect 2824 15719 2859 15723
rect 2893 15719 2928 15723
rect 2962 15719 2996 15723
rect 2275 15689 2307 15719
rect 2347 15689 2376 15719
rect 2419 15689 2445 15719
rect 2491 15689 2514 15719
rect 2563 15689 2583 15719
rect 2635 15689 2652 15719
rect 2707 15689 2721 15719
rect 2779 15689 2790 15719
rect 2851 15689 2859 15719
rect 2923 15689 2928 15719
rect 2995 15689 2996 15719
rect 3030 15719 3064 15723
rect 3098 15719 3132 15723
rect 3166 15719 3200 15723
rect 3234 15719 3268 15723
rect 3302 15719 3336 15723
rect 3370 15719 3404 15723
rect 3438 15719 3472 15723
rect 3506 15719 3540 15723
rect 3030 15689 3033 15719
rect 3098 15689 3105 15719
rect 3166 15689 3177 15719
rect 3234 15689 3249 15719
rect 3302 15689 3321 15719
rect 3370 15689 3393 15719
rect 3438 15689 3465 15719
rect 3506 15689 3537 15719
rect 3574 15689 3608 15723
rect 3654 15703 3676 15723
rect 3726 15703 3744 15723
rect 3798 15703 3812 15723
rect 3870 15703 3880 15723
rect 3942 15703 3948 15723
rect 4014 15703 4016 15723
rect 3642 15689 3676 15703
rect 3710 15689 3744 15703
rect 3778 15689 3812 15703
rect 3846 15689 3880 15703
rect 3914 15689 3948 15703
rect 3982 15689 4016 15703
rect 4050 15703 4052 15723
rect 4118 15703 4124 15723
rect 4186 15703 4196 15723
rect 4254 15703 4268 15723
rect 4322 15703 4340 15723
rect 4390 15703 4412 15723
rect 4458 15703 4484 15723
rect 4526 15703 4557 15723
rect 4050 15689 4084 15703
rect 4118 15689 4152 15703
rect 4186 15689 4220 15703
rect 4254 15689 4288 15703
rect 4322 15689 4356 15703
rect 4390 15689 4424 15703
rect 4458 15689 4492 15703
rect 4526 15689 4560 15703
rect 4594 15689 4628 15723
rect 4664 15703 4696 15723
rect 4737 15703 4764 15723
rect 4810 15703 4832 15723
rect 4883 15703 4900 15723
rect 4956 15703 4968 15723
rect 5029 15703 5036 15723
rect 5102 15703 5104 15723
rect 4662 15689 4696 15703
rect 4730 15689 4764 15703
rect 4798 15689 4832 15703
rect 4866 15689 4900 15703
rect 4934 15689 4968 15703
rect 5002 15689 5036 15703
rect 5070 15689 5104 15703
rect 5138 15703 5141 15723
rect 5206 15703 5214 15723
rect 5274 15703 5287 15723
rect 5342 15703 5360 15723
rect 5138 15689 5172 15703
rect 5206 15689 5240 15703
rect 5274 15689 5308 15703
rect 5342 15689 5376 15703
rect 5410 15689 5444 15723
rect 5478 15689 5512 15723
rect 5546 15689 5580 15723
rect 5614 15689 5648 15723
rect 5682 15689 5716 15723
rect 5750 15689 5784 15723
rect 5818 15689 5852 15723
rect 5886 15689 5920 15723
rect 5954 15689 5988 15723
rect 6022 15689 6056 15723
rect 6090 15689 6124 15723
rect 6158 15689 6192 15723
rect 6226 15689 6260 15723
rect 6294 15689 6328 15723
rect 6362 15689 6396 15723
rect 6430 15689 6464 15723
rect 6498 15689 6532 15723
rect 6566 15689 6600 15723
rect 6634 15689 6668 15723
rect 6702 15689 6736 15723
rect 6770 15689 6804 15723
rect 6838 15689 6872 15723
rect 6906 15689 6940 15723
rect 6974 15689 7008 15723
rect 7042 15689 7076 15723
rect 7110 15689 7144 15723
rect 7178 15689 7212 15723
rect 7246 15689 7280 15723
rect 7314 15689 7348 15723
rect 7382 15689 7416 15723
rect 7450 15689 7484 15723
rect 7518 15689 7552 15723
rect 7586 15689 7620 15723
rect 7654 15689 7688 15723
rect 7722 15689 7756 15723
rect 7790 15689 7824 15723
rect 7858 15689 7892 15723
rect 7926 15689 7960 15723
rect 7994 15689 8028 15723
rect 8062 15689 8096 15723
rect 8130 15689 8164 15723
rect 8198 15689 8232 15723
rect 8266 15689 8300 15723
rect 8334 15689 8368 15723
rect 8402 15689 8436 15723
rect 8470 15689 8504 15723
rect 8538 15689 8572 15723
rect 8606 15689 8640 15723
rect 8674 15689 8708 15723
rect 8742 15689 8776 15723
rect 8810 15689 8844 15723
rect 8878 15689 8912 15723
rect 8946 15689 8980 15723
rect 9014 15689 9048 15723
rect 9082 15689 9116 15723
rect 9150 15689 9184 15723
rect 9218 15689 9252 15723
rect 9286 15689 9320 15723
rect 9354 15689 9388 15723
rect 9422 15689 9456 15723
rect 9490 15689 9524 15723
rect 9558 15689 9592 15723
rect 9626 15689 9660 15723
rect 9694 15689 9728 15723
rect 9762 15689 9796 15723
rect 9830 15689 9864 15723
rect 9898 15689 9932 15723
rect 9966 15689 10000 15723
rect 10034 15689 10068 15723
rect 10102 15689 10136 15723
rect 10170 15689 10204 15723
rect 10238 15689 10272 15723
rect 10306 15689 10340 15723
rect 10374 15689 10408 15723
rect 10442 15689 10476 15723
rect 10510 15689 10544 15723
rect 10578 15689 10612 15723
rect 10646 15689 10680 15723
rect 10714 15689 10748 15723
rect 10782 15689 10816 15723
rect 10850 15689 10884 15723
rect 10918 15689 10952 15723
rect 10986 15689 11020 15723
rect 11054 15689 11088 15723
rect 11122 15689 11156 15723
rect 11190 15689 11224 15723
rect 11258 15689 11292 15723
rect 11326 15689 11360 15723
rect 11394 15689 11428 15723
rect 11462 15689 11496 15723
rect 11530 15689 11564 15723
rect 11598 15689 11632 15723
rect 11666 15689 11700 15723
rect 11734 15689 11768 15723
rect 11802 15689 11836 15723
rect 11870 15689 11904 15723
rect 11938 15689 11972 15723
rect 12006 15689 12040 15723
rect 12074 15689 12108 15723
rect 12142 15689 12176 15723
rect 12210 15689 12244 15723
rect 12278 15689 12312 15723
rect 12346 15689 12380 15723
rect 12414 15689 12448 15723
rect 12482 15689 12516 15723
rect 12550 15689 12584 15723
rect 12618 15689 12652 15723
rect 12686 15689 12720 15723
rect 12754 15689 12788 15723
rect 12822 15689 12856 15723
rect 12890 15689 12924 15723
rect 12958 15689 12992 15723
rect 13026 15689 13060 15723
rect 13094 15689 13128 15723
rect 13162 15689 13196 15723
rect 13230 15689 13264 15723
rect 13298 15689 13332 15723
rect 13366 15689 13400 15723
rect 13434 15689 13468 15723
rect 13502 15689 13536 15723
rect 13570 15689 13604 15723
rect 13638 15689 13672 15723
rect 13706 15689 13740 15723
rect 13774 15689 13808 15723
rect 13842 15689 13876 15723
rect 13910 15689 13944 15723
rect 13978 15689 14012 15723
rect 14046 15689 14080 15723
rect 14114 15689 14148 15723
rect 14182 15689 14216 15723
rect 14250 15689 14284 15723
rect 14318 15689 14352 15723
rect 14386 15710 14420 15723
rect 14454 15710 14492 15744
rect 14526 15710 14564 15744
rect 14598 15710 14636 15744
rect 14670 15710 14708 15744
rect 14742 15710 14780 15744
rect 14814 15710 14852 15744
rect 14886 15710 14924 15744
rect 14958 15710 14996 15744
rect 15030 15710 15068 15744
rect 15102 15710 15106 15744
rect 14386 15689 15106 15710
rect 1410 15685 1449 15689
rect 1483 15685 1521 15689
rect 1555 15685 1593 15689
rect 1627 15685 1665 15689
rect 1699 15685 1737 15689
rect 1771 15685 1809 15689
rect 1843 15685 1881 15689
rect 1915 15685 1953 15689
rect 1987 15685 2025 15689
rect 2059 15685 2097 15689
rect 2131 15685 2169 15689
rect 2203 15685 2241 15689
rect 2275 15685 2313 15689
rect 2347 15685 2385 15689
rect 2419 15685 2457 15689
rect 2491 15685 2529 15689
rect 2563 15685 2601 15689
rect 2635 15685 2673 15689
rect 2707 15685 2745 15689
rect 2779 15685 2817 15689
rect 2851 15685 2889 15689
rect 2923 15685 2961 15689
rect 2995 15685 3033 15689
rect 3067 15685 3105 15689
rect 3139 15685 3177 15689
rect 3211 15685 3249 15689
rect 3283 15685 3321 15689
rect 3355 15685 3393 15689
rect 3427 15685 3465 15689
rect 3499 15685 3537 15689
rect 3571 15685 15106 15689
rect 205 15683 15106 15685
rect 67 15675 15106 15683
rect 67 15673 14420 15675
rect 67 15639 68 15673
rect 102 15639 139 15673
rect 173 15639 210 15673
rect 244 15639 281 15673
rect 315 15639 352 15673
rect 386 15651 14420 15673
rect 386 15647 12660 15651
rect 386 15639 5396 15647
rect 66 15605 69 15639
rect 103 15605 153 15639
rect 187 15605 237 15639
rect 271 15605 321 15639
rect 355 15605 405 15639
rect 439 15616 5396 15639
rect 439 15605 481 15616
rect 66 15604 481 15605
rect 66 15570 68 15604
rect 102 15570 139 15604
rect 173 15570 210 15604
rect 244 15570 281 15604
rect 315 15570 352 15604
rect 386 15583 481 15604
rect 515 15613 5396 15616
rect 5430 15617 12660 15647
rect 12694 15617 12730 15651
rect 12764 15617 12800 15651
rect 12834 15617 12869 15651
rect 12903 15617 12938 15651
rect 12972 15617 13007 15651
rect 13041 15617 13076 15651
rect 13110 15617 13145 15651
rect 13179 15617 13214 15651
rect 13248 15617 13283 15651
rect 13317 15617 13352 15651
rect 13386 15617 13421 15651
rect 13455 15617 13490 15651
rect 13524 15617 13559 15651
rect 13593 15617 13628 15651
rect 13662 15617 13697 15651
rect 13731 15617 13766 15651
rect 13800 15617 13835 15651
rect 13869 15617 13904 15651
rect 13938 15617 13973 15651
rect 14007 15617 14042 15651
rect 14076 15617 14111 15651
rect 14145 15617 14180 15651
rect 14214 15617 14249 15651
rect 14283 15617 14318 15651
rect 14352 15641 14420 15651
rect 14454 15641 14492 15675
rect 14526 15641 14564 15675
rect 14598 15641 14636 15675
rect 14670 15641 14708 15675
rect 14742 15641 14780 15675
rect 14814 15641 14852 15675
rect 14886 15641 14924 15675
rect 14958 15641 14996 15675
rect 15030 15641 15068 15675
rect 15102 15641 15106 15675
rect 14352 15617 15106 15641
rect 5430 15613 15106 15617
rect 515 15607 15106 15613
rect 515 15583 594 15607
rect 386 15570 420 15583
rect 66 15562 420 15570
rect 454 15582 481 15583
rect 66 15535 69 15562
rect 103 15535 153 15562
rect 187 15535 237 15562
rect 271 15535 321 15562
rect 355 15535 405 15562
rect 454 15549 488 15582
rect 522 15573 594 15583
rect 628 15573 663 15607
rect 697 15573 732 15607
rect 766 15573 801 15607
rect 835 15573 870 15607
rect 904 15573 939 15607
rect 973 15573 1008 15607
rect 1042 15573 1077 15607
rect 1111 15573 1146 15607
rect 1180 15573 1215 15607
rect 1249 15573 1284 15607
rect 1318 15573 1353 15607
rect 1387 15573 1422 15607
rect 1456 15573 1491 15607
rect 1525 15573 1560 15607
rect 1594 15573 1629 15607
rect 1663 15573 1698 15607
rect 1732 15573 1767 15607
rect 1801 15573 1836 15607
rect 1870 15573 1904 15607
rect 1938 15573 1972 15607
rect 2006 15573 2040 15607
rect 2074 15573 2108 15607
rect 2142 15573 2176 15607
rect 2210 15573 2244 15607
rect 2278 15573 2312 15607
rect 2346 15573 2380 15607
rect 2414 15573 2448 15607
rect 2482 15573 2516 15607
rect 2550 15573 2584 15607
rect 2618 15573 2652 15607
rect 2686 15573 2720 15607
rect 2754 15573 2788 15607
rect 2822 15573 2856 15607
rect 2890 15573 2924 15607
rect 2958 15573 2992 15607
rect 3026 15573 3060 15607
rect 3094 15573 3128 15607
rect 3162 15573 3196 15607
rect 3230 15573 3264 15607
rect 3298 15573 3332 15607
rect 3366 15573 3400 15607
rect 3434 15573 3468 15607
rect 3502 15573 3536 15607
rect 3570 15573 3604 15607
rect 3638 15573 3672 15607
rect 3706 15573 3740 15607
rect 3774 15573 3808 15607
rect 3842 15573 3876 15607
rect 3910 15573 3944 15607
rect 3978 15573 4012 15607
rect 4046 15573 4080 15607
rect 4114 15573 4148 15607
rect 4182 15573 4216 15607
rect 4250 15573 4284 15607
rect 4318 15573 4352 15607
rect 4386 15573 4420 15607
rect 4454 15573 4488 15607
rect 4522 15573 4556 15607
rect 4590 15573 4624 15607
rect 4658 15573 4692 15607
rect 4726 15573 4760 15607
rect 4794 15573 4828 15607
rect 4862 15573 4896 15607
rect 4930 15573 4964 15607
rect 4998 15573 5032 15607
rect 5066 15573 5100 15607
rect 5134 15573 5168 15607
rect 5202 15573 5236 15607
rect 5270 15573 5304 15607
rect 5338 15573 5372 15607
rect 5406 15573 5430 15607
rect 66 15501 68 15535
rect 103 15528 139 15535
rect 187 15528 210 15535
rect 271 15528 281 15535
rect 102 15501 139 15528
rect 173 15501 210 15528
rect 244 15501 281 15528
rect 315 15528 321 15535
rect 386 15528 405 15535
rect 439 15541 522 15549
rect 439 15528 481 15541
rect 315 15501 352 15528
rect 386 15514 481 15528
rect 515 15514 522 15541
rect 5396 15569 5430 15573
rect 386 15501 420 15514
rect 66 15485 420 15501
rect 454 15507 481 15514
rect 66 15466 69 15485
rect 103 15466 153 15485
rect 187 15466 237 15485
rect 271 15466 321 15485
rect 355 15466 405 15485
rect 454 15480 488 15507
rect 66 15432 68 15466
rect 103 15451 139 15466
rect 187 15451 210 15466
rect 271 15451 281 15466
rect 102 15432 139 15451
rect 173 15432 210 15451
rect 244 15432 281 15451
rect 315 15451 321 15466
rect 386 15451 405 15466
rect 439 15466 522 15480
rect 439 15451 481 15466
rect 315 15432 352 15451
rect 386 15445 481 15451
rect 515 15445 522 15466
rect 386 15432 420 15445
rect 66 15411 420 15432
rect 454 15432 481 15445
rect 454 15411 488 15432
rect 66 15408 522 15411
rect 66 15397 69 15408
rect 103 15397 153 15408
rect 187 15397 237 15408
rect 271 15397 321 15408
rect 355 15397 405 15408
rect 66 15363 68 15397
rect 103 15374 139 15397
rect 187 15374 210 15397
rect 271 15374 281 15397
rect 102 15363 139 15374
rect 173 15363 210 15374
rect 244 15363 281 15374
rect 315 15374 321 15397
rect 386 15374 405 15397
rect 439 15391 522 15408
rect 439 15375 481 15391
rect 515 15375 522 15391
rect 315 15363 352 15374
rect 386 15363 420 15374
rect 66 15341 420 15363
rect 454 15357 481 15375
rect 454 15341 488 15357
rect 66 15331 522 15341
rect 66 15328 69 15331
rect 103 15328 153 15331
rect 187 15328 237 15331
rect 271 15328 321 15331
rect 355 15328 405 15331
rect 66 15294 68 15328
rect 103 15297 139 15328
rect 187 15297 210 15328
rect 271 15297 281 15328
rect 102 15294 139 15297
rect 173 15294 210 15297
rect 244 15294 281 15297
rect 315 15297 321 15328
rect 386 15297 405 15328
rect 439 15316 522 15331
rect 439 15305 481 15316
rect 515 15305 522 15316
rect 315 15294 352 15297
rect 386 15294 420 15297
rect 66 15271 420 15294
rect 454 15282 481 15305
rect 454 15271 488 15282
rect 66 15259 522 15271
rect 66 15225 68 15259
rect 102 15254 139 15259
rect 173 15254 210 15259
rect 244 15254 281 15259
rect 103 15225 139 15254
rect 187 15225 210 15254
rect 271 15225 281 15254
rect 315 15254 352 15259
rect 386 15254 522 15259
rect 315 15225 321 15254
rect 386 15225 405 15254
rect 439 15241 522 15254
rect 439 15235 481 15241
rect 515 15235 522 15241
rect 66 15220 69 15225
rect 103 15220 153 15225
rect 187 15220 237 15225
rect 271 15220 321 15225
rect 355 15220 405 15225
rect 66 15201 420 15220
rect 454 15207 481 15235
rect 454 15201 488 15207
rect 66 15190 522 15201
rect 66 15156 68 15190
rect 102 15177 139 15190
rect 173 15177 210 15190
rect 244 15177 281 15190
rect 103 15156 139 15177
rect 187 15156 210 15177
rect 271 15156 281 15177
rect 315 15177 352 15190
rect 386 15177 522 15190
rect 315 15156 321 15177
rect 386 15156 405 15177
rect 439 15166 522 15177
rect 439 15165 481 15166
rect 515 15165 522 15166
rect 66 15143 69 15156
rect 103 15143 153 15156
rect 187 15143 237 15156
rect 271 15143 321 15156
rect 355 15143 405 15156
rect 66 15131 420 15143
rect 454 15132 481 15165
rect 454 15131 488 15132
rect 66 15121 522 15131
rect 66 15087 68 15121
rect 102 15100 139 15121
rect 173 15100 210 15121
rect 244 15100 281 15121
rect 103 15087 139 15100
rect 187 15087 210 15100
rect 271 15087 281 15100
rect 315 15100 352 15121
rect 386 15100 522 15121
rect 315 15087 321 15100
rect 386 15087 405 15100
rect 439 15095 522 15100
rect 66 15066 69 15087
rect 103 15066 153 15087
rect 187 15066 237 15087
rect 271 15066 321 15087
rect 355 15066 405 15087
rect 454 15091 488 15095
rect 66 15061 420 15066
rect 454 15061 481 15091
rect 66 15057 481 15061
rect 515 15057 522 15061
rect 66 15052 522 15057
rect 66 15018 68 15052
rect 102 15022 139 15052
rect 173 15022 210 15052
rect 244 15022 281 15052
rect 103 15018 139 15022
rect 187 15018 210 15022
rect 271 15018 281 15022
rect 315 15022 352 15052
rect 386 15025 522 15052
rect 386 15022 420 15025
rect 315 15018 321 15022
rect 386 15018 405 15022
rect 66 14988 69 15018
rect 103 14988 153 15018
rect 187 14988 237 15018
rect 271 14988 321 15018
rect 355 14988 405 15018
rect 454 15016 488 15025
rect 454 14991 481 15016
rect 439 14988 481 14991
rect 66 14983 481 14988
rect 66 14949 68 14983
rect 102 14949 139 14983
rect 173 14949 210 14983
rect 244 14949 281 14983
rect 315 14949 352 14983
rect 386 14982 481 14983
rect 515 14982 522 14991
rect 386 14955 522 14982
rect 386 14949 420 14955
rect 66 14944 420 14949
rect 66 14914 69 14944
rect 103 14914 153 14944
rect 187 14914 237 14944
rect 271 14914 321 14944
rect 355 14914 405 14944
rect 454 14941 488 14955
rect 454 14921 481 14941
rect 66 14880 68 14914
rect 103 14910 139 14914
rect 187 14910 210 14914
rect 271 14910 281 14914
rect 102 14880 139 14910
rect 173 14880 210 14910
rect 244 14880 281 14910
rect 315 14910 321 14914
rect 386 14910 405 14914
rect 439 14910 481 14921
rect 315 14880 352 14910
rect 386 14907 481 14910
rect 515 14907 522 14921
rect 386 14885 522 14907
rect 386 14880 420 14885
rect 66 14866 420 14880
rect 454 14867 488 14885
rect 574 15508 5344 15521
rect 574 15474 694 15508
rect 728 15474 766 15508
rect 800 15474 838 15508
rect 872 15474 910 15508
rect 944 15474 982 15508
rect 1016 15474 1054 15508
rect 1088 15474 1126 15508
rect 1160 15474 1198 15508
rect 1232 15474 1270 15508
rect 1304 15474 1342 15508
rect 1376 15474 1414 15508
rect 1448 15474 1486 15508
rect 1520 15474 1558 15508
rect 1592 15474 1630 15508
rect 1664 15474 1702 15508
rect 1736 15474 1774 15508
rect 1808 15474 1846 15508
rect 1880 15474 1918 15508
rect 1952 15474 1990 15508
rect 2024 15474 2062 15508
rect 2096 15474 2134 15508
rect 2168 15474 2206 15508
rect 2240 15474 2278 15508
rect 2312 15474 2350 15508
rect 2384 15474 2422 15508
rect 2456 15474 2494 15508
rect 2528 15474 2566 15508
rect 2600 15474 2638 15508
rect 2672 15474 2710 15508
rect 2744 15474 2782 15508
rect 2816 15474 2854 15508
rect 2888 15474 2926 15508
rect 2960 15474 2998 15508
rect 3032 15474 3070 15508
rect 3104 15474 3142 15508
rect 3176 15474 3214 15508
rect 3248 15474 3286 15508
rect 3320 15474 3358 15508
rect 3392 15474 3430 15508
rect 3464 15474 3502 15508
rect 3536 15474 3574 15508
rect 3608 15474 3646 15508
rect 3680 15474 3718 15508
rect 3752 15474 3790 15508
rect 3824 15474 3862 15508
rect 3896 15474 3935 15508
rect 3969 15504 5344 15508
rect 3969 15474 4017 15504
rect 574 15470 4017 15474
rect 4051 15470 4094 15504
rect 4128 15470 4171 15504
rect 4205 15470 4248 15504
rect 4282 15470 4325 15504
rect 4359 15470 4402 15504
rect 4436 15470 4479 15504
rect 4513 15470 4556 15504
rect 4590 15470 4632 15504
rect 4666 15470 4708 15504
rect 4742 15470 4784 15504
rect 4818 15470 4860 15504
rect 4894 15470 4936 15504
rect 4970 15470 5012 15504
rect 5046 15470 5088 15504
rect 5122 15470 5164 15504
rect 5198 15470 5344 15504
rect 574 15444 5344 15470
rect 574 15436 5228 15444
rect 574 15402 622 15436
rect 656 15421 5228 15436
rect 656 15402 698 15421
rect 732 15420 767 15421
rect 801 15420 836 15421
rect 870 15420 905 15421
rect 939 15420 974 15421
rect 1008 15420 1043 15421
rect 1077 15420 1112 15421
rect 574 15387 698 15402
rect 744 15387 767 15420
rect 817 15387 836 15420
rect 890 15387 905 15420
rect 963 15387 974 15420
rect 1036 15387 1043 15420
rect 1109 15387 1112 15420
rect 1146 15420 1181 15421
rect 1215 15420 1250 15421
rect 1284 15420 1319 15421
rect 1353 15420 1388 15421
rect 1422 15420 1457 15421
rect 1491 15420 1526 15421
rect 1560 15420 1595 15421
rect 1629 15420 1664 15421
rect 1698 15420 1733 15421
rect 1146 15387 1148 15420
rect 1215 15387 1221 15420
rect 1284 15387 1294 15420
rect 1353 15387 1367 15420
rect 1422 15387 1440 15420
rect 1491 15387 1513 15420
rect 1560 15387 1586 15420
rect 1629 15387 1659 15420
rect 1698 15387 1732 15420
rect 1767 15387 1802 15421
rect 1836 15420 1871 15421
rect 1905 15420 1940 15421
rect 1974 15420 2009 15421
rect 2043 15420 2078 15421
rect 2112 15420 2147 15421
rect 2181 15420 2216 15421
rect 2250 15420 2285 15421
rect 2319 15420 2354 15421
rect 1839 15387 1871 15420
rect 1912 15387 1940 15420
rect 1985 15387 2009 15420
rect 2058 15387 2078 15420
rect 2131 15387 2147 15420
rect 2204 15387 2216 15420
rect 2277 15387 2285 15420
rect 2350 15387 2354 15420
rect 2388 15420 2423 15421
rect 2388 15387 2389 15420
rect 574 15386 710 15387
rect 744 15386 783 15387
rect 817 15386 856 15387
rect 890 15386 929 15387
rect 963 15386 1002 15387
rect 1036 15386 1075 15387
rect 1109 15386 1148 15387
rect 1182 15386 1221 15387
rect 1255 15386 1294 15387
rect 1328 15386 1367 15387
rect 1401 15386 1440 15387
rect 1474 15386 1513 15387
rect 1547 15386 1586 15387
rect 1620 15386 1659 15387
rect 1693 15386 1732 15387
rect 1766 15386 1805 15387
rect 1839 15386 1878 15387
rect 1912 15386 1951 15387
rect 1985 15386 2024 15387
rect 2058 15386 2097 15387
rect 2131 15386 2170 15387
rect 2204 15386 2243 15387
rect 2277 15386 2316 15387
rect 2350 15386 2389 15387
rect 2457 15420 2492 15421
rect 2526 15420 2561 15421
rect 2595 15420 2630 15421
rect 2664 15420 2699 15421
rect 2733 15420 2768 15421
rect 2802 15420 2837 15421
rect 2871 15420 2906 15421
rect 2940 15420 2975 15421
rect 2457 15387 2462 15420
rect 2526 15387 2535 15420
rect 2595 15387 2608 15420
rect 2664 15387 2681 15420
rect 2733 15387 2754 15420
rect 2802 15387 2827 15420
rect 2871 15387 2900 15420
rect 2940 15387 2973 15420
rect 3009 15387 3044 15421
rect 3078 15420 3113 15421
rect 3147 15420 3182 15421
rect 3216 15420 3251 15421
rect 3285 15420 3320 15421
rect 3354 15420 3389 15421
rect 3423 15420 3458 15421
rect 3492 15420 3527 15421
rect 3081 15387 3113 15420
rect 3155 15387 3182 15420
rect 3229 15387 3251 15420
rect 3303 15387 3320 15420
rect 3377 15387 3389 15420
rect 3451 15387 3458 15420
rect 3525 15387 3527 15420
rect 3561 15420 3596 15421
rect 3630 15420 3665 15421
rect 3699 15420 3734 15421
rect 3768 15420 3803 15421
rect 3837 15420 3872 15421
rect 3906 15420 3941 15421
rect 3561 15387 3565 15420
rect 3630 15387 3639 15420
rect 3699 15387 3713 15420
rect 3768 15387 3787 15420
rect 3837 15387 3861 15420
rect 3906 15387 3935 15420
rect 3975 15387 4010 15421
rect 4044 15387 4079 15421
rect 4113 15387 4148 15421
rect 4182 15391 4217 15421
rect 4182 15387 4211 15391
rect 4251 15387 4286 15421
rect 4320 15391 4355 15421
rect 4389 15391 4424 15421
rect 4458 15391 4493 15421
rect 4527 15391 4562 15421
rect 4596 15391 4631 15421
rect 4321 15387 4355 15391
rect 4397 15387 4424 15391
rect 4473 15387 4493 15391
rect 4549 15387 4562 15391
rect 4625 15387 4631 15391
rect 4665 15391 4700 15421
rect 4734 15391 4769 15421
rect 4803 15391 4838 15421
rect 4872 15391 4907 15421
rect 4941 15391 4976 15421
rect 5010 15391 5045 15421
rect 4665 15387 4667 15391
rect 4734 15387 4743 15391
rect 4803 15387 4819 15391
rect 4872 15387 4894 15391
rect 4941 15387 4969 15391
rect 5010 15387 5044 15391
rect 5079 15387 5114 15421
rect 5148 15410 5228 15421
rect 5262 15410 5344 15444
rect 5148 15397 5344 15410
rect 5148 15387 5208 15397
rect 2423 15386 2462 15387
rect 2496 15386 2535 15387
rect 2569 15386 2608 15387
rect 2642 15386 2681 15387
rect 2715 15386 2754 15387
rect 2788 15386 2827 15387
rect 2861 15386 2900 15387
rect 2934 15386 2973 15387
rect 3007 15386 3047 15387
rect 3081 15386 3121 15387
rect 3155 15386 3195 15387
rect 3229 15386 3269 15387
rect 3303 15386 3343 15387
rect 3377 15386 3417 15387
rect 3451 15386 3491 15387
rect 3525 15386 3565 15387
rect 3599 15386 3639 15387
rect 3673 15386 3713 15387
rect 3747 15386 3787 15387
rect 3821 15386 3861 15387
rect 3895 15386 3935 15387
rect 3969 15386 4211 15387
rect 574 15362 4211 15386
rect 574 15328 622 15362
rect 656 15357 4211 15362
rect 4245 15357 4287 15387
rect 4321 15357 4363 15387
rect 4397 15357 4439 15387
rect 4473 15357 4515 15387
rect 4549 15357 4591 15387
rect 4625 15357 4667 15387
rect 4701 15357 4743 15387
rect 4777 15357 4819 15387
rect 4853 15357 4894 15387
rect 4928 15357 4969 15387
rect 5003 15357 5044 15387
rect 5078 15363 5208 15387
rect 5242 15372 5344 15397
rect 5078 15357 5228 15363
rect 656 15337 744 15357
rect 656 15328 710 15337
rect 574 15323 710 15328
rect 574 15289 674 15323
rect 708 15303 710 15323
rect 5178 15338 5228 15357
rect 5262 15338 5344 15372
rect 708 15289 744 15303
rect 574 15288 744 15289
rect 574 15254 622 15288
rect 656 15254 744 15288
rect 574 15252 710 15254
rect 574 15218 674 15252
rect 708 15220 710 15252
rect 708 15218 744 15220
rect 574 15214 744 15218
rect 574 15180 622 15214
rect 656 15181 744 15214
rect 778 15271 794 15305
rect 828 15271 862 15305
rect 921 15271 930 15305
rect 993 15271 998 15305
rect 1065 15271 1066 15305
rect 1100 15271 1103 15305
rect 1168 15271 1175 15305
rect 1236 15271 1247 15305
rect 1304 15271 1319 15305
rect 1372 15271 1391 15305
rect 1440 15271 1463 15305
rect 1508 15271 1535 15305
rect 1576 15271 1607 15305
rect 1644 15271 1678 15305
rect 1713 15271 1751 15305
rect 1785 15271 1823 15305
rect 1857 15271 1895 15305
rect 1929 15271 1962 15305
rect 2001 15271 2030 15305
rect 2073 15271 2098 15305
rect 2145 15271 2166 15305
rect 2217 15271 2234 15305
rect 2290 15271 2302 15305
rect 2363 15271 2370 15305
rect 2436 15271 2438 15305
rect 2472 15271 2483 15305
rect 2540 15271 2555 15305
rect 2608 15271 2627 15305
rect 2676 15271 2699 15305
rect 2744 15271 2771 15305
rect 2812 15271 2843 15305
rect 2880 15271 2915 15305
rect 2949 15271 2987 15305
rect 3021 15271 3059 15305
rect 3117 15271 3131 15305
rect 3185 15271 3204 15305
rect 3253 15271 3277 15305
rect 3321 15271 3350 15305
rect 3389 15271 3423 15305
rect 3457 15271 3491 15305
rect 3530 15271 3559 15305
rect 3603 15271 3627 15305
rect 3676 15271 3695 15305
rect 3749 15271 3763 15305
rect 3822 15271 3831 15305
rect 3895 15271 3899 15305
rect 3933 15271 3934 15305
rect 4001 15271 4007 15305
rect 4041 15271 4080 15305
rect 4114 15271 4204 15305
rect 4238 15271 4272 15305
rect 4306 15271 4340 15305
rect 4374 15271 4408 15305
rect 4442 15271 4476 15305
rect 4510 15271 4544 15305
rect 4578 15271 4612 15305
rect 4646 15271 4680 15305
rect 4714 15271 4748 15305
rect 4782 15271 4816 15305
rect 4850 15271 4884 15305
rect 4918 15271 4952 15305
rect 4986 15271 5020 15305
rect 5054 15271 5088 15305
rect 5122 15271 5138 15305
rect 778 15237 5138 15271
rect 778 15204 1764 15237
rect 4145 15204 5138 15237
rect 5178 15300 5344 15338
rect 5178 15284 5228 15300
rect 5178 15250 5208 15284
rect 5262 15266 5344 15300
rect 5242 15250 5344 15266
rect 5178 15228 5344 15250
rect 656 15180 674 15181
rect 574 15147 674 15180
rect 708 15171 744 15181
rect 708 15147 710 15171
rect 574 15140 710 15147
rect 574 15106 622 15140
rect 656 15137 710 15140
rect 1804 15169 1820 15203
rect 1866 15169 1906 15203
rect 1940 15169 1980 15203
rect 2014 15169 2054 15203
rect 2088 15169 2128 15203
rect 2162 15169 2202 15203
rect 2236 15169 2276 15203
rect 2310 15169 2350 15203
rect 2384 15169 2424 15203
rect 2458 15169 2498 15203
rect 2532 15169 2572 15203
rect 2606 15169 2646 15203
rect 2680 15169 2720 15203
rect 2754 15169 2794 15203
rect 2828 15169 2868 15203
rect 2902 15169 2939 15203
rect 2976 15169 3016 15203
rect 3050 15169 3090 15203
rect 3124 15169 3164 15203
rect 3198 15169 3238 15203
rect 3272 15169 3312 15203
rect 3346 15169 3386 15203
rect 3420 15169 3460 15203
rect 3494 15169 3534 15203
rect 3568 15169 3607 15203
rect 3641 15169 3680 15203
rect 3714 15169 3753 15203
rect 3787 15169 3826 15203
rect 3860 15169 3899 15203
rect 3933 15169 3972 15203
rect 4006 15169 4045 15203
rect 4094 15169 4110 15203
rect 5178 15194 5228 15228
rect 5262 15194 5344 15228
rect 5178 15156 5344 15194
rect 5178 15152 5228 15156
rect 744 15137 1764 15152
rect 656 15129 1764 15137
rect 4145 15150 5228 15152
rect 4145 15136 5208 15150
rect 4145 15129 4211 15136
rect 4245 15129 4287 15136
rect 4321 15129 4363 15136
rect 4397 15129 4439 15136
rect 4473 15129 4515 15136
rect 4549 15129 4591 15136
rect 4625 15129 4667 15136
rect 4701 15129 4743 15136
rect 4777 15129 4819 15136
rect 4853 15129 4894 15136
rect 4928 15129 4969 15136
rect 5003 15129 5044 15136
rect 5078 15129 5208 15136
rect 656 15109 794 15129
rect 656 15106 674 15109
rect 574 15075 674 15106
rect 708 15095 794 15109
rect 828 15095 862 15129
rect 896 15095 930 15129
rect 964 15095 998 15129
rect 1032 15095 1066 15129
rect 1100 15095 1134 15129
rect 1168 15095 1202 15129
rect 1236 15095 1270 15129
rect 1304 15095 1338 15129
rect 1372 15095 1406 15129
rect 1440 15095 1474 15129
rect 1508 15095 1542 15129
rect 1576 15095 1610 15129
rect 1644 15095 1678 15129
rect 1712 15095 1962 15129
rect 1996 15095 2030 15129
rect 2064 15095 2098 15129
rect 2132 15095 2166 15129
rect 2200 15095 2234 15129
rect 2268 15095 2302 15129
rect 2336 15095 2370 15129
rect 2404 15095 2438 15129
rect 2472 15095 2506 15129
rect 2540 15095 2574 15129
rect 2608 15095 2642 15129
rect 2676 15095 2710 15129
rect 2744 15095 2778 15129
rect 2812 15095 2846 15129
rect 2880 15095 3083 15129
rect 3117 15095 3151 15129
rect 3185 15095 3219 15129
rect 3253 15095 3287 15129
rect 3321 15095 3355 15129
rect 3389 15095 3423 15129
rect 3457 15095 3491 15129
rect 3525 15095 3559 15129
rect 3593 15095 3627 15129
rect 3661 15095 3695 15129
rect 3729 15095 3763 15129
rect 3797 15095 3831 15129
rect 3865 15095 3899 15129
rect 3933 15095 3967 15129
rect 4001 15095 4204 15129
rect 4245 15102 4272 15129
rect 4321 15102 4340 15129
rect 4397 15102 4408 15129
rect 4473 15102 4476 15129
rect 4238 15095 4272 15102
rect 4306 15095 4340 15102
rect 4374 15095 4408 15102
rect 4442 15095 4476 15102
rect 4510 15102 4515 15129
rect 4578 15102 4591 15129
rect 4646 15102 4667 15129
rect 4714 15102 4743 15129
rect 4510 15095 4544 15102
rect 4578 15095 4612 15102
rect 4646 15095 4680 15102
rect 4714 15095 4748 15102
rect 4782 15095 4816 15129
rect 4853 15102 4884 15129
rect 4928 15102 4952 15129
rect 5003 15102 5020 15129
rect 5078 15102 5088 15129
rect 4850 15095 4884 15102
rect 4918 15095 4952 15102
rect 4986 15095 5020 15102
rect 5054 15095 5088 15102
rect 5122 15116 5208 15129
rect 5262 15122 5344 15156
rect 5242 15116 5344 15122
rect 5122 15095 5344 15116
rect 708 15089 5344 15095
rect 708 15075 710 15089
rect 574 15066 710 15075
rect 574 15032 622 15066
rect 656 15055 710 15066
rect 744 15055 5344 15089
rect 656 15037 5344 15055
rect 656 15032 674 15037
rect 574 15003 674 15032
rect 708 15024 5344 15037
rect 708 15013 2465 15024
rect 2499 15013 2538 15024
rect 2572 15013 2611 15024
rect 2645 15013 2684 15024
rect 2718 15013 2757 15024
rect 2791 15013 2830 15024
rect 2864 15013 2903 15024
rect 2937 15013 2976 15024
rect 3010 15013 3049 15024
rect 3083 15013 3122 15024
rect 3156 15013 3195 15024
rect 3229 15013 3268 15024
rect 3302 15013 3341 15024
rect 3375 15013 3414 15024
rect 3448 15013 3487 15024
rect 3521 15013 3560 15024
rect 3594 15013 3633 15024
rect 3667 15013 3706 15024
rect 3740 15013 3779 15024
rect 3813 15013 3852 15024
rect 3886 15013 3925 15024
rect 3959 15013 3998 15024
rect 4032 15013 4071 15024
rect 4105 15013 4144 15024
rect 4178 15013 4217 15024
rect 4251 15013 4290 15024
rect 4324 15013 4363 15024
rect 4397 15013 4436 15024
rect 4470 15013 4509 15024
rect 4543 15013 4582 15024
rect 4616 15013 4655 15024
rect 4689 15013 4728 15024
rect 4762 15013 4801 15024
rect 4835 15013 4874 15024
rect 708 15007 768 15013
rect 802 15007 837 15013
rect 871 15007 906 15013
rect 940 15007 975 15013
rect 1009 15007 1044 15013
rect 1078 15007 1113 15013
rect 708 15003 710 15007
rect 574 14992 710 15003
rect 574 14958 622 14992
rect 656 14973 710 14992
rect 744 14979 768 15007
rect 817 14979 837 15007
rect 890 14979 906 15007
rect 963 14979 975 15007
rect 1036 14979 1044 15007
rect 1109 14979 1113 15007
rect 1147 15007 1182 15013
rect 1147 14979 1148 15007
rect 744 14973 783 14979
rect 817 14973 856 14979
rect 890 14973 929 14979
rect 963 14973 1002 14979
rect 1036 14973 1075 14979
rect 1109 14973 1148 14979
rect 1216 15007 1251 15013
rect 1285 15007 1320 15013
rect 1354 15007 1389 15013
rect 1423 15007 1458 15013
rect 1492 15007 1527 15013
rect 1561 15007 1596 15013
rect 1630 15007 1665 15013
rect 1699 15007 1734 15013
rect 1216 14979 1221 15007
rect 1285 14979 1294 15007
rect 1354 14979 1367 15007
rect 1423 14979 1440 15007
rect 1492 14979 1513 15007
rect 1561 14979 1586 15007
rect 1630 14979 1659 15007
rect 1699 14979 1732 15007
rect 1768 14979 1803 15013
rect 1837 15007 1872 15013
rect 1906 15007 1941 15013
rect 1975 15007 2010 15013
rect 2044 15007 2079 15013
rect 2113 15007 2148 15013
rect 2182 15007 2217 15013
rect 2251 15007 2286 15013
rect 2320 15007 2355 15013
rect 1839 14979 1872 15007
rect 1912 14979 1941 15007
rect 1984 14979 2010 15007
rect 2056 14979 2079 15007
rect 2128 14979 2148 15007
rect 2200 14979 2217 15007
rect 2272 14979 2286 15007
rect 2344 14979 2355 15007
rect 2389 14979 2424 15013
rect 2458 14990 2465 15013
rect 2527 14990 2538 15013
rect 2596 14990 2611 15013
rect 2665 14990 2684 15013
rect 2734 14990 2757 15013
rect 2803 14990 2830 15013
rect 2872 14990 2903 15013
rect 2458 14979 2493 14990
rect 2527 14979 2562 14990
rect 2596 14979 2631 14990
rect 2665 14979 2700 14990
rect 2734 14979 2769 14990
rect 2803 14979 2838 14990
rect 2872 14979 2907 14990
rect 2941 14979 2976 15013
rect 3010 14979 3045 15013
rect 3083 14990 3114 15013
rect 3156 14990 3183 15013
rect 3229 14990 3252 15013
rect 3302 14990 3321 15013
rect 3375 14990 3390 15013
rect 3448 14990 3459 15013
rect 3521 14990 3528 15013
rect 3594 14990 3597 15013
rect 3079 14979 3114 14990
rect 3148 14979 3183 14990
rect 3217 14979 3252 14990
rect 3286 14979 3321 14990
rect 3355 14979 3390 14990
rect 3424 14979 3459 14990
rect 3493 14979 3528 14990
rect 3562 14979 3597 14990
rect 3631 14990 3633 15013
rect 3700 14990 3706 15013
rect 3769 14990 3779 15013
rect 3838 14990 3852 15013
rect 3907 14990 3925 15013
rect 3976 14990 3998 15013
rect 4045 14990 4071 15013
rect 4114 14990 4144 15013
rect 4183 14990 4217 15013
rect 3631 14979 3666 14990
rect 3700 14979 3735 14990
rect 3769 14979 3804 14990
rect 3838 14979 3873 14990
rect 3907 14979 3942 14990
rect 3976 14979 4011 14990
rect 4045 14979 4080 14990
rect 4114 14979 4149 14990
rect 4183 14979 4218 14990
rect 4252 14979 4287 15013
rect 4324 14990 4356 15013
rect 4397 14990 4425 15013
rect 4470 14990 4494 15013
rect 4543 14990 4563 15013
rect 4616 14990 4632 15013
rect 4689 14990 4701 15013
rect 4762 14990 4770 15013
rect 4835 14990 4839 15013
rect 4321 14979 4356 14990
rect 4390 14979 4425 14990
rect 4459 14979 4494 14990
rect 4528 14979 4563 14990
rect 4597 14979 4632 14990
rect 4666 14979 4701 14990
rect 4735 14979 4770 14990
rect 4804 14979 4839 14990
rect 4873 14990 4874 15013
rect 4908 15013 4947 15024
rect 4981 15013 5020 15024
rect 5054 15013 5094 15024
rect 5128 15013 5168 15024
rect 5202 15013 5344 15024
rect 4873 14979 4908 14990
rect 4942 14990 4947 15013
rect 5011 14990 5020 15013
rect 5080 14990 5094 15013
rect 5149 14990 5168 15013
rect 4942 14979 4977 14990
rect 5011 14979 5046 14990
rect 5080 14979 5115 14990
rect 5149 14979 5184 14990
rect 5218 14979 5344 15013
rect 1182 14973 1221 14979
rect 1255 14973 1294 14979
rect 1328 14973 1367 14979
rect 1401 14973 1440 14979
rect 1474 14973 1513 14979
rect 1547 14973 1586 14979
rect 1620 14973 1659 14979
rect 1693 14973 1732 14979
rect 1766 14973 1805 14979
rect 1839 14973 1878 14979
rect 1912 14973 1950 14979
rect 1984 14973 2022 14979
rect 2056 14973 2094 14979
rect 2128 14973 2166 14979
rect 2200 14973 2238 14979
rect 2272 14973 2310 14979
rect 2344 14973 5344 14979
rect 656 14958 5344 14973
rect 574 14919 5344 14958
rect 574 14885 694 14919
rect 728 14885 768 14919
rect 802 14885 842 14919
rect 876 14885 916 14919
rect 950 14885 990 14919
rect 1024 14885 1064 14919
rect 1098 14885 1138 14919
rect 1172 14885 1212 14919
rect 1246 14885 1286 14919
rect 1320 14885 1360 14919
rect 1394 14885 1434 14919
rect 1468 14885 1507 14919
rect 1541 14885 1580 14919
rect 1614 14885 1653 14919
rect 1687 14885 1726 14919
rect 1760 14885 1799 14919
rect 1833 14885 1872 14919
rect 1906 14885 1945 14919
rect 1979 14885 2018 14919
rect 2052 14885 2091 14919
rect 2125 14885 2164 14919
rect 2198 14885 2237 14919
rect 2271 14885 2310 14919
rect 2344 14885 5344 14919
rect 574 14879 5344 14885
rect 5396 15491 5430 15535
rect 5396 15413 5430 15457
rect 5396 15335 5430 15379
rect 5396 15257 5430 15301
rect 5396 15179 5430 15223
rect 5396 15101 5430 15145
rect 5396 15023 5430 15067
rect 5396 14945 5430 14989
rect 66 14845 69 14866
rect 103 14845 153 14866
rect 187 14845 237 14866
rect 271 14845 321 14866
rect 355 14845 405 14866
rect 454 14851 481 14867
rect 66 14832 68 14845
rect 103 14832 139 14845
rect 187 14832 210 14845
rect 271 14832 281 14845
rect 67 14811 68 14832
rect 102 14811 139 14832
rect 173 14811 210 14832
rect 244 14811 281 14832
rect 315 14832 321 14845
rect 386 14832 405 14845
rect 439 14833 481 14851
rect 515 14833 522 14851
rect 439 14832 522 14833
rect 315 14811 352 14832
rect 386 14827 522 14832
rect 5396 14867 5430 14911
rect 5396 14827 5430 14833
rect 386 14811 5430 14827
rect 67 14793 5430 14811
rect 12580 15606 15106 15607
rect 12580 15581 14420 15606
rect 12580 15547 12660 15581
rect 12694 15547 12730 15581
rect 12764 15547 12800 15581
rect 12834 15547 12869 15581
rect 12903 15547 12938 15581
rect 12972 15547 13007 15581
rect 13041 15547 13076 15581
rect 13110 15547 13145 15581
rect 13179 15547 13214 15581
rect 13248 15547 13283 15581
rect 13317 15547 13352 15581
rect 13386 15547 13421 15581
rect 13455 15547 13490 15581
rect 13524 15547 13559 15581
rect 13593 15547 13628 15581
rect 13662 15547 13697 15581
rect 13731 15547 13766 15581
rect 13800 15547 13835 15581
rect 13869 15547 13904 15581
rect 13938 15547 13973 15581
rect 14007 15547 14042 15581
rect 14076 15547 14111 15581
rect 14145 15547 14180 15581
rect 14214 15547 14249 15581
rect 14283 15547 14318 15581
rect 14352 15572 14420 15581
rect 14454 15572 14492 15606
rect 14526 15572 14564 15606
rect 14598 15572 14636 15606
rect 14670 15572 14708 15606
rect 14742 15572 14780 15606
rect 14814 15572 14852 15606
rect 14886 15572 14924 15606
rect 14958 15572 14996 15606
rect 15030 15572 15068 15606
rect 15102 15572 15106 15606
rect 14352 15547 15106 15572
rect 12580 15537 15106 15547
rect 12580 15511 14420 15537
rect 12580 15477 12660 15511
rect 12694 15477 12730 15511
rect 12764 15477 12800 15511
rect 12834 15477 12869 15511
rect 12903 15477 12938 15511
rect 12972 15477 13007 15511
rect 13041 15477 13076 15511
rect 13110 15477 13145 15511
rect 13179 15477 13214 15511
rect 13248 15477 13283 15511
rect 13317 15477 13352 15511
rect 13386 15477 13421 15511
rect 13455 15477 13490 15511
rect 13524 15477 13559 15511
rect 13593 15477 13628 15511
rect 13662 15477 13697 15511
rect 13731 15477 13766 15511
rect 13800 15477 13835 15511
rect 13869 15477 13904 15511
rect 13938 15477 13973 15511
rect 14007 15477 14042 15511
rect 14076 15477 14111 15511
rect 14145 15477 14180 15511
rect 14214 15477 14249 15511
rect 14283 15477 14318 15511
rect 14352 15503 14420 15511
rect 14454 15503 14492 15537
rect 14526 15503 14564 15537
rect 14598 15503 14636 15537
rect 14670 15503 14708 15537
rect 14742 15503 14780 15537
rect 14814 15503 14852 15537
rect 14886 15503 14924 15537
rect 14958 15503 14996 15537
rect 15030 15503 15068 15537
rect 15102 15503 15106 15537
rect 14352 15477 15106 15503
rect 12580 15468 15106 15477
rect 12580 15464 14420 15468
rect 14454 15464 14492 15468
rect 14526 15464 14564 15468
rect 14598 15464 14636 15468
rect 14670 15464 14708 15468
rect 14742 15464 14780 15468
rect 14814 15464 14852 15468
rect 12580 15441 12860 15464
rect 12894 15441 12934 15464
rect 12968 15441 13008 15464
rect 13042 15441 13082 15464
rect 13116 15441 13156 15464
rect 13190 15441 13230 15464
rect 13264 15441 13304 15464
rect 13338 15441 13378 15464
rect 13412 15441 13452 15464
rect 13486 15441 13526 15464
rect 13560 15441 13600 15464
rect 13634 15441 13674 15464
rect 13708 15441 13748 15464
rect 13782 15441 13822 15464
rect 13856 15441 13896 15464
rect 13930 15441 13970 15464
rect 14004 15441 14044 15464
rect 14078 15441 14118 15464
rect 14152 15441 14191 15464
rect 14225 15441 14264 15464
rect 14298 15441 14337 15464
rect 12580 15407 12660 15441
rect 12694 15407 12730 15441
rect 12764 15407 12800 15441
rect 12834 15430 12860 15441
rect 12903 15430 12934 15441
rect 12834 15407 12869 15430
rect 12903 15407 12938 15430
rect 12972 15407 13007 15441
rect 13042 15430 13076 15441
rect 13116 15430 13145 15441
rect 13190 15430 13214 15441
rect 13264 15430 13283 15441
rect 13338 15430 13352 15441
rect 13412 15430 13421 15441
rect 13486 15430 13490 15441
rect 13041 15407 13076 15430
rect 13110 15407 13145 15430
rect 13179 15407 13214 15430
rect 13248 15407 13283 15430
rect 13317 15407 13352 15430
rect 13386 15407 13421 15430
rect 13455 15407 13490 15430
rect 13524 15430 13526 15441
rect 13593 15430 13600 15441
rect 13662 15430 13674 15441
rect 13731 15430 13748 15441
rect 13800 15430 13822 15441
rect 13869 15430 13896 15441
rect 13938 15430 13970 15441
rect 13524 15407 13559 15430
rect 13593 15407 13628 15430
rect 13662 15407 13697 15430
rect 13731 15407 13766 15430
rect 13800 15407 13835 15430
rect 13869 15407 13904 15430
rect 13938 15407 13973 15430
rect 14007 15407 14042 15441
rect 14078 15430 14111 15441
rect 14152 15430 14180 15441
rect 14225 15430 14249 15441
rect 14298 15430 14318 15441
rect 14371 15430 14410 15464
rect 14454 15434 14483 15464
rect 14526 15434 14556 15464
rect 14598 15434 14629 15464
rect 14670 15434 14702 15464
rect 14742 15434 14775 15464
rect 14814 15434 14848 15464
rect 14886 15434 14924 15468
rect 14958 15434 14996 15468
rect 15030 15434 15068 15468
rect 15102 15434 15106 15468
rect 14444 15430 14483 15434
rect 14517 15430 14556 15434
rect 14590 15430 14629 15434
rect 14663 15430 14702 15434
rect 14736 15430 14775 15434
rect 14809 15430 14848 15434
rect 14882 15430 15106 15434
rect 14076 15407 14111 15430
rect 14145 15407 14180 15430
rect 14214 15407 14249 15430
rect 14283 15407 14318 15430
rect 14352 15407 15106 15430
rect 12580 15399 15106 15407
rect 12580 15382 14420 15399
rect 14454 15382 14492 15399
rect 14526 15382 14564 15399
rect 14598 15382 14636 15399
rect 14670 15382 14708 15399
rect 14742 15382 14780 15399
rect 14814 15382 14852 15399
rect 12580 15371 12860 15382
rect 12894 15371 12934 15382
rect 12968 15371 13008 15382
rect 13042 15371 13082 15382
rect 13116 15371 13156 15382
rect 13190 15371 13230 15382
rect 13264 15371 13304 15382
rect 13338 15371 13378 15382
rect 13412 15371 13452 15382
rect 13486 15371 13526 15382
rect 13560 15371 13600 15382
rect 13634 15371 13674 15382
rect 13708 15371 13748 15382
rect 13782 15371 13822 15382
rect 13856 15371 13896 15382
rect 13930 15371 13970 15382
rect 14004 15371 14044 15382
rect 14078 15371 14118 15382
rect 14152 15371 14191 15382
rect 14225 15371 14264 15382
rect 14298 15371 14337 15382
rect 12580 15337 12660 15371
rect 12694 15337 12730 15371
rect 12764 15337 12800 15371
rect 12834 15348 12860 15371
rect 12903 15348 12934 15371
rect 12834 15337 12869 15348
rect 12903 15337 12938 15348
rect 12972 15337 13007 15371
rect 13042 15348 13076 15371
rect 13116 15348 13145 15371
rect 13190 15348 13214 15371
rect 13264 15348 13283 15371
rect 13338 15348 13352 15371
rect 13412 15348 13421 15371
rect 13486 15348 13490 15371
rect 13041 15337 13076 15348
rect 13110 15337 13145 15348
rect 13179 15337 13214 15348
rect 13248 15337 13283 15348
rect 13317 15337 13352 15348
rect 13386 15337 13421 15348
rect 13455 15337 13490 15348
rect 13524 15348 13526 15371
rect 13593 15348 13600 15371
rect 13662 15348 13674 15371
rect 13731 15348 13748 15371
rect 13800 15348 13822 15371
rect 13869 15348 13896 15371
rect 13938 15348 13970 15371
rect 13524 15337 13559 15348
rect 13593 15337 13628 15348
rect 13662 15337 13697 15348
rect 13731 15337 13766 15348
rect 13800 15337 13835 15348
rect 13869 15337 13904 15348
rect 13938 15337 13973 15348
rect 14007 15337 14042 15371
rect 14078 15348 14111 15371
rect 14152 15348 14180 15371
rect 14225 15348 14249 15371
rect 14298 15348 14318 15371
rect 14371 15348 14410 15382
rect 14454 15365 14483 15382
rect 14526 15365 14556 15382
rect 14598 15365 14629 15382
rect 14670 15365 14702 15382
rect 14742 15365 14775 15382
rect 14814 15365 14848 15382
rect 14886 15365 14924 15399
rect 14958 15365 14996 15399
rect 15030 15365 15068 15399
rect 15102 15365 15106 15399
rect 14444 15348 14483 15365
rect 14517 15348 14556 15365
rect 14590 15348 14629 15365
rect 14663 15348 14702 15365
rect 14736 15348 14775 15365
rect 14809 15348 14848 15365
rect 14882 15348 15106 15365
rect 14076 15337 14111 15348
rect 14145 15337 14180 15348
rect 14214 15337 14249 15348
rect 14283 15337 14318 15348
rect 14352 15337 15106 15348
rect 12580 15330 15106 15337
rect 12580 15301 14420 15330
rect 12580 15267 12660 15301
rect 12694 15267 12730 15301
rect 12764 15267 12800 15301
rect 12834 15300 12869 15301
rect 12903 15300 12938 15301
rect 12834 15267 12860 15300
rect 12903 15267 12934 15300
rect 12972 15267 13007 15301
rect 13041 15300 13076 15301
rect 13110 15300 13145 15301
rect 13179 15300 13214 15301
rect 13248 15300 13283 15301
rect 13317 15300 13352 15301
rect 13386 15300 13421 15301
rect 13455 15300 13490 15301
rect 13042 15267 13076 15300
rect 13116 15267 13145 15300
rect 13190 15267 13214 15300
rect 13264 15267 13283 15300
rect 13338 15267 13352 15300
rect 13412 15267 13421 15300
rect 13486 15267 13490 15300
rect 13524 15300 13559 15301
rect 13593 15300 13628 15301
rect 13662 15300 13697 15301
rect 13731 15300 13766 15301
rect 13800 15300 13835 15301
rect 13869 15300 13904 15301
rect 13938 15300 13973 15301
rect 13524 15267 13526 15300
rect 13593 15267 13600 15300
rect 13662 15267 13674 15300
rect 13731 15267 13748 15300
rect 13800 15267 13822 15300
rect 13869 15267 13896 15300
rect 13938 15267 13970 15300
rect 14007 15267 14042 15301
rect 14076 15300 14111 15301
rect 14145 15300 14180 15301
rect 14214 15300 14249 15301
rect 14283 15300 14318 15301
rect 14352 15300 14420 15301
rect 14454 15300 14492 15330
rect 14526 15300 14564 15330
rect 14598 15300 14636 15330
rect 14670 15300 14708 15330
rect 14742 15300 14780 15330
rect 14814 15300 14852 15330
rect 14078 15267 14111 15300
rect 14152 15267 14180 15300
rect 14225 15267 14249 15300
rect 14298 15267 14318 15300
rect 12580 15266 12860 15267
rect 12894 15266 12934 15267
rect 12968 15266 13008 15267
rect 13042 15266 13082 15267
rect 13116 15266 13156 15267
rect 13190 15266 13230 15267
rect 13264 15266 13304 15267
rect 13338 15266 13378 15267
rect 13412 15266 13452 15267
rect 13486 15266 13526 15267
rect 13560 15266 13600 15267
rect 13634 15266 13674 15267
rect 13708 15266 13748 15267
rect 13782 15266 13822 15267
rect 13856 15266 13896 15267
rect 13930 15266 13970 15267
rect 14004 15266 14044 15267
rect 14078 15266 14118 15267
rect 14152 15266 14191 15267
rect 14225 15266 14264 15267
rect 14298 15266 14337 15267
rect 14371 15266 14410 15300
rect 14454 15296 14483 15300
rect 14526 15296 14556 15300
rect 14598 15296 14629 15300
rect 14670 15296 14702 15300
rect 14742 15296 14775 15300
rect 14814 15296 14848 15300
rect 14886 15296 14924 15330
rect 14958 15296 14996 15330
rect 15030 15296 15068 15330
rect 15102 15296 15106 15330
rect 14444 15266 14483 15296
rect 14517 15266 14556 15296
rect 14590 15266 14629 15296
rect 14663 15266 14702 15296
rect 14736 15266 14775 15296
rect 14809 15266 14848 15296
rect 14882 15266 15106 15296
rect 12580 15261 15106 15266
rect 12580 15231 14420 15261
rect 12580 15197 12660 15231
rect 12694 15197 12730 15231
rect 12764 15197 12800 15231
rect 12834 15218 12869 15231
rect 12903 15218 12938 15231
rect 12834 15197 12860 15218
rect 12903 15197 12934 15218
rect 12972 15197 13007 15231
rect 13041 15218 13076 15231
rect 13110 15218 13145 15231
rect 13179 15218 13214 15231
rect 13248 15218 13283 15231
rect 13317 15218 13352 15231
rect 13386 15218 13421 15231
rect 13455 15218 13490 15231
rect 13042 15197 13076 15218
rect 13116 15197 13145 15218
rect 13190 15197 13214 15218
rect 13264 15197 13283 15218
rect 13338 15197 13352 15218
rect 13412 15197 13421 15218
rect 13486 15197 13490 15218
rect 13524 15218 13559 15231
rect 13593 15218 13628 15231
rect 13662 15218 13697 15231
rect 13731 15218 13766 15231
rect 13800 15218 13835 15231
rect 13869 15218 13904 15231
rect 13938 15218 13973 15231
rect 13524 15197 13526 15218
rect 13593 15197 13600 15218
rect 13662 15197 13674 15218
rect 13731 15197 13748 15218
rect 13800 15197 13822 15218
rect 13869 15197 13896 15218
rect 13938 15197 13970 15218
rect 14007 15197 14042 15231
rect 14076 15218 14111 15231
rect 14145 15218 14180 15231
rect 14214 15218 14249 15231
rect 14283 15218 14318 15231
rect 14352 15227 14420 15231
rect 14454 15227 14492 15261
rect 14526 15227 14564 15261
rect 14598 15227 14636 15261
rect 14670 15227 14708 15261
rect 14742 15227 14780 15261
rect 14814 15227 14852 15261
rect 14886 15227 14924 15261
rect 14958 15227 14996 15261
rect 15030 15227 15068 15261
rect 15102 15227 15106 15261
rect 14352 15218 15106 15227
rect 14078 15197 14111 15218
rect 14152 15197 14180 15218
rect 14225 15197 14249 15218
rect 14298 15197 14318 15218
rect 12580 15184 12860 15197
rect 12894 15184 12934 15197
rect 12968 15184 13008 15197
rect 13042 15184 13082 15197
rect 13116 15184 13156 15197
rect 13190 15184 13230 15197
rect 13264 15184 13304 15197
rect 13338 15184 13378 15197
rect 13412 15184 13452 15197
rect 13486 15184 13526 15197
rect 13560 15184 13600 15197
rect 13634 15184 13674 15197
rect 13708 15184 13748 15197
rect 13782 15184 13822 15197
rect 13856 15184 13896 15197
rect 13930 15184 13970 15197
rect 14004 15184 14044 15197
rect 14078 15184 14118 15197
rect 14152 15184 14191 15197
rect 14225 15184 14264 15197
rect 14298 15184 14337 15197
rect 14371 15184 14410 15218
rect 14444 15192 14483 15218
rect 14517 15192 14556 15218
rect 14590 15192 14629 15218
rect 14663 15192 14702 15218
rect 14736 15192 14775 15218
rect 14809 15192 14848 15218
rect 14882 15192 15106 15218
rect 14454 15184 14483 15192
rect 14526 15184 14556 15192
rect 14598 15184 14629 15192
rect 14670 15184 14702 15192
rect 14742 15184 14775 15192
rect 14814 15184 14848 15192
rect 12580 15161 14420 15184
rect 12580 15127 12660 15161
rect 12694 15127 12730 15161
rect 12764 15127 12800 15161
rect 12834 15136 12869 15161
rect 12903 15136 12938 15161
rect 12834 15127 12860 15136
rect 12903 15127 12934 15136
rect 12972 15127 13007 15161
rect 13041 15136 13076 15161
rect 13110 15136 13145 15161
rect 13179 15136 13214 15161
rect 13248 15136 13283 15161
rect 13317 15136 13352 15161
rect 13386 15136 13421 15161
rect 13455 15136 13490 15161
rect 13042 15127 13076 15136
rect 13116 15127 13145 15136
rect 13190 15127 13214 15136
rect 13264 15127 13283 15136
rect 13338 15127 13352 15136
rect 13412 15127 13421 15136
rect 13486 15127 13490 15136
rect 13524 15136 13559 15161
rect 13593 15136 13628 15161
rect 13662 15136 13697 15161
rect 13731 15136 13766 15161
rect 13800 15136 13835 15161
rect 13869 15136 13904 15161
rect 13938 15136 13973 15161
rect 13524 15127 13526 15136
rect 13593 15127 13600 15136
rect 13662 15127 13674 15136
rect 13731 15127 13748 15136
rect 13800 15127 13822 15136
rect 13869 15127 13896 15136
rect 13938 15127 13970 15136
rect 14007 15127 14042 15161
rect 14076 15136 14111 15161
rect 14145 15136 14180 15161
rect 14214 15136 14249 15161
rect 14283 15136 14318 15161
rect 14352 15158 14420 15161
rect 14454 15158 14492 15184
rect 14526 15158 14564 15184
rect 14598 15158 14636 15184
rect 14670 15158 14708 15184
rect 14742 15158 14780 15184
rect 14814 15158 14852 15184
rect 14886 15158 14924 15192
rect 14958 15158 14996 15192
rect 15030 15158 15068 15192
rect 15102 15158 15106 15192
rect 14352 15136 15106 15158
rect 14078 15127 14111 15136
rect 14152 15127 14180 15136
rect 14225 15127 14249 15136
rect 14298 15127 14318 15136
rect 12580 15102 12860 15127
rect 12894 15102 12934 15127
rect 12968 15102 13008 15127
rect 13042 15102 13082 15127
rect 13116 15102 13156 15127
rect 13190 15102 13230 15127
rect 13264 15102 13304 15127
rect 13338 15102 13378 15127
rect 13412 15102 13452 15127
rect 13486 15102 13526 15127
rect 13560 15102 13600 15127
rect 13634 15102 13674 15127
rect 13708 15102 13748 15127
rect 13782 15102 13822 15127
rect 13856 15102 13896 15127
rect 13930 15102 13970 15127
rect 14004 15102 14044 15127
rect 14078 15102 14118 15127
rect 14152 15102 14191 15127
rect 14225 15102 14264 15127
rect 14298 15102 14337 15127
rect 14371 15102 14410 15136
rect 14444 15123 14483 15136
rect 14517 15123 14556 15136
rect 14590 15123 14629 15136
rect 14663 15123 14702 15136
rect 14736 15123 14775 15136
rect 14809 15123 14848 15136
rect 14882 15123 15106 15136
rect 14454 15102 14483 15123
rect 14526 15102 14556 15123
rect 14598 15102 14629 15123
rect 14670 15102 14702 15123
rect 14742 15102 14775 15123
rect 14814 15102 14848 15123
rect 12580 15091 14420 15102
rect 12580 15057 12660 15091
rect 12694 15057 12730 15091
rect 12764 15057 12800 15091
rect 12834 15057 12869 15091
rect 12903 15057 12938 15091
rect 12972 15057 13007 15091
rect 13041 15057 13076 15091
rect 13110 15057 13145 15091
rect 13179 15057 13214 15091
rect 13248 15057 13283 15091
rect 13317 15057 13352 15091
rect 13386 15057 13421 15091
rect 13455 15057 13490 15091
rect 13524 15057 13559 15091
rect 13593 15057 13628 15091
rect 13662 15057 13697 15091
rect 13731 15057 13766 15091
rect 13800 15057 13835 15091
rect 13869 15057 13904 15091
rect 13938 15057 13973 15091
rect 14007 15057 14042 15091
rect 14076 15057 14111 15091
rect 14145 15057 14180 15091
rect 14214 15057 14249 15091
rect 14283 15057 14318 15091
rect 14352 15089 14420 15091
rect 14454 15089 14492 15102
rect 14526 15089 14564 15102
rect 14598 15089 14636 15102
rect 14670 15089 14708 15102
rect 14742 15089 14780 15102
rect 14814 15089 14852 15102
rect 14886 15089 14924 15123
rect 14958 15089 14996 15123
rect 15030 15089 15068 15123
rect 15102 15089 15106 15123
rect 14352 15057 15106 15089
rect 12580 15054 15106 15057
rect 12580 15021 12860 15054
rect 12894 15021 12934 15054
rect 12968 15021 13008 15054
rect 13042 15021 13082 15054
rect 13116 15021 13156 15054
rect 13190 15021 13230 15054
rect 13264 15021 13304 15054
rect 13338 15021 13378 15054
rect 13412 15021 13452 15054
rect 13486 15021 13526 15054
rect 13560 15021 13600 15054
rect 13634 15021 13674 15054
rect 13708 15021 13748 15054
rect 13782 15021 13822 15054
rect 13856 15021 13896 15054
rect 13930 15021 13970 15054
rect 14004 15021 14044 15054
rect 14078 15021 14118 15054
rect 14152 15021 14191 15054
rect 14225 15021 14264 15054
rect 14298 15021 14337 15054
rect 12580 14987 12660 15021
rect 12694 14987 12730 15021
rect 12764 14987 12800 15021
rect 12834 15020 12860 15021
rect 12903 15020 12934 15021
rect 12834 14987 12869 15020
rect 12903 14987 12938 15020
rect 12972 14987 13007 15021
rect 13042 15020 13076 15021
rect 13116 15020 13145 15021
rect 13190 15020 13214 15021
rect 13264 15020 13283 15021
rect 13338 15020 13352 15021
rect 13412 15020 13421 15021
rect 13486 15020 13490 15021
rect 13041 14987 13076 15020
rect 13110 14987 13145 15020
rect 13179 14987 13214 15020
rect 13248 14987 13283 15020
rect 13317 14987 13352 15020
rect 13386 14987 13421 15020
rect 13455 14987 13490 15020
rect 13524 15020 13526 15021
rect 13593 15020 13600 15021
rect 13662 15020 13674 15021
rect 13731 15020 13748 15021
rect 13800 15020 13822 15021
rect 13869 15020 13896 15021
rect 13938 15020 13970 15021
rect 13524 14987 13559 15020
rect 13593 14987 13628 15020
rect 13662 14987 13697 15020
rect 13731 14987 13766 15020
rect 13800 14987 13835 15020
rect 13869 14987 13904 15020
rect 13938 14987 13973 15020
rect 14007 14987 14042 15021
rect 14078 15020 14111 15021
rect 14152 15020 14180 15021
rect 14225 15020 14249 15021
rect 14298 15020 14318 15021
rect 14371 15020 14410 15054
rect 14454 15020 14483 15054
rect 14526 15020 14556 15054
rect 14598 15020 14629 15054
rect 14670 15020 14702 15054
rect 14742 15020 14775 15054
rect 14814 15020 14848 15054
rect 14886 15020 14924 15054
rect 14958 15020 14996 15054
rect 15030 15020 15068 15054
rect 15102 15020 15106 15054
rect 14076 14987 14111 15020
rect 14145 14987 14180 15020
rect 14214 14987 14249 15020
rect 14283 14987 14318 15020
rect 14352 14987 15106 15020
rect 12580 14985 15106 14987
rect 12580 14972 14420 14985
rect 14454 14972 14492 14985
rect 14526 14972 14564 14985
rect 14598 14972 14636 14985
rect 14670 14972 14708 14985
rect 14742 14972 14780 14985
rect 14814 14972 14852 14985
rect 12580 14951 12860 14972
rect 12894 14951 12934 14972
rect 12968 14951 13008 14972
rect 13042 14951 13082 14972
rect 13116 14951 13156 14972
rect 13190 14951 13230 14972
rect 13264 14951 13304 14972
rect 13338 14951 13378 14972
rect 13412 14951 13452 14972
rect 13486 14951 13526 14972
rect 13560 14951 13600 14972
rect 13634 14951 13674 14972
rect 13708 14951 13748 14972
rect 13782 14951 13822 14972
rect 13856 14951 13896 14972
rect 13930 14951 13970 14972
rect 14004 14951 14044 14972
rect 14078 14951 14118 14972
rect 14152 14951 14191 14972
rect 14225 14951 14264 14972
rect 14298 14951 14337 14972
rect 12580 14917 12660 14951
rect 12694 14917 12730 14951
rect 12764 14917 12800 14951
rect 12834 14938 12860 14951
rect 12903 14938 12934 14951
rect 12834 14917 12869 14938
rect 12903 14917 12938 14938
rect 12972 14917 13007 14951
rect 13042 14938 13076 14951
rect 13116 14938 13145 14951
rect 13190 14938 13214 14951
rect 13264 14938 13283 14951
rect 13338 14938 13352 14951
rect 13412 14938 13421 14951
rect 13486 14938 13490 14951
rect 13041 14917 13076 14938
rect 13110 14917 13145 14938
rect 13179 14917 13214 14938
rect 13248 14917 13283 14938
rect 13317 14917 13352 14938
rect 13386 14917 13421 14938
rect 13455 14917 13490 14938
rect 13524 14938 13526 14951
rect 13593 14938 13600 14951
rect 13662 14938 13674 14951
rect 13731 14938 13748 14951
rect 13800 14938 13822 14951
rect 13869 14938 13896 14951
rect 13938 14938 13970 14951
rect 13524 14917 13559 14938
rect 13593 14917 13628 14938
rect 13662 14917 13697 14938
rect 13731 14917 13766 14938
rect 13800 14917 13835 14938
rect 13869 14917 13904 14938
rect 13938 14917 13973 14938
rect 14007 14917 14042 14951
rect 14078 14938 14111 14951
rect 14152 14938 14180 14951
rect 14225 14938 14249 14951
rect 14298 14938 14318 14951
rect 14371 14938 14410 14972
rect 14454 14951 14483 14972
rect 14526 14951 14556 14972
rect 14598 14951 14629 14972
rect 14670 14951 14702 14972
rect 14742 14951 14775 14972
rect 14814 14951 14848 14972
rect 14886 14951 14924 14985
rect 14958 14951 14996 14985
rect 15030 14951 15068 14985
rect 15102 14951 15106 14985
rect 14444 14938 14483 14951
rect 14517 14938 14556 14951
rect 14590 14938 14629 14951
rect 14663 14938 14702 14951
rect 14736 14938 14775 14951
rect 14809 14938 14848 14951
rect 14882 14938 15106 14951
rect 14076 14917 14111 14938
rect 14145 14917 14180 14938
rect 14214 14917 14249 14938
rect 14283 14917 14318 14938
rect 14352 14917 15106 14938
rect 12580 14916 15106 14917
rect 12580 14882 14420 14916
rect 14454 14882 14492 14916
rect 14526 14882 14564 14916
rect 14598 14882 14636 14916
rect 14670 14882 14708 14916
rect 14742 14882 14780 14916
rect 14814 14882 14852 14916
rect 14886 14882 14924 14916
rect 14958 14882 14996 14916
rect 15030 14882 15068 14916
rect 15102 14882 15106 14916
rect 12580 14881 15106 14882
rect 12580 14847 12660 14881
rect 12694 14847 12730 14881
rect 12764 14847 12800 14881
rect 12834 14847 12869 14881
rect 12903 14847 12938 14881
rect 12972 14847 13007 14881
rect 13041 14847 13076 14881
rect 13110 14847 13145 14881
rect 13179 14847 13214 14881
rect 13248 14847 13283 14881
rect 13317 14847 13352 14881
rect 13386 14847 13421 14881
rect 13455 14847 13490 14881
rect 13524 14847 13559 14881
rect 13593 14847 13628 14881
rect 13662 14847 13697 14881
rect 13731 14847 13766 14881
rect 13800 14847 13835 14881
rect 13869 14847 13904 14881
rect 13938 14847 13973 14881
rect 14007 14847 14042 14881
rect 14076 14847 14111 14881
rect 14145 14847 14180 14881
rect 14214 14847 14249 14881
rect 14283 14847 14318 14881
rect 14352 14847 15106 14881
rect 12580 14813 14420 14847
rect 14454 14813 14492 14847
rect 14526 14813 14564 14847
rect 14598 14813 14636 14847
rect 14670 14813 14708 14847
rect 14742 14813 14780 14847
rect 14814 14813 14852 14847
rect 14886 14813 14924 14847
rect 14958 14813 14996 14847
rect 15030 14813 15068 14847
rect 15102 14813 15106 14847
rect 12580 14793 15106 14813
rect 67 14777 15106 14793
rect 773 10499 787 14137
rect 14337 10499 14351 14137
rect -947 9680 15117 9685
rect -947 9647 -723 9680
rect -947 9613 -932 9647
rect -898 9613 -864 9647
rect -830 9613 -796 9647
rect -762 9646 -723 9647
rect -689 9646 -654 9680
rect -620 9646 -585 9680
rect -551 9646 -516 9680
rect -482 9646 -447 9680
rect -413 9646 -378 9680
rect -344 9646 -309 9680
rect -275 9646 -240 9680
rect -206 9646 -171 9680
rect -137 9646 -102 9680
rect -68 9646 -33 9680
rect -762 9613 -33 9646
rect -947 9612 -33 9613
rect -947 9578 -723 9612
rect -689 9578 -654 9612
rect -620 9578 -585 9612
rect -551 9578 -516 9612
rect -482 9578 -447 9612
rect -413 9578 -378 9612
rect -344 9578 -309 9612
rect -275 9578 -240 9612
rect -206 9578 -171 9612
rect -137 9578 -102 9612
rect -68 9578 -33 9612
rect -947 9571 -33 9578
rect -947 9537 -932 9571
rect -898 9537 -864 9571
rect -830 9537 -796 9571
rect -762 9544 -33 9571
rect -762 9537 -723 9544
rect -947 9510 -723 9537
rect -689 9510 -654 9544
rect -620 9510 -585 9544
rect -551 9510 -516 9544
rect -482 9514 -447 9544
rect -450 9510 -447 9514
rect -413 9514 -378 9544
rect -344 9514 -309 9544
rect -275 9514 -240 9544
rect -206 9514 -171 9544
rect -137 9514 -102 9544
rect -68 9514 -33 9544
rect 14893 9647 15117 9680
rect 14893 9613 14932 9647
rect 14966 9613 15000 9647
rect 15034 9613 15068 9647
rect 15102 9613 15117 9647
rect 14893 9571 15117 9613
rect 14893 9537 14932 9571
rect 14966 9537 15000 9571
rect 15034 9537 15068 9571
rect 15102 9537 15117 9571
rect -413 9510 -411 9514
rect -344 9510 -338 9514
rect -275 9510 -265 9514
rect -206 9510 -192 9514
rect -137 9510 -119 9514
rect -68 9510 -46 9514
rect -947 9495 -484 9510
rect -947 9461 -932 9495
rect -898 9461 -864 9495
rect -830 9461 -796 9495
rect -762 9480 -484 9495
rect -450 9480 -411 9510
rect -377 9480 -338 9510
rect -304 9480 -265 9510
rect -231 9480 -192 9510
rect -158 9480 -119 9510
rect -85 9480 -46 9510
rect 14893 9495 15117 9537
rect -762 9476 -33 9480
rect -762 9461 -723 9476
rect -947 9442 -723 9461
rect -689 9442 -654 9476
rect -620 9442 -585 9476
rect -551 9442 -516 9476
rect -482 9442 -447 9476
rect -413 9442 -378 9476
rect -344 9442 -309 9476
rect -275 9442 -240 9476
rect -206 9442 -171 9476
rect -137 9442 -102 9476
rect -68 9442 -33 9476
rect -947 9428 -33 9442
rect 14893 9461 14932 9495
rect 14966 9461 15000 9495
rect 15034 9461 15068 9495
rect 15102 9461 15117 9495
rect -947 9418 -484 9428
rect -947 9384 -932 9418
rect -898 9384 -864 9418
rect -830 9384 -796 9418
rect -762 9408 -484 9418
rect -450 9408 -411 9428
rect -377 9408 -338 9428
rect -304 9408 -265 9428
rect -231 9408 -192 9428
rect -158 9408 -119 9428
rect -85 9408 -46 9428
rect -762 9384 -723 9408
rect -947 9374 -723 9384
rect -689 9374 -654 9408
rect -620 9374 -585 9408
rect -551 9374 -516 9408
rect -450 9394 -447 9408
rect -482 9374 -447 9394
rect -413 9394 -411 9408
rect -344 9394 -338 9408
rect -275 9394 -265 9408
rect -206 9394 -192 9408
rect -137 9394 -119 9408
rect -68 9394 -46 9408
rect 14893 9418 15117 9461
rect -413 9374 -378 9394
rect -344 9374 -309 9394
rect -275 9374 -240 9394
rect -206 9374 -171 9394
rect -137 9374 -102 9394
rect -68 9374 -33 9394
rect -947 9342 -33 9374
rect 14893 9384 14932 9418
rect 14966 9384 15000 9418
rect 15034 9384 15068 9418
rect 15102 9384 15117 9418
rect -947 9341 -484 9342
rect -947 9307 -932 9341
rect -898 9307 -864 9341
rect -830 9307 -796 9341
rect -762 9340 -484 9341
rect -450 9340 -411 9342
rect -377 9340 -338 9342
rect -304 9340 -265 9342
rect -231 9340 -192 9342
rect -158 9340 -119 9342
rect -85 9340 -46 9342
rect -762 9307 -723 9340
rect -947 9306 -723 9307
rect -689 9306 -654 9340
rect -620 9306 -585 9340
rect -551 9306 -516 9340
rect -450 9308 -447 9340
rect -482 9306 -447 9308
rect -413 9308 -411 9340
rect -344 9308 -338 9340
rect -275 9308 -265 9340
rect -206 9308 -192 9340
rect -137 9308 -119 9340
rect -68 9308 -46 9340
rect 14893 9341 15117 9384
rect -413 9306 -378 9308
rect -344 9306 -309 9308
rect -275 9306 -240 9308
rect -206 9306 -171 9308
rect -137 9306 -102 9308
rect -68 9306 -33 9308
rect -947 9272 -33 9306
rect -947 9264 -723 9272
rect -947 9230 -932 9264
rect -898 9230 -864 9264
rect -830 9230 -796 9264
rect -762 9238 -723 9264
rect -689 9238 -654 9272
rect -620 9238 -585 9272
rect -551 9238 -516 9272
rect -482 9256 -447 9272
rect -450 9238 -447 9256
rect -413 9256 -378 9272
rect -344 9256 -309 9272
rect -275 9256 -240 9272
rect -206 9256 -171 9272
rect -137 9256 -102 9272
rect -68 9256 -33 9272
rect 14893 9307 14932 9341
rect 14966 9307 15000 9341
rect 15034 9307 15068 9341
rect 15102 9307 15117 9341
rect 14893 9264 15117 9307
rect -413 9238 -411 9256
rect -344 9238 -338 9256
rect -275 9238 -265 9256
rect -206 9238 -192 9256
rect -137 9238 -119 9256
rect -68 9238 -46 9256
rect -762 9230 -484 9238
rect -947 9222 -484 9230
rect -450 9222 -411 9238
rect -377 9222 -338 9238
rect -304 9222 -265 9238
rect -231 9222 -192 9238
rect -158 9222 -119 9238
rect -85 9222 -46 9238
rect 14893 9230 14932 9264
rect 14966 9230 15000 9264
rect 15034 9230 15068 9264
rect 15102 9230 15117 9264
rect -947 9204 -33 9222
rect -947 9187 -723 9204
rect -947 9153 -932 9187
rect -898 9153 -864 9187
rect -830 9153 -796 9187
rect -762 9170 -723 9187
rect -689 9170 -654 9204
rect -620 9170 -585 9204
rect -551 9170 -516 9204
rect -482 9170 -447 9204
rect -413 9170 -378 9204
rect -344 9170 -309 9204
rect -275 9170 -240 9204
rect -206 9170 -171 9204
rect -137 9170 -102 9204
rect -68 9170 -33 9204
rect 14893 9187 15117 9230
rect -762 9153 -484 9170
rect -947 9136 -484 9153
rect -450 9136 -411 9170
rect -377 9136 -338 9170
rect -304 9136 -265 9170
rect -231 9136 -192 9170
rect -158 9136 -119 9170
rect -85 9136 -46 9170
rect 14893 9153 14932 9187
rect 14966 9153 15000 9187
rect 15034 9153 15068 9187
rect 15102 9153 15117 9187
rect -947 9110 -723 9136
rect -947 9076 -932 9110
rect -898 9076 -864 9110
rect -830 9076 -796 9110
rect -762 9102 -723 9110
rect -689 9102 -654 9136
rect -620 9102 -585 9136
rect -551 9102 -516 9136
rect -482 9102 -447 9136
rect -413 9102 -378 9136
rect -344 9102 -309 9136
rect -275 9102 -240 9136
rect -206 9102 -171 9136
rect -137 9102 -102 9136
rect -68 9102 -33 9136
rect -762 9076 -33 9102
rect -947 9068 -33 9076
rect -947 9034 -723 9068
rect -689 9034 -654 9068
rect -620 9034 -585 9068
rect -551 9034 -516 9068
rect -482 9034 -447 9068
rect -413 9034 -378 9068
rect -344 9034 -309 9068
rect -275 9034 -240 9068
rect -206 9034 -171 9068
rect -137 9034 -102 9068
rect -68 9034 -33 9068
rect -947 9033 -33 9034
rect -947 8999 -932 9033
rect -898 8999 -864 9033
rect -830 8999 -796 9033
rect -762 9000 -33 9033
rect -762 8999 -723 9000
rect -947 8966 -723 8999
rect -689 8966 -654 9000
rect -620 8966 -585 9000
rect -551 8966 -516 9000
rect -482 8966 -447 9000
rect -413 8966 -378 9000
rect -344 8966 -309 9000
rect -275 8966 -240 9000
rect -206 8966 -171 9000
rect -137 8966 -102 9000
rect -68 8966 -33 9000
rect 14893 9110 15117 9153
rect 14893 9076 14932 9110
rect 14966 9076 15000 9110
rect 15034 9076 15068 9110
rect 15102 9076 15117 9110
rect 14893 9033 15117 9076
rect 14893 8999 14932 9033
rect 14966 8999 15000 9033
rect 15034 8999 15068 9033
rect 15102 8999 15117 9033
rect 14893 8966 15117 8999
rect -947 8961 15117 8966
rect 8367 8808 15102 8809
rect 42 8774 15102 8808
rect 42 8740 68 8774
rect 102 8740 138 8774
rect 172 8740 208 8774
rect 242 8753 278 8774
rect 312 8753 348 8774
rect 382 8753 418 8774
rect 452 8753 488 8774
rect 522 8753 558 8774
rect 592 8753 628 8774
rect 662 8753 698 8774
rect 732 8753 768 8774
rect 802 8753 838 8774
rect 242 8740 248 8753
rect 312 8740 322 8753
rect 382 8740 396 8753
rect 452 8740 470 8753
rect 522 8740 544 8753
rect 592 8740 618 8753
rect 662 8740 691 8753
rect 732 8740 764 8753
rect 802 8740 837 8753
rect 872 8740 908 8774
rect 942 8760 978 8774
rect 1012 8760 1048 8774
rect 1082 8760 1118 8774
rect 1152 8760 1188 8774
rect 1222 8760 1258 8774
rect 1292 8760 1328 8774
rect 1362 8760 1398 8774
rect 1432 8760 1467 8774
rect 1501 8760 1536 8774
rect 1570 8760 1605 8774
rect 1639 8760 1674 8774
rect 1708 8760 1743 8774
rect 1777 8760 1812 8774
rect 946 8740 978 8760
rect 1018 8740 1048 8760
rect 1090 8740 1118 8760
rect 1162 8740 1188 8760
rect 1234 8740 1258 8760
rect 1306 8740 1328 8760
rect 1378 8740 1398 8760
rect 1450 8740 1467 8760
rect 1522 8740 1536 8760
rect 1594 8740 1605 8760
rect 1666 8740 1674 8760
rect 1738 8740 1743 8760
rect 1810 8740 1812 8760
rect 1846 8760 1881 8774
rect 1915 8760 1950 8774
rect 1984 8760 2019 8774
rect 2053 8760 2088 8774
rect 2122 8760 2157 8774
rect 1846 8740 1849 8760
rect 1915 8740 1922 8760
rect 1984 8740 1995 8760
rect 2053 8740 2068 8760
rect 2122 8740 2141 8760
rect 2191 8740 2226 8774
rect 2260 8753 2295 8774
rect 2329 8753 2364 8774
rect 2398 8753 2433 8774
rect 2467 8753 2502 8774
rect 2261 8740 2295 8753
rect 2340 8740 2364 8753
rect 2419 8740 2433 8753
rect 2498 8740 2502 8753
rect 2536 8753 2571 8774
rect 2605 8753 2640 8774
rect 2674 8753 2709 8774
rect 2743 8753 2778 8774
rect 2536 8740 2543 8753
rect 2605 8740 2621 8753
rect 2674 8740 2699 8753
rect 2743 8740 2777 8753
rect 2812 8740 2847 8774
rect 2881 8773 15102 8774
rect 2881 8770 8393 8773
rect 2881 8753 2933 8770
rect 42 8719 248 8740
rect 282 8719 322 8740
rect 356 8719 396 8740
rect 430 8719 470 8740
rect 504 8719 544 8740
rect 578 8719 618 8740
rect 652 8719 691 8740
rect 725 8719 764 8740
rect 798 8719 837 8740
rect 871 8726 912 8740
rect 946 8726 984 8740
rect 1018 8726 1056 8740
rect 1090 8726 1128 8740
rect 1162 8726 1200 8740
rect 1234 8726 1272 8740
rect 1306 8726 1344 8740
rect 1378 8726 1416 8740
rect 1450 8726 1488 8740
rect 1522 8726 1560 8740
rect 1594 8726 1632 8740
rect 1666 8726 1704 8740
rect 1738 8726 1776 8740
rect 1810 8726 1849 8740
rect 1883 8726 1922 8740
rect 1956 8726 1995 8740
rect 2029 8726 2068 8740
rect 2102 8726 2141 8740
rect 2175 8726 2227 8740
rect 871 8719 2227 8726
rect 2261 8719 2306 8740
rect 2340 8719 2385 8740
rect 2419 8719 2464 8740
rect 2498 8719 2543 8740
rect 2577 8719 2621 8740
rect 2655 8719 2699 8740
rect 2733 8719 2777 8740
rect 2811 8719 2855 8740
rect 2889 8719 2933 8753
rect 2967 8736 3002 8770
rect 3036 8753 3071 8770
rect 3045 8736 3071 8753
rect 3105 8736 3139 8770
rect 3173 8736 3207 8770
rect 3241 8736 3275 8770
rect 3309 8736 3343 8770
rect 3377 8736 3411 8770
rect 3445 8760 3479 8770
rect 3445 8736 3477 8760
rect 3513 8736 3547 8770
rect 3581 8760 3615 8770
rect 3649 8760 3683 8770
rect 3717 8760 3751 8770
rect 3785 8760 3819 8770
rect 3853 8760 3887 8770
rect 3921 8760 3955 8770
rect 3989 8760 4023 8770
rect 3584 8736 3615 8760
rect 3657 8736 3683 8760
rect 3730 8736 3751 8760
rect 3803 8736 3819 8760
rect 3876 8736 3887 8760
rect 3949 8736 3955 8760
rect 4022 8736 4023 8760
rect 4057 8760 4091 8770
rect 4125 8760 4159 8770
rect 4193 8760 4227 8770
rect 4261 8760 4295 8770
rect 4329 8760 4363 8770
rect 4397 8760 4431 8770
rect 4057 8736 4061 8760
rect 4125 8736 4134 8760
rect 4193 8736 4207 8760
rect 4261 8736 4280 8760
rect 4329 8736 4353 8760
rect 4397 8736 4426 8760
rect 4465 8736 4499 8770
rect 4533 8736 4567 8770
rect 4601 8760 4635 8770
rect 4669 8760 4703 8770
rect 4737 8760 4771 8770
rect 4805 8760 4839 8770
rect 4873 8760 4907 8770
rect 4941 8760 4975 8770
rect 4606 8736 4635 8760
rect 4679 8736 4703 8760
rect 4752 8736 4771 8760
rect 4825 8736 4839 8760
rect 4898 8736 4907 8760
rect 4971 8736 4975 8760
rect 5009 8760 5043 8770
rect 5077 8760 5111 8770
rect 5145 8760 5179 8770
rect 5213 8760 5247 8770
rect 5281 8760 5315 8770
rect 5349 8760 5383 8770
rect 5417 8760 5451 8770
rect 5009 8736 5010 8760
rect 5077 8736 5083 8760
rect 5145 8736 5156 8760
rect 5213 8736 5229 8760
rect 5281 8736 5302 8760
rect 5349 8736 5375 8760
rect 5417 8736 5448 8760
rect 5485 8736 5519 8770
rect 5553 8760 5587 8770
rect 5621 8760 5655 8770
rect 5689 8760 5723 8770
rect 5757 8760 5791 8770
rect 5825 8760 5859 8770
rect 5893 8760 5927 8770
rect 5961 8760 5995 8770
rect 5555 8736 5587 8760
rect 5628 8736 5655 8760
rect 5701 8736 5723 8760
rect 5774 8736 5791 8760
rect 5847 8736 5859 8760
rect 5920 8736 5927 8760
rect 5993 8736 5995 8760
rect 6029 8760 6063 8770
rect 6097 8760 6131 8770
rect 6165 8760 6199 8770
rect 6233 8760 6267 8770
rect 6301 8760 6335 8770
rect 6369 8760 6403 8770
rect 6437 8760 6471 8770
rect 6029 8736 6032 8760
rect 6097 8736 6105 8760
rect 6165 8736 6178 8760
rect 6233 8736 6251 8760
rect 6301 8736 6324 8760
rect 6369 8736 6397 8760
rect 6437 8736 6470 8760
rect 6505 8736 6539 8770
rect 6573 8760 6607 8770
rect 6641 8760 6675 8770
rect 6709 8760 6743 8770
rect 6777 8760 6811 8770
rect 6845 8760 6879 8770
rect 6913 8760 6947 8770
rect 6577 8736 6607 8760
rect 6650 8736 6675 8760
rect 6723 8736 6743 8760
rect 6796 8736 6811 8760
rect 6869 8736 6879 8760
rect 6942 8736 6947 8760
rect 6981 8760 7015 8770
rect 2967 8719 3011 8736
rect 3045 8726 3477 8736
rect 3511 8726 3550 8736
rect 3584 8726 3623 8736
rect 3657 8726 3696 8736
rect 3730 8726 3769 8736
rect 3803 8726 3842 8736
rect 3876 8726 3915 8736
rect 3949 8726 3988 8736
rect 4022 8726 4061 8736
rect 4095 8726 4134 8736
rect 4168 8726 4207 8736
rect 4241 8726 4280 8736
rect 4314 8726 4353 8736
rect 4387 8726 4426 8736
rect 4460 8726 4499 8736
rect 4533 8726 4572 8736
rect 4606 8726 4645 8736
rect 4679 8726 4718 8736
rect 4752 8726 4791 8736
rect 4825 8726 4864 8736
rect 4898 8726 4937 8736
rect 4971 8726 5010 8736
rect 5044 8726 5083 8736
rect 5117 8726 5156 8736
rect 5190 8726 5229 8736
rect 5263 8726 5302 8736
rect 5336 8726 5375 8736
rect 5409 8726 5448 8736
rect 5482 8726 5521 8736
rect 5555 8726 5594 8736
rect 5628 8726 5667 8736
rect 5701 8726 5740 8736
rect 5774 8726 5813 8736
rect 5847 8726 5886 8736
rect 5920 8726 5959 8736
rect 5993 8726 6032 8736
rect 6066 8726 6105 8736
rect 6139 8726 6178 8736
rect 6212 8726 6251 8736
rect 6285 8726 6324 8736
rect 6358 8726 6397 8736
rect 6431 8726 6470 8736
rect 6504 8726 6543 8736
rect 6577 8726 6616 8736
rect 6650 8726 6689 8736
rect 6723 8726 6762 8736
rect 6796 8726 6835 8736
rect 6869 8726 6908 8736
rect 6942 8726 6981 8736
rect 7049 8760 7083 8770
rect 7117 8760 7151 8770
rect 7185 8760 7219 8770
rect 7253 8760 7287 8770
rect 7321 8760 7355 8770
rect 7389 8760 7423 8770
rect 7049 8736 7054 8760
rect 7117 8736 7127 8760
rect 7185 8736 7200 8760
rect 7253 8736 7273 8760
rect 7321 8736 7346 8760
rect 7389 8736 7419 8760
rect 7457 8736 7491 8770
rect 7525 8760 7559 8770
rect 7593 8760 7627 8770
rect 7661 8760 7695 8770
rect 7729 8760 7763 8770
rect 7797 8760 7831 8770
rect 7865 8760 7899 8770
rect 7933 8760 7967 8770
rect 7526 8736 7559 8760
rect 7599 8736 7627 8760
rect 7672 8736 7695 8760
rect 7745 8736 7763 8760
rect 7818 8736 7831 8760
rect 7891 8736 7899 8760
rect 7964 8736 7967 8760
rect 8001 8760 8035 8770
rect 8069 8760 8103 8770
rect 8137 8760 8171 8770
rect 8205 8760 8239 8770
rect 8273 8760 8307 8770
rect 8341 8760 8393 8770
rect 8427 8760 8462 8773
rect 8496 8760 8531 8773
rect 8565 8760 8600 8773
rect 8634 8760 8669 8773
rect 8703 8760 8738 8773
rect 8772 8760 8807 8773
rect 8841 8760 8876 8773
rect 8910 8760 8945 8773
rect 8979 8760 9014 8773
rect 8001 8736 8003 8760
rect 8069 8736 8075 8760
rect 8137 8736 8147 8760
rect 8205 8736 8219 8760
rect 8273 8736 8291 8760
rect 8341 8736 8363 8760
rect 8427 8739 8435 8760
rect 8496 8739 8507 8760
rect 8565 8739 8579 8760
rect 8634 8739 8651 8760
rect 8703 8739 8723 8760
rect 8772 8739 8795 8760
rect 8841 8739 8867 8760
rect 8910 8739 8939 8760
rect 8979 8739 9011 8760
rect 9048 8739 9083 8773
rect 9117 8739 9152 8773
rect 9186 8760 9220 8773
rect 9254 8760 9288 8773
rect 9322 8760 9356 8773
rect 9390 8760 9424 8773
rect 9458 8760 9492 8773
rect 9526 8760 9560 8773
rect 9594 8760 9628 8773
rect 9662 8760 9696 8773
rect 9189 8739 9220 8760
rect 9261 8739 9288 8760
rect 9333 8739 9356 8760
rect 9405 8739 9424 8760
rect 9477 8739 9492 8760
rect 9549 8739 9560 8760
rect 9621 8739 9628 8760
rect 9693 8739 9696 8760
rect 9730 8760 9764 8773
rect 9798 8760 9832 8773
rect 9866 8760 9900 8773
rect 9934 8760 9968 8773
rect 10002 8760 10036 8773
rect 10070 8760 10104 8773
rect 10138 8760 10172 8773
rect 10206 8760 10240 8773
rect 10274 8760 10308 8773
rect 9730 8739 9731 8760
rect 9798 8739 9803 8760
rect 9866 8739 9875 8760
rect 9934 8739 9947 8760
rect 10002 8739 10019 8760
rect 10070 8739 10091 8760
rect 10138 8739 10163 8760
rect 10206 8739 10235 8760
rect 10274 8739 10307 8760
rect 10342 8739 10376 8773
rect 10410 8760 10444 8773
rect 10478 8760 10512 8773
rect 10546 8760 10580 8773
rect 10614 8760 10648 8773
rect 10682 8760 10716 8773
rect 10750 8760 10784 8773
rect 10818 8760 10852 8773
rect 10886 8760 10920 8773
rect 10413 8739 10444 8760
rect 10485 8739 10512 8760
rect 10557 8739 10580 8760
rect 10629 8739 10648 8760
rect 10701 8739 10716 8760
rect 10773 8739 10784 8760
rect 10845 8739 10852 8760
rect 10917 8739 10920 8760
rect 10954 8760 10988 8773
rect 11022 8760 11056 8773
rect 11090 8760 11124 8773
rect 11158 8760 11192 8773
rect 11226 8760 11260 8773
rect 11294 8760 11328 8773
rect 11362 8760 11396 8773
rect 11430 8760 11464 8773
rect 11498 8760 11532 8773
rect 10954 8739 10955 8760
rect 11022 8739 11027 8760
rect 11090 8739 11099 8760
rect 11158 8739 11171 8760
rect 11226 8739 11243 8760
rect 11294 8739 11315 8760
rect 11362 8739 11387 8760
rect 11430 8739 11459 8760
rect 11498 8739 11531 8760
rect 11566 8739 11600 8773
rect 11634 8760 11668 8773
rect 11702 8760 11736 8773
rect 11770 8760 11804 8773
rect 11838 8760 11872 8773
rect 11906 8760 11940 8773
rect 11974 8760 12008 8773
rect 12042 8760 12076 8773
rect 12110 8760 12144 8773
rect 11637 8739 11668 8760
rect 11709 8739 11736 8760
rect 11781 8739 11804 8760
rect 11853 8739 11872 8760
rect 11925 8739 11940 8760
rect 11997 8739 12008 8760
rect 12069 8739 12076 8760
rect 12141 8739 12144 8760
rect 12178 8760 12212 8773
rect 12246 8760 12280 8773
rect 12314 8760 12348 8773
rect 12382 8760 12416 8773
rect 12450 8760 12484 8773
rect 12518 8760 12552 8773
rect 12586 8760 12620 8773
rect 12654 8760 12688 8773
rect 12722 8760 12756 8773
rect 12178 8739 12179 8760
rect 12246 8739 12251 8760
rect 12314 8739 12323 8760
rect 12382 8739 12395 8760
rect 12450 8739 12467 8760
rect 12518 8739 12539 8760
rect 12586 8739 12611 8760
rect 12654 8739 12683 8760
rect 12722 8739 12755 8760
rect 12790 8739 12824 8773
rect 12858 8760 12892 8773
rect 12926 8760 12960 8773
rect 12994 8760 13028 8773
rect 13062 8760 13096 8773
rect 13130 8760 13164 8773
rect 13198 8760 13232 8773
rect 13266 8760 13300 8773
rect 13334 8760 13368 8773
rect 12861 8739 12892 8760
rect 12933 8739 12960 8760
rect 13005 8739 13028 8760
rect 13077 8739 13096 8760
rect 13149 8739 13164 8760
rect 13221 8739 13232 8760
rect 13293 8739 13300 8760
rect 13365 8739 13368 8760
rect 13402 8760 13436 8773
rect 13470 8760 13504 8773
rect 13538 8760 13572 8773
rect 13606 8760 13640 8773
rect 13674 8760 13708 8773
rect 13742 8760 13776 8773
rect 13810 8760 13844 8773
rect 13878 8760 13912 8773
rect 13946 8760 13980 8773
rect 13402 8739 13403 8760
rect 13470 8739 13475 8760
rect 13538 8739 13547 8760
rect 13606 8739 13619 8760
rect 13674 8739 13691 8760
rect 13742 8739 13763 8760
rect 13810 8739 13835 8760
rect 13878 8739 13907 8760
rect 13946 8739 13979 8760
rect 14014 8739 14048 8773
rect 14082 8760 14116 8773
rect 14150 8760 14184 8773
rect 14218 8760 14252 8773
rect 14286 8760 14320 8773
rect 14354 8760 14388 8773
rect 14422 8760 14456 8773
rect 14490 8760 14524 8773
rect 14558 8760 14592 8773
rect 14085 8739 14116 8760
rect 14157 8739 14184 8760
rect 14229 8739 14252 8760
rect 14301 8739 14320 8760
rect 14373 8739 14388 8760
rect 14445 8739 14456 8760
rect 14517 8739 14524 8760
rect 14589 8739 14592 8760
rect 14626 8760 14660 8773
rect 14694 8760 14728 8773
rect 14762 8760 14796 8773
rect 14830 8760 14864 8773
rect 14626 8739 14627 8760
rect 14694 8739 14699 8760
rect 14762 8739 14771 8760
rect 14830 8739 14843 8760
rect 14898 8739 15102 8773
rect 7015 8726 7054 8736
rect 7088 8726 7127 8736
rect 7161 8726 7200 8736
rect 7234 8726 7273 8736
rect 7307 8726 7346 8736
rect 7380 8726 7419 8736
rect 7453 8726 7492 8736
rect 7526 8726 7565 8736
rect 7599 8726 7638 8736
rect 7672 8726 7711 8736
rect 7745 8726 7784 8736
rect 7818 8726 7857 8736
rect 7891 8726 7930 8736
rect 7964 8726 8003 8736
rect 8037 8726 8075 8736
rect 8109 8726 8147 8736
rect 8181 8726 8219 8736
rect 8253 8726 8291 8736
rect 8325 8726 8363 8736
rect 8397 8726 8435 8739
rect 8469 8726 8507 8739
rect 8541 8726 8579 8739
rect 8613 8726 8651 8739
rect 8685 8726 8723 8739
rect 8757 8726 8795 8739
rect 8829 8726 8867 8739
rect 8901 8726 8939 8739
rect 8973 8726 9011 8739
rect 9045 8726 9083 8739
rect 9117 8726 9155 8739
rect 9189 8726 9227 8739
rect 9261 8726 9299 8739
rect 9333 8726 9371 8739
rect 9405 8726 9443 8739
rect 9477 8726 9515 8739
rect 9549 8726 9587 8739
rect 9621 8726 9659 8739
rect 9693 8726 9731 8739
rect 9765 8726 9803 8739
rect 9837 8726 9875 8739
rect 9909 8726 9947 8739
rect 9981 8726 10019 8739
rect 10053 8726 10091 8739
rect 10125 8726 10163 8739
rect 10197 8726 10235 8739
rect 10269 8726 10307 8739
rect 10341 8726 10379 8739
rect 10413 8726 10451 8739
rect 10485 8726 10523 8739
rect 10557 8726 10595 8739
rect 10629 8726 10667 8739
rect 10701 8726 10739 8739
rect 10773 8726 10811 8739
rect 10845 8726 10883 8739
rect 10917 8726 10955 8739
rect 10989 8726 11027 8739
rect 11061 8726 11099 8739
rect 11133 8726 11171 8739
rect 11205 8726 11243 8739
rect 11277 8726 11315 8739
rect 11349 8726 11387 8739
rect 11421 8726 11459 8739
rect 11493 8726 11531 8739
rect 11565 8726 11603 8739
rect 11637 8726 11675 8739
rect 11709 8726 11747 8739
rect 11781 8726 11819 8739
rect 11853 8726 11891 8739
rect 11925 8726 11963 8739
rect 11997 8726 12035 8739
rect 12069 8726 12107 8739
rect 12141 8726 12179 8739
rect 12213 8726 12251 8739
rect 12285 8726 12323 8739
rect 12357 8726 12395 8739
rect 12429 8726 12467 8739
rect 12501 8726 12539 8739
rect 12573 8726 12611 8739
rect 12645 8726 12683 8739
rect 12717 8726 12755 8739
rect 12789 8726 12827 8739
rect 12861 8726 12899 8739
rect 12933 8726 12971 8739
rect 13005 8726 13043 8739
rect 13077 8726 13115 8739
rect 13149 8726 13187 8739
rect 13221 8726 13259 8739
rect 13293 8726 13331 8739
rect 13365 8726 13403 8739
rect 13437 8726 13475 8739
rect 13509 8726 13547 8739
rect 13581 8726 13619 8739
rect 13653 8726 13691 8739
rect 13725 8726 13763 8739
rect 13797 8726 13835 8739
rect 13869 8726 13907 8739
rect 13941 8726 13979 8739
rect 14013 8726 14051 8739
rect 14085 8726 14123 8739
rect 14157 8726 14195 8739
rect 14229 8726 14267 8739
rect 14301 8726 14339 8739
rect 14373 8726 14411 8739
rect 14445 8726 14483 8739
rect 14517 8726 14555 8739
rect 14589 8726 14627 8739
rect 14661 8726 14699 8739
rect 14733 8726 14771 8739
rect 14805 8726 14843 8739
rect 14877 8726 15102 8739
rect 3045 8721 15102 8726
rect 3045 8719 14932 8721
rect 42 8700 14932 8719
rect 42 8666 68 8700
rect 102 8666 138 8700
rect 172 8666 208 8700
rect 242 8666 278 8700
rect 312 8666 348 8700
rect 382 8666 418 8700
rect 452 8666 488 8700
rect 522 8666 558 8700
rect 592 8666 628 8700
rect 662 8666 698 8700
rect 732 8666 768 8700
rect 802 8666 838 8700
rect 872 8666 908 8700
rect 942 8666 978 8700
rect 1012 8666 1048 8700
rect 1082 8666 1118 8700
rect 1152 8666 1188 8700
rect 1222 8666 1258 8700
rect 1292 8666 1328 8700
rect 1362 8666 1398 8700
rect 1432 8666 1467 8700
rect 1501 8666 1536 8700
rect 1570 8666 1605 8700
rect 1639 8666 1674 8700
rect 1708 8666 1743 8700
rect 1777 8666 1812 8700
rect 1846 8666 1881 8700
rect 1915 8666 1950 8700
rect 1984 8666 2019 8700
rect 2053 8666 2088 8700
rect 2122 8666 2157 8700
rect 2191 8666 2226 8700
rect 2260 8666 2295 8700
rect 2329 8666 2364 8700
rect 2398 8666 2433 8700
rect 2467 8666 2502 8700
rect 2536 8666 2571 8700
rect 2605 8666 2640 8700
rect 2674 8666 2709 8700
rect 2743 8666 2778 8700
rect 2812 8666 2847 8700
rect 2881 8666 2933 8700
rect 2967 8666 3002 8700
rect 3036 8666 3071 8700
rect 3105 8666 3139 8700
rect 3173 8666 3207 8700
rect 3241 8666 3275 8700
rect 3309 8666 3343 8700
rect 3377 8666 3411 8700
rect 3445 8666 3479 8700
rect 3513 8666 3547 8700
rect 3581 8666 3615 8700
rect 3649 8666 3683 8700
rect 3717 8666 3751 8700
rect 3785 8666 3819 8700
rect 3853 8666 3887 8700
rect 3921 8666 3955 8700
rect 3989 8666 4023 8700
rect 4057 8666 4091 8700
rect 4125 8666 4159 8700
rect 4193 8666 4227 8700
rect 4261 8666 4295 8700
rect 4329 8666 4363 8700
rect 4397 8666 4431 8700
rect 4465 8666 4499 8700
rect 4533 8666 4567 8700
rect 4601 8666 4635 8700
rect 4669 8666 4703 8700
rect 4737 8666 4771 8700
rect 4805 8666 4839 8700
rect 4873 8666 4907 8700
rect 4941 8666 4975 8700
rect 5009 8666 5043 8700
rect 5077 8666 5111 8700
rect 5145 8666 5179 8700
rect 5213 8666 5247 8700
rect 5281 8666 5315 8700
rect 5349 8666 5383 8700
rect 5417 8666 5451 8700
rect 5485 8666 5519 8700
rect 5553 8666 5587 8700
rect 5621 8666 5655 8700
rect 5689 8666 5723 8700
rect 5757 8666 5791 8700
rect 5825 8666 5859 8700
rect 5893 8666 5927 8700
rect 5961 8666 5995 8700
rect 6029 8666 6063 8700
rect 6097 8666 6131 8700
rect 6165 8666 6199 8700
rect 6233 8666 6267 8700
rect 6301 8666 6335 8700
rect 6369 8666 6403 8700
rect 6437 8666 6471 8700
rect 6505 8666 6539 8700
rect 6573 8666 6607 8700
rect 6641 8666 6675 8700
rect 6709 8666 6743 8700
rect 6777 8666 6811 8700
rect 6845 8666 6879 8700
rect 6913 8666 6947 8700
rect 6981 8666 7015 8700
rect 7049 8666 7083 8700
rect 7117 8666 7151 8700
rect 7185 8666 7219 8700
rect 7253 8666 7287 8700
rect 7321 8666 7355 8700
rect 7389 8666 7423 8700
rect 7457 8666 7491 8700
rect 7525 8666 7559 8700
rect 7593 8666 7627 8700
rect 7661 8666 7695 8700
rect 7729 8666 7763 8700
rect 7797 8666 7831 8700
rect 7865 8666 7899 8700
rect 7933 8666 7967 8700
rect 8001 8666 8035 8700
rect 8069 8666 8103 8700
rect 8137 8666 8171 8700
rect 8205 8666 8239 8700
rect 8273 8666 8307 8700
rect 8341 8693 14932 8700
rect 8341 8666 8393 8693
rect 42 8659 8393 8666
rect 8427 8659 8462 8693
rect 8496 8659 8531 8693
rect 8565 8659 8600 8693
rect 8634 8659 8669 8693
rect 8703 8659 8738 8693
rect 8772 8659 8807 8693
rect 8841 8659 8876 8693
rect 8910 8659 8945 8693
rect 8979 8659 9014 8693
rect 9048 8659 9083 8693
rect 9117 8659 9152 8693
rect 9186 8659 9220 8693
rect 9254 8659 9288 8693
rect 9322 8659 9356 8693
rect 9390 8659 9424 8693
rect 9458 8659 9492 8693
rect 9526 8659 9560 8693
rect 9594 8659 9628 8693
rect 9662 8659 9696 8693
rect 9730 8659 9764 8693
rect 9798 8659 9832 8693
rect 9866 8659 9900 8693
rect 9934 8659 9968 8693
rect 10002 8659 10036 8693
rect 10070 8659 10104 8693
rect 10138 8659 10172 8693
rect 10206 8659 10240 8693
rect 10274 8659 10308 8693
rect 10342 8659 10376 8693
rect 10410 8659 10444 8693
rect 10478 8659 10512 8693
rect 10546 8659 10580 8693
rect 10614 8659 10648 8693
rect 10682 8659 10716 8693
rect 10750 8659 10784 8693
rect 10818 8659 10852 8693
rect 10886 8659 10920 8693
rect 10954 8659 10988 8693
rect 11022 8659 11056 8693
rect 11090 8659 11124 8693
rect 11158 8659 11192 8693
rect 11226 8659 11260 8693
rect 11294 8659 11328 8693
rect 11362 8659 11396 8693
rect 11430 8659 11464 8693
rect 11498 8659 11532 8693
rect 11566 8659 11600 8693
rect 11634 8659 11668 8693
rect 11702 8659 11736 8693
rect 11770 8659 11804 8693
rect 11838 8659 11872 8693
rect 11906 8659 11940 8693
rect 11974 8659 12008 8693
rect 12042 8659 12076 8693
rect 12110 8659 12144 8693
rect 12178 8659 12212 8693
rect 12246 8659 12280 8693
rect 12314 8659 12348 8693
rect 12382 8659 12416 8693
rect 12450 8659 12484 8693
rect 12518 8659 12552 8693
rect 12586 8659 12620 8693
rect 12654 8659 12688 8693
rect 12722 8659 12756 8693
rect 12790 8659 12824 8693
rect 12858 8659 12892 8693
rect 12926 8659 12960 8693
rect 12994 8659 13028 8693
rect 13062 8659 13096 8693
rect 13130 8659 13164 8693
rect 13198 8659 13232 8693
rect 13266 8659 13300 8693
rect 13334 8659 13368 8693
rect 13402 8659 13436 8693
rect 13470 8659 13504 8693
rect 13538 8659 13572 8693
rect 13606 8659 13640 8693
rect 13674 8659 13708 8693
rect 13742 8659 13776 8693
rect 13810 8659 13844 8693
rect 13878 8659 13912 8693
rect 13946 8659 13980 8693
rect 14014 8659 14048 8693
rect 14082 8659 14116 8693
rect 14150 8659 14184 8693
rect 14218 8659 14252 8693
rect 14286 8659 14320 8693
rect 14354 8659 14388 8693
rect 14422 8659 14456 8693
rect 14490 8659 14524 8693
rect 14558 8659 14592 8693
rect 14626 8659 14660 8693
rect 14694 8659 14728 8693
rect 14762 8659 14796 8693
rect 14830 8659 14864 8693
rect 14898 8687 14932 8693
rect 14966 8687 15000 8721
rect 15034 8687 15068 8721
rect 14898 8659 15102 8687
rect 42 8649 15102 8659
rect 42 8636 14932 8649
rect 42 8626 912 8636
rect 946 8626 984 8636
rect 1018 8626 1056 8636
rect 1090 8626 1128 8636
rect 1162 8626 1200 8636
rect 1234 8626 1272 8636
rect 1306 8626 1344 8636
rect 1378 8626 1416 8636
rect 1450 8626 1488 8636
rect 1522 8626 1560 8636
rect 1594 8626 1632 8636
rect 1666 8626 1704 8636
rect 1738 8626 1776 8636
rect 1810 8626 1849 8636
rect 1883 8626 1922 8636
rect 1956 8626 1995 8636
rect 2029 8626 2068 8636
rect 2102 8626 2141 8636
rect 2175 8630 3477 8636
rect 3511 8630 3550 8636
rect 3584 8630 3623 8636
rect 3657 8630 3696 8636
rect 3730 8630 3769 8636
rect 3803 8630 3842 8636
rect 3876 8630 3915 8636
rect 3949 8630 3988 8636
rect 4022 8630 4061 8636
rect 4095 8630 4134 8636
rect 4168 8630 4207 8636
rect 4241 8630 4280 8636
rect 4314 8630 4353 8636
rect 4387 8630 4426 8636
rect 4460 8630 4499 8636
rect 4533 8630 4572 8636
rect 4606 8630 4645 8636
rect 4679 8630 4718 8636
rect 4752 8630 4791 8636
rect 4825 8630 4864 8636
rect 4898 8630 4937 8636
rect 4971 8630 5010 8636
rect 5044 8630 5083 8636
rect 5117 8630 5156 8636
rect 5190 8630 5229 8636
rect 5263 8630 5302 8636
rect 5336 8630 5375 8636
rect 5409 8630 5448 8636
rect 5482 8630 5521 8636
rect 5555 8630 5594 8636
rect 5628 8630 5667 8636
rect 5701 8630 5740 8636
rect 5774 8630 5813 8636
rect 5847 8630 5886 8636
rect 5920 8630 5959 8636
rect 5993 8630 6032 8636
rect 6066 8630 6105 8636
rect 6139 8630 6178 8636
rect 6212 8630 6251 8636
rect 6285 8630 6324 8636
rect 6358 8630 6397 8636
rect 6431 8630 6470 8636
rect 6504 8630 6543 8636
rect 6577 8630 6616 8636
rect 6650 8630 6689 8636
rect 6723 8630 6762 8636
rect 6796 8630 6835 8636
rect 6869 8630 6908 8636
rect 6942 8630 6981 8636
rect 2175 8626 2933 8630
rect 42 8592 68 8626
rect 102 8592 138 8626
rect 172 8592 208 8626
rect 242 8592 278 8626
rect 312 8592 348 8626
rect 382 8592 418 8626
rect 452 8592 488 8626
rect 522 8592 558 8626
rect 592 8592 628 8626
rect 662 8592 698 8626
rect 732 8592 768 8626
rect 802 8592 838 8626
rect 872 8592 908 8626
rect 946 8602 978 8626
rect 1018 8602 1048 8626
rect 1090 8602 1118 8626
rect 1162 8602 1188 8626
rect 1234 8602 1258 8626
rect 1306 8602 1328 8626
rect 1378 8602 1398 8626
rect 1450 8602 1467 8626
rect 1522 8602 1536 8626
rect 1594 8602 1605 8626
rect 1666 8602 1674 8626
rect 1738 8602 1743 8626
rect 1810 8602 1812 8626
rect 942 8592 978 8602
rect 1012 8592 1048 8602
rect 1082 8592 1118 8602
rect 1152 8592 1188 8602
rect 1222 8592 1258 8602
rect 1292 8592 1328 8602
rect 1362 8592 1398 8602
rect 1432 8592 1467 8602
rect 1501 8592 1536 8602
rect 1570 8592 1605 8602
rect 1639 8592 1674 8602
rect 1708 8592 1743 8602
rect 1777 8592 1812 8602
rect 1846 8602 1849 8626
rect 1915 8602 1922 8626
rect 1984 8602 1995 8626
rect 2053 8602 2068 8626
rect 2122 8602 2141 8626
rect 1846 8592 1881 8602
rect 1915 8592 1950 8602
rect 1984 8592 2019 8602
rect 2053 8592 2088 8602
rect 2122 8592 2157 8602
rect 2191 8592 2226 8626
rect 2260 8592 2295 8626
rect 2329 8592 2364 8626
rect 2398 8592 2433 8626
rect 2467 8592 2502 8626
rect 2536 8592 2571 8626
rect 2605 8592 2640 8626
rect 2674 8592 2709 8626
rect 2743 8592 2778 8626
rect 2812 8592 2847 8626
rect 2881 8596 2933 8626
rect 2967 8596 3002 8630
rect 3036 8596 3071 8630
rect 3105 8596 3139 8630
rect 3173 8596 3207 8630
rect 3241 8596 3275 8630
rect 3309 8596 3343 8630
rect 3377 8596 3411 8630
rect 3445 8602 3477 8630
rect 3445 8596 3479 8602
rect 3513 8596 3547 8630
rect 3584 8602 3615 8630
rect 3657 8602 3683 8630
rect 3730 8602 3751 8630
rect 3803 8602 3819 8630
rect 3876 8602 3887 8630
rect 3949 8602 3955 8630
rect 4022 8602 4023 8630
rect 3581 8596 3615 8602
rect 3649 8596 3683 8602
rect 3717 8596 3751 8602
rect 3785 8596 3819 8602
rect 3853 8596 3887 8602
rect 3921 8596 3955 8602
rect 3989 8596 4023 8602
rect 4057 8602 4061 8630
rect 4125 8602 4134 8630
rect 4193 8602 4207 8630
rect 4261 8602 4280 8630
rect 4329 8602 4353 8630
rect 4397 8602 4426 8630
rect 4057 8596 4091 8602
rect 4125 8596 4159 8602
rect 4193 8596 4227 8602
rect 4261 8596 4295 8602
rect 4329 8596 4363 8602
rect 4397 8596 4431 8602
rect 4465 8596 4499 8630
rect 4533 8596 4567 8630
rect 4606 8602 4635 8630
rect 4679 8602 4703 8630
rect 4752 8602 4771 8630
rect 4825 8602 4839 8630
rect 4898 8602 4907 8630
rect 4971 8602 4975 8630
rect 4601 8596 4635 8602
rect 4669 8596 4703 8602
rect 4737 8596 4771 8602
rect 4805 8596 4839 8602
rect 4873 8596 4907 8602
rect 4941 8596 4975 8602
rect 5009 8602 5010 8630
rect 5077 8602 5083 8630
rect 5145 8602 5156 8630
rect 5213 8602 5229 8630
rect 5281 8602 5302 8630
rect 5349 8602 5375 8630
rect 5417 8602 5448 8630
rect 5009 8596 5043 8602
rect 5077 8596 5111 8602
rect 5145 8596 5179 8602
rect 5213 8596 5247 8602
rect 5281 8596 5315 8602
rect 5349 8596 5383 8602
rect 5417 8596 5451 8602
rect 5485 8596 5519 8630
rect 5555 8602 5587 8630
rect 5628 8602 5655 8630
rect 5701 8602 5723 8630
rect 5774 8602 5791 8630
rect 5847 8602 5859 8630
rect 5920 8602 5927 8630
rect 5993 8602 5995 8630
rect 5553 8596 5587 8602
rect 5621 8596 5655 8602
rect 5689 8596 5723 8602
rect 5757 8596 5791 8602
rect 5825 8596 5859 8602
rect 5893 8596 5927 8602
rect 5961 8596 5995 8602
rect 6029 8602 6032 8630
rect 6097 8602 6105 8630
rect 6165 8602 6178 8630
rect 6233 8602 6251 8630
rect 6301 8602 6324 8630
rect 6369 8602 6397 8630
rect 6437 8602 6470 8630
rect 6029 8596 6063 8602
rect 6097 8596 6131 8602
rect 6165 8596 6199 8602
rect 6233 8596 6267 8602
rect 6301 8596 6335 8602
rect 6369 8596 6403 8602
rect 6437 8596 6471 8602
rect 6505 8596 6539 8630
rect 6577 8602 6607 8630
rect 6650 8602 6675 8630
rect 6723 8602 6743 8630
rect 6796 8602 6811 8630
rect 6869 8602 6879 8630
rect 6942 8602 6947 8630
rect 6573 8596 6607 8602
rect 6641 8596 6675 8602
rect 6709 8596 6743 8602
rect 6777 8596 6811 8602
rect 6845 8596 6879 8602
rect 6913 8596 6947 8602
rect 7015 8630 7054 8636
rect 7088 8630 7127 8636
rect 7161 8630 7200 8636
rect 7234 8630 7273 8636
rect 7307 8630 7346 8636
rect 7380 8630 7419 8636
rect 7453 8630 7492 8636
rect 7526 8630 7565 8636
rect 7599 8630 7638 8636
rect 7672 8630 7711 8636
rect 7745 8630 7784 8636
rect 7818 8630 7857 8636
rect 7891 8630 7930 8636
rect 7964 8630 8003 8636
rect 8037 8630 8075 8636
rect 8109 8630 8147 8636
rect 8181 8630 8219 8636
rect 8253 8630 8291 8636
rect 8325 8630 8363 8636
rect 6981 8596 7015 8602
rect 7049 8602 7054 8630
rect 7117 8602 7127 8630
rect 7185 8602 7200 8630
rect 7253 8602 7273 8630
rect 7321 8602 7346 8630
rect 7389 8602 7419 8630
rect 7049 8596 7083 8602
rect 7117 8596 7151 8602
rect 7185 8596 7219 8602
rect 7253 8596 7287 8602
rect 7321 8596 7355 8602
rect 7389 8596 7423 8602
rect 7457 8596 7491 8630
rect 7526 8602 7559 8630
rect 7599 8602 7627 8630
rect 7672 8602 7695 8630
rect 7745 8602 7763 8630
rect 7818 8602 7831 8630
rect 7891 8602 7899 8630
rect 7964 8602 7967 8630
rect 7525 8596 7559 8602
rect 7593 8596 7627 8602
rect 7661 8596 7695 8602
rect 7729 8596 7763 8602
rect 7797 8596 7831 8602
rect 7865 8596 7899 8602
rect 7933 8596 7967 8602
rect 8001 8602 8003 8630
rect 8069 8602 8075 8630
rect 8137 8602 8147 8630
rect 8205 8602 8219 8630
rect 8273 8602 8291 8630
rect 8341 8602 8363 8630
rect 8397 8613 8435 8636
rect 8469 8613 8507 8636
rect 8541 8613 8579 8636
rect 8613 8613 8651 8636
rect 8685 8613 8723 8636
rect 8757 8613 8795 8636
rect 8829 8613 8867 8636
rect 8901 8613 8939 8636
rect 8973 8613 9011 8636
rect 9045 8613 9083 8636
rect 9117 8613 9155 8636
rect 9189 8613 9227 8636
rect 9261 8613 9299 8636
rect 9333 8613 9371 8636
rect 9405 8613 9443 8636
rect 9477 8613 9515 8636
rect 9549 8613 9587 8636
rect 9621 8613 9659 8636
rect 9693 8613 9731 8636
rect 9765 8613 9803 8636
rect 9837 8613 9875 8636
rect 9909 8613 9947 8636
rect 9981 8613 10019 8636
rect 10053 8613 10091 8636
rect 10125 8613 10163 8636
rect 10197 8613 10235 8636
rect 10269 8613 10307 8636
rect 10341 8613 10379 8636
rect 10413 8613 10451 8636
rect 10485 8613 10523 8636
rect 10557 8613 10595 8636
rect 10629 8613 10667 8636
rect 10701 8613 10739 8636
rect 10773 8613 10811 8636
rect 10845 8613 10883 8636
rect 10917 8613 10955 8636
rect 10989 8613 11027 8636
rect 11061 8613 11099 8636
rect 11133 8613 11171 8636
rect 11205 8613 11243 8636
rect 11277 8613 11315 8636
rect 11349 8613 11387 8636
rect 11421 8613 11459 8636
rect 11493 8613 11531 8636
rect 11565 8613 11603 8636
rect 11637 8613 11675 8636
rect 11709 8613 11747 8636
rect 11781 8613 11819 8636
rect 11853 8613 11891 8636
rect 11925 8613 11963 8636
rect 11997 8613 12035 8636
rect 12069 8613 12107 8636
rect 12141 8613 12179 8636
rect 12213 8613 12251 8636
rect 12285 8613 12323 8636
rect 12357 8613 12395 8636
rect 12429 8613 12467 8636
rect 12501 8613 12539 8636
rect 12573 8613 12611 8636
rect 12645 8613 12683 8636
rect 12717 8613 12755 8636
rect 12789 8613 12827 8636
rect 12861 8613 12899 8636
rect 12933 8613 12971 8636
rect 13005 8613 13043 8636
rect 13077 8613 13115 8636
rect 13149 8613 13187 8636
rect 13221 8613 13259 8636
rect 13293 8613 13331 8636
rect 13365 8613 13403 8636
rect 13437 8613 13475 8636
rect 13509 8613 13547 8636
rect 13581 8613 13619 8636
rect 13653 8613 13691 8636
rect 13725 8613 13763 8636
rect 13797 8613 13835 8636
rect 13869 8613 13907 8636
rect 13941 8613 13979 8636
rect 14013 8613 14051 8636
rect 14085 8613 14123 8636
rect 14157 8613 14195 8636
rect 14229 8613 14267 8636
rect 14301 8613 14339 8636
rect 14373 8613 14411 8636
rect 14445 8613 14483 8636
rect 14517 8613 14555 8636
rect 14589 8613 14627 8636
rect 14661 8613 14699 8636
rect 14733 8613 14771 8636
rect 14805 8613 14843 8636
rect 14877 8615 14932 8636
rect 14966 8615 15000 8649
rect 15034 8615 15068 8649
rect 14877 8613 15102 8615
rect 8427 8602 8435 8613
rect 8496 8602 8507 8613
rect 8565 8602 8579 8613
rect 8634 8602 8651 8613
rect 8703 8602 8723 8613
rect 8772 8602 8795 8613
rect 8841 8602 8867 8613
rect 8910 8602 8939 8613
rect 8979 8602 9011 8613
rect 8001 8596 8035 8602
rect 8069 8596 8103 8602
rect 8137 8596 8171 8602
rect 8205 8596 8239 8602
rect 8273 8596 8307 8602
rect 8341 8596 8393 8602
rect 2881 8592 8393 8596
rect 42 8579 8393 8592
rect 8427 8579 8462 8602
rect 8496 8579 8531 8602
rect 8565 8579 8600 8602
rect 8634 8579 8669 8602
rect 8703 8579 8738 8602
rect 8772 8579 8807 8602
rect 8841 8579 8876 8602
rect 8910 8579 8945 8602
rect 8979 8579 9014 8602
rect 9048 8579 9083 8613
rect 9117 8579 9152 8613
rect 9189 8602 9220 8613
rect 9261 8602 9288 8613
rect 9333 8602 9356 8613
rect 9405 8602 9424 8613
rect 9477 8602 9492 8613
rect 9549 8602 9560 8613
rect 9621 8602 9628 8613
rect 9693 8602 9696 8613
rect 9186 8579 9220 8602
rect 9254 8579 9288 8602
rect 9322 8579 9356 8602
rect 9390 8579 9424 8602
rect 9458 8579 9492 8602
rect 9526 8579 9560 8602
rect 9594 8579 9628 8602
rect 9662 8579 9696 8602
rect 9730 8602 9731 8613
rect 9798 8602 9803 8613
rect 9866 8602 9875 8613
rect 9934 8602 9947 8613
rect 10002 8602 10019 8613
rect 10070 8602 10091 8613
rect 10138 8602 10163 8613
rect 10206 8602 10235 8613
rect 10274 8602 10307 8613
rect 9730 8579 9764 8602
rect 9798 8579 9832 8602
rect 9866 8579 9900 8602
rect 9934 8579 9968 8602
rect 10002 8579 10036 8602
rect 10070 8579 10104 8602
rect 10138 8579 10172 8602
rect 10206 8579 10240 8602
rect 10274 8579 10308 8602
rect 10342 8579 10376 8613
rect 10413 8602 10444 8613
rect 10485 8602 10512 8613
rect 10557 8602 10580 8613
rect 10629 8602 10648 8613
rect 10701 8602 10716 8613
rect 10773 8602 10784 8613
rect 10845 8602 10852 8613
rect 10917 8602 10920 8613
rect 10410 8579 10444 8602
rect 10478 8579 10512 8602
rect 10546 8579 10580 8602
rect 10614 8579 10648 8602
rect 10682 8579 10716 8602
rect 10750 8579 10784 8602
rect 10818 8579 10852 8602
rect 10886 8579 10920 8602
rect 10954 8602 10955 8613
rect 11022 8602 11027 8613
rect 11090 8602 11099 8613
rect 11158 8602 11171 8613
rect 11226 8602 11243 8613
rect 11294 8602 11315 8613
rect 11362 8602 11387 8613
rect 11430 8602 11459 8613
rect 11498 8602 11531 8613
rect 10954 8579 10988 8602
rect 11022 8579 11056 8602
rect 11090 8579 11124 8602
rect 11158 8579 11192 8602
rect 11226 8579 11260 8602
rect 11294 8579 11328 8602
rect 11362 8579 11396 8602
rect 11430 8579 11464 8602
rect 11498 8579 11532 8602
rect 11566 8579 11600 8613
rect 11637 8602 11668 8613
rect 11709 8602 11736 8613
rect 11781 8602 11804 8613
rect 11853 8602 11872 8613
rect 11925 8602 11940 8613
rect 11997 8602 12008 8613
rect 12069 8602 12076 8613
rect 12141 8602 12144 8613
rect 11634 8579 11668 8602
rect 11702 8579 11736 8602
rect 11770 8579 11804 8602
rect 11838 8579 11872 8602
rect 11906 8579 11940 8602
rect 11974 8579 12008 8602
rect 12042 8579 12076 8602
rect 12110 8579 12144 8602
rect 12178 8602 12179 8613
rect 12246 8602 12251 8613
rect 12314 8602 12323 8613
rect 12382 8602 12395 8613
rect 12450 8602 12467 8613
rect 12518 8602 12539 8613
rect 12586 8602 12611 8613
rect 12654 8602 12683 8613
rect 12722 8602 12755 8613
rect 12178 8579 12212 8602
rect 12246 8579 12280 8602
rect 12314 8579 12348 8602
rect 12382 8579 12416 8602
rect 12450 8579 12484 8602
rect 12518 8579 12552 8602
rect 12586 8579 12620 8602
rect 12654 8579 12688 8602
rect 12722 8579 12756 8602
rect 12790 8579 12824 8613
rect 12861 8602 12892 8613
rect 12933 8602 12960 8613
rect 13005 8602 13028 8613
rect 13077 8602 13096 8613
rect 13149 8602 13164 8613
rect 13221 8602 13232 8613
rect 13293 8602 13300 8613
rect 13365 8602 13368 8613
rect 12858 8579 12892 8602
rect 12926 8579 12960 8602
rect 12994 8579 13028 8602
rect 13062 8579 13096 8602
rect 13130 8579 13164 8602
rect 13198 8579 13232 8602
rect 13266 8579 13300 8602
rect 13334 8579 13368 8602
rect 13402 8602 13403 8613
rect 13470 8602 13475 8613
rect 13538 8602 13547 8613
rect 13606 8602 13619 8613
rect 13674 8602 13691 8613
rect 13742 8602 13763 8613
rect 13810 8602 13835 8613
rect 13878 8602 13907 8613
rect 13946 8602 13979 8613
rect 13402 8579 13436 8602
rect 13470 8579 13504 8602
rect 13538 8579 13572 8602
rect 13606 8579 13640 8602
rect 13674 8579 13708 8602
rect 13742 8579 13776 8602
rect 13810 8579 13844 8602
rect 13878 8579 13912 8602
rect 13946 8579 13980 8602
rect 14014 8579 14048 8613
rect 14085 8602 14116 8613
rect 14157 8602 14184 8613
rect 14229 8602 14252 8613
rect 14301 8602 14320 8613
rect 14373 8602 14388 8613
rect 14445 8602 14456 8613
rect 14517 8602 14524 8613
rect 14589 8602 14592 8613
rect 14082 8579 14116 8602
rect 14150 8579 14184 8602
rect 14218 8579 14252 8602
rect 14286 8579 14320 8602
rect 14354 8579 14388 8602
rect 14422 8579 14456 8602
rect 14490 8579 14524 8602
rect 14558 8579 14592 8602
rect 14626 8602 14627 8613
rect 14694 8602 14699 8613
rect 14762 8602 14771 8613
rect 14830 8602 14843 8613
rect 14626 8579 14660 8602
rect 14694 8579 14728 8602
rect 14762 8579 14796 8602
rect 14830 8579 14864 8602
rect 14898 8579 15102 8613
rect 42 8577 15102 8579
rect 42 8560 14932 8577
rect 42 8552 2933 8560
rect 42 8518 68 8552
rect 102 8518 138 8552
rect 172 8518 208 8552
rect 242 8518 278 8552
rect 312 8518 348 8552
rect 382 8518 418 8552
rect 452 8518 488 8552
rect 522 8518 558 8552
rect 592 8518 628 8552
rect 662 8518 698 8552
rect 732 8518 768 8552
rect 802 8518 838 8552
rect 872 8518 908 8552
rect 942 8518 978 8552
rect 1012 8518 1048 8552
rect 1082 8518 1118 8552
rect 1152 8518 1188 8552
rect 1222 8518 1258 8552
rect 1292 8518 1328 8552
rect 1362 8518 1398 8552
rect 1432 8518 1467 8552
rect 1501 8518 1536 8552
rect 1570 8518 1605 8552
rect 1639 8518 1674 8552
rect 1708 8518 1743 8552
rect 1777 8518 1812 8552
rect 1846 8518 1881 8552
rect 1915 8518 1950 8552
rect 1984 8518 2019 8552
rect 2053 8518 2088 8552
rect 2122 8518 2157 8552
rect 2191 8518 2226 8552
rect 2260 8518 2295 8552
rect 2329 8518 2364 8552
rect 2398 8518 2433 8552
rect 2467 8518 2502 8552
rect 2536 8518 2571 8552
rect 2605 8518 2640 8552
rect 2674 8518 2709 8552
rect 2743 8518 2778 8552
rect 2812 8518 2847 8552
rect 2881 8526 2933 8552
rect 2967 8526 3002 8560
rect 3036 8526 3071 8560
rect 3105 8526 3139 8560
rect 3173 8526 3207 8560
rect 3241 8526 3275 8560
rect 3309 8526 3343 8560
rect 3377 8526 3411 8560
rect 3445 8526 3479 8560
rect 3513 8526 3547 8560
rect 3581 8526 3615 8560
rect 3649 8526 3683 8560
rect 3717 8526 3751 8560
rect 3785 8526 3819 8560
rect 3853 8526 3887 8560
rect 3921 8526 3955 8560
rect 3989 8526 4023 8560
rect 4057 8526 4091 8560
rect 4125 8526 4159 8560
rect 4193 8526 4227 8560
rect 4261 8526 4295 8560
rect 4329 8526 4363 8560
rect 4397 8526 4431 8560
rect 4465 8526 4499 8560
rect 4533 8526 4567 8560
rect 4601 8526 4635 8560
rect 4669 8526 4703 8560
rect 4737 8526 4771 8560
rect 4805 8526 4839 8560
rect 4873 8526 4907 8560
rect 4941 8526 4975 8560
rect 5009 8526 5043 8560
rect 5077 8526 5111 8560
rect 5145 8526 5179 8560
rect 5213 8526 5247 8560
rect 5281 8526 5315 8560
rect 5349 8526 5383 8560
rect 5417 8526 5451 8560
rect 5485 8526 5519 8560
rect 5553 8526 5587 8560
rect 5621 8526 5655 8560
rect 5689 8526 5723 8560
rect 5757 8526 5791 8560
rect 5825 8526 5859 8560
rect 5893 8526 5927 8560
rect 5961 8526 5995 8560
rect 6029 8526 6063 8560
rect 6097 8526 6131 8560
rect 6165 8526 6199 8560
rect 6233 8526 6267 8560
rect 6301 8526 6335 8560
rect 6369 8526 6403 8560
rect 6437 8526 6471 8560
rect 6505 8526 6539 8560
rect 6573 8526 6607 8560
rect 6641 8526 6675 8560
rect 6709 8526 6743 8560
rect 6777 8526 6811 8560
rect 6845 8526 6879 8560
rect 6913 8526 6947 8560
rect 6981 8526 7015 8560
rect 7049 8526 7083 8560
rect 7117 8526 7151 8560
rect 7185 8526 7219 8560
rect 7253 8526 7287 8560
rect 7321 8526 7355 8560
rect 7389 8526 7423 8560
rect 7457 8526 7491 8560
rect 7525 8526 7559 8560
rect 7593 8526 7627 8560
rect 7661 8526 7695 8560
rect 7729 8526 7763 8560
rect 7797 8526 7831 8560
rect 7865 8526 7899 8560
rect 7933 8526 7967 8560
rect 8001 8526 8035 8560
rect 8069 8526 8103 8560
rect 8137 8526 8171 8560
rect 8205 8526 8239 8560
rect 8273 8526 8307 8560
rect 8341 8546 14932 8560
rect 8341 8533 13992 8546
rect 14026 8533 14076 8546
rect 14110 8543 14932 8546
rect 14966 8543 15000 8577
rect 15034 8543 15068 8577
rect 14110 8533 15102 8543
rect 8341 8526 8393 8533
rect 2881 8518 8393 8526
rect 42 8499 8393 8518
rect 8427 8499 8462 8533
rect 8496 8499 8531 8533
rect 8565 8499 8600 8533
rect 8634 8499 8669 8533
rect 8703 8499 8738 8533
rect 8772 8499 8807 8533
rect 8841 8499 8876 8533
rect 8910 8499 8945 8533
rect 8979 8499 9014 8533
rect 9048 8499 9083 8533
rect 9117 8499 9152 8533
rect 9186 8499 9220 8533
rect 9254 8499 9288 8533
rect 9322 8499 9356 8533
rect 9390 8499 9424 8533
rect 9458 8499 9492 8533
rect 9526 8499 9560 8533
rect 9594 8499 9628 8533
rect 9662 8499 9696 8533
rect 9730 8499 9764 8533
rect 9798 8499 9832 8533
rect 9866 8499 9900 8533
rect 9934 8499 9968 8533
rect 10002 8499 10036 8533
rect 10070 8499 10104 8533
rect 10138 8499 10172 8533
rect 10206 8499 10240 8533
rect 10274 8499 10308 8533
rect 10342 8499 10376 8533
rect 10410 8499 10444 8533
rect 10478 8499 10512 8533
rect 10546 8499 10580 8533
rect 10614 8499 10648 8533
rect 10682 8499 10716 8533
rect 10750 8499 10784 8533
rect 10818 8499 10852 8533
rect 10886 8499 10920 8533
rect 10954 8499 10988 8533
rect 11022 8499 11056 8533
rect 11090 8499 11124 8533
rect 11158 8499 11192 8533
rect 11226 8499 11260 8533
rect 11294 8499 11328 8533
rect 11362 8499 11396 8533
rect 11430 8499 11464 8533
rect 11498 8499 11532 8533
rect 11566 8499 11600 8533
rect 11634 8499 11668 8533
rect 11702 8499 11736 8533
rect 11770 8499 11804 8533
rect 11838 8499 11872 8533
rect 11906 8499 11940 8533
rect 11974 8499 12008 8533
rect 12042 8499 12076 8533
rect 12110 8499 12144 8533
rect 12178 8499 12212 8533
rect 12246 8499 12280 8533
rect 12314 8499 12348 8533
rect 12382 8499 12416 8533
rect 12450 8499 12484 8533
rect 12518 8499 12552 8533
rect 12586 8499 12620 8533
rect 12654 8499 12688 8533
rect 12722 8499 12756 8533
rect 12790 8499 12824 8533
rect 12858 8499 12892 8533
rect 12926 8499 12960 8533
rect 12994 8499 13028 8533
rect 13062 8499 13096 8533
rect 13130 8499 13164 8533
rect 13198 8499 13232 8533
rect 13266 8499 13300 8533
rect 13334 8499 13368 8533
rect 13402 8499 13436 8533
rect 13470 8499 13504 8533
rect 13538 8499 13572 8533
rect 13606 8499 13640 8533
rect 13674 8499 13708 8533
rect 13742 8499 13776 8533
rect 13810 8499 13844 8533
rect 13878 8499 13912 8533
rect 13946 8499 13980 8533
rect 14026 8512 14048 8533
rect 14110 8512 14116 8533
rect 14014 8499 14048 8512
rect 14082 8499 14116 8512
rect 14150 8499 14184 8533
rect 14218 8512 14252 8533
rect 14286 8512 14320 8533
rect 14354 8512 14388 8533
rect 14422 8512 14456 8533
rect 14490 8512 14524 8533
rect 14219 8499 14252 8512
rect 14291 8499 14320 8512
rect 14363 8499 14388 8512
rect 14435 8499 14456 8512
rect 14507 8499 14524 8512
rect 14558 8499 14592 8533
rect 14626 8499 14660 8533
rect 14694 8499 14728 8533
rect 14762 8499 14796 8533
rect 14830 8499 14864 8533
rect 14898 8505 15102 8533
rect 14898 8499 14932 8505
rect 42 8490 14185 8499
rect 42 8484 2933 8490
rect 34 8460 136 8484
rect 34 8426 68 8460
rect 102 8426 136 8460
rect 34 8392 136 8426
rect 34 8358 68 8392
rect 102 8358 136 8392
rect 2907 8456 2933 8484
rect 2967 8456 3002 8490
rect 3036 8456 3071 8490
rect 3105 8456 3139 8490
rect 3173 8456 3207 8490
rect 3241 8456 3275 8490
rect 3309 8456 3343 8490
rect 3377 8456 3411 8490
rect 3445 8456 3479 8490
rect 3513 8456 3547 8490
rect 3581 8456 3615 8490
rect 3649 8456 3683 8490
rect 3717 8456 3751 8490
rect 3785 8456 3819 8490
rect 3853 8456 3887 8490
rect 3921 8456 3955 8490
rect 3989 8456 4023 8490
rect 4057 8456 4091 8490
rect 4125 8456 4159 8490
rect 4193 8456 4227 8490
rect 4261 8456 4295 8490
rect 4329 8456 4363 8490
rect 4397 8456 4431 8490
rect 4465 8456 4499 8490
rect 4533 8456 4567 8490
rect 4601 8456 4635 8490
rect 4669 8456 4703 8490
rect 4737 8456 4771 8490
rect 4805 8456 4839 8490
rect 4873 8456 4907 8490
rect 4941 8456 4975 8490
rect 5009 8456 5043 8490
rect 5077 8456 5111 8490
rect 5145 8456 5179 8490
rect 5213 8456 5247 8490
rect 5281 8456 5315 8490
rect 5349 8456 5383 8490
rect 5417 8456 5451 8490
rect 5485 8456 5519 8490
rect 5553 8456 5587 8490
rect 5621 8456 5655 8490
rect 5689 8456 5723 8490
rect 5757 8456 5791 8490
rect 5825 8456 5859 8490
rect 5893 8456 5927 8490
rect 5961 8456 5995 8490
rect 6029 8456 6063 8490
rect 6097 8456 6131 8490
rect 6165 8456 6199 8490
rect 6233 8456 6267 8490
rect 6301 8456 6335 8490
rect 6369 8456 6403 8490
rect 6437 8456 6471 8490
rect 6505 8456 6539 8490
rect 6573 8456 6607 8490
rect 6641 8456 6675 8490
rect 6709 8456 6743 8490
rect 6777 8456 6811 8490
rect 6845 8456 6879 8490
rect 6913 8456 6947 8490
rect 6981 8456 7015 8490
rect 7049 8456 7083 8490
rect 7117 8456 7151 8490
rect 7185 8456 7219 8490
rect 7253 8456 7287 8490
rect 7321 8456 7355 8490
rect 7389 8456 7423 8490
rect 7457 8456 7491 8490
rect 7525 8456 7559 8490
rect 7593 8456 7627 8490
rect 7661 8456 7695 8490
rect 7729 8456 7763 8490
rect 7797 8456 7831 8490
rect 7865 8456 7899 8490
rect 7933 8456 7967 8490
rect 8001 8456 8035 8490
rect 8069 8456 8103 8490
rect 8137 8456 8171 8490
rect 8205 8456 8239 8490
rect 8273 8456 8307 8490
rect 8341 8478 14185 8490
rect 14219 8478 14257 8499
rect 14291 8478 14329 8499
rect 14363 8478 14401 8499
rect 14435 8478 14473 8499
rect 14507 8478 14932 8499
rect 8341 8474 14932 8478
rect 8341 8456 13992 8474
rect 2907 8453 13992 8456
rect 14026 8453 14076 8474
rect 14110 8471 14932 8474
rect 14966 8471 15000 8505
rect 15034 8471 15068 8505
rect 14110 8462 15102 8471
rect 14110 8453 14614 8462
rect 14648 8453 14692 8462
rect 14726 8453 14770 8462
rect 14804 8453 14848 8462
rect 14882 8453 14926 8462
rect 2907 8420 8393 8453
rect 2907 8386 2933 8420
rect 2967 8386 3002 8420
rect 3036 8386 3071 8420
rect 3105 8386 3139 8420
rect 3173 8386 3207 8420
rect 3241 8386 3275 8420
rect 3309 8386 3343 8420
rect 3377 8386 3411 8420
rect 3445 8386 3479 8420
rect 3513 8386 3547 8420
rect 3581 8386 3615 8420
rect 3649 8386 3683 8420
rect 3717 8386 3751 8420
rect 3785 8386 3819 8420
rect 3853 8386 3887 8420
rect 3921 8386 3955 8420
rect 3989 8386 4023 8420
rect 4057 8386 4091 8420
rect 4125 8386 4159 8420
rect 4193 8386 4227 8420
rect 4261 8386 4295 8420
rect 4329 8386 4363 8420
rect 4397 8386 4431 8420
rect 4465 8386 4499 8420
rect 4533 8386 4567 8420
rect 4601 8386 4635 8420
rect 4669 8386 4703 8420
rect 4737 8386 4771 8420
rect 4805 8386 4839 8420
rect 4873 8386 4907 8420
rect 4941 8386 4975 8420
rect 5009 8386 5043 8420
rect 5077 8386 5111 8420
rect 5145 8386 5179 8420
rect 5213 8386 5247 8420
rect 5281 8386 5315 8420
rect 5349 8386 5383 8420
rect 5417 8386 5451 8420
rect 5485 8386 5519 8420
rect 5553 8386 5587 8420
rect 5621 8386 5655 8420
rect 5689 8386 5723 8420
rect 5757 8386 5791 8420
rect 5825 8386 5859 8420
rect 5893 8386 5927 8420
rect 5961 8386 5995 8420
rect 6029 8386 6063 8420
rect 6097 8386 6131 8420
rect 6165 8386 6199 8420
rect 6233 8386 6267 8420
rect 6301 8386 6335 8420
rect 6369 8386 6403 8420
rect 6437 8386 6471 8420
rect 6505 8386 6539 8420
rect 6573 8386 6607 8420
rect 6641 8386 6675 8420
rect 6709 8386 6743 8420
rect 6777 8386 6811 8420
rect 6845 8386 6879 8420
rect 6913 8386 6947 8420
rect 6981 8386 7015 8420
rect 7049 8386 7083 8420
rect 7117 8386 7151 8420
rect 7185 8386 7219 8420
rect 7253 8386 7287 8420
rect 7321 8386 7355 8420
rect 7389 8386 7423 8420
rect 7457 8386 7491 8420
rect 7525 8386 7559 8420
rect 7593 8386 7627 8420
rect 7661 8386 7695 8420
rect 7729 8386 7763 8420
rect 7797 8386 7831 8420
rect 7865 8386 7899 8420
rect 7933 8386 7967 8420
rect 8001 8386 8035 8420
rect 8069 8386 8103 8420
rect 8137 8386 8171 8420
rect 8205 8386 8239 8420
rect 8273 8386 8307 8420
rect 8341 8419 8393 8420
rect 8427 8419 8462 8453
rect 8496 8419 8531 8453
rect 8565 8419 8600 8453
rect 8634 8419 8669 8453
rect 8703 8419 8738 8453
rect 8772 8419 8807 8453
rect 8841 8419 8876 8453
rect 8910 8419 8945 8453
rect 8979 8419 9014 8453
rect 9048 8419 9083 8453
rect 9117 8419 9152 8453
rect 9186 8419 9220 8453
rect 9254 8419 9288 8453
rect 9322 8419 9356 8453
rect 9390 8419 9424 8453
rect 9458 8419 9492 8453
rect 9526 8419 9560 8453
rect 9594 8419 9628 8453
rect 9662 8419 9696 8453
rect 9730 8419 9764 8453
rect 9798 8419 9832 8453
rect 9866 8419 9900 8453
rect 9934 8419 9968 8453
rect 10002 8419 10036 8453
rect 10070 8419 10104 8453
rect 10138 8419 10172 8453
rect 10206 8419 10240 8453
rect 10274 8419 10308 8453
rect 10342 8419 10376 8453
rect 10410 8419 10444 8453
rect 10478 8419 10512 8453
rect 10546 8419 10580 8453
rect 10614 8419 10648 8453
rect 10682 8419 10716 8453
rect 10750 8419 10784 8453
rect 10818 8419 10852 8453
rect 10886 8419 10920 8453
rect 10954 8419 10988 8453
rect 11022 8419 11056 8453
rect 11090 8419 11124 8453
rect 11158 8419 11192 8453
rect 11226 8419 11260 8453
rect 11294 8419 11328 8453
rect 11362 8419 11396 8453
rect 11430 8419 11464 8453
rect 11498 8419 11532 8453
rect 11566 8419 11600 8453
rect 11634 8419 11668 8453
rect 11702 8419 11736 8453
rect 11770 8419 11804 8453
rect 11838 8419 11872 8453
rect 11906 8419 11940 8453
rect 11974 8419 12008 8453
rect 12042 8419 12076 8453
rect 12110 8419 12144 8453
rect 12178 8419 12212 8453
rect 12246 8419 12280 8453
rect 12314 8419 12348 8453
rect 12382 8419 12416 8453
rect 12450 8419 12484 8453
rect 12518 8419 12552 8453
rect 12586 8419 12620 8453
rect 12654 8419 12688 8453
rect 12722 8419 12756 8453
rect 12790 8419 12824 8453
rect 12858 8419 12892 8453
rect 12926 8419 12960 8453
rect 12994 8419 13028 8453
rect 13062 8419 13096 8453
rect 13130 8419 13164 8453
rect 13198 8419 13232 8453
rect 13266 8419 13300 8453
rect 13334 8419 13368 8453
rect 13402 8419 13436 8453
rect 13470 8419 13504 8453
rect 13538 8419 13572 8453
rect 13606 8419 13640 8453
rect 13674 8419 13708 8453
rect 13742 8419 13776 8453
rect 13810 8419 13844 8453
rect 13878 8419 13912 8453
rect 13946 8419 13980 8453
rect 14026 8440 14048 8453
rect 14110 8440 14116 8453
rect 14014 8419 14048 8440
rect 14082 8419 14116 8440
rect 14150 8419 14184 8453
rect 14218 8435 14252 8453
rect 14286 8435 14320 8453
rect 14354 8435 14388 8453
rect 14422 8435 14456 8453
rect 14490 8435 14524 8453
rect 14219 8419 14252 8435
rect 14291 8419 14320 8435
rect 14363 8419 14388 8435
rect 14435 8419 14456 8435
rect 14507 8419 14524 8435
rect 14558 8419 14592 8453
rect 14648 8428 14660 8453
rect 14726 8428 14728 8453
rect 14626 8419 14660 8428
rect 14694 8419 14728 8428
rect 14762 8428 14770 8453
rect 14830 8428 14848 8453
rect 14898 8428 14926 8453
rect 14960 8433 15004 8462
rect 15038 8433 15102 8462
rect 14762 8419 14796 8428
rect 14830 8419 14864 8428
rect 14898 8419 14932 8428
rect 8341 8401 14185 8419
rect 14219 8401 14257 8419
rect 14291 8401 14329 8419
rect 14363 8401 14401 8419
rect 14435 8401 14473 8419
rect 14507 8401 14932 8419
rect 8341 8386 13992 8401
rect 2907 8383 13992 8386
rect 34 8324 136 8358
rect 34 8290 68 8324
rect 102 8290 136 8324
rect 235 8361 437 8371
rect 2445 8361 2647 8371
rect 235 8355 438 8361
rect 235 8321 248 8355
rect 285 8321 319 8355
rect 354 8321 387 8355
rect 426 8321 438 8355
rect 235 8315 438 8321
rect 2444 8355 2647 8361
rect 2444 8321 2456 8355
rect 2495 8321 2528 8355
rect 2563 8321 2597 8355
rect 2634 8321 2647 8355
rect 235 8305 437 8315
rect 34 8256 136 8290
rect 34 8222 68 8256
rect 102 8222 136 8256
rect 2444 8247 2647 8321
rect 2907 8350 8367 8383
rect 2907 8316 2933 8350
rect 2967 8316 3002 8350
rect 3036 8316 3071 8350
rect 3105 8316 3139 8350
rect 3173 8316 3207 8350
rect 3241 8316 3275 8350
rect 3309 8316 3343 8350
rect 3377 8316 3411 8350
rect 3445 8316 3479 8350
rect 3513 8316 3547 8350
rect 3581 8316 3615 8350
rect 3649 8316 3683 8350
rect 3717 8316 3751 8350
rect 3785 8316 3819 8350
rect 3853 8316 3887 8350
rect 3921 8316 3955 8350
rect 3989 8316 4023 8350
rect 4057 8316 4091 8350
rect 4125 8316 4159 8350
rect 4193 8316 4227 8350
rect 4261 8316 4295 8350
rect 4329 8316 4363 8350
rect 4397 8316 4431 8350
rect 4465 8316 4499 8350
rect 4533 8316 4567 8350
rect 4601 8316 4635 8350
rect 4669 8316 4703 8350
rect 4737 8316 4771 8350
rect 4805 8316 4839 8350
rect 4873 8316 4907 8350
rect 4941 8316 4975 8350
rect 5009 8316 5043 8350
rect 5077 8316 5111 8350
rect 5145 8316 5179 8350
rect 5213 8316 5247 8350
rect 5281 8316 5315 8350
rect 5349 8316 5383 8350
rect 5417 8316 5451 8350
rect 5485 8316 5519 8350
rect 5553 8316 5587 8350
rect 5621 8316 5655 8350
rect 5689 8316 5723 8350
rect 5757 8316 5791 8350
rect 5825 8316 5859 8350
rect 5893 8316 5927 8350
rect 5961 8316 5995 8350
rect 6029 8316 6063 8350
rect 6097 8316 6131 8350
rect 6165 8316 6199 8350
rect 6233 8316 6267 8350
rect 6301 8316 6335 8350
rect 6369 8316 6403 8350
rect 6437 8316 6471 8350
rect 6505 8316 6539 8350
rect 6573 8316 6607 8350
rect 6641 8316 6675 8350
rect 6709 8316 6743 8350
rect 6777 8316 6811 8350
rect 6845 8316 6879 8350
rect 6913 8316 6947 8350
rect 6981 8316 7015 8350
rect 7049 8316 7083 8350
rect 7117 8316 7151 8350
rect 7185 8316 7219 8350
rect 7253 8316 7287 8350
rect 7321 8316 7355 8350
rect 7389 8316 7423 8350
rect 7457 8316 7491 8350
rect 7525 8316 7559 8350
rect 7593 8316 7627 8350
rect 7661 8316 7695 8350
rect 7729 8316 7763 8350
rect 7797 8316 7831 8350
rect 7865 8316 7899 8350
rect 7933 8316 7967 8350
rect 8001 8316 8035 8350
rect 8069 8316 8103 8350
rect 8137 8316 8171 8350
rect 8205 8316 8239 8350
rect 8273 8316 8307 8350
rect 8341 8316 8367 8350
rect 2907 8280 8367 8316
rect 34 8192 136 8222
rect 2907 8246 2933 8280
rect 2967 8246 3002 8280
rect 3036 8246 3071 8280
rect 3105 8246 3139 8280
rect 3173 8246 3207 8280
rect 3241 8246 3275 8280
rect 3309 8246 3343 8280
rect 3377 8246 3411 8280
rect 3445 8246 3479 8280
rect 3513 8246 3547 8280
rect 3581 8246 3615 8280
rect 3649 8246 3683 8280
rect 3717 8246 3751 8280
rect 3785 8246 3819 8280
rect 3853 8246 3887 8280
rect 3921 8246 3955 8280
rect 3989 8246 4023 8280
rect 4057 8246 4091 8280
rect 4125 8246 4159 8280
rect 4193 8246 4227 8280
rect 4261 8246 4295 8280
rect 4329 8246 4363 8280
rect 4397 8246 4431 8280
rect 4465 8246 4499 8280
rect 4533 8246 4567 8280
rect 4601 8246 4635 8280
rect 4669 8246 4703 8280
rect 4737 8246 4771 8280
rect 4805 8246 4839 8280
rect 4873 8246 4907 8280
rect 4941 8246 4975 8280
rect 5009 8246 5043 8280
rect 5077 8246 5111 8280
rect 5145 8246 5179 8280
rect 5213 8246 5247 8280
rect 5281 8246 5315 8280
rect 5349 8246 5383 8280
rect 5417 8246 5451 8280
rect 5485 8246 5519 8280
rect 5553 8246 5587 8280
rect 5621 8246 5655 8280
rect 5689 8246 5723 8280
rect 5757 8246 5791 8280
rect 5825 8246 5859 8280
rect 5893 8246 5927 8280
rect 5961 8246 5995 8280
rect 6029 8246 6063 8280
rect 6097 8246 6131 8280
rect 6165 8246 6199 8280
rect 6233 8246 6267 8280
rect 6301 8246 6335 8280
rect 6369 8246 6403 8280
rect 6437 8246 6471 8280
rect 6505 8246 6539 8280
rect 6573 8246 6607 8280
rect 6641 8246 6675 8280
rect 6709 8246 6743 8280
rect 6777 8246 6811 8280
rect 6845 8246 6879 8280
rect 6913 8246 6947 8280
rect 6981 8246 7015 8280
rect 7049 8246 7083 8280
rect 7117 8246 7151 8280
rect 7185 8246 7219 8280
rect 7253 8246 7287 8280
rect 7321 8246 7355 8280
rect 7389 8246 7423 8280
rect 7457 8246 7491 8280
rect 7525 8246 7559 8280
rect 7593 8246 7627 8280
rect 7661 8246 7695 8280
rect 7729 8246 7763 8280
rect 7797 8246 7831 8280
rect 7865 8246 7899 8280
rect 7933 8246 7967 8280
rect 8001 8246 8035 8280
rect 8069 8246 8103 8280
rect 8137 8246 8171 8280
rect 8205 8246 8239 8280
rect 8273 8246 8307 8280
rect 8341 8246 8367 8280
rect 13506 8367 13992 8383
rect 14026 8367 14076 8401
rect 14110 8399 14932 8401
rect 14966 8399 15000 8433
rect 15038 8428 15068 8433
rect 15034 8399 15068 8428
rect 14110 8388 15102 8399
rect 14110 8367 14614 8388
rect 13506 8358 14614 8367
rect 13506 8357 14185 8358
rect 14219 8357 14257 8358
rect 14291 8357 14329 8358
rect 14363 8357 14401 8358
rect 14435 8357 14473 8358
rect 14507 8357 14614 8358
rect 14648 8357 14692 8388
rect 14726 8357 14770 8388
rect 14804 8357 14848 8388
rect 14882 8357 14926 8388
rect 14960 8361 15004 8388
rect 15038 8361 15102 8388
rect 13506 8323 13532 8357
rect 13566 8323 13603 8357
rect 13637 8323 13674 8357
rect 13708 8323 13744 8357
rect 13778 8323 13814 8357
rect 13848 8323 13884 8357
rect 13918 8323 13954 8357
rect 13988 8323 14024 8357
rect 14058 8323 14094 8357
rect 14128 8323 14164 8357
rect 14219 8324 14234 8357
rect 14291 8324 14304 8357
rect 14363 8324 14374 8357
rect 14435 8324 14444 8357
rect 14507 8324 14514 8357
rect 14198 8323 14234 8324
rect 14268 8323 14304 8324
rect 14338 8323 14374 8324
rect 14408 8323 14444 8324
rect 14478 8323 14514 8324
rect 14548 8323 14584 8357
rect 14648 8354 14654 8357
rect 14618 8323 14654 8354
rect 14688 8354 14692 8357
rect 14758 8354 14770 8357
rect 14828 8354 14848 8357
rect 14898 8354 14926 8357
rect 14688 8323 14724 8354
rect 14758 8323 14794 8354
rect 14828 8323 14864 8354
rect 14898 8327 14932 8354
rect 14966 8327 15000 8361
rect 15038 8354 15068 8361
rect 15034 8327 15068 8354
rect 14898 8323 15102 8327
rect 13506 8314 15102 8323
rect 13506 8283 14614 8314
rect 14648 8283 14692 8314
rect 14726 8283 14770 8314
rect 14804 8283 14848 8314
rect 14882 8283 14926 8314
rect 14960 8289 15004 8314
rect 15038 8289 15102 8314
rect 2907 8210 8367 8246
rect 2907 8192 2933 8210
rect 42 8176 2933 8192
rect 2967 8176 3002 8210
rect 3036 8176 3071 8210
rect 3105 8176 3139 8210
rect 3173 8176 3207 8210
rect 3241 8176 3275 8210
rect 3309 8176 3343 8210
rect 3377 8176 3411 8210
rect 3445 8176 3479 8210
rect 3513 8176 3547 8210
rect 3581 8176 3615 8210
rect 3649 8176 3683 8210
rect 3717 8176 3751 8210
rect 3785 8176 3819 8210
rect 3853 8176 3887 8210
rect 3921 8176 3955 8210
rect 3989 8176 4023 8210
rect 4057 8176 4091 8210
rect 4125 8176 4159 8210
rect 4193 8176 4227 8210
rect 4261 8176 4295 8210
rect 4329 8176 4363 8210
rect 4397 8176 4431 8210
rect 4465 8176 4499 8210
rect 4533 8176 4567 8210
rect 4601 8176 4635 8210
rect 4669 8176 4703 8210
rect 4737 8176 4771 8210
rect 4805 8176 4839 8210
rect 4873 8176 4907 8210
rect 4941 8176 4975 8210
rect 5009 8176 5043 8210
rect 5077 8176 5111 8210
rect 5145 8176 5179 8210
rect 5213 8176 5247 8210
rect 5281 8176 5315 8210
rect 5349 8176 5383 8210
rect 5417 8176 5451 8210
rect 5485 8176 5519 8210
rect 5553 8176 5587 8210
rect 5621 8176 5655 8210
rect 5689 8176 5723 8210
rect 5757 8176 5791 8210
rect 5825 8176 5859 8210
rect 5893 8176 5927 8210
rect 5961 8176 5995 8210
rect 6029 8176 6063 8210
rect 6097 8176 6131 8210
rect 6165 8176 6199 8210
rect 6233 8176 6267 8210
rect 6301 8176 6335 8210
rect 6369 8176 6403 8210
rect 6437 8176 6471 8210
rect 6505 8176 6539 8210
rect 6573 8176 6607 8210
rect 6641 8176 6675 8210
rect 6709 8176 6743 8210
rect 6777 8176 6811 8210
rect 6845 8176 6879 8210
rect 6913 8176 6947 8210
rect 6981 8176 7015 8210
rect 7049 8176 7083 8210
rect 7117 8176 7151 8210
rect 7185 8176 7219 8210
rect 7253 8176 7287 8210
rect 7321 8176 7355 8210
rect 7389 8176 7423 8210
rect 7457 8176 7491 8210
rect 7525 8176 7559 8210
rect 7593 8176 7627 8210
rect 7661 8176 7695 8210
rect 7729 8176 7763 8210
rect 7797 8176 7831 8210
rect 7865 8176 7899 8210
rect 7933 8176 7967 8210
rect 8001 8176 8035 8210
rect 8069 8176 8103 8210
rect 8137 8176 8171 8210
rect 8205 8176 8239 8210
rect 8273 8176 8307 8210
rect 8341 8176 8367 8210
rect 42 8157 8367 8176
rect 42 8123 68 8157
rect 102 8123 138 8157
rect 172 8123 208 8157
rect 242 8123 278 8157
rect 312 8123 348 8157
rect 382 8123 418 8157
rect 452 8123 488 8157
rect 522 8123 558 8157
rect 592 8123 628 8157
rect 662 8123 698 8157
rect 732 8123 768 8157
rect 802 8123 838 8157
rect 872 8123 908 8157
rect 942 8123 978 8157
rect 1012 8123 1048 8157
rect 1082 8123 1118 8157
rect 1152 8123 1188 8157
rect 1222 8123 1258 8157
rect 1292 8123 1328 8157
rect 1362 8123 1398 8157
rect 1432 8123 1467 8157
rect 1501 8123 1536 8157
rect 1570 8123 1605 8157
rect 1639 8123 1674 8157
rect 1708 8123 1743 8157
rect 1777 8123 1812 8157
rect 1846 8123 1881 8157
rect 1915 8123 1950 8157
rect 1984 8123 2019 8157
rect 2053 8123 2088 8157
rect 2122 8123 2157 8157
rect 2191 8123 2226 8157
rect 2260 8123 2295 8157
rect 2329 8123 2364 8157
rect 2398 8123 2433 8157
rect 2467 8123 2502 8157
rect 2536 8123 2571 8157
rect 2605 8123 2640 8157
rect 2674 8123 2709 8157
rect 2743 8123 2778 8157
rect 2812 8123 2847 8157
rect 2881 8140 8367 8157
rect 2881 8123 2933 8140
rect 42 8106 2933 8123
rect 2967 8106 3002 8140
rect 3036 8106 3071 8140
rect 3105 8106 3139 8140
rect 3173 8106 3207 8140
rect 3241 8106 3275 8140
rect 3309 8106 3343 8140
rect 3377 8106 3411 8140
rect 3445 8106 3479 8140
rect 3513 8106 3547 8140
rect 3581 8106 3615 8140
rect 3649 8106 3683 8140
rect 3717 8106 3751 8140
rect 3785 8106 3819 8140
rect 3853 8106 3887 8140
rect 3921 8106 3955 8140
rect 3989 8106 4023 8140
rect 4057 8106 4091 8140
rect 4125 8106 4159 8140
rect 4193 8106 4227 8140
rect 4261 8106 4295 8140
rect 4329 8106 4363 8140
rect 4397 8106 4431 8140
rect 4465 8106 4499 8140
rect 4533 8106 4567 8140
rect 4601 8106 4635 8140
rect 4669 8106 4703 8140
rect 4737 8106 4771 8140
rect 4805 8106 4839 8140
rect 4873 8106 4907 8140
rect 4941 8106 4975 8140
rect 5009 8106 5043 8140
rect 5077 8106 5111 8140
rect 5145 8106 5179 8140
rect 5213 8106 5247 8140
rect 5281 8106 5315 8140
rect 5349 8106 5383 8140
rect 5417 8106 5451 8140
rect 5485 8106 5519 8140
rect 5553 8106 5587 8140
rect 5621 8106 5655 8140
rect 5689 8106 5723 8140
rect 5757 8106 5791 8140
rect 5825 8106 5859 8140
rect 5893 8106 5927 8140
rect 5961 8106 5995 8140
rect 6029 8106 6063 8140
rect 6097 8106 6131 8140
rect 6165 8106 6199 8140
rect 6233 8106 6267 8140
rect 6301 8106 6335 8140
rect 6369 8106 6403 8140
rect 6437 8106 6471 8140
rect 6505 8106 6539 8140
rect 6573 8106 6607 8140
rect 6641 8106 6675 8140
rect 6709 8106 6743 8140
rect 6777 8106 6811 8140
rect 6845 8106 6879 8140
rect 6913 8106 6947 8140
rect 6981 8106 7015 8140
rect 7049 8106 7083 8140
rect 7117 8106 7151 8140
rect 7185 8106 7219 8140
rect 7253 8106 7287 8140
rect 7321 8106 7355 8140
rect 7389 8106 7423 8140
rect 7457 8106 7491 8140
rect 7525 8106 7559 8140
rect 7593 8106 7627 8140
rect 7661 8106 7695 8140
rect 7729 8106 7763 8140
rect 7797 8106 7831 8140
rect 7865 8106 7899 8140
rect 7933 8106 7967 8140
rect 8001 8106 8035 8140
rect 8069 8106 8103 8140
rect 8137 8106 8171 8140
rect 8205 8106 8239 8140
rect 8273 8106 8307 8140
rect 8341 8106 8367 8140
rect 42 8082 8367 8106
rect 42 8048 68 8082
rect 102 8048 138 8082
rect 172 8048 208 8082
rect 242 8048 278 8082
rect 312 8048 348 8082
rect 382 8048 418 8082
rect 452 8048 488 8082
rect 522 8048 558 8082
rect 592 8048 628 8082
rect 662 8048 698 8082
rect 732 8048 768 8082
rect 802 8048 838 8082
rect 872 8048 908 8082
rect 942 8048 978 8082
rect 1012 8048 1048 8082
rect 1082 8048 1118 8082
rect 1152 8048 1188 8082
rect 1222 8048 1258 8082
rect 1292 8048 1328 8082
rect 1362 8048 1398 8082
rect 1432 8048 1467 8082
rect 1501 8048 1536 8082
rect 1570 8048 1605 8082
rect 1639 8048 1674 8082
rect 1708 8048 1743 8082
rect 1777 8048 1812 8082
rect 1846 8048 1881 8082
rect 1915 8048 1950 8082
rect 1984 8048 2019 8082
rect 2053 8048 2088 8082
rect 2122 8048 2157 8082
rect 2191 8048 2226 8082
rect 2260 8048 2295 8082
rect 2329 8048 2364 8082
rect 2398 8048 2433 8082
rect 2467 8048 2502 8082
rect 2536 8048 2571 8082
rect 2605 8048 2640 8082
rect 2674 8048 2709 8082
rect 2743 8048 2778 8082
rect 2812 8048 2847 8082
rect 2881 8070 8367 8082
rect 2881 8048 2933 8070
rect 42 8036 2933 8048
rect 2967 8036 3002 8070
rect 3036 8036 3071 8070
rect 3105 8036 3139 8070
rect 3173 8036 3207 8070
rect 3241 8036 3275 8070
rect 3309 8036 3343 8070
rect 3377 8036 3411 8070
rect 3445 8036 3479 8070
rect 3513 8036 3547 8070
rect 3581 8036 3615 8070
rect 3649 8036 3683 8070
rect 3717 8036 3751 8070
rect 3785 8036 3819 8070
rect 3853 8036 3887 8070
rect 3921 8036 3955 8070
rect 3989 8036 4023 8070
rect 4057 8036 4091 8070
rect 4125 8036 4159 8070
rect 4193 8036 4227 8070
rect 4261 8036 4295 8070
rect 4329 8036 4363 8070
rect 4397 8036 4431 8070
rect 4465 8036 4499 8070
rect 4533 8036 4567 8070
rect 4601 8036 4635 8070
rect 4669 8036 4703 8070
rect 4737 8036 4771 8070
rect 4805 8036 4839 8070
rect 4873 8036 4907 8070
rect 4941 8036 4975 8070
rect 5009 8036 5043 8070
rect 5077 8036 5111 8070
rect 5145 8036 5179 8070
rect 5213 8036 5247 8070
rect 5281 8036 5315 8070
rect 5349 8036 5383 8070
rect 5417 8036 5451 8070
rect 5485 8036 5519 8070
rect 5553 8036 5587 8070
rect 5621 8036 5655 8070
rect 5689 8036 5723 8070
rect 5757 8036 5791 8070
rect 5825 8036 5859 8070
rect 5893 8036 5927 8070
rect 5961 8036 5995 8070
rect 6029 8036 6063 8070
rect 6097 8036 6131 8070
rect 6165 8036 6199 8070
rect 6233 8036 6267 8070
rect 6301 8036 6335 8070
rect 6369 8036 6403 8070
rect 6437 8036 6471 8070
rect 6505 8036 6539 8070
rect 6573 8036 6607 8070
rect 6641 8036 6675 8070
rect 6709 8036 6743 8070
rect 6777 8036 6811 8070
rect 6845 8036 6879 8070
rect 6913 8036 6947 8070
rect 6981 8036 7015 8070
rect 7049 8036 7083 8070
rect 7117 8036 7151 8070
rect 7185 8036 7219 8070
rect 7253 8036 7287 8070
rect 7321 8036 7355 8070
rect 7389 8036 7423 8070
rect 7457 8036 7491 8070
rect 7525 8036 7559 8070
rect 7593 8036 7627 8070
rect 7661 8036 7695 8070
rect 7729 8036 7763 8070
rect 7797 8036 7831 8070
rect 7865 8036 7899 8070
rect 7933 8036 7967 8070
rect 8001 8036 8035 8070
rect 8069 8036 8103 8070
rect 8137 8036 8171 8070
rect 8205 8036 8239 8070
rect 8273 8036 8307 8070
rect 8341 8036 8367 8070
rect 42 8007 8367 8036
rect 42 7973 68 8007
rect 102 7973 138 8007
rect 172 7973 208 8007
rect 242 7973 278 8007
rect 312 7973 348 8007
rect 382 7973 418 8007
rect 452 7973 488 8007
rect 522 7973 558 8007
rect 592 7973 628 8007
rect 662 7973 698 8007
rect 732 7973 768 8007
rect 802 7973 838 8007
rect 872 7973 908 8007
rect 942 7973 978 8007
rect 1012 7973 1048 8007
rect 1082 7973 1118 8007
rect 1152 7973 1188 8007
rect 1222 7973 1258 8007
rect 1292 7973 1328 8007
rect 1362 7973 1398 8007
rect 1432 7973 1467 8007
rect 1501 7973 1536 8007
rect 1570 7973 1605 8007
rect 1639 7973 1674 8007
rect 1708 7973 1743 8007
rect 1777 7973 1812 8007
rect 1846 7973 1881 8007
rect 1915 7973 1950 8007
rect 1984 7973 2019 8007
rect 2053 7973 2088 8007
rect 2122 7973 2157 8007
rect 2191 7973 2226 8007
rect 2260 7973 2295 8007
rect 2329 7973 2364 8007
rect 2398 7973 2433 8007
rect 2467 7973 2502 8007
rect 2536 7973 2571 8007
rect 2605 7973 2640 8007
rect 2674 7973 2709 8007
rect 2743 7973 2778 8007
rect 2812 7973 2847 8007
rect 2881 8000 8367 8007
rect 2881 7973 2933 8000
rect 42 7966 2933 7973
rect 2967 7966 3002 8000
rect 3036 7966 3071 8000
rect 3105 7966 3139 8000
rect 3173 7966 3207 8000
rect 3241 7966 3275 8000
rect 3309 7966 3343 8000
rect 3377 7966 3411 8000
rect 3445 7966 3479 8000
rect 3513 7966 3547 8000
rect 3581 7966 3615 8000
rect 3649 7966 3683 8000
rect 3717 7966 3751 8000
rect 3785 7966 3819 8000
rect 3853 7966 3887 8000
rect 3921 7966 3955 8000
rect 3989 7966 4023 8000
rect 4057 7966 4091 8000
rect 4125 7966 4159 8000
rect 4193 7966 4227 8000
rect 4261 7966 4295 8000
rect 4329 7966 4363 8000
rect 4397 7966 4431 8000
rect 4465 7966 4499 8000
rect 4533 7966 4567 8000
rect 4601 7966 4635 8000
rect 4669 7966 4703 8000
rect 4737 7966 4771 8000
rect 4805 7966 4839 8000
rect 4873 7966 4907 8000
rect 4941 7966 4975 8000
rect 5009 7966 5043 8000
rect 5077 7966 5111 8000
rect 5145 7966 5179 8000
rect 5213 7966 5247 8000
rect 5281 7966 5315 8000
rect 5349 7966 5383 8000
rect 5417 7966 5451 8000
rect 5485 7966 5519 8000
rect 5553 7966 5587 8000
rect 5621 7966 5655 8000
rect 5689 7966 5723 8000
rect 5757 7966 5791 8000
rect 5825 7966 5859 8000
rect 5893 7966 5927 8000
rect 5961 7966 5995 8000
rect 6029 7966 6063 8000
rect 6097 7966 6131 8000
rect 6165 7966 6199 8000
rect 6233 7966 6267 8000
rect 6301 7966 6335 8000
rect 6369 7966 6403 8000
rect 6437 7966 6471 8000
rect 6505 7966 6539 8000
rect 6573 7966 6607 8000
rect 6641 7966 6675 8000
rect 6709 7966 6743 8000
rect 6777 7966 6811 8000
rect 6845 7966 6879 8000
rect 6913 7966 6947 8000
rect 6981 7966 7015 8000
rect 7049 7966 7083 8000
rect 7117 7966 7151 8000
rect 7185 7966 7219 8000
rect 7253 7966 7287 8000
rect 7321 7966 7355 8000
rect 7389 7966 7423 8000
rect 7457 7966 7491 8000
rect 7525 7966 7559 8000
rect 7593 7966 7627 8000
rect 7661 7966 7695 8000
rect 7729 7966 7763 8000
rect 7797 7966 7831 8000
rect 7865 7966 7899 8000
rect 7933 7966 7967 8000
rect 8001 7966 8035 8000
rect 8069 7966 8103 8000
rect 8137 7966 8171 8000
rect 8205 7966 8239 8000
rect 8273 7966 8307 8000
rect 8341 7966 8367 8000
rect 42 7932 8367 7966
rect 42 7898 68 7932
rect 102 7898 138 7932
rect 172 7898 208 7932
rect 242 7898 278 7932
rect 312 7898 348 7932
rect 382 7898 418 7932
rect 452 7898 488 7932
rect 522 7898 558 7932
rect 592 7898 628 7932
rect 662 7898 698 7932
rect 732 7898 768 7932
rect 802 7898 838 7932
rect 872 7898 908 7932
rect 942 7898 978 7932
rect 1012 7898 1048 7932
rect 1082 7898 1118 7932
rect 1152 7898 1188 7932
rect 1222 7898 1258 7932
rect 1292 7898 1328 7932
rect 1362 7898 1398 7932
rect 1432 7898 1467 7932
rect 1501 7898 1536 7932
rect 1570 7898 1605 7932
rect 1639 7898 1674 7932
rect 1708 7898 1743 7932
rect 1777 7898 1812 7932
rect 1846 7898 1881 7932
rect 1915 7898 1950 7932
rect 1984 7898 2019 7932
rect 2053 7898 2088 7932
rect 2122 7898 2157 7932
rect 2191 7898 2226 7932
rect 2260 7898 2295 7932
rect 2329 7898 2364 7932
rect 2398 7898 2433 7932
rect 2467 7898 2502 7932
rect 2536 7898 2571 7932
rect 2605 7898 2640 7932
rect 2674 7898 2709 7932
rect 2743 7898 2778 7932
rect 2812 7898 2847 7932
rect 2881 7930 8367 7932
rect 2881 7898 2933 7930
rect 42 7896 2933 7898
rect 2967 7896 3002 7930
rect 3036 7896 3071 7930
rect 3105 7896 3139 7930
rect 3173 7896 3207 7930
rect 3241 7896 3275 7930
rect 3309 7896 3343 7930
rect 3377 7896 3411 7930
rect 3445 7896 3479 7930
rect 3513 7896 3547 7930
rect 3581 7896 3615 7930
rect 3649 7896 3683 7930
rect 3717 7896 3751 7930
rect 3785 7896 3819 7930
rect 3853 7896 3887 7930
rect 3921 7896 3955 7930
rect 3989 7896 4023 7930
rect 4057 7896 4091 7930
rect 4125 7896 4159 7930
rect 4193 7896 4227 7930
rect 4261 7896 4295 7930
rect 4329 7896 4363 7930
rect 4397 7896 4431 7930
rect 4465 7896 4499 7930
rect 4533 7896 4567 7930
rect 4601 7896 4635 7930
rect 4669 7896 4703 7930
rect 4737 7896 4771 7930
rect 4805 7896 4839 7930
rect 4873 7896 4907 7930
rect 4941 7896 4975 7930
rect 5009 7896 5043 7930
rect 5077 7896 5111 7930
rect 5145 7896 5179 7930
rect 5213 7896 5247 7930
rect 5281 7896 5315 7930
rect 5349 7896 5383 7930
rect 5417 7896 5451 7930
rect 5485 7896 5519 7930
rect 5553 7896 5587 7930
rect 5621 7896 5655 7930
rect 5689 7896 5723 7930
rect 5757 7896 5791 7930
rect 5825 7896 5859 7930
rect 5893 7896 5927 7930
rect 5961 7896 5995 7930
rect 6029 7896 6063 7930
rect 6097 7896 6131 7930
rect 6165 7896 6199 7930
rect 6233 7896 6267 7930
rect 6301 7896 6335 7930
rect 6369 7896 6403 7930
rect 6437 7896 6471 7930
rect 6505 7896 6539 7930
rect 6573 7896 6607 7930
rect 6641 7896 6675 7930
rect 6709 7896 6743 7930
rect 6777 7896 6811 7930
rect 6845 7896 6879 7930
rect 6913 7896 6947 7930
rect 6981 7896 7015 7930
rect 7049 7896 7083 7930
rect 7117 7896 7151 7930
rect 7185 7896 7219 7930
rect 7253 7896 7287 7930
rect 7321 7896 7355 7930
rect 7389 7896 7423 7930
rect 7457 7896 7491 7930
rect 7525 7896 7559 7930
rect 7593 7896 7627 7930
rect 7661 7896 7695 7930
rect 7729 7896 7763 7930
rect 7797 7896 7831 7930
rect 7865 7896 7899 7930
rect 7933 7896 7967 7930
rect 8001 7896 8035 7930
rect 8069 7896 8103 7930
rect 8137 7896 8171 7930
rect 8205 7896 8239 7930
rect 8273 7896 8307 7930
rect 8341 7896 8367 7930
rect 8494 8254 8628 8255
rect 8494 7932 8509 8254
rect 8615 7932 8628 8254
rect 8494 7917 8628 7932
rect 9596 8247 9714 8255
rect 9630 8239 9678 8247
rect 9712 8239 9714 8247
rect 9596 8144 9612 8213
rect 9596 8041 9612 8110
rect 9596 7933 9612 8007
rect 9596 7917 9714 7933
rect 10314 8247 10430 8255
rect 10348 8239 10396 8247
rect 10416 8144 10430 8213
rect 10416 8041 10430 8110
rect 10416 7933 10430 8007
rect 10314 7917 10430 7933
rect 10800 8254 10934 8255
rect 10800 8220 10804 8254
rect 10838 8239 10898 8254
rect 10932 8220 10934 8254
rect 10800 8179 10816 8220
rect 10918 8179 10934 8220
rect 10800 8145 10804 8179
rect 10932 8145 10934 8179
rect 10800 8104 10816 8145
rect 10918 8104 10934 8145
rect 10800 8070 10804 8104
rect 10932 8070 10934 8104
rect 10800 8028 10816 8070
rect 10918 8028 10934 8070
rect 10800 7994 10804 8028
rect 10932 7994 10934 8028
rect 10800 7952 10816 7994
rect 10918 7952 10934 7994
rect 10800 7918 10804 7952
rect 10838 7918 10898 7933
rect 10932 7918 10934 7952
rect 10800 7917 10934 7918
rect 13506 8249 13532 8283
rect 13566 8249 13603 8283
rect 13637 8249 13674 8283
rect 13708 8249 13744 8283
rect 13778 8249 13814 8283
rect 13848 8249 13884 8283
rect 13918 8249 13954 8283
rect 13988 8249 14024 8283
rect 14058 8249 14094 8283
rect 14128 8249 14164 8283
rect 14198 8280 14234 8283
rect 14268 8280 14304 8283
rect 14338 8280 14374 8283
rect 14408 8280 14444 8283
rect 14478 8280 14514 8283
rect 14219 8249 14234 8280
rect 14291 8249 14304 8280
rect 14363 8249 14374 8280
rect 14435 8249 14444 8280
rect 14507 8249 14514 8280
rect 14548 8249 14584 8283
rect 14648 8280 14654 8283
rect 14618 8249 14654 8280
rect 14688 8280 14692 8283
rect 14758 8280 14770 8283
rect 14828 8280 14848 8283
rect 14898 8280 14926 8283
rect 14688 8249 14724 8280
rect 14758 8249 14794 8280
rect 14828 8249 14864 8280
rect 14898 8255 14932 8280
rect 14966 8255 15000 8289
rect 15038 8280 15068 8289
rect 15034 8255 15068 8280
rect 14898 8249 15102 8255
rect 13506 8246 14185 8249
rect 14219 8246 14257 8249
rect 14291 8246 14329 8249
rect 14363 8246 14401 8249
rect 14435 8246 14473 8249
rect 14507 8246 15102 8249
rect 13506 8240 15102 8246
rect 13506 8209 14614 8240
rect 14648 8209 14692 8240
rect 14726 8209 14770 8240
rect 14804 8209 14848 8240
rect 14882 8209 14926 8240
rect 14960 8217 15004 8240
rect 15038 8217 15102 8240
rect 13506 8175 13532 8209
rect 13566 8175 13603 8209
rect 13637 8175 13674 8209
rect 13708 8175 13744 8209
rect 13778 8175 13814 8209
rect 13848 8175 13884 8209
rect 13918 8175 13954 8209
rect 13988 8175 14024 8209
rect 14058 8175 14094 8209
rect 14128 8175 14164 8209
rect 14198 8202 14234 8209
rect 14268 8202 14304 8209
rect 14338 8202 14374 8209
rect 14408 8202 14444 8209
rect 14478 8202 14514 8209
rect 14219 8175 14234 8202
rect 14291 8175 14304 8202
rect 14363 8175 14374 8202
rect 14435 8175 14444 8202
rect 14507 8175 14514 8202
rect 14548 8175 14584 8209
rect 14648 8206 14654 8209
rect 14618 8175 14654 8206
rect 14688 8206 14692 8209
rect 14758 8206 14770 8209
rect 14828 8206 14848 8209
rect 14898 8206 14926 8209
rect 14688 8175 14724 8206
rect 14758 8175 14794 8206
rect 14828 8175 14864 8206
rect 14898 8183 14932 8206
rect 14966 8183 15000 8217
rect 15038 8206 15068 8217
rect 15034 8183 15068 8206
rect 14898 8175 15102 8183
rect 13506 8168 14185 8175
rect 14219 8168 14257 8175
rect 14291 8168 14329 8175
rect 14363 8168 14401 8175
rect 14435 8168 14473 8175
rect 14507 8168 15102 8175
rect 13506 8166 15102 8168
rect 13506 8135 14614 8166
rect 14648 8135 14692 8166
rect 14726 8135 14770 8166
rect 14804 8135 14848 8166
rect 14882 8135 14926 8166
rect 14960 8145 15004 8166
rect 15038 8145 15102 8166
rect 13506 8101 13532 8135
rect 13566 8101 13603 8135
rect 13637 8101 13674 8135
rect 13708 8101 13744 8135
rect 13778 8101 13814 8135
rect 13848 8101 13884 8135
rect 13918 8101 13954 8135
rect 13988 8101 14024 8135
rect 14058 8101 14094 8135
rect 14128 8101 14164 8135
rect 14198 8101 14234 8135
rect 14268 8101 14304 8135
rect 14338 8101 14374 8135
rect 14408 8115 14444 8135
rect 14478 8115 14514 8135
rect 14408 8101 14431 8115
rect 14478 8101 14511 8115
rect 14548 8101 14584 8135
rect 14648 8132 14654 8135
rect 14618 8101 14654 8132
rect 14688 8132 14692 8135
rect 14758 8132 14770 8135
rect 14828 8132 14848 8135
rect 14898 8132 14926 8135
rect 14688 8101 14724 8132
rect 14758 8101 14794 8132
rect 14828 8101 14864 8132
rect 14898 8111 14932 8132
rect 14966 8111 15000 8145
rect 15038 8132 15068 8145
rect 15034 8111 15068 8132
rect 14898 8101 15102 8111
rect 13506 8081 14431 8101
rect 14465 8081 14511 8101
rect 14545 8092 15102 8101
rect 14545 8081 14614 8092
rect 13506 8061 14614 8081
rect 14648 8061 14692 8092
rect 14726 8061 14770 8092
rect 14804 8061 14848 8092
rect 14882 8061 14926 8092
rect 14960 8073 15004 8092
rect 15038 8073 15102 8092
rect 13506 8027 13532 8061
rect 13566 8027 13603 8061
rect 13637 8027 13674 8061
rect 13708 8027 13744 8061
rect 13778 8027 13814 8061
rect 13848 8027 13884 8061
rect 13918 8027 13954 8061
rect 13988 8027 14024 8061
rect 14058 8027 14094 8061
rect 14128 8027 14164 8061
rect 14198 8027 14234 8061
rect 14268 8027 14304 8061
rect 14338 8027 14374 8061
rect 14408 8033 14444 8061
rect 14478 8033 14514 8061
rect 14408 8027 14431 8033
rect 14478 8027 14511 8033
rect 14548 8027 14584 8061
rect 14648 8058 14654 8061
rect 14618 8027 14654 8058
rect 14688 8058 14692 8061
rect 14758 8058 14770 8061
rect 14828 8058 14848 8061
rect 14898 8058 14926 8061
rect 14688 8027 14724 8058
rect 14758 8027 14794 8058
rect 14828 8027 14864 8058
rect 14898 8039 14932 8058
rect 14966 8039 15000 8073
rect 15038 8058 15068 8073
rect 15034 8039 15068 8058
rect 14898 8027 15102 8039
rect 13506 7999 14431 8027
rect 14465 7999 14511 8027
rect 14545 8018 15102 8027
rect 14545 7999 14614 8018
rect 13506 7987 14614 7999
rect 14648 7987 14692 8018
rect 14726 7987 14770 8018
rect 14804 7987 14848 8018
rect 14882 7987 14926 8018
rect 14960 8001 15004 8018
rect 15038 8001 15102 8018
rect 13506 7953 13532 7987
rect 13566 7953 13603 7987
rect 13637 7953 13674 7987
rect 13708 7953 13744 7987
rect 13778 7953 13814 7987
rect 13848 7953 13884 7987
rect 13918 7953 13954 7987
rect 13988 7953 14024 7987
rect 14058 7953 14094 7987
rect 14128 7953 14164 7987
rect 14198 7953 14234 7987
rect 14268 7953 14304 7987
rect 14338 7953 14374 7987
rect 14408 7953 14444 7987
rect 14478 7953 14514 7987
rect 14548 7953 14584 7987
rect 14648 7984 14654 7987
rect 14618 7953 14654 7984
rect 14688 7984 14692 7987
rect 14758 7984 14770 7987
rect 14828 7984 14848 7987
rect 14898 7984 14926 7987
rect 14688 7953 14724 7984
rect 14758 7953 14794 7984
rect 14828 7953 14864 7984
rect 14898 7967 14932 7984
rect 14966 7967 15000 8001
rect 15038 7984 15068 8001
rect 15034 7967 15068 7984
rect 14898 7953 15102 7967
rect 13506 7950 15102 7953
rect 42 7860 8367 7896
rect 42 7857 2933 7860
rect 42 7823 68 7857
rect 102 7823 138 7857
rect 172 7823 208 7857
rect 242 7823 278 7857
rect 312 7823 348 7857
rect 382 7823 418 7857
rect 452 7823 488 7857
rect 522 7823 558 7857
rect 592 7823 628 7857
rect 662 7823 698 7857
rect 732 7823 768 7857
rect 802 7823 838 7857
rect 872 7823 908 7857
rect 942 7823 978 7857
rect 1012 7823 1048 7857
rect 1082 7823 1118 7857
rect 1152 7823 1188 7857
rect 1222 7823 1258 7857
rect 1292 7823 1328 7857
rect 1362 7823 1398 7857
rect 1432 7823 1467 7857
rect 1501 7823 1536 7857
rect 1570 7823 1605 7857
rect 1639 7823 1674 7857
rect 1708 7823 1743 7857
rect 1777 7823 1812 7857
rect 1846 7823 1881 7857
rect 1915 7823 1950 7857
rect 1984 7823 2019 7857
rect 2053 7823 2088 7857
rect 2122 7823 2157 7857
rect 2191 7823 2226 7857
rect 2260 7823 2295 7857
rect 2329 7823 2364 7857
rect 2398 7823 2433 7857
rect 2467 7823 2502 7857
rect 2536 7823 2571 7857
rect 2605 7823 2640 7857
rect 2674 7823 2709 7857
rect 2743 7823 2778 7857
rect 2812 7823 2847 7857
rect 2881 7826 2933 7857
rect 2967 7826 3002 7860
rect 3036 7826 3071 7860
rect 3105 7826 3139 7860
rect 3173 7826 3207 7860
rect 3241 7826 3275 7860
rect 3309 7826 3343 7860
rect 3377 7826 3411 7860
rect 3445 7826 3479 7860
rect 3513 7826 3547 7860
rect 3581 7826 3615 7860
rect 3649 7826 3683 7860
rect 3717 7826 3751 7860
rect 3785 7826 3819 7860
rect 3853 7826 3887 7860
rect 3921 7826 3955 7860
rect 3989 7826 4023 7860
rect 4057 7826 4091 7860
rect 4125 7826 4159 7860
rect 4193 7826 4227 7860
rect 4261 7826 4295 7860
rect 4329 7826 4363 7860
rect 4397 7826 4431 7860
rect 4465 7826 4499 7860
rect 4533 7826 4567 7860
rect 4601 7826 4635 7860
rect 4669 7826 4703 7860
rect 4737 7826 4771 7860
rect 4805 7826 4839 7860
rect 4873 7826 4907 7860
rect 4941 7826 4975 7860
rect 5009 7826 5043 7860
rect 5077 7826 5111 7860
rect 5145 7826 5179 7860
rect 5213 7826 5247 7860
rect 5281 7826 5315 7860
rect 5349 7826 5383 7860
rect 5417 7826 5451 7860
rect 5485 7826 5519 7860
rect 5553 7826 5587 7860
rect 5621 7826 5655 7860
rect 5689 7826 5723 7860
rect 5757 7826 5791 7860
rect 5825 7826 5859 7860
rect 5893 7826 5927 7860
rect 5961 7826 5995 7860
rect 6029 7826 6063 7860
rect 6097 7826 6131 7860
rect 6165 7826 6199 7860
rect 6233 7826 6267 7860
rect 6301 7826 6335 7860
rect 6369 7826 6403 7860
rect 6437 7826 6471 7860
rect 6505 7826 6539 7860
rect 6573 7826 6607 7860
rect 6641 7826 6675 7860
rect 6709 7826 6743 7860
rect 6777 7826 6811 7860
rect 6845 7826 6879 7860
rect 6913 7826 6947 7860
rect 6981 7826 7015 7860
rect 7049 7826 7083 7860
rect 7117 7826 7151 7860
rect 7185 7826 7219 7860
rect 7253 7826 7287 7860
rect 7321 7826 7355 7860
rect 7389 7826 7423 7860
rect 7457 7826 7491 7860
rect 7525 7826 7559 7860
rect 7593 7826 7627 7860
rect 7661 7826 7695 7860
rect 7729 7826 7763 7860
rect 7797 7826 7831 7860
rect 7865 7826 7899 7860
rect 7933 7826 7967 7860
rect 8001 7826 8035 7860
rect 8069 7826 8103 7860
rect 8137 7826 8171 7860
rect 8205 7826 8239 7860
rect 8273 7826 8307 7860
rect 8341 7826 8367 7860
rect 2881 7823 8367 7826
rect 42 7788 8367 7823
rect 13506 7916 14431 7950
rect 14465 7916 14511 7950
rect 14545 7944 15102 7950
rect 14545 7916 14614 7944
rect 13506 7913 14614 7916
rect 14648 7913 14692 7944
rect 14726 7913 14770 7944
rect 14804 7913 14848 7944
rect 14882 7913 14926 7944
rect 14960 7929 15004 7944
rect 15038 7929 15102 7944
rect 13506 7879 13532 7913
rect 13566 7879 13603 7913
rect 13637 7879 13674 7913
rect 13708 7879 13744 7913
rect 13778 7879 13814 7913
rect 13848 7879 13884 7913
rect 13918 7879 13954 7913
rect 13988 7879 14024 7913
rect 14058 7879 14094 7913
rect 14128 7879 14164 7913
rect 14198 7879 14234 7913
rect 14268 7879 14304 7913
rect 14338 7879 14374 7913
rect 14408 7879 14444 7913
rect 14478 7879 14514 7913
rect 14548 7879 14584 7913
rect 14648 7910 14654 7913
rect 14618 7879 14654 7910
rect 14688 7910 14692 7913
rect 14758 7910 14770 7913
rect 14828 7910 14848 7913
rect 14898 7910 14926 7913
rect 14688 7879 14724 7910
rect 14758 7879 14794 7910
rect 14828 7879 14864 7910
rect 14898 7895 14932 7910
rect 14966 7895 15000 7929
rect 15038 7910 15068 7929
rect 15034 7895 15068 7910
rect 14898 7879 15102 7895
rect 13506 7870 15102 7879
rect 13506 7839 14614 7870
rect 14648 7839 14692 7870
rect 14726 7839 14770 7870
rect 14804 7839 14848 7870
rect 14882 7839 14926 7870
rect 14960 7857 15004 7870
rect 15038 7857 15102 7870
rect 13506 7805 13532 7839
rect 13566 7805 13603 7839
rect 13637 7805 13674 7839
rect 13708 7805 13744 7839
rect 13778 7805 13814 7839
rect 13848 7805 13884 7839
rect 13918 7805 13954 7839
rect 13988 7805 14024 7839
rect 14058 7805 14094 7839
rect 14128 7805 14164 7839
rect 14198 7805 14234 7839
rect 14268 7805 14304 7839
rect 14338 7805 14374 7839
rect 14408 7805 14444 7839
rect 14478 7805 14514 7839
rect 14548 7805 14584 7839
rect 14648 7836 14654 7839
rect 14618 7805 14654 7836
rect 14688 7836 14692 7839
rect 14758 7836 14770 7839
rect 14828 7836 14848 7839
rect 14898 7836 14926 7839
rect 14688 7805 14724 7836
rect 14758 7805 14794 7836
rect 14828 7805 14864 7836
rect 14898 7823 14932 7836
rect 14966 7823 15000 7857
rect 15038 7836 15068 7857
rect 15034 7823 15068 7836
rect 14898 7805 15102 7823
rect 13506 7796 15102 7805
rect 13506 7788 14614 7796
rect 42 7762 14614 7788
rect 14648 7762 14692 7796
rect 14726 7762 14770 7796
rect 14804 7762 14848 7796
rect 14882 7762 14926 7796
rect 14960 7785 15004 7796
rect 15038 7785 15102 7796
rect 42 7751 14932 7762
rect 14966 7751 15000 7785
rect 15038 7762 15068 7785
rect 15034 7751 15068 7762
rect 42 7749 15102 7751
rect 42 7715 68 7749
rect 102 7715 137 7749
rect 171 7715 206 7749
rect 240 7715 275 7749
rect 309 7715 344 7749
rect 378 7715 413 7749
rect 447 7715 482 7749
rect 516 7715 551 7749
rect 585 7715 620 7749
rect 654 7715 689 7749
rect 723 7715 758 7749
rect 792 7715 827 7749
rect 861 7715 896 7749
rect 930 7715 965 7749
rect 999 7715 1034 7749
rect 1068 7715 1103 7749
rect 1137 7715 1172 7749
rect 1206 7715 1241 7749
rect 1275 7715 1310 7749
rect 1344 7715 1379 7749
rect 1413 7715 1448 7749
rect 1482 7715 1517 7749
rect 1551 7715 1586 7749
rect 1620 7715 1655 7749
rect 1689 7715 1724 7749
rect 1758 7715 1793 7749
rect 1827 7715 1862 7749
rect 1896 7715 1931 7749
rect 1965 7715 2000 7749
rect 2034 7715 2069 7749
rect 2103 7715 2138 7749
rect 2172 7715 2207 7749
rect 2241 7715 2276 7749
rect 2310 7715 2345 7749
rect 2379 7715 2414 7749
rect 2448 7715 2483 7749
rect 2517 7715 2552 7749
rect 2586 7715 2621 7749
rect 2655 7715 2690 7749
rect 2724 7715 2759 7749
rect 2793 7715 2828 7749
rect 2862 7715 2896 7749
rect 2930 7715 2964 7749
rect 2998 7715 3032 7749
rect 3066 7715 3100 7749
rect 3134 7715 3168 7749
rect 3202 7715 3236 7749
rect 3270 7715 3304 7749
rect 3338 7715 3372 7749
rect 3406 7715 3440 7749
rect 3474 7715 3508 7749
rect 3542 7715 3576 7749
rect 3610 7715 3644 7749
rect 3678 7715 3712 7749
rect 3746 7715 3780 7749
rect 3814 7715 3848 7749
rect 3882 7715 3916 7749
rect 3950 7715 3984 7749
rect 4018 7715 4052 7749
rect 4086 7715 4120 7749
rect 4154 7715 4188 7749
rect 4222 7715 4256 7749
rect 4290 7715 4324 7749
rect 4358 7715 4392 7749
rect 4426 7715 4460 7749
rect 4494 7715 4528 7749
rect 4562 7715 4596 7749
rect 4630 7715 4664 7749
rect 4698 7715 4732 7749
rect 4766 7715 4800 7749
rect 4834 7715 4868 7749
rect 4902 7715 4936 7749
rect 4970 7715 5004 7749
rect 5038 7715 5072 7749
rect 5106 7715 5140 7749
rect 5174 7715 5208 7749
rect 5242 7715 5276 7749
rect 5310 7715 5344 7749
rect 5378 7715 5412 7749
rect 5446 7715 5480 7749
rect 5514 7715 5548 7749
rect 5582 7715 5616 7749
rect 5650 7715 5684 7749
rect 5718 7715 5752 7749
rect 5786 7715 5820 7749
rect 5854 7715 5888 7749
rect 5922 7715 5956 7749
rect 5990 7715 6024 7749
rect 6058 7715 6092 7749
rect 6126 7715 6160 7749
rect 6194 7715 6228 7749
rect 6262 7715 6296 7749
rect 6330 7715 6364 7749
rect 6398 7715 6432 7749
rect 6466 7715 6500 7749
rect 6534 7715 6568 7749
rect 6602 7715 6636 7749
rect 6670 7715 6704 7749
rect 6738 7715 6772 7749
rect 6806 7715 6840 7749
rect 6874 7715 6908 7749
rect 6942 7715 6976 7749
rect 7010 7715 7044 7749
rect 7078 7715 7112 7749
rect 7146 7715 7180 7749
rect 7214 7715 7248 7749
rect 7282 7715 7316 7749
rect 7350 7715 7384 7749
rect 7418 7715 7452 7749
rect 7486 7715 7520 7749
rect 7554 7715 7588 7749
rect 7622 7715 7656 7749
rect 7690 7715 7724 7749
rect 7758 7715 7792 7749
rect 7826 7715 7860 7749
rect 7894 7715 7928 7749
rect 7962 7715 7996 7749
rect 8030 7715 8064 7749
rect 8098 7715 8132 7749
rect 8166 7715 8200 7749
rect 8234 7715 8268 7749
rect 8302 7715 8336 7749
rect 8370 7715 8404 7749
rect 8438 7715 8472 7749
rect 8506 7715 8540 7749
rect 8574 7715 8608 7749
rect 8642 7715 8676 7749
rect 8710 7715 8744 7749
rect 8778 7715 8812 7749
rect 8846 7715 8880 7749
rect 8914 7715 8948 7749
rect 8982 7715 9016 7749
rect 9050 7715 9084 7749
rect 9118 7715 9152 7749
rect 9186 7715 9220 7749
rect 9254 7715 9288 7749
rect 9322 7715 9356 7749
rect 9390 7715 9424 7749
rect 9458 7715 9492 7749
rect 9526 7715 9560 7749
rect 9594 7715 9628 7749
rect 9662 7715 9696 7749
rect 9730 7715 9764 7749
rect 9798 7715 9832 7749
rect 9866 7715 9900 7749
rect 9934 7715 9968 7749
rect 10002 7715 10036 7749
rect 10070 7715 10104 7749
rect 10138 7715 10172 7749
rect 10206 7715 10240 7749
rect 10274 7715 10308 7749
rect 10342 7715 10376 7749
rect 10410 7715 10444 7749
rect 10478 7715 10512 7749
rect 10546 7715 10580 7749
rect 10614 7715 10648 7749
rect 10682 7715 10716 7749
rect 10750 7715 10784 7749
rect 10818 7715 10852 7749
rect 10886 7715 10920 7749
rect 10954 7715 10988 7749
rect 11022 7715 11056 7749
rect 11090 7715 11124 7749
rect 11158 7715 11192 7749
rect 11226 7715 11260 7749
rect 11294 7715 11328 7749
rect 11362 7715 11396 7749
rect 11430 7715 11464 7749
rect 11498 7715 11532 7749
rect 11566 7715 11600 7749
rect 11634 7715 11668 7749
rect 11702 7715 11736 7749
rect 11770 7715 11804 7749
rect 11838 7715 11872 7749
rect 11906 7715 11940 7749
rect 11974 7715 12008 7749
rect 12042 7715 12076 7749
rect 12110 7715 12144 7749
rect 12178 7715 12212 7749
rect 12246 7715 12280 7749
rect 12314 7715 12348 7749
rect 12382 7715 12416 7749
rect 12450 7715 12484 7749
rect 12518 7715 12552 7749
rect 12586 7715 12620 7749
rect 12654 7715 12688 7749
rect 12722 7715 12756 7749
rect 12790 7715 12824 7749
rect 12858 7715 12892 7749
rect 12926 7715 12960 7749
rect 12994 7715 13028 7749
rect 13062 7715 13096 7749
rect 13130 7715 13164 7749
rect 13198 7715 13232 7749
rect 13266 7715 13300 7749
rect 13334 7715 13368 7749
rect 13402 7715 13436 7749
rect 13470 7715 13504 7749
rect 13538 7715 13572 7749
rect 13606 7715 13640 7749
rect 13674 7715 13708 7749
rect 13742 7715 13776 7749
rect 13810 7715 13844 7749
rect 13878 7715 13912 7749
rect 13946 7715 13980 7749
rect 14014 7715 14048 7749
rect 14082 7715 14116 7749
rect 14150 7715 14184 7749
rect 14218 7715 14252 7749
rect 14286 7715 14320 7749
rect 14354 7715 14388 7749
rect 14422 7715 14456 7749
rect 14490 7715 14524 7749
rect 14558 7715 14592 7749
rect 14626 7722 14660 7749
rect 14694 7722 14728 7749
rect 14648 7715 14660 7722
rect 14726 7715 14728 7722
rect 14762 7722 14796 7749
rect 14830 7722 14864 7749
rect 14898 7722 15102 7749
rect 14762 7715 14770 7722
rect 14830 7715 14848 7722
rect 14898 7715 14926 7722
rect 42 7688 14614 7715
rect 14648 7688 14692 7715
rect 14726 7688 14770 7715
rect 14804 7688 14848 7715
rect 14882 7688 14926 7715
rect 14960 7713 15004 7722
rect 15038 7713 15102 7722
rect 42 7679 14932 7688
rect 14966 7679 15000 7713
rect 15038 7688 15068 7713
rect 15034 7679 15068 7688
rect 42 7677 15102 7679
rect 34 7676 15102 7677
rect 34 7642 2733 7676
rect 34 7608 68 7642
rect 102 7608 137 7642
rect 171 7608 206 7642
rect 240 7608 275 7642
rect 309 7608 344 7642
rect 378 7608 413 7642
rect 447 7608 482 7642
rect 516 7608 551 7642
rect 585 7608 620 7642
rect 654 7608 689 7642
rect 723 7608 758 7642
rect 792 7608 827 7642
rect 861 7608 896 7642
rect 930 7608 965 7642
rect 999 7608 1033 7642
rect 1067 7608 1101 7642
rect 1135 7608 1169 7642
rect 1203 7608 1237 7642
rect 1271 7608 1305 7642
rect 1339 7608 1373 7642
rect 1407 7608 1441 7642
rect 1475 7608 1509 7642
rect 1543 7608 1577 7642
rect 1611 7608 1645 7642
rect 1679 7608 1713 7642
rect 1747 7608 1781 7642
rect 1815 7608 1849 7642
rect 1883 7608 1917 7642
rect 1951 7608 1985 7642
rect 2019 7608 2053 7642
rect 2087 7608 2121 7642
rect 2155 7608 2189 7642
rect 2223 7608 2257 7642
rect 2291 7608 2325 7642
rect 2359 7608 2393 7642
rect 2427 7608 2461 7642
rect 2495 7608 2529 7642
rect 2563 7608 2597 7642
rect 2631 7608 2665 7642
rect 2699 7608 2733 7642
rect 34 7570 2733 7608
rect 34 7536 68 7570
rect 102 7536 137 7570
rect 171 7536 206 7570
rect 240 7536 275 7570
rect 309 7536 344 7570
rect 378 7536 413 7570
rect 447 7536 482 7570
rect 516 7536 551 7570
rect 585 7536 620 7570
rect 654 7536 689 7570
rect 723 7536 758 7570
rect 792 7536 827 7570
rect 861 7536 896 7570
rect 930 7536 965 7570
rect 999 7536 1033 7570
rect 1067 7536 1101 7570
rect 1135 7536 1169 7570
rect 1203 7536 1237 7570
rect 1271 7536 1305 7570
rect 1339 7536 1373 7570
rect 1407 7536 1441 7570
rect 1475 7536 1509 7570
rect 1543 7536 1577 7570
rect 1611 7536 1645 7570
rect 1679 7536 1713 7570
rect 1747 7536 1781 7570
rect 1815 7536 1849 7570
rect 1883 7536 1917 7570
rect 1951 7536 1985 7570
rect 2019 7536 2053 7570
rect 2087 7536 2121 7570
rect 2155 7536 2189 7570
rect 2223 7536 2257 7570
rect 2291 7536 2325 7570
rect 2359 7536 2393 7570
rect 2427 7536 2461 7570
rect 2495 7536 2529 7570
rect 2563 7536 2597 7570
rect 2631 7536 2665 7570
rect 2699 7536 2733 7570
rect 34 7498 2733 7536
rect 34 7464 68 7498
rect 102 7464 137 7498
rect 171 7464 206 7498
rect 240 7464 275 7498
rect 309 7464 344 7498
rect 378 7464 413 7498
rect 447 7464 482 7498
rect 516 7464 551 7498
rect 585 7464 620 7498
rect 654 7464 689 7498
rect 723 7464 758 7498
rect 792 7464 827 7498
rect 861 7464 896 7498
rect 930 7464 965 7498
rect 999 7464 1033 7498
rect 1067 7464 1101 7498
rect 1135 7464 1169 7498
rect 1203 7464 1237 7498
rect 1271 7464 1305 7498
rect 1339 7464 1373 7498
rect 1407 7464 1441 7498
rect 1475 7464 1509 7498
rect 1543 7464 1577 7498
rect 1611 7464 1645 7498
rect 1679 7464 1713 7498
rect 1747 7464 1781 7498
rect 1815 7464 1849 7498
rect 1883 7464 1917 7498
rect 1951 7464 1985 7498
rect 2019 7464 2053 7498
rect 2087 7464 2121 7498
rect 2155 7464 2189 7498
rect 2223 7464 2257 7498
rect 2291 7464 2325 7498
rect 2359 7464 2393 7498
rect 2427 7464 2461 7498
rect 2495 7464 2529 7498
rect 2563 7464 2597 7498
rect 2631 7464 2665 7498
rect 2699 7464 2733 7498
rect 34 7426 2733 7464
rect 34 7392 68 7426
rect 102 7392 137 7426
rect 171 7392 206 7426
rect 240 7392 275 7426
rect 309 7392 344 7426
rect 378 7392 413 7426
rect 447 7392 482 7426
rect 516 7392 551 7426
rect 585 7392 620 7426
rect 654 7392 689 7426
rect 723 7392 758 7426
rect 792 7392 827 7426
rect 861 7392 896 7426
rect 930 7392 965 7426
rect 999 7392 1033 7426
rect 1067 7392 1101 7426
rect 1135 7392 1169 7426
rect 1203 7392 1237 7426
rect 1271 7392 1305 7426
rect 1339 7392 1373 7426
rect 1407 7392 1441 7426
rect 1475 7392 1509 7426
rect 1543 7392 1577 7426
rect 1611 7392 1645 7426
rect 1679 7392 1713 7426
rect 1747 7392 1781 7426
rect 1815 7392 1849 7426
rect 1883 7392 1917 7426
rect 1951 7392 1985 7426
rect 2019 7392 2053 7426
rect 2087 7392 2121 7426
rect 2155 7392 2189 7426
rect 2223 7392 2257 7426
rect 2291 7392 2325 7426
rect 2359 7392 2393 7426
rect 2427 7392 2461 7426
rect 2495 7392 2529 7426
rect 2563 7392 2597 7426
rect 2631 7392 2665 7426
rect 2699 7392 2733 7426
rect 34 7381 2733 7392
rect 12498 7648 15102 7676
rect 12498 7640 14614 7648
rect 14648 7640 14692 7648
rect 14726 7640 14770 7648
rect 14804 7640 14848 7648
rect 14882 7640 14926 7648
rect 14960 7641 15004 7648
rect 15038 7641 15102 7648
rect 12498 7606 12524 7640
rect 12558 7606 12593 7640
rect 12627 7606 12662 7640
rect 12696 7606 12731 7640
rect 12765 7606 12800 7640
rect 12834 7606 12869 7640
rect 12903 7606 12938 7640
rect 12972 7606 13007 7640
rect 13041 7606 13076 7640
rect 13110 7606 13145 7640
rect 13179 7606 13214 7640
rect 13248 7606 13283 7640
rect 13317 7606 13352 7640
rect 13386 7606 13421 7640
rect 13455 7606 13490 7640
rect 13524 7606 13559 7640
rect 13593 7606 13628 7640
rect 13662 7606 13697 7640
rect 13731 7606 13766 7640
rect 13800 7606 13835 7640
rect 13869 7606 13904 7640
rect 13938 7606 13973 7640
rect 14007 7606 14042 7640
rect 14076 7606 14111 7640
rect 14145 7606 14180 7640
rect 14214 7606 14249 7640
rect 14283 7606 14318 7640
rect 14352 7606 14387 7640
rect 14421 7606 14456 7640
rect 14490 7606 14524 7640
rect 14558 7606 14592 7640
rect 14648 7614 14660 7640
rect 14726 7614 14728 7640
rect 14626 7606 14660 7614
rect 14694 7606 14728 7614
rect 14762 7614 14770 7640
rect 14830 7614 14848 7640
rect 14898 7614 14926 7640
rect 14762 7606 14796 7614
rect 14830 7606 14864 7614
rect 14898 7607 14932 7614
rect 14966 7607 15000 7641
rect 15038 7614 15068 7641
rect 15034 7607 15068 7614
rect 14898 7606 15102 7607
rect 12498 7574 15102 7606
rect 12498 7556 14614 7574
rect 14648 7556 14692 7574
rect 14726 7556 14770 7574
rect 14804 7556 14848 7574
rect 14882 7556 14926 7574
rect 14960 7569 15004 7574
rect 15038 7569 15102 7574
rect 12498 7522 12524 7556
rect 12558 7522 12593 7556
rect 12627 7522 12662 7556
rect 12696 7522 12731 7556
rect 12765 7522 12800 7556
rect 12834 7522 12869 7556
rect 12903 7522 12938 7556
rect 12972 7522 13007 7556
rect 13041 7522 13076 7556
rect 13110 7522 13145 7556
rect 13179 7522 13214 7556
rect 13248 7522 13283 7556
rect 13317 7522 13352 7556
rect 13386 7522 13421 7556
rect 13455 7522 13490 7556
rect 13524 7522 13559 7556
rect 13593 7522 13628 7556
rect 13662 7522 13697 7556
rect 13731 7522 13766 7556
rect 13800 7522 13835 7556
rect 13869 7522 13904 7556
rect 13938 7522 13973 7556
rect 14007 7522 14042 7556
rect 14076 7522 14111 7556
rect 14145 7522 14180 7556
rect 14214 7522 14249 7556
rect 14283 7522 14318 7556
rect 14352 7522 14387 7556
rect 14421 7522 14456 7556
rect 14490 7522 14524 7556
rect 14558 7522 14592 7556
rect 14648 7540 14660 7556
rect 14726 7540 14728 7556
rect 14626 7522 14660 7540
rect 14694 7522 14728 7540
rect 14762 7540 14770 7556
rect 14830 7540 14848 7556
rect 14898 7540 14926 7556
rect 14762 7522 14796 7540
rect 14830 7522 14864 7540
rect 14898 7535 14932 7540
rect 14966 7535 15000 7569
rect 15038 7540 15068 7569
rect 15034 7535 15068 7540
rect 14898 7522 15102 7535
rect 12498 7499 15102 7522
rect 12498 7472 14614 7499
rect 14648 7472 14692 7499
rect 14726 7472 14770 7499
rect 14804 7472 14848 7499
rect 14882 7472 14926 7499
rect 14960 7497 15004 7499
rect 15038 7497 15102 7499
rect 12498 7438 12524 7472
rect 12558 7438 12593 7472
rect 12627 7438 12662 7472
rect 12696 7438 12731 7472
rect 12765 7438 12800 7472
rect 12834 7438 12869 7472
rect 12903 7438 12938 7472
rect 12972 7438 13007 7472
rect 13041 7438 13076 7472
rect 13110 7438 13145 7472
rect 13179 7438 13214 7472
rect 13248 7438 13283 7472
rect 13317 7438 13352 7472
rect 13386 7438 13421 7472
rect 13455 7438 13490 7472
rect 13524 7438 13559 7472
rect 13593 7438 13628 7472
rect 13662 7438 13697 7472
rect 13731 7438 13766 7472
rect 13800 7438 13835 7472
rect 13869 7438 13904 7472
rect 13938 7438 13973 7472
rect 14007 7438 14042 7472
rect 14076 7438 14111 7472
rect 14145 7438 14180 7472
rect 14214 7438 14249 7472
rect 14283 7438 14318 7472
rect 14352 7438 14387 7472
rect 14421 7438 14456 7472
rect 14490 7438 14524 7472
rect 14558 7438 14592 7472
rect 14648 7465 14660 7472
rect 14726 7465 14728 7472
rect 14626 7438 14660 7465
rect 14694 7438 14728 7465
rect 14762 7465 14770 7472
rect 14830 7465 14848 7472
rect 14898 7465 14926 7472
rect 14762 7438 14796 7465
rect 14830 7438 14864 7465
rect 14898 7463 14932 7465
rect 14966 7463 15000 7497
rect 15038 7465 15068 7497
rect 15034 7463 15068 7465
rect 14898 7438 15102 7463
rect 12498 7425 15102 7438
rect 12498 7424 14932 7425
rect 12498 7390 14614 7424
rect 14648 7390 14692 7424
rect 14726 7390 14770 7424
rect 14804 7390 14848 7424
rect 14882 7390 14926 7424
rect 14966 7391 15000 7425
rect 15034 7424 15068 7425
rect 15038 7391 15068 7424
rect 14960 7390 15004 7391
rect 15038 7390 15102 7391
rect 12498 7388 15102 7390
rect 25 7374 7756 7381
rect 25 7340 57 7374
rect 91 7354 132 7374
rect 166 7354 207 7374
rect 241 7354 282 7374
rect 316 7354 357 7374
rect 391 7354 432 7374
rect 466 7354 507 7374
rect 541 7354 582 7374
rect 616 7354 657 7374
rect 691 7354 732 7374
rect 766 7354 807 7374
rect 841 7354 882 7374
rect 916 7354 957 7374
rect 991 7354 1032 7374
rect 1066 7354 1107 7374
rect 1141 7354 1182 7374
rect 1216 7354 1256 7374
rect 1290 7354 1330 7374
rect 1364 7354 7756 7374
rect 102 7340 132 7354
rect 25 7320 68 7340
rect 102 7320 137 7340
rect 171 7320 206 7354
rect 241 7340 275 7354
rect 316 7340 344 7354
rect 391 7340 413 7354
rect 466 7340 482 7354
rect 541 7340 551 7354
rect 616 7340 620 7354
rect 240 7320 275 7340
rect 309 7320 344 7340
rect 378 7320 413 7340
rect 447 7320 482 7340
rect 516 7320 551 7340
rect 585 7320 620 7340
rect 654 7340 657 7354
rect 723 7340 732 7354
rect 792 7340 807 7354
rect 861 7340 882 7354
rect 930 7340 957 7354
rect 999 7340 1032 7354
rect 654 7320 689 7340
rect 723 7320 758 7340
rect 792 7320 827 7340
rect 861 7320 896 7340
rect 930 7320 965 7340
rect 999 7320 1033 7340
rect 1067 7320 1101 7354
rect 1141 7340 1169 7354
rect 1216 7340 1237 7354
rect 1290 7340 1305 7354
rect 1364 7340 1373 7354
rect 1135 7320 1169 7340
rect 1203 7320 1237 7340
rect 1271 7320 1305 7340
rect 1339 7320 1373 7340
rect 1407 7320 1441 7354
rect 1475 7320 1509 7354
rect 1543 7320 1577 7354
rect 1611 7320 1645 7354
rect 1679 7320 1713 7354
rect 1747 7320 1781 7354
rect 1815 7320 1849 7354
rect 1883 7320 1917 7354
rect 1951 7320 1985 7354
rect 2019 7320 2053 7354
rect 2087 7320 2121 7354
rect 2155 7320 2189 7354
rect 2223 7320 2257 7354
rect 2291 7320 2325 7354
rect 2359 7320 2393 7354
rect 2427 7320 2461 7354
rect 2495 7320 2529 7354
rect 2563 7320 2597 7354
rect 2631 7320 2665 7354
rect 2699 7320 7756 7354
rect 25 7290 7756 7320
rect 12498 7354 12524 7388
rect 12558 7354 12593 7388
rect 12627 7354 12662 7388
rect 12696 7354 12731 7388
rect 12765 7354 12800 7388
rect 12834 7354 12869 7388
rect 12903 7354 12938 7388
rect 12972 7354 13007 7388
rect 13041 7354 13076 7388
rect 13110 7354 13145 7388
rect 13179 7354 13214 7388
rect 13248 7354 13283 7388
rect 13317 7354 13352 7388
rect 13386 7354 13421 7388
rect 13455 7354 13490 7388
rect 13524 7354 13559 7388
rect 13593 7354 13628 7388
rect 13662 7354 13697 7388
rect 13731 7354 13766 7388
rect 13800 7354 13835 7388
rect 13869 7354 13904 7388
rect 13938 7354 13973 7388
rect 14007 7354 14042 7388
rect 14076 7354 14111 7388
rect 14145 7354 14180 7388
rect 14214 7354 14249 7388
rect 14283 7354 14318 7388
rect 14352 7354 14387 7388
rect 14421 7354 14456 7388
rect 14490 7354 14524 7388
rect 14558 7354 14592 7388
rect 14626 7354 14660 7388
rect 14694 7354 14728 7388
rect 14762 7354 14796 7388
rect 14830 7354 14864 7388
rect 14898 7354 15102 7388
rect 12498 7353 15102 7354
rect 12498 7349 14932 7353
rect 12498 7317 14614 7349
rect 25 7256 57 7290
rect 91 7282 132 7290
rect 166 7282 207 7290
rect 241 7282 282 7290
rect 316 7282 357 7290
rect 391 7282 432 7290
rect 466 7282 507 7290
rect 541 7282 582 7290
rect 616 7282 657 7290
rect 691 7282 732 7290
rect 766 7282 807 7290
rect 841 7282 882 7290
rect 916 7282 957 7290
rect 991 7282 1032 7290
rect 1066 7282 1107 7290
rect 1141 7282 1182 7290
rect 1216 7282 1256 7290
rect 1290 7282 1330 7290
rect 1364 7282 7756 7290
rect 102 7256 132 7282
rect 25 7248 68 7256
rect 102 7248 137 7256
rect 171 7248 206 7282
rect 241 7256 275 7282
rect 316 7256 344 7282
rect 391 7256 413 7282
rect 466 7256 482 7282
rect 541 7256 551 7282
rect 616 7256 620 7282
rect 240 7248 275 7256
rect 309 7248 344 7256
rect 378 7248 413 7256
rect 447 7248 482 7256
rect 516 7248 551 7256
rect 585 7248 620 7256
rect 654 7256 657 7282
rect 723 7256 732 7282
rect 792 7256 807 7282
rect 861 7256 882 7282
rect 930 7256 957 7282
rect 999 7256 1032 7282
rect 654 7248 689 7256
rect 723 7248 758 7256
rect 792 7248 827 7256
rect 861 7248 896 7256
rect 930 7248 965 7256
rect 999 7248 1033 7256
rect 1067 7248 1101 7282
rect 1141 7256 1169 7282
rect 1216 7256 1237 7282
rect 1290 7256 1305 7282
rect 1364 7256 1373 7282
rect 1135 7248 1169 7256
rect 1203 7248 1237 7256
rect 1271 7248 1305 7256
rect 1339 7248 1373 7256
rect 1407 7248 1441 7282
rect 1475 7248 1509 7282
rect 1543 7248 1577 7282
rect 1611 7248 1645 7282
rect 1679 7248 1713 7282
rect 1747 7248 1781 7282
rect 1815 7248 1849 7282
rect 1883 7248 1917 7282
rect 1951 7248 1985 7282
rect 2019 7248 2053 7282
rect 2087 7248 2121 7282
rect 2155 7248 2189 7282
rect 2223 7248 2257 7282
rect 2291 7248 2325 7282
rect 2359 7248 2393 7282
rect 2427 7248 2461 7282
rect 2495 7248 2529 7282
rect 2563 7248 2597 7282
rect 2631 7248 2665 7282
rect 2699 7248 7756 7282
rect 25 7220 7756 7248
rect 25 7210 1431 7220
rect 1465 7210 1504 7220
rect 1538 7210 1577 7220
rect 1611 7210 1650 7220
rect 1684 7210 1723 7220
rect 1757 7210 1796 7220
rect 1830 7210 1869 7220
rect 1903 7210 1942 7220
rect 1976 7210 2015 7220
rect 2049 7210 2088 7220
rect 2122 7210 2161 7220
rect 2195 7210 2234 7220
rect 2268 7210 2307 7220
rect 2341 7210 2380 7220
rect 2414 7210 2453 7220
rect 2487 7210 2526 7220
rect 2560 7210 2599 7220
rect 2633 7210 2672 7220
rect 25 7206 68 7210
rect 102 7206 137 7210
rect 25 7172 57 7206
rect 102 7176 132 7206
rect 171 7176 206 7210
rect 240 7206 275 7210
rect 309 7206 344 7210
rect 378 7206 413 7210
rect 447 7206 482 7210
rect 516 7206 551 7210
rect 585 7206 620 7210
rect 241 7176 275 7206
rect 316 7176 344 7206
rect 391 7176 413 7206
rect 466 7176 482 7206
rect 541 7176 551 7206
rect 616 7176 620 7206
rect 654 7206 689 7210
rect 723 7206 758 7210
rect 792 7206 827 7210
rect 861 7206 896 7210
rect 930 7206 965 7210
rect 999 7206 1033 7210
rect 654 7176 657 7206
rect 723 7176 732 7206
rect 792 7176 807 7206
rect 861 7176 882 7206
rect 930 7176 957 7206
rect 999 7176 1032 7206
rect 1067 7176 1101 7210
rect 1135 7206 1169 7210
rect 1203 7206 1237 7210
rect 1271 7206 1305 7210
rect 1339 7206 1373 7210
rect 1141 7176 1169 7206
rect 1216 7176 1237 7206
rect 1290 7176 1305 7206
rect 1364 7176 1373 7206
rect 1407 7186 1431 7210
rect 1475 7186 1504 7210
rect 1407 7176 1441 7186
rect 1475 7176 1509 7186
rect 1543 7176 1577 7210
rect 1611 7176 1645 7210
rect 1684 7186 1713 7210
rect 1757 7186 1781 7210
rect 1830 7186 1849 7210
rect 1903 7186 1917 7210
rect 1976 7186 1985 7210
rect 2049 7186 2053 7210
rect 1679 7176 1713 7186
rect 1747 7176 1781 7186
rect 1815 7176 1849 7186
rect 1883 7176 1917 7186
rect 1951 7176 1985 7186
rect 2019 7176 2053 7186
rect 2087 7186 2088 7210
rect 2155 7186 2161 7210
rect 2223 7186 2234 7210
rect 2291 7186 2307 7210
rect 2359 7186 2380 7210
rect 2427 7186 2453 7210
rect 2495 7186 2526 7210
rect 2087 7176 2121 7186
rect 2155 7176 2189 7186
rect 2223 7176 2257 7186
rect 2291 7176 2325 7186
rect 2359 7176 2393 7186
rect 2427 7176 2461 7186
rect 2495 7176 2529 7186
rect 2563 7176 2597 7210
rect 2633 7186 2665 7210
rect 2706 7186 2745 7220
rect 2779 7186 2818 7220
rect 2852 7186 2891 7220
rect 2925 7186 2964 7220
rect 2998 7186 3037 7220
rect 3071 7186 3110 7220
rect 3144 7186 3183 7220
rect 3217 7186 3256 7220
rect 3290 7186 3329 7220
rect 3363 7186 3402 7220
rect 3436 7186 3475 7220
rect 3509 7186 3548 7220
rect 3582 7186 3621 7220
rect 3655 7186 3694 7220
rect 3728 7186 3767 7220
rect 3801 7186 3840 7220
rect 3874 7186 3913 7220
rect 3947 7186 3986 7220
rect 4020 7186 4059 7220
rect 4093 7186 4132 7220
rect 4166 7186 4205 7220
rect 4239 7186 4278 7220
rect 4312 7186 4351 7220
rect 4385 7186 4424 7220
rect 4458 7186 4497 7220
rect 4531 7186 4570 7220
rect 4604 7186 4643 7220
rect 4677 7186 4716 7220
rect 4750 7186 4789 7220
rect 4823 7186 4862 7220
rect 4896 7186 4935 7220
rect 4969 7186 5008 7220
rect 5042 7186 5081 7220
rect 5115 7186 5154 7220
rect 5188 7186 5227 7220
rect 5261 7186 5300 7220
rect 5334 7186 5373 7220
rect 5407 7186 5446 7220
rect 5480 7186 5519 7220
rect 5553 7186 5592 7220
rect 5626 7186 5665 7220
rect 5699 7186 5738 7220
rect 5772 7186 5811 7220
rect 5845 7186 5884 7220
rect 5918 7186 5957 7220
rect 5991 7186 6030 7220
rect 6064 7186 6103 7220
rect 6137 7186 6176 7220
rect 6210 7186 6249 7220
rect 6283 7186 6322 7220
rect 6356 7186 6395 7220
rect 6429 7186 6468 7220
rect 6502 7186 6540 7220
rect 6574 7186 6612 7220
rect 6646 7186 6684 7220
rect 6718 7186 6756 7220
rect 6790 7186 6828 7220
rect 6862 7186 6900 7220
rect 6934 7186 6972 7220
rect 7006 7186 7044 7220
rect 7078 7186 7116 7220
rect 7150 7186 7756 7220
rect 2631 7176 2665 7186
rect 2699 7176 7756 7186
rect 91 7172 132 7176
rect 166 7172 207 7176
rect 241 7172 282 7176
rect 316 7172 357 7176
rect 391 7172 432 7176
rect 466 7172 507 7176
rect 541 7172 582 7176
rect 616 7172 657 7176
rect 691 7172 732 7176
rect 766 7172 807 7176
rect 841 7172 882 7176
rect 916 7172 957 7176
rect 991 7172 1032 7176
rect 1066 7172 1107 7176
rect 1141 7172 1182 7176
rect 1216 7172 1256 7176
rect 1290 7172 1330 7176
rect 1364 7172 7756 7176
rect 25 7138 7756 7172
rect 25 7122 68 7138
rect 102 7122 137 7138
rect 25 7088 57 7122
rect 102 7104 132 7122
rect 171 7104 206 7138
rect 240 7122 275 7138
rect 309 7122 344 7138
rect 378 7122 413 7138
rect 447 7122 482 7138
rect 516 7122 551 7138
rect 585 7122 620 7138
rect 241 7104 275 7122
rect 316 7104 344 7122
rect 391 7104 413 7122
rect 466 7104 482 7122
rect 541 7104 551 7122
rect 616 7104 620 7122
rect 654 7122 689 7138
rect 723 7122 758 7138
rect 792 7122 827 7138
rect 861 7122 896 7138
rect 930 7122 965 7138
rect 999 7122 1033 7138
rect 654 7104 657 7122
rect 723 7104 732 7122
rect 792 7104 807 7122
rect 861 7104 882 7122
rect 930 7104 957 7122
rect 999 7104 1032 7122
rect 1067 7104 1101 7138
rect 1135 7122 1169 7138
rect 1203 7122 1237 7138
rect 1271 7122 1305 7138
rect 1339 7122 1373 7138
rect 1141 7104 1169 7122
rect 1216 7104 1237 7122
rect 1290 7104 1305 7122
rect 1364 7104 1373 7122
rect 1407 7104 1441 7138
rect 1475 7104 1509 7138
rect 1543 7104 1577 7138
rect 1611 7104 1645 7138
rect 1679 7104 1713 7138
rect 1747 7104 1781 7138
rect 1815 7104 1849 7138
rect 1883 7104 1917 7138
rect 1951 7104 1985 7138
rect 2019 7104 2053 7138
rect 2087 7104 2121 7138
rect 2155 7104 2189 7138
rect 2223 7104 2257 7138
rect 2291 7104 2325 7138
rect 2359 7104 2393 7138
rect 2427 7104 2461 7138
rect 2495 7104 2529 7138
rect 2563 7104 2597 7138
rect 2631 7104 2665 7138
rect 2699 7104 7756 7138
rect 91 7088 132 7104
rect 166 7088 207 7104
rect 241 7088 282 7104
rect 316 7088 357 7104
rect 391 7088 432 7104
rect 466 7088 507 7104
rect 541 7088 582 7104
rect 616 7088 657 7104
rect 691 7088 732 7104
rect 766 7088 807 7104
rect 841 7088 882 7104
rect 916 7088 957 7104
rect 991 7088 1032 7104
rect 1066 7088 1107 7104
rect 1141 7088 1182 7104
rect 1216 7088 1256 7104
rect 1290 7088 1330 7104
rect 1364 7088 7756 7104
rect 25 7066 7756 7088
rect 25 7038 68 7066
rect 102 7038 137 7066
rect 25 7004 57 7038
rect 102 7032 132 7038
rect 171 7032 206 7066
rect 240 7038 275 7066
rect 309 7038 344 7066
rect 378 7038 413 7066
rect 447 7038 482 7066
rect 516 7038 551 7066
rect 585 7038 620 7066
rect 241 7032 275 7038
rect 316 7032 344 7038
rect 391 7032 413 7038
rect 466 7032 482 7038
rect 541 7032 551 7038
rect 616 7032 620 7038
rect 654 7038 689 7066
rect 723 7038 758 7066
rect 792 7038 827 7066
rect 861 7038 896 7066
rect 930 7038 965 7066
rect 999 7038 1033 7066
rect 654 7032 657 7038
rect 723 7032 732 7038
rect 792 7032 807 7038
rect 861 7032 882 7038
rect 930 7032 957 7038
rect 999 7032 1032 7038
rect 1067 7032 1101 7066
rect 1135 7038 1169 7066
rect 1203 7038 1237 7066
rect 1271 7038 1305 7066
rect 1339 7038 1373 7066
rect 1141 7032 1169 7038
rect 1216 7032 1237 7038
rect 1290 7032 1305 7038
rect 1364 7032 1373 7038
rect 1407 7032 1441 7066
rect 1475 7032 1509 7066
rect 1543 7032 1577 7066
rect 1611 7032 1645 7066
rect 1679 7032 1713 7066
rect 1747 7032 1781 7066
rect 1815 7032 1849 7066
rect 1883 7032 1917 7066
rect 1951 7032 1985 7066
rect 2019 7032 2053 7066
rect 2087 7032 2121 7066
rect 2155 7032 2189 7066
rect 2223 7032 2257 7066
rect 2291 7032 2325 7066
rect 2359 7032 2393 7066
rect 2427 7032 2461 7066
rect 2495 7032 2529 7066
rect 2563 7032 2597 7066
rect 2631 7032 2665 7066
rect 2699 7047 7756 7066
rect 2699 7032 2757 7047
rect 91 7004 132 7032
rect 166 7004 207 7032
rect 241 7004 282 7032
rect 316 7004 357 7032
rect 391 7004 432 7032
rect 466 7004 507 7032
rect 541 7004 582 7032
rect 616 7004 657 7032
rect 691 7004 732 7032
rect 766 7004 807 7032
rect 841 7004 882 7032
rect 916 7004 957 7032
rect 991 7004 1032 7032
rect 1066 7004 1107 7032
rect 1141 7004 1182 7032
rect 1216 7004 1256 7032
rect 1290 7004 1330 7032
rect 1364 7013 2757 7032
rect 2791 7013 2825 7047
rect 2859 7013 2893 7047
rect 2927 7013 2961 7047
rect 2995 7013 3029 7047
rect 3063 7013 3097 7047
rect 3131 7013 3165 7047
rect 3199 7013 3233 7047
rect 3267 7013 3301 7047
rect 3335 7013 3369 7047
rect 3403 7013 3437 7047
rect 3471 7013 3505 7047
rect 3539 7013 3573 7047
rect 3607 7013 3641 7047
rect 3675 7013 3709 7047
rect 3743 7013 3777 7047
rect 3811 7013 3845 7047
rect 3879 7013 3913 7047
rect 3947 7013 3981 7047
rect 4015 7013 4049 7047
rect 4083 7013 4117 7047
rect 4151 7013 4185 7047
rect 4219 7013 4253 7047
rect 4287 7013 4321 7047
rect 4355 7013 4389 7047
rect 4423 7013 4457 7047
rect 4491 7013 4525 7047
rect 4559 7013 4593 7047
rect 4627 7013 4661 7047
rect 4695 7013 4729 7047
rect 4763 7013 4797 7047
rect 4831 7013 4865 7047
rect 4899 7013 4933 7047
rect 4967 7013 5001 7047
rect 5035 7013 5069 7047
rect 5103 7013 5137 7047
rect 5171 7013 5205 7047
rect 5239 7013 5273 7047
rect 5307 7013 5341 7047
rect 5375 7013 5409 7047
rect 5443 7013 5477 7047
rect 5511 7013 5545 7047
rect 5579 7013 5613 7047
rect 5647 7013 5681 7047
rect 5715 7013 5749 7047
rect 5783 7013 5817 7047
rect 5851 7013 5885 7047
rect 5919 7013 5953 7047
rect 5987 7013 6021 7047
rect 6055 7013 6089 7047
rect 6123 7013 6157 7047
rect 6191 7013 6225 7047
rect 6259 7013 6293 7047
rect 6327 7013 6361 7047
rect 6395 7013 6429 7047
rect 6463 7013 6497 7047
rect 6531 7013 6565 7047
rect 6599 7013 6633 7047
rect 6667 7013 6701 7047
rect 6735 7013 6769 7047
rect 6803 7013 6837 7047
rect 6871 7013 6905 7047
rect 6939 7013 6973 7047
rect 7007 7013 7041 7047
rect 7075 7013 7109 7047
rect 7143 7013 7177 7047
rect 7211 7013 7245 7047
rect 7279 7013 7313 7047
rect 7347 7013 7381 7047
rect 7415 7013 7449 7047
rect 7483 7013 7517 7047
rect 7551 7013 7585 7047
rect 7619 7013 7653 7047
rect 7687 7013 7756 7047
rect 1364 7004 7756 7013
rect 25 6997 7756 7004
rect 7183 6957 7756 6997
rect 8184 7315 14614 7317
rect 14648 7315 14692 7349
rect 14726 7315 14770 7349
rect 14804 7315 14848 7349
rect 14882 7315 14926 7349
rect 14966 7319 15000 7353
rect 15034 7349 15068 7353
rect 15038 7319 15068 7349
rect 14960 7315 15004 7319
rect 15038 7315 15102 7319
rect 8184 7282 15102 7315
rect 8184 7248 8210 7282
rect 8244 7248 8279 7282
rect 8313 7248 8348 7282
rect 8382 7248 8417 7282
rect 8451 7248 8486 7282
rect 8520 7248 8555 7282
rect 8589 7248 8624 7282
rect 8658 7248 8693 7282
rect 8727 7248 8762 7282
rect 8796 7248 8831 7282
rect 8865 7248 8900 7282
rect 8934 7248 8969 7282
rect 9003 7248 9038 7282
rect 9072 7248 9107 7282
rect 9141 7248 9176 7282
rect 9210 7248 9245 7282
rect 9279 7248 9314 7282
rect 9348 7248 9383 7282
rect 9417 7248 9452 7282
rect 9486 7248 9521 7282
rect 9555 7248 9590 7282
rect 9624 7248 9659 7282
rect 9693 7248 9728 7282
rect 9762 7248 9797 7282
rect 9831 7248 9866 7282
rect 9900 7248 9935 7282
rect 9969 7248 10004 7282
rect 10038 7248 10073 7282
rect 10107 7248 10142 7282
rect 10176 7248 10211 7282
rect 10245 7248 10280 7282
rect 10314 7248 10349 7282
rect 10383 7248 10418 7282
rect 10452 7248 10487 7282
rect 10521 7248 10556 7282
rect 10590 7248 10625 7282
rect 10659 7248 10694 7282
rect 10728 7248 10763 7282
rect 10797 7248 10832 7282
rect 10866 7248 10901 7282
rect 10935 7248 10970 7282
rect 11004 7248 11039 7282
rect 11073 7248 11108 7282
rect 11142 7248 11177 7282
rect 11211 7248 11246 7282
rect 11280 7248 11315 7282
rect 11349 7248 11384 7282
rect 11418 7248 11453 7282
rect 11487 7248 11522 7282
rect 11556 7248 11591 7282
rect 11625 7248 11660 7282
rect 11694 7248 11729 7282
rect 11763 7248 11798 7282
rect 11832 7248 11867 7282
rect 11901 7248 11936 7282
rect 11970 7248 12005 7282
rect 12039 7248 12074 7282
rect 12108 7248 12143 7282
rect 12177 7248 12212 7282
rect 12246 7248 12280 7282
rect 12314 7248 12348 7282
rect 12382 7248 12416 7282
rect 12450 7248 12484 7282
rect 12518 7248 12552 7282
rect 12586 7248 12620 7282
rect 12654 7248 12688 7282
rect 12722 7248 12756 7282
rect 12790 7248 12824 7282
rect 12858 7248 12892 7282
rect 12926 7248 12960 7282
rect 12994 7248 13028 7282
rect 13062 7248 13096 7282
rect 13130 7248 13164 7282
rect 13198 7248 13232 7282
rect 13266 7248 13300 7282
rect 13334 7248 13368 7282
rect 13402 7248 13436 7282
rect 13470 7248 13504 7282
rect 13538 7248 13572 7282
rect 13606 7248 13640 7282
rect 13674 7248 13708 7282
rect 13742 7248 13776 7282
rect 13810 7248 13844 7282
rect 13878 7248 13912 7282
rect 13946 7248 13980 7282
rect 14014 7248 14048 7282
rect 14082 7248 14116 7282
rect 14150 7248 14184 7282
rect 14218 7248 14252 7282
rect 14286 7248 14320 7282
rect 14354 7248 14388 7282
rect 14422 7248 14456 7282
rect 14490 7248 14524 7282
rect 14558 7248 14592 7282
rect 14626 7274 14660 7282
rect 14694 7274 14728 7282
rect 14648 7248 14660 7274
rect 14726 7248 14728 7274
rect 14762 7274 14796 7282
rect 14830 7274 14864 7282
rect 14898 7281 15102 7282
rect 14898 7274 14932 7281
rect 14762 7248 14770 7274
rect 14830 7248 14848 7274
rect 14898 7248 14926 7274
rect 8184 7240 14614 7248
rect 14648 7240 14692 7248
rect 14726 7240 14770 7248
rect 14804 7240 14848 7248
rect 14882 7240 14926 7248
rect 14966 7247 15000 7281
rect 15034 7274 15068 7281
rect 15038 7247 15068 7274
rect 14960 7240 15004 7247
rect 15038 7240 15102 7247
rect 8184 7210 15102 7240
rect 8184 7176 8210 7210
rect 8244 7176 8279 7210
rect 8313 7176 8348 7210
rect 8382 7176 8417 7210
rect 8451 7176 8486 7210
rect 8520 7176 8555 7210
rect 8589 7176 8624 7210
rect 8658 7176 8693 7210
rect 8727 7176 8762 7210
rect 8796 7176 8831 7210
rect 8865 7176 8900 7210
rect 8934 7176 8969 7210
rect 9003 7176 9038 7210
rect 9072 7176 9107 7210
rect 9141 7176 9176 7210
rect 9210 7176 9245 7210
rect 9279 7176 9314 7210
rect 9348 7176 9383 7210
rect 9417 7176 9452 7210
rect 9486 7176 9521 7210
rect 9555 7176 9590 7210
rect 9624 7176 9659 7210
rect 9693 7176 9728 7210
rect 9762 7176 9797 7210
rect 9831 7176 9866 7210
rect 9900 7176 9935 7210
rect 9969 7176 10004 7210
rect 10038 7176 10073 7210
rect 10107 7176 10142 7210
rect 10176 7176 10211 7210
rect 10245 7176 10280 7210
rect 10314 7176 10349 7210
rect 10383 7176 10418 7210
rect 10452 7176 10487 7210
rect 10521 7176 10556 7210
rect 10590 7176 10625 7210
rect 10659 7176 10694 7210
rect 10728 7176 10763 7210
rect 10797 7176 10832 7210
rect 10866 7176 10901 7210
rect 10935 7176 10970 7210
rect 11004 7176 11039 7210
rect 11073 7176 11108 7210
rect 11142 7176 11177 7210
rect 11211 7176 11246 7210
rect 11280 7176 11315 7210
rect 11349 7176 11384 7210
rect 11418 7176 11453 7210
rect 11487 7176 11522 7210
rect 11556 7176 11591 7210
rect 11625 7176 11660 7210
rect 11694 7176 11729 7210
rect 11763 7176 11798 7210
rect 11832 7176 11867 7210
rect 11901 7176 11936 7210
rect 11970 7176 12005 7210
rect 12039 7176 12074 7210
rect 12108 7176 12143 7210
rect 12177 7176 12212 7210
rect 12246 7176 12280 7210
rect 12314 7176 12348 7210
rect 12382 7176 12416 7210
rect 12450 7176 12484 7210
rect 12518 7176 12552 7210
rect 12586 7176 12620 7210
rect 12654 7176 12688 7210
rect 12722 7176 12756 7210
rect 12790 7176 12824 7210
rect 12858 7176 12892 7210
rect 12926 7176 12960 7210
rect 12994 7176 13028 7210
rect 13062 7176 13096 7210
rect 13130 7176 13164 7210
rect 13198 7176 13232 7210
rect 13266 7176 13300 7210
rect 13334 7176 13368 7210
rect 13402 7176 13436 7210
rect 13470 7176 13504 7210
rect 13538 7176 13572 7210
rect 13606 7176 13640 7210
rect 13674 7176 13708 7210
rect 13742 7176 13776 7210
rect 13810 7176 13844 7210
rect 13878 7176 13912 7210
rect 13946 7176 13980 7210
rect 14014 7176 14048 7210
rect 14082 7176 14116 7210
rect 14150 7176 14184 7210
rect 14218 7176 14252 7210
rect 14286 7176 14320 7210
rect 14354 7176 14388 7210
rect 14422 7176 14456 7210
rect 14490 7176 14524 7210
rect 14558 7176 14592 7210
rect 14626 7199 14660 7210
rect 14694 7199 14728 7210
rect 14648 7176 14660 7199
rect 14726 7176 14728 7199
rect 14762 7199 14796 7210
rect 14830 7199 14864 7210
rect 14898 7209 15102 7210
rect 14898 7199 14932 7209
rect 14762 7176 14770 7199
rect 14830 7176 14848 7199
rect 14898 7176 14926 7199
rect 8184 7165 14614 7176
rect 14648 7165 14692 7176
rect 14726 7165 14770 7176
rect 14804 7165 14848 7176
rect 14882 7165 14926 7176
rect 14966 7175 15000 7209
rect 15034 7199 15068 7209
rect 15038 7175 15068 7199
rect 14960 7165 15004 7175
rect 15038 7165 15102 7175
rect 8184 7138 15102 7165
rect 8184 7104 8210 7138
rect 8244 7104 8279 7138
rect 8313 7104 8348 7138
rect 8382 7104 8417 7138
rect 8451 7104 8486 7138
rect 8520 7104 8555 7138
rect 8589 7104 8624 7138
rect 8658 7104 8693 7138
rect 8727 7104 8762 7138
rect 8796 7104 8831 7138
rect 8865 7104 8900 7138
rect 8934 7104 8969 7138
rect 9003 7104 9038 7138
rect 9072 7104 9107 7138
rect 9141 7104 9176 7138
rect 9210 7104 9245 7138
rect 9279 7104 9314 7138
rect 9348 7104 9383 7138
rect 9417 7104 9452 7138
rect 9486 7104 9521 7138
rect 9555 7104 9590 7138
rect 9624 7104 9659 7138
rect 9693 7104 9728 7138
rect 9762 7104 9797 7138
rect 9831 7104 9866 7138
rect 9900 7104 9935 7138
rect 9969 7104 10004 7138
rect 10038 7104 10073 7138
rect 10107 7104 10142 7138
rect 10176 7104 10211 7138
rect 10245 7104 10280 7138
rect 10314 7104 10349 7138
rect 10383 7104 10418 7138
rect 10452 7104 10487 7138
rect 10521 7104 10556 7138
rect 10590 7104 10625 7138
rect 10659 7104 10694 7138
rect 10728 7104 10763 7138
rect 10797 7104 10832 7138
rect 10866 7104 10901 7138
rect 10935 7104 10970 7138
rect 11004 7104 11039 7138
rect 11073 7104 11108 7138
rect 11142 7104 11177 7138
rect 11211 7104 11246 7138
rect 11280 7104 11315 7138
rect 11349 7104 11384 7138
rect 11418 7104 11453 7138
rect 11487 7104 11522 7138
rect 11556 7104 11591 7138
rect 11625 7104 11660 7138
rect 11694 7104 11729 7138
rect 11763 7104 11798 7138
rect 11832 7104 11867 7138
rect 11901 7104 11936 7138
rect 11970 7104 12005 7138
rect 12039 7104 12074 7138
rect 12108 7104 12143 7138
rect 12177 7104 12212 7138
rect 12246 7104 12280 7138
rect 12314 7104 12348 7138
rect 12382 7104 12416 7138
rect 12450 7104 12484 7138
rect 12518 7104 12552 7138
rect 12586 7104 12620 7138
rect 12654 7104 12688 7138
rect 12722 7104 12756 7138
rect 12790 7104 12824 7138
rect 12858 7104 12892 7138
rect 12926 7104 12960 7138
rect 12994 7104 13028 7138
rect 13062 7104 13096 7138
rect 13130 7104 13164 7138
rect 13198 7104 13232 7138
rect 13266 7104 13300 7138
rect 13334 7104 13368 7138
rect 13402 7104 13436 7138
rect 13470 7104 13504 7138
rect 13538 7104 13572 7138
rect 13606 7104 13640 7138
rect 13674 7104 13708 7138
rect 13742 7104 13776 7138
rect 13810 7104 13844 7138
rect 13878 7104 13912 7138
rect 13946 7104 13980 7138
rect 14014 7104 14048 7138
rect 14082 7104 14116 7138
rect 14150 7104 14184 7138
rect 14218 7104 14252 7138
rect 14286 7104 14320 7138
rect 14354 7104 14388 7138
rect 14422 7104 14456 7138
rect 14490 7104 14524 7138
rect 14558 7104 14592 7138
rect 14626 7124 14660 7138
rect 14694 7124 14728 7138
rect 14648 7104 14660 7124
rect 14726 7104 14728 7124
rect 14762 7124 14796 7138
rect 14830 7124 14864 7138
rect 14898 7137 15102 7138
rect 14898 7124 14932 7137
rect 14762 7104 14770 7124
rect 14830 7104 14848 7124
rect 14898 7104 14926 7124
rect 8184 7090 14614 7104
rect 14648 7090 14692 7104
rect 14726 7090 14770 7104
rect 14804 7090 14848 7104
rect 14882 7090 14926 7104
rect 14966 7103 15000 7137
rect 15034 7124 15068 7137
rect 15038 7103 15068 7124
rect 14960 7090 15004 7103
rect 15038 7090 15102 7103
rect 8184 7066 15102 7090
rect 8184 7032 8210 7066
rect 8244 7032 8279 7066
rect 8313 7032 8348 7066
rect 8382 7032 8417 7066
rect 8451 7032 8486 7066
rect 8520 7032 8555 7066
rect 8589 7032 8624 7066
rect 8658 7032 8693 7066
rect 8727 7032 8762 7066
rect 8796 7032 8831 7066
rect 8865 7032 8900 7066
rect 8934 7032 8969 7066
rect 9003 7032 9038 7066
rect 9072 7032 9107 7066
rect 9141 7032 9176 7066
rect 9210 7032 9245 7066
rect 9279 7032 9314 7066
rect 9348 7032 9383 7066
rect 9417 7032 9452 7066
rect 9486 7032 9521 7066
rect 9555 7032 9590 7066
rect 9624 7032 9659 7066
rect 9693 7032 9728 7066
rect 9762 7032 9797 7066
rect 9831 7032 9866 7066
rect 9900 7032 9935 7066
rect 9969 7032 10004 7066
rect 10038 7032 10073 7066
rect 10107 7032 10142 7066
rect 10176 7032 10211 7066
rect 10245 7032 10280 7066
rect 10314 7032 10349 7066
rect 10383 7032 10418 7066
rect 10452 7032 10487 7066
rect 10521 7032 10556 7066
rect 10590 7032 10625 7066
rect 10659 7032 10694 7066
rect 10728 7032 10763 7066
rect 10797 7032 10832 7066
rect 10866 7032 10901 7066
rect 10935 7032 10970 7066
rect 11004 7032 11039 7066
rect 11073 7032 11108 7066
rect 11142 7032 11177 7066
rect 11211 7032 11246 7066
rect 11280 7032 11315 7066
rect 11349 7032 11384 7066
rect 11418 7032 11453 7066
rect 11487 7032 11522 7066
rect 11556 7032 11591 7066
rect 11625 7032 11660 7066
rect 11694 7032 11729 7066
rect 11763 7032 11798 7066
rect 11832 7032 11867 7066
rect 11901 7032 11936 7066
rect 11970 7032 12005 7066
rect 12039 7032 12074 7066
rect 12108 7032 12143 7066
rect 12177 7032 12212 7066
rect 12246 7032 12280 7066
rect 12314 7032 12348 7066
rect 12382 7032 12416 7066
rect 12450 7032 12484 7066
rect 12518 7032 12552 7066
rect 12586 7032 12620 7066
rect 12654 7032 12688 7066
rect 12722 7032 12756 7066
rect 12790 7032 12824 7066
rect 12858 7032 12892 7066
rect 12926 7032 12960 7066
rect 12994 7032 13028 7066
rect 13062 7032 13096 7066
rect 13130 7032 13164 7066
rect 13198 7032 13232 7066
rect 13266 7032 13300 7066
rect 13334 7032 13368 7066
rect 13402 7032 13436 7066
rect 13470 7032 13504 7066
rect 13538 7032 13572 7066
rect 13606 7032 13640 7066
rect 13674 7032 13708 7066
rect 13742 7032 13776 7066
rect 13810 7032 13844 7066
rect 13878 7032 13912 7066
rect 13946 7032 13980 7066
rect 14014 7032 14048 7066
rect 14082 7032 14116 7066
rect 14150 7032 14184 7066
rect 14218 7032 14252 7066
rect 14286 7032 14320 7066
rect 14354 7032 14388 7066
rect 14422 7032 14456 7066
rect 14490 7032 14524 7066
rect 14558 7032 14592 7066
rect 14626 7032 14660 7066
rect 14694 7032 14728 7066
rect 14762 7032 14796 7066
rect 14830 7032 14864 7066
rect 14898 7065 15102 7066
rect 14898 7032 14932 7065
rect 8184 7031 14932 7032
rect 14966 7031 15000 7065
rect 15034 7031 15068 7065
rect 8184 6997 15102 7031
rect 8184 6957 8488 6997
rect 44 6809 68 6843
rect 102 6809 137 6843
rect 171 6809 206 6843
rect 240 6809 275 6843
rect 309 6809 344 6843
rect 378 6809 413 6843
rect 447 6809 482 6843
rect 516 6809 551 6843
rect 585 6809 620 6843
rect 654 6809 689 6843
rect 723 6809 758 6843
rect 792 6809 827 6843
rect 861 6809 896 6843
rect 930 6809 965 6843
rect 999 6809 1034 6843
rect 1068 6809 1103 6843
rect 1137 6809 1172 6843
rect 1206 6809 1241 6843
rect 1275 6809 1310 6843
rect 1344 6809 1379 6843
rect 1413 6809 1448 6843
rect 1482 6809 1517 6843
rect 1551 6809 1586 6843
rect 1620 6809 1655 6843
rect 1689 6809 1724 6843
rect 1758 6809 1793 6843
rect 1827 6809 1862 6843
rect 1896 6809 1931 6843
rect 1965 6809 2000 6843
rect 2034 6809 2069 6843
rect 2103 6809 2138 6843
rect 2172 6809 2207 6843
rect 2241 6809 2276 6843
rect 2310 6809 2345 6843
rect 2379 6809 2414 6843
rect 2448 6809 2483 6843
rect 2517 6809 2552 6843
rect 2586 6809 2621 6843
rect 2655 6809 2690 6843
rect 2724 6809 2759 6843
rect 2793 6809 2828 6843
rect 2862 6809 2897 6843
rect 2931 6809 2966 6843
rect 3000 6809 3035 6843
rect 3069 6809 3104 6843
rect 3138 6809 3173 6843
rect 3207 6809 3242 6843
rect 3276 6809 3310 6843
rect 3344 6809 3378 6843
rect 3412 6809 3446 6843
rect 3480 6809 3514 6843
rect 3548 6809 3582 6843
rect 3616 6809 3650 6843
rect 3684 6809 3718 6843
rect 3752 6809 3786 6843
rect 3820 6809 3854 6843
rect 3888 6809 3922 6843
rect 3956 6809 3990 6843
rect 4024 6809 4058 6843
rect 4092 6809 4126 6843
rect 4160 6809 4194 6843
rect 4228 6809 4262 6843
rect 4296 6809 4330 6843
rect 4364 6809 4398 6843
rect 4432 6809 4466 6843
rect 4500 6809 4534 6843
rect 4568 6809 4602 6843
rect 4636 6809 4670 6843
rect 4704 6809 4738 6843
rect 4772 6809 4806 6843
rect 4840 6809 4874 6843
rect 4908 6809 4942 6843
rect 4976 6809 5010 6843
rect 5044 6809 5078 6843
rect 5112 6809 5146 6843
rect 5180 6809 5214 6843
rect 5248 6809 5282 6843
rect 5316 6809 5350 6843
rect 5384 6809 5418 6843
rect 5452 6809 5486 6843
rect 5520 6809 5554 6843
rect 5588 6809 5622 6843
rect 5656 6809 5690 6843
rect 5724 6809 5758 6843
rect 5792 6809 5826 6843
rect 5860 6809 5894 6843
rect 5928 6809 5962 6843
rect 5996 6809 6030 6843
rect 6064 6809 6098 6843
rect 6132 6809 6166 6843
rect 6200 6809 6234 6843
rect 6268 6809 6302 6843
rect 6336 6809 6370 6843
rect 6404 6809 6438 6843
rect 6472 6809 6506 6843
rect 6540 6809 6574 6843
rect 6608 6809 6642 6843
rect 6676 6809 6710 6843
rect 6744 6809 6778 6843
rect 6812 6809 6846 6843
rect 6880 6809 6914 6843
rect 6948 6809 6982 6843
rect 7016 6809 7050 6843
rect 7084 6809 7108 6843
rect 44 6756 7108 6809
rect 44 6722 68 6756
rect 102 6722 137 6756
rect 171 6722 206 6756
rect 240 6722 275 6756
rect 309 6722 344 6756
rect 378 6722 413 6756
rect 447 6722 482 6756
rect 516 6722 551 6756
rect 585 6722 620 6756
rect 654 6722 689 6756
rect 723 6722 758 6756
rect 792 6722 827 6756
rect 861 6722 896 6756
rect 930 6722 965 6756
rect 999 6722 1034 6756
rect 1068 6722 1103 6756
rect 1137 6722 1172 6756
rect 1206 6722 1241 6756
rect 1275 6722 1310 6756
rect 1344 6722 1379 6756
rect 1413 6722 1448 6756
rect 1482 6722 1517 6756
rect 1551 6722 1586 6756
rect 1620 6722 1655 6756
rect 1689 6722 1724 6756
rect 1758 6722 1793 6756
rect 1827 6722 1862 6756
rect 1896 6722 1931 6756
rect 1965 6722 2000 6756
rect 2034 6722 2069 6756
rect 2103 6722 2138 6756
rect 2172 6722 2207 6756
rect 2241 6722 2276 6756
rect 2310 6722 2345 6756
rect 2379 6722 2414 6756
rect 2448 6722 2483 6756
rect 2517 6722 2552 6756
rect 2586 6722 2621 6756
rect 2655 6722 2690 6756
rect 2724 6722 2759 6756
rect 2793 6722 2828 6756
rect 2862 6722 2897 6756
rect 2931 6722 2966 6756
rect 3000 6722 3035 6756
rect 3069 6722 3104 6756
rect 3138 6722 3173 6756
rect 3207 6722 3242 6756
rect 3276 6722 3310 6756
rect 3344 6722 3378 6756
rect 3412 6722 3446 6756
rect 3480 6722 3514 6756
rect 3548 6722 3582 6756
rect 3616 6722 3650 6756
rect 3684 6722 3718 6756
rect 3752 6722 3786 6756
rect 3820 6722 3854 6756
rect 3888 6722 3922 6756
rect 3956 6722 3990 6756
rect 4024 6722 4058 6756
rect 4092 6722 4126 6756
rect 4160 6722 4194 6756
rect 4228 6722 4262 6756
rect 4296 6722 4330 6756
rect 4364 6722 4398 6756
rect 4432 6722 4466 6756
rect 4500 6722 4534 6756
rect 4568 6722 4602 6756
rect 4636 6722 4670 6756
rect 4704 6722 4738 6756
rect 4772 6722 4806 6756
rect 4840 6722 4874 6756
rect 4908 6722 4942 6756
rect 4976 6722 5010 6756
rect 5044 6722 5078 6756
rect 5112 6722 5146 6756
rect 5180 6722 5214 6756
rect 5248 6722 5282 6756
rect 5316 6722 5350 6756
rect 5384 6722 5418 6756
rect 5452 6722 5486 6756
rect 5520 6722 5554 6756
rect 5588 6722 5622 6756
rect 5656 6722 5690 6756
rect 5724 6722 5758 6756
rect 5792 6722 5826 6756
rect 5860 6722 5894 6756
rect 5928 6722 5962 6756
rect 5996 6722 6030 6756
rect 6064 6722 6098 6756
rect 6132 6722 6166 6756
rect 6200 6722 6234 6756
rect 6268 6722 6302 6756
rect 6336 6722 6370 6756
rect 6404 6722 6438 6756
rect 6472 6722 6506 6756
rect 6540 6722 6574 6756
rect 6608 6722 6642 6756
rect 6676 6722 6710 6756
rect 6744 6722 6778 6756
rect 6812 6722 6846 6756
rect 6880 6722 6914 6756
rect 6948 6722 6982 6756
rect 7016 6722 7050 6756
rect 7084 6722 7108 6756
rect 7183 6739 8488 6957
rect 12493 6809 12517 6843
rect 12551 6809 12586 6843
rect 12620 6809 12655 6843
rect 12689 6809 12724 6843
rect 12758 6809 12793 6843
rect 12827 6809 12862 6843
rect 12896 6809 12931 6843
rect 12965 6809 13000 6843
rect 13034 6809 13069 6843
rect 13103 6809 13138 6843
rect 13172 6809 13207 6843
rect 13241 6809 13276 6843
rect 13310 6809 13345 6843
rect 13379 6809 13414 6843
rect 13448 6809 13483 6843
rect 13517 6809 13552 6843
rect 13586 6809 13621 6843
rect 13655 6809 13690 6843
rect 13724 6809 13759 6843
rect 13793 6809 13828 6843
rect 13862 6809 13897 6843
rect 13931 6809 13966 6843
rect 14000 6809 14035 6843
rect 14069 6809 14104 6843
rect 14138 6809 14173 6843
rect 14207 6809 14242 6843
rect 14276 6809 14311 6843
rect 14345 6809 14380 6843
rect 14414 6809 14449 6843
rect 14483 6809 14518 6843
rect 14552 6809 14587 6843
rect 14621 6809 14655 6843
rect 14689 6809 14723 6843
rect 14757 6809 14791 6843
rect 14825 6809 14859 6843
rect 14893 6825 15117 6843
rect 14893 6809 15068 6825
rect 12493 6805 15068 6809
rect 12493 6771 14932 6805
rect 14966 6771 15000 6805
rect 15034 6771 15068 6805
rect 15102 6771 15117 6825
rect 12493 6756 15117 6771
rect 44 6669 7108 6722
rect 44 6635 68 6669
rect 102 6635 137 6669
rect 171 6635 206 6669
rect 240 6635 275 6669
rect 309 6635 344 6669
rect 378 6635 413 6669
rect 447 6635 482 6669
rect 516 6635 551 6669
rect 585 6635 620 6669
rect 654 6635 689 6669
rect 723 6635 758 6669
rect 792 6635 827 6669
rect 861 6635 896 6669
rect 930 6635 965 6669
rect 999 6635 1034 6669
rect 1068 6635 1103 6669
rect 1137 6635 1172 6669
rect 1206 6635 1241 6669
rect 1275 6635 1310 6669
rect 1344 6635 1379 6669
rect 1413 6635 1448 6669
rect 1482 6635 1517 6669
rect 1551 6635 1586 6669
rect 1620 6635 1655 6669
rect 1689 6635 1724 6669
rect 1758 6635 1793 6669
rect 1827 6635 1862 6669
rect 1896 6635 1931 6669
rect 1965 6635 2000 6669
rect 2034 6635 2069 6669
rect 2103 6635 2138 6669
rect 2172 6635 2207 6669
rect 2241 6635 2276 6669
rect 2310 6635 2345 6669
rect 2379 6635 2414 6669
rect 2448 6635 2483 6669
rect 2517 6635 2552 6669
rect 2586 6635 2621 6669
rect 2655 6635 2690 6669
rect 2724 6635 2759 6669
rect 2793 6635 2828 6669
rect 2862 6635 2897 6669
rect 2931 6635 2966 6669
rect 3000 6635 3035 6669
rect 3069 6635 3104 6669
rect 3138 6635 3173 6669
rect 3207 6635 3242 6669
rect 3276 6635 3310 6669
rect 3344 6635 3378 6669
rect 3412 6635 3446 6669
rect 3480 6635 3514 6669
rect 3548 6635 3582 6669
rect 3616 6635 3650 6669
rect 3684 6635 3718 6669
rect 3752 6635 3786 6669
rect 3820 6635 3854 6669
rect 3888 6635 3922 6669
rect 3956 6635 3990 6669
rect 4024 6635 4058 6669
rect 4092 6635 4126 6669
rect 4160 6635 4194 6669
rect 4228 6635 4262 6669
rect 4296 6635 4330 6669
rect 4364 6635 4398 6669
rect 4432 6635 4466 6669
rect 4500 6635 4534 6669
rect 4568 6635 4602 6669
rect 4636 6635 4670 6669
rect 4704 6635 4738 6669
rect 4772 6635 4806 6669
rect 4840 6635 4874 6669
rect 4908 6635 4942 6669
rect 4976 6635 5010 6669
rect 5044 6635 5078 6669
rect 5112 6635 5146 6669
rect 5180 6635 5214 6669
rect 5248 6635 5282 6669
rect 5316 6635 5350 6669
rect 5384 6635 5418 6669
rect 5452 6635 5486 6669
rect 5520 6635 5554 6669
rect 5588 6635 5622 6669
rect 5656 6635 5690 6669
rect 5724 6635 5758 6669
rect 5792 6635 5826 6669
rect 5860 6635 5894 6669
rect 5928 6635 5962 6669
rect 5996 6635 6030 6669
rect 6064 6635 6098 6669
rect 6132 6635 6166 6669
rect 6200 6635 6234 6669
rect 6268 6635 6302 6669
rect 6336 6635 6370 6669
rect 6404 6635 6438 6669
rect 6472 6635 6506 6669
rect 6540 6635 6574 6669
rect 6608 6635 6642 6669
rect 6676 6635 6710 6669
rect 6744 6635 6778 6669
rect 6812 6635 6846 6669
rect 6880 6635 6914 6669
rect 6948 6635 6982 6669
rect 7016 6635 7050 6669
rect 7084 6635 7108 6669
rect 12493 6722 12517 6756
rect 12551 6722 12586 6756
rect 12620 6722 12655 6756
rect 12689 6722 12724 6756
rect 12758 6722 12793 6756
rect 12827 6722 12862 6756
rect 12896 6722 12931 6756
rect 12965 6722 13000 6756
rect 13034 6722 13069 6756
rect 13103 6722 13138 6756
rect 13172 6722 13207 6756
rect 13241 6722 13276 6756
rect 13310 6722 13345 6756
rect 13379 6722 13414 6756
rect 13448 6722 13483 6756
rect 13517 6722 13552 6756
rect 13586 6722 13621 6756
rect 13655 6722 13690 6756
rect 13724 6722 13759 6756
rect 13793 6722 13828 6756
rect 13862 6722 13897 6756
rect 13931 6722 13966 6756
rect 14000 6722 14035 6756
rect 14069 6722 14104 6756
rect 14138 6722 14173 6756
rect 14207 6722 14242 6756
rect 14276 6722 14311 6756
rect 14345 6722 14380 6756
rect 14414 6722 14449 6756
rect 14483 6722 14518 6756
rect 14552 6722 14587 6756
rect 14621 6722 14655 6756
rect 14689 6722 14723 6756
rect 14757 6722 14791 6756
rect 14825 6722 14859 6756
rect 14893 6753 15117 6756
rect 14893 6731 15068 6753
rect 14893 6722 14932 6731
rect 12493 6697 14932 6722
rect 14966 6697 15000 6731
rect 15034 6697 15068 6731
rect 15102 6697 15117 6753
rect 12493 6681 15117 6697
rect 12493 6669 15068 6681
rect 12493 6635 12517 6669
rect 12551 6635 12586 6669
rect 12620 6635 12655 6669
rect 12689 6635 12724 6669
rect 12758 6635 12793 6669
rect 12827 6635 12862 6669
rect 12896 6635 12931 6669
rect 12965 6635 13000 6669
rect 13034 6635 13069 6669
rect 13103 6635 13138 6669
rect 13172 6635 13207 6669
rect 13241 6635 13276 6669
rect 13310 6635 13345 6669
rect 13379 6635 13414 6669
rect 13448 6635 13483 6669
rect 13517 6635 13552 6669
rect 13586 6635 13621 6669
rect 13655 6635 13690 6669
rect 13724 6635 13759 6669
rect 13793 6635 13828 6669
rect 13862 6635 13897 6669
rect 13931 6635 13966 6669
rect 14000 6635 14035 6669
rect 14069 6635 14104 6669
rect 14138 6635 14173 6669
rect 14207 6635 14242 6669
rect 14276 6635 14311 6669
rect 14345 6635 14380 6669
rect 14414 6635 14449 6669
rect 14483 6635 14518 6669
rect 14552 6635 14587 6669
rect 14621 6635 14655 6669
rect 14689 6635 14723 6669
rect 14757 6635 14791 6669
rect 14825 6635 14859 6669
rect 14893 6657 15068 6669
rect 14893 6635 14932 6657
rect 44 6623 14932 6635
rect 14966 6623 15000 6657
rect 15034 6623 15068 6657
rect 15102 6623 15117 6681
rect 44 6609 15117 6623
rect 44 6583 15068 6609
rect 44 6582 14932 6583
rect 44 6548 68 6582
rect 102 6548 137 6582
rect 171 6548 206 6582
rect 240 6548 275 6582
rect 309 6548 344 6582
rect 378 6548 413 6582
rect 447 6548 482 6582
rect 516 6548 551 6582
rect 585 6548 620 6582
rect 654 6548 689 6582
rect 723 6548 758 6582
rect 792 6548 827 6582
rect 861 6548 896 6582
rect 930 6548 965 6582
rect 999 6548 1034 6582
rect 1068 6548 1103 6582
rect 1137 6548 1172 6582
rect 1206 6548 1241 6582
rect 1275 6548 1310 6582
rect 1344 6548 1379 6582
rect 1413 6548 1448 6582
rect 1482 6548 1517 6582
rect 1551 6548 1586 6582
rect 1620 6548 1655 6582
rect 1689 6548 1724 6582
rect 1758 6548 1793 6582
rect 1827 6548 1862 6582
rect 1896 6548 1931 6582
rect 1965 6548 2000 6582
rect 2034 6548 2069 6582
rect 2103 6548 2138 6582
rect 2172 6548 2207 6582
rect 2241 6548 2276 6582
rect 2310 6548 2345 6582
rect 2379 6548 2414 6582
rect 2448 6548 2483 6582
rect 2517 6548 2551 6582
rect 2585 6548 2619 6582
rect 2653 6548 2687 6582
rect 2721 6548 2755 6582
rect 2789 6548 2823 6582
rect 2857 6548 2891 6582
rect 2925 6548 2959 6582
rect 2993 6548 3027 6582
rect 3061 6548 3095 6582
rect 3129 6548 3163 6582
rect 3197 6548 3231 6582
rect 3265 6548 3299 6582
rect 3333 6548 3367 6582
rect 3401 6548 3435 6582
rect 3469 6548 3503 6582
rect 3537 6548 3571 6582
rect 3605 6548 3639 6582
rect 3673 6548 3707 6582
rect 3741 6548 3775 6582
rect 3809 6548 3843 6582
rect 3877 6548 3911 6582
rect 3945 6548 3979 6582
rect 4013 6548 4047 6582
rect 4081 6548 4115 6582
rect 4149 6548 4183 6582
rect 4217 6548 4251 6582
rect 4285 6548 4319 6582
rect 4353 6548 4387 6582
rect 4421 6548 4455 6582
rect 4489 6548 4523 6582
rect 4557 6548 4591 6582
rect 4625 6548 4659 6582
rect 4693 6548 4727 6582
rect 4761 6548 4795 6582
rect 4829 6548 4863 6582
rect 4897 6548 4931 6582
rect 4965 6548 4999 6582
rect 5033 6548 5067 6582
rect 5101 6548 5135 6582
rect 5169 6548 5203 6582
rect 5237 6548 5271 6582
rect 5305 6548 5339 6582
rect 5373 6548 5407 6582
rect 5441 6548 5475 6582
rect 5509 6548 5543 6582
rect 5577 6548 5611 6582
rect 5645 6548 5679 6582
rect 5713 6548 5747 6582
rect 5781 6548 5815 6582
rect 5849 6548 5883 6582
rect 5917 6548 5951 6582
rect 5985 6548 6019 6582
rect 6053 6548 6087 6582
rect 6121 6548 6155 6582
rect 6189 6548 6223 6582
rect 6257 6548 6291 6582
rect 6325 6548 6359 6582
rect 6393 6548 6427 6582
rect 6461 6548 6495 6582
rect 6529 6548 6563 6582
rect 6597 6548 6631 6582
rect 6665 6548 6699 6582
rect 6733 6548 6767 6582
rect 6801 6548 6835 6582
rect 6869 6548 6903 6582
rect 6937 6548 6971 6582
rect 7005 6548 7039 6582
rect 7073 6548 7107 6582
rect 7141 6548 7175 6582
rect 7209 6548 7243 6582
rect 7277 6548 7311 6582
rect 7345 6548 7379 6582
rect 7413 6548 7447 6582
rect 7481 6548 7515 6582
rect 7549 6548 7583 6582
rect 7617 6548 7651 6582
rect 7685 6548 7719 6582
rect 7753 6548 7787 6582
rect 7821 6548 7855 6582
rect 7889 6548 7923 6582
rect 7957 6548 7991 6582
rect 8025 6548 8059 6582
rect 8093 6548 8127 6582
rect 8161 6548 8195 6582
rect 8229 6548 8263 6582
rect 8297 6548 8331 6582
rect 8365 6548 8399 6582
rect 8433 6548 8467 6582
rect 8501 6548 8535 6582
rect 8569 6548 8603 6582
rect 8637 6548 8671 6582
rect 8705 6548 8739 6582
rect 8773 6548 8807 6582
rect 8841 6548 8875 6582
rect 8909 6548 8943 6582
rect 8977 6548 9011 6582
rect 9045 6548 9079 6582
rect 9113 6548 9147 6582
rect 9181 6548 9215 6582
rect 9249 6548 9283 6582
rect 9317 6548 9351 6582
rect 9385 6548 9419 6582
rect 9453 6548 9487 6582
rect 9521 6548 9555 6582
rect 9589 6548 9623 6582
rect 9657 6548 9691 6582
rect 9725 6548 9759 6582
rect 9793 6548 9827 6582
rect 9861 6548 9895 6582
rect 9929 6548 9963 6582
rect 9997 6548 10031 6582
rect 10065 6548 10099 6582
rect 10133 6548 10167 6582
rect 10201 6548 10235 6582
rect 10269 6548 10303 6582
rect 10337 6548 10371 6582
rect 10405 6548 10439 6582
rect 10473 6548 10507 6582
rect 10541 6548 10575 6582
rect 10609 6548 10643 6582
rect 10677 6548 10711 6582
rect 10745 6548 10779 6582
rect 10813 6548 10847 6582
rect 10881 6548 10915 6582
rect 10949 6548 10983 6582
rect 11017 6548 11051 6582
rect 11085 6548 11119 6582
rect 11153 6548 11187 6582
rect 11221 6548 11255 6582
rect 11289 6548 11323 6582
rect 11357 6548 11391 6582
rect 11425 6548 11459 6582
rect 11493 6548 11527 6582
rect 11561 6548 11595 6582
rect 11629 6548 11663 6582
rect 11697 6548 11731 6582
rect 11765 6548 11799 6582
rect 11833 6548 11867 6582
rect 11901 6548 11935 6582
rect 11969 6548 12003 6582
rect 12037 6548 12071 6582
rect 12105 6548 12139 6582
rect 12173 6548 12207 6582
rect 12241 6548 12275 6582
rect 12309 6548 12343 6582
rect 12377 6548 12411 6582
rect 12445 6548 12479 6582
rect 12513 6548 12547 6582
rect 12581 6548 12615 6582
rect 12649 6548 12683 6582
rect 12717 6548 12751 6582
rect 12785 6548 12819 6582
rect 12853 6548 12887 6582
rect 12921 6548 12955 6582
rect 12989 6548 13023 6582
rect 13057 6548 13091 6582
rect 13125 6548 13159 6582
rect 13193 6548 13227 6582
rect 13261 6548 13295 6582
rect 13329 6548 13363 6582
rect 13397 6548 13431 6582
rect 13465 6548 13499 6582
rect 13533 6548 13567 6582
rect 13601 6548 13635 6582
rect 13669 6548 13703 6582
rect 13737 6548 13771 6582
rect 13805 6548 13839 6582
rect 13873 6548 13907 6582
rect 13941 6548 13975 6582
rect 14009 6548 14043 6582
rect 14077 6548 14111 6582
rect 14145 6548 14179 6582
rect 14213 6548 14247 6582
rect 14281 6548 14315 6582
rect 14349 6548 14383 6582
rect 14417 6548 14451 6582
rect 14485 6548 14519 6582
rect 14553 6548 14587 6582
rect 14621 6548 14655 6582
rect 14689 6548 14723 6582
rect 14757 6548 14791 6582
rect 14825 6548 14859 6582
rect 14893 6549 14932 6582
rect 14966 6549 15000 6583
rect 15034 6549 15068 6583
rect 15102 6549 15117 6609
rect 14893 6548 15117 6549
rect 44 6537 15117 6548
rect 44 6509 15068 6537
rect 44 6508 14932 6509
rect 44 6474 68 6508
rect 102 6474 137 6508
rect 171 6474 206 6508
rect 240 6474 275 6508
rect 309 6474 344 6508
rect 378 6474 413 6508
rect 447 6474 482 6508
rect 516 6474 551 6508
rect 585 6474 620 6508
rect 654 6474 689 6508
rect 723 6474 758 6508
rect 792 6474 827 6508
rect 861 6474 896 6508
rect 930 6474 965 6508
rect 999 6474 1034 6508
rect 1068 6474 1103 6508
rect 1137 6474 1172 6508
rect 1206 6474 1241 6508
rect 1275 6474 1310 6508
rect 1344 6474 1379 6508
rect 1413 6474 1448 6508
rect 1482 6474 1517 6508
rect 1551 6474 1586 6508
rect 1620 6474 1655 6508
rect 1689 6474 1724 6508
rect 1758 6474 1793 6508
rect 1827 6474 1862 6508
rect 1896 6474 1931 6508
rect 1965 6474 2000 6508
rect 2034 6474 2069 6508
rect 2103 6474 2138 6508
rect 2172 6474 2207 6508
rect 2241 6474 2276 6508
rect 2310 6474 2345 6508
rect 2379 6474 2414 6508
rect 2448 6474 2483 6508
rect 2517 6474 2551 6508
rect 2585 6474 2619 6508
rect 2653 6474 2687 6508
rect 2721 6474 2755 6508
rect 2789 6474 2823 6508
rect 2857 6474 2891 6508
rect 2925 6474 2959 6508
rect 2993 6474 3027 6508
rect 3061 6474 3095 6508
rect 3129 6474 3163 6508
rect 3197 6474 3231 6508
rect 3265 6474 3299 6508
rect 3333 6474 3367 6508
rect 3401 6474 3435 6508
rect 3469 6474 3503 6508
rect 3537 6474 3571 6508
rect 3605 6474 3639 6508
rect 3673 6474 3707 6508
rect 3741 6474 3775 6508
rect 3809 6474 3843 6508
rect 3877 6474 3911 6508
rect 3945 6474 3979 6508
rect 4013 6474 4047 6508
rect 4081 6474 4115 6508
rect 4149 6474 4183 6508
rect 4217 6474 4251 6508
rect 4285 6474 4319 6508
rect 4353 6474 4387 6508
rect 4421 6474 4455 6508
rect 4489 6474 4523 6508
rect 4557 6474 4591 6508
rect 4625 6474 4659 6508
rect 4693 6474 4727 6508
rect 4761 6474 4795 6508
rect 4829 6474 4863 6508
rect 4897 6474 4931 6508
rect 4965 6474 4999 6508
rect 5033 6474 5067 6508
rect 5101 6474 5135 6508
rect 5169 6474 5203 6508
rect 5237 6474 5271 6508
rect 5305 6474 5339 6508
rect 5373 6474 5407 6508
rect 5441 6474 5475 6508
rect 5509 6474 5543 6508
rect 5577 6474 5611 6508
rect 5645 6474 5679 6508
rect 5713 6474 5747 6508
rect 5781 6474 5815 6508
rect 5849 6474 5883 6508
rect 5917 6474 5951 6508
rect 5985 6474 6019 6508
rect 6053 6474 6087 6508
rect 6121 6474 6155 6508
rect 6189 6474 6223 6508
rect 6257 6474 6291 6508
rect 6325 6474 6359 6508
rect 6393 6474 6427 6508
rect 6461 6474 6495 6508
rect 6529 6474 6563 6508
rect 6597 6474 6631 6508
rect 6665 6474 6699 6508
rect 6733 6474 6767 6508
rect 6801 6474 6835 6508
rect 6869 6474 6903 6508
rect 6937 6474 6971 6508
rect 7005 6474 7039 6508
rect 7073 6474 7107 6508
rect 7141 6474 7175 6508
rect 7209 6474 7243 6508
rect 7277 6474 7311 6508
rect 7345 6474 7379 6508
rect 7413 6474 7447 6508
rect 7481 6474 7515 6508
rect 7549 6474 7583 6508
rect 7617 6474 7651 6508
rect 7685 6474 7719 6508
rect 7753 6474 7787 6508
rect 7821 6474 7855 6508
rect 7889 6474 7923 6508
rect 7957 6474 7991 6508
rect 8025 6474 8059 6508
rect 8093 6474 8127 6508
rect 8161 6474 8195 6508
rect 8229 6474 8263 6508
rect 8297 6474 8331 6508
rect 8365 6474 8399 6508
rect 8433 6474 8467 6508
rect 8501 6474 8535 6508
rect 8569 6474 8603 6508
rect 8637 6474 8671 6508
rect 8705 6474 8739 6508
rect 8773 6474 8807 6508
rect 8841 6474 8875 6508
rect 8909 6474 8943 6508
rect 8977 6474 9011 6508
rect 9045 6474 9079 6508
rect 9113 6474 9147 6508
rect 9181 6474 9215 6508
rect 9249 6474 9283 6508
rect 9317 6474 9351 6508
rect 9385 6474 9419 6508
rect 9453 6474 9487 6508
rect 9521 6474 9555 6508
rect 9589 6474 9623 6508
rect 9657 6474 9691 6508
rect 9725 6474 9759 6508
rect 9793 6474 9827 6508
rect 9861 6474 9895 6508
rect 9929 6474 9963 6508
rect 9997 6474 10031 6508
rect 10065 6474 10099 6508
rect 10133 6474 10167 6508
rect 10201 6474 10235 6508
rect 10269 6474 10303 6508
rect 10337 6474 10371 6508
rect 10405 6474 10439 6508
rect 10473 6474 10507 6508
rect 10541 6474 10575 6508
rect 10609 6474 10643 6508
rect 10677 6474 10711 6508
rect 10745 6474 10779 6508
rect 10813 6474 10847 6508
rect 10881 6474 10915 6508
rect 10949 6474 10983 6508
rect 11017 6474 11051 6508
rect 11085 6474 11119 6508
rect 11153 6474 11187 6508
rect 11221 6474 11255 6508
rect 11289 6474 11323 6508
rect 11357 6474 11391 6508
rect 11425 6474 11459 6508
rect 11493 6474 11527 6508
rect 11561 6474 11595 6508
rect 11629 6474 11663 6508
rect 11697 6474 11731 6508
rect 11765 6474 11799 6508
rect 11833 6474 11867 6508
rect 11901 6474 11935 6508
rect 11969 6474 12003 6508
rect 12037 6474 12071 6508
rect 12105 6474 12139 6508
rect 12173 6474 12207 6508
rect 12241 6474 12275 6508
rect 12309 6474 12343 6508
rect 12377 6474 12411 6508
rect 12445 6474 12479 6508
rect 12513 6474 12547 6508
rect 12581 6474 12615 6508
rect 12649 6474 12683 6508
rect 12717 6474 12751 6508
rect 12785 6474 12819 6508
rect 12853 6474 12887 6508
rect 12921 6474 12955 6508
rect 12989 6474 13023 6508
rect 13057 6474 13091 6508
rect 13125 6474 13159 6508
rect 13193 6474 13227 6508
rect 13261 6474 13295 6508
rect 13329 6474 13363 6508
rect 13397 6474 13431 6508
rect 13465 6474 13499 6508
rect 13533 6474 13567 6508
rect 13601 6474 13635 6508
rect 13669 6474 13703 6508
rect 13737 6474 13771 6508
rect 13805 6474 13839 6508
rect 13873 6474 13907 6508
rect 13941 6474 13975 6508
rect 14009 6474 14043 6508
rect 14077 6474 14111 6508
rect 14145 6474 14179 6508
rect 14213 6474 14247 6508
rect 14281 6474 14315 6508
rect 14349 6474 14383 6508
rect 14417 6474 14451 6508
rect 14485 6474 14519 6508
rect 14553 6474 14587 6508
rect 14621 6474 14655 6508
rect 14689 6474 14723 6508
rect 14757 6474 14791 6508
rect 14825 6474 14859 6508
rect 14893 6475 14932 6508
rect 14966 6475 15000 6509
rect 15034 6475 15068 6509
rect 15102 6475 15117 6537
rect 14893 6474 15117 6475
rect 44 6465 15117 6474
rect 44 6439 15068 6465
rect 44 6400 68 6439
rect 102 6434 141 6439
rect 175 6434 214 6439
rect 248 6434 287 6439
rect 321 6434 360 6439
rect 394 6434 433 6439
rect 467 6434 506 6439
rect 540 6434 579 6439
rect 613 6434 652 6439
rect 686 6434 725 6439
rect 759 6434 798 6439
rect 832 6434 871 6439
rect 905 6434 944 6439
rect 978 6434 1017 6439
rect 1051 6434 1090 6439
rect 15020 6435 15068 6439
rect 102 6400 137 6434
rect 175 6405 206 6434
rect 248 6405 275 6434
rect 321 6405 344 6434
rect 394 6405 413 6434
rect 467 6405 482 6434
rect 540 6405 551 6434
rect 613 6405 620 6434
rect 686 6405 689 6434
rect 171 6400 206 6405
rect 240 6400 275 6405
rect 309 6400 344 6405
rect 378 6400 413 6405
rect 447 6400 482 6405
rect 516 6400 551 6405
rect 585 6400 620 6405
rect 654 6400 689 6405
rect 723 6405 725 6434
rect 792 6405 798 6434
rect 861 6405 871 6434
rect 930 6405 944 6434
rect 999 6405 1017 6434
rect 723 6400 758 6405
rect 792 6400 827 6405
rect 861 6400 896 6405
rect 930 6400 965 6405
rect 999 6400 1034 6405
rect 1068 6400 1090 6434
rect 15034 6401 15068 6435
rect 15102 6401 15117 6465
rect 44 6367 1090 6400
rect 44 6326 68 6367
rect 102 6360 141 6367
rect 175 6360 214 6367
rect 248 6360 287 6367
rect 321 6360 360 6367
rect 394 6360 433 6367
rect 467 6360 506 6367
rect 540 6360 579 6367
rect 613 6360 652 6367
rect 686 6360 725 6367
rect 759 6360 798 6367
rect 832 6360 871 6367
rect 905 6360 944 6367
rect 978 6360 1017 6367
rect 1051 6360 1090 6367
rect 15020 6393 15117 6401
rect 15020 6360 15068 6393
rect 102 6326 137 6360
rect 175 6333 206 6360
rect 248 6333 275 6360
rect 321 6333 344 6360
rect 394 6333 413 6360
rect 467 6333 482 6360
rect 540 6333 551 6360
rect 613 6333 620 6360
rect 686 6333 689 6360
rect 171 6326 206 6333
rect 240 6326 275 6333
rect 309 6326 344 6333
rect 378 6326 413 6333
rect 447 6326 482 6333
rect 516 6326 551 6333
rect 585 6326 620 6333
rect 654 6326 689 6333
rect 723 6333 725 6360
rect 792 6333 798 6360
rect 861 6333 871 6360
rect 930 6333 944 6360
rect 999 6333 1017 6360
rect 723 6326 758 6333
rect 792 6326 827 6333
rect 861 6326 896 6333
rect 930 6326 965 6333
rect 999 6326 1034 6333
rect 1068 6326 1090 6360
rect 15034 6326 15068 6360
rect 15102 6326 15117 6393
rect 44 6295 1090 6326
rect 44 6252 68 6295
rect 102 6286 141 6295
rect 175 6286 214 6295
rect 248 6286 287 6295
rect 321 6286 360 6295
rect 394 6286 433 6295
rect 467 6286 506 6295
rect 540 6286 579 6295
rect 613 6286 652 6295
rect 686 6286 725 6295
rect 759 6286 798 6295
rect 832 6286 871 6295
rect 905 6286 944 6295
rect 978 6286 1017 6295
rect 1051 6286 1090 6295
rect 15020 6321 15117 6326
rect 15020 6287 15068 6321
rect 15102 6287 15117 6321
rect 102 6252 137 6286
rect 175 6261 206 6286
rect 248 6261 275 6286
rect 321 6261 344 6286
rect 394 6261 413 6286
rect 467 6261 482 6286
rect 540 6261 551 6286
rect 613 6261 620 6286
rect 686 6261 689 6286
rect 171 6252 206 6261
rect 240 6252 275 6261
rect 309 6252 344 6261
rect 378 6252 413 6261
rect 447 6252 482 6261
rect 516 6252 551 6261
rect 585 6252 620 6261
rect 654 6252 689 6261
rect 723 6261 725 6286
rect 792 6261 798 6286
rect 861 6261 871 6286
rect 930 6261 944 6286
rect 999 6261 1017 6286
rect 723 6252 758 6261
rect 792 6252 827 6261
rect 861 6252 896 6261
rect 930 6252 965 6261
rect 999 6252 1034 6261
rect 1068 6252 1090 6286
rect 15020 6285 15117 6287
rect 44 6223 1090 6252
rect 15034 6251 15068 6285
rect 15102 6251 15117 6285
rect 44 6178 68 6223
rect 102 6212 141 6223
rect 175 6212 214 6223
rect 248 6212 287 6223
rect 321 6212 360 6223
rect 394 6212 433 6223
rect 467 6212 506 6223
rect 540 6212 579 6223
rect 613 6212 652 6223
rect 686 6212 725 6223
rect 759 6212 798 6223
rect 832 6212 871 6223
rect 905 6212 944 6223
rect 978 6212 1017 6223
rect 1051 6212 1090 6223
rect 15020 6249 15117 6251
rect 15020 6215 15068 6249
rect 15102 6215 15117 6249
rect 102 6178 137 6212
rect 175 6189 206 6212
rect 248 6189 275 6212
rect 321 6189 344 6212
rect 394 6189 413 6212
rect 467 6189 482 6212
rect 540 6189 551 6212
rect 613 6189 620 6212
rect 686 6189 689 6212
rect 171 6178 206 6189
rect 240 6178 275 6189
rect 309 6178 344 6189
rect 378 6178 413 6189
rect 447 6178 482 6189
rect 516 6178 551 6189
rect 585 6178 620 6189
rect 654 6178 689 6189
rect 723 6189 725 6212
rect 792 6189 798 6212
rect 861 6189 871 6212
rect 930 6189 944 6212
rect 999 6189 1017 6212
rect 723 6178 758 6189
rect 792 6178 827 6189
rect 861 6178 896 6189
rect 930 6178 965 6189
rect 999 6178 1034 6189
rect 1068 6178 1090 6212
rect 15020 6210 15117 6215
rect 44 6151 1090 6178
rect 15034 6176 15068 6210
rect 44 6104 68 6151
rect 102 6138 141 6151
rect 175 6138 214 6151
rect 248 6138 287 6151
rect 321 6138 360 6151
rect 394 6138 433 6151
rect 467 6138 506 6151
rect 540 6138 579 6151
rect 613 6138 652 6151
rect 686 6138 725 6151
rect 759 6138 798 6151
rect 832 6138 871 6151
rect 905 6138 944 6151
rect 978 6138 1017 6151
rect 1051 6138 1090 6151
rect 15020 6143 15068 6176
rect 15102 6143 15117 6210
rect 102 6104 137 6138
rect 175 6117 206 6138
rect 248 6117 275 6138
rect 321 6117 344 6138
rect 394 6117 413 6138
rect 467 6117 482 6138
rect 540 6117 551 6138
rect 613 6117 620 6138
rect 686 6117 689 6138
rect 171 6104 206 6117
rect 240 6104 275 6117
rect 309 6104 344 6117
rect 378 6104 413 6117
rect 447 6104 482 6117
rect 516 6104 551 6117
rect 585 6104 620 6117
rect 654 6104 689 6117
rect 723 6117 725 6138
rect 792 6117 798 6138
rect 861 6117 871 6138
rect 930 6117 944 6138
rect 999 6117 1017 6138
rect 1068 6117 1090 6138
rect 15020 6135 15117 6143
rect 723 6104 758 6117
rect 792 6104 827 6117
rect 861 6104 896 6117
rect 930 6104 965 6117
rect 999 6104 1034 6117
rect 1068 6104 1103 6117
rect 1137 6104 1172 6117
rect 1206 6104 1241 6117
rect 1275 6104 1310 6117
rect 1344 6104 1379 6117
rect 1413 6104 1448 6117
rect 1482 6104 1517 6117
rect 1551 6104 1586 6117
rect 1620 6104 1655 6117
rect 1689 6104 1724 6117
rect 1758 6104 1793 6117
rect 1827 6104 1862 6117
rect 1896 6104 1931 6117
rect 1965 6104 2000 6117
rect 2034 6104 2069 6117
rect 2103 6104 2138 6117
rect 2172 6104 2207 6117
rect 2241 6104 2276 6117
rect 2310 6104 2345 6117
rect 2379 6104 2414 6117
rect 2448 6104 2483 6117
rect 2517 6104 2551 6117
rect 2585 6104 2619 6117
rect 2653 6104 2687 6117
rect 2721 6104 2755 6117
rect 2789 6104 2823 6117
rect 2857 6104 2891 6117
rect 2925 6104 2959 6117
rect 2993 6104 3027 6117
rect 3061 6104 3095 6117
rect 3129 6104 3163 6117
rect 3197 6104 3231 6117
rect 3265 6104 3299 6117
rect 3333 6104 3367 6117
rect 3401 6104 3435 6117
rect 3469 6104 3503 6117
rect 3537 6104 3571 6117
rect 3605 6104 3639 6117
rect 3673 6104 3707 6117
rect 3741 6104 3775 6117
rect 3809 6104 3843 6117
rect 3877 6104 3911 6117
rect 3945 6104 3979 6117
rect 4013 6104 4047 6117
rect 4081 6104 4115 6117
rect 4149 6104 4183 6117
rect 4217 6104 4251 6117
rect 4285 6104 4319 6117
rect 4353 6104 4387 6117
rect 4421 6104 4455 6117
rect 4489 6104 4523 6117
rect 4557 6104 4591 6117
rect 4625 6104 4659 6117
rect 4693 6104 4727 6117
rect 4761 6104 4795 6117
rect 4829 6104 4863 6117
rect 4897 6104 4931 6117
rect 4965 6104 4999 6117
rect 5033 6104 5067 6117
rect 5101 6104 5135 6117
rect 5169 6104 5203 6117
rect 5237 6104 5271 6117
rect 5305 6104 5339 6117
rect 5373 6104 5407 6117
rect 5441 6104 5475 6117
rect 5509 6104 5543 6117
rect 5577 6104 5611 6117
rect 5645 6104 5679 6117
rect 5713 6104 5747 6117
rect 5781 6104 5815 6117
rect 5849 6104 5883 6117
rect 5917 6104 5951 6117
rect 5985 6104 6019 6117
rect 6053 6104 6087 6117
rect 6121 6104 6155 6117
rect 6189 6104 6223 6117
rect 6257 6104 6291 6117
rect 6325 6104 6359 6117
rect 6393 6104 6427 6117
rect 6461 6104 6495 6117
rect 6529 6104 6563 6117
rect 6597 6104 6631 6117
rect 6665 6104 6699 6117
rect 6733 6104 6767 6117
rect 6801 6104 6835 6117
rect 6869 6104 6903 6117
rect 6937 6104 6971 6117
rect 7005 6104 7039 6117
rect 7073 6104 7107 6117
rect 7141 6104 7175 6117
rect 7209 6104 7243 6117
rect 7277 6104 7311 6117
rect 7345 6104 7379 6117
rect 7413 6104 7447 6117
rect 7481 6104 7515 6117
rect 7549 6104 7583 6117
rect 7617 6104 7651 6117
rect 7685 6104 7719 6117
rect 7753 6104 7787 6117
rect 7821 6104 7855 6117
rect 7889 6104 7923 6117
rect 7957 6104 7991 6117
rect 8025 6104 8059 6117
rect 8093 6104 8127 6117
rect 8161 6104 8195 6117
rect 8229 6104 8263 6117
rect 8297 6104 8331 6117
rect 8365 6104 8399 6117
rect 8433 6104 8467 6117
rect 8501 6104 8535 6117
rect 8569 6104 8603 6117
rect 8637 6104 8671 6117
rect 8705 6104 8739 6117
rect 8773 6104 8807 6117
rect 8841 6104 8875 6117
rect 8909 6104 8943 6117
rect 8977 6104 9011 6117
rect 9045 6104 9079 6117
rect 9113 6104 9147 6117
rect 9181 6104 9215 6117
rect 9249 6104 9283 6117
rect 9317 6104 9351 6117
rect 9385 6104 9419 6117
rect 9453 6104 9487 6117
rect 9521 6104 9555 6117
rect 9589 6104 9623 6117
rect 9657 6104 9691 6117
rect 9725 6104 9759 6117
rect 9793 6104 9827 6117
rect 9861 6104 9895 6117
rect 9929 6104 9963 6117
rect 9997 6104 10031 6117
rect 10065 6104 10099 6117
rect 10133 6104 10167 6117
rect 10201 6104 10235 6117
rect 10269 6104 10303 6117
rect 10337 6104 10371 6117
rect 10405 6104 10439 6117
rect 10473 6104 10507 6117
rect 10541 6104 10575 6117
rect 10609 6104 10643 6117
rect 10677 6104 10711 6117
rect 10745 6104 10779 6117
rect 10813 6104 10847 6117
rect 10881 6104 10915 6117
rect 10949 6104 10983 6117
rect 11017 6104 11051 6117
rect 11085 6104 11119 6117
rect 11153 6104 11187 6117
rect 11221 6104 11255 6117
rect 11289 6104 11323 6117
rect 11357 6104 11391 6117
rect 11425 6104 11459 6117
rect 11493 6104 11527 6117
rect 11561 6104 11595 6117
rect 11629 6104 11663 6117
rect 11697 6104 11731 6117
rect 11765 6104 11799 6117
rect 11833 6104 11867 6117
rect 11901 6104 11935 6117
rect 11969 6104 12003 6117
rect 12037 6104 12071 6117
rect 12105 6104 12139 6117
rect 12173 6104 12207 6117
rect 12241 6104 12275 6117
rect 12309 6104 12343 6117
rect 12377 6104 12411 6117
rect 12445 6104 12479 6117
rect 12513 6104 12547 6117
rect 12581 6104 12615 6117
rect 12649 6104 12683 6117
rect 12717 6104 12751 6117
rect 12785 6104 12819 6117
rect 12853 6104 12887 6117
rect 12921 6104 12955 6117
rect 12989 6104 13023 6117
rect 13057 6104 13091 6117
rect 13125 6104 13159 6117
rect 13193 6104 13227 6117
rect 13261 6104 13295 6117
rect 13329 6104 13363 6117
rect 13397 6104 13431 6117
rect 13465 6104 13499 6117
rect 13533 6104 13567 6117
rect 13601 6104 13635 6117
rect 13669 6104 13703 6117
rect 13737 6104 13771 6117
rect 13805 6104 13839 6117
rect 13873 6104 13907 6117
rect 13941 6104 13975 6117
rect 14009 6104 14043 6117
rect 14077 6104 14111 6117
rect 14145 6104 14179 6117
rect 14213 6104 14247 6117
rect 14281 6104 14315 6117
rect 14349 6104 14383 6117
rect 14417 6104 14451 6117
rect 14485 6104 14519 6117
rect 14553 6104 14587 6117
rect 14621 6104 14655 6117
rect 14689 6104 14723 6117
rect 14757 6104 14791 6117
rect 14825 6104 14859 6117
rect 14893 6104 14932 6117
rect 44 6101 14932 6104
rect 14966 6101 15000 6117
rect 15034 6101 15068 6135
rect 44 6071 15068 6101
rect 15102 6071 15117 6135
rect 44 6060 15117 6071
rect 44 6051 14932 6060
rect 14917 6026 14932 6051
rect 14966 6026 15000 6060
rect 15034 6026 15068 6060
rect 14917 5999 15068 6026
rect 15102 5999 15117 6060
rect 14917 5988 15117 5999
rect 14977 5961 15117 5988
rect 14977 5954 15068 5961
rect 14977 4628 15000 5954
rect 15102 4628 15117 5961
rect 14977 4593 15117 4628
rect 14977 4559 15000 4593
rect 15034 4559 15068 4593
rect 15102 4559 15117 4593
rect 14977 4524 15117 4559
rect 14977 4490 15000 4524
rect 15034 4490 15068 4524
rect 14977 4487 15068 4490
rect 15102 4487 15117 4524
rect 14977 4455 15117 4487
rect 14977 4421 15000 4455
rect 15034 4421 15068 4455
rect 14977 4415 15068 4421
rect 15102 4415 15117 4455
rect 14977 4386 15117 4415
rect 14977 4352 15000 4386
rect 15034 4352 15068 4386
rect 14977 4343 15068 4352
rect 15102 4343 15117 4386
rect 14977 4317 15117 4343
rect 14977 4283 15000 4317
rect 15034 4283 15068 4317
rect 14977 4271 15068 4283
rect 15102 4271 15117 4317
rect 14977 4248 15117 4271
rect 14977 4214 15000 4248
rect 15034 4214 15068 4248
rect 14977 4199 15068 4214
rect 15102 4199 15117 4248
rect 14977 4179 15117 4199
rect 14977 4145 15000 4179
rect 15034 4145 15068 4179
rect 14977 4127 15068 4145
rect 15102 4127 15117 4179
rect 14977 4110 15117 4127
rect 14977 4076 15000 4110
rect 15034 4076 15068 4110
rect 14977 4055 15068 4076
rect 15102 4055 15117 4110
rect 14977 4041 15117 4055
rect 14977 4007 15000 4041
rect 15034 4007 15068 4041
rect 14977 3983 15068 4007
rect 15102 3983 15117 4041
rect 14977 3972 15117 3983
rect 14977 3938 15000 3972
rect 15034 3938 15068 3972
rect 14977 3911 15068 3938
rect 15102 3911 15117 3972
rect 14977 3903 15117 3911
rect 14977 3869 15000 3903
rect 15034 3869 15068 3903
rect 14977 3839 15068 3869
rect 15102 3839 15117 3903
rect 14977 3834 15117 3839
rect 14977 3800 15000 3834
rect 15034 3800 15068 3834
rect 14977 3767 15068 3800
rect 15102 3767 15117 3834
rect 14977 3765 15117 3767
rect 14977 3731 15000 3765
rect 15034 3731 15068 3765
rect 15102 3731 15117 3765
rect 14977 3729 15117 3731
rect 14977 3696 15068 3729
rect 14977 3662 15000 3696
rect 15034 3662 15068 3696
rect 15102 3662 15117 3729
rect 14977 3657 15117 3662
rect 14977 3627 15068 3657
rect 14977 3593 15000 3627
rect 15034 3593 15068 3627
rect 15102 3593 15117 3657
rect 14977 3585 15117 3593
rect 14977 3558 15068 3585
rect 14977 3524 15000 3558
rect 15034 3524 15068 3558
rect 15102 3524 15117 3585
rect 14977 3513 15117 3524
rect 14977 3489 15068 3513
rect 14977 3455 15000 3489
rect 15034 3455 15068 3489
rect 15102 3455 15117 3513
rect 14977 3441 15117 3455
rect 14977 3420 15068 3441
rect 14977 3386 15000 3420
rect 15034 3386 15068 3420
rect 15102 3386 15117 3441
rect 14977 3369 15117 3386
rect 14977 3351 15068 3369
rect 14977 3317 15000 3351
rect 15034 3317 15068 3351
rect 15102 3317 15117 3369
rect 14977 3297 15117 3317
rect 14977 3282 15068 3297
rect 14977 3248 15000 3282
rect 15034 3248 15068 3282
rect 15102 3248 15117 3297
rect 14977 3225 15117 3248
rect 14977 3213 15068 3225
rect 14977 3179 15000 3213
rect 15034 3179 15068 3213
rect 15102 3179 15117 3225
rect 14977 3153 15117 3179
rect 14977 3144 15068 3153
rect 14977 3110 15000 3144
rect 15034 3110 15068 3144
rect 15102 3110 15117 3153
rect 14977 3081 15117 3110
rect 14977 3075 15068 3081
rect 14977 3041 15000 3075
rect 15034 3041 15068 3075
rect 15102 3041 15117 3081
rect 14977 3009 15117 3041
rect 14977 3006 15068 3009
rect 14977 2972 15000 3006
rect 15034 2972 15068 3006
rect 15102 2972 15117 3009
rect 14977 2937 15117 2972
rect 14977 2903 15000 2937
rect 15034 2903 15068 2937
rect 15102 2903 15117 2937
rect 14977 2868 15117 2903
rect 14977 2834 15000 2868
rect 15034 2834 15068 2868
rect 14977 2831 15068 2834
rect 15102 2831 15117 2868
rect 14977 2799 15117 2831
rect 14977 2765 15000 2799
rect 15034 2765 15068 2799
rect 14977 2759 15068 2765
rect 15102 2759 15117 2799
rect 14977 2730 15117 2759
rect 14977 2696 15000 2730
rect 15034 2696 15068 2730
rect 14977 2687 15068 2696
rect 15102 2687 15117 2730
rect 14977 2661 15117 2687
rect 14977 2627 15000 2661
rect 15034 2627 15068 2661
rect 14977 2615 15068 2627
rect 15102 2615 15117 2661
rect 14977 2592 15117 2615
rect 14977 2558 15000 2592
rect 15034 2558 15068 2592
rect 14977 2543 15068 2558
rect 15102 2543 15117 2592
rect 14977 2523 15117 2543
rect 14977 2489 15000 2523
rect 15034 2489 15068 2523
rect 14977 2471 15068 2489
rect 15102 2471 15117 2523
rect 14977 2454 15117 2471
rect 14977 2420 15000 2454
rect 15034 2420 15068 2454
rect 14977 2399 15068 2420
rect 15102 2399 15117 2454
rect 14977 2385 15117 2399
rect 14977 2351 15000 2385
rect 15034 2351 15068 2385
rect 14977 2327 15068 2351
rect 15102 2327 15117 2385
rect 14977 2316 15117 2327
rect 14977 2282 15000 2316
rect 15034 2282 15068 2316
rect 14977 2255 15068 2282
rect 15102 2255 15117 2316
rect 14977 2247 15117 2255
rect 14977 2213 15000 2247
rect 15034 2213 15068 2247
rect 14977 2183 15068 2213
rect 15102 2183 15117 2247
rect 14977 2178 15117 2183
rect 14977 2144 15000 2178
rect 15034 2144 15068 2178
rect 14977 2111 15068 2144
rect 15102 2111 15117 2178
rect 14977 2109 15117 2111
rect 14977 2075 15000 2109
rect 15034 2075 15068 2109
rect 15102 2075 15117 2109
rect 14977 2073 15117 2075
rect 14977 2040 15068 2073
rect 14977 2006 15000 2040
rect 15034 2006 15068 2040
rect 15102 2006 15117 2073
rect 14977 2001 15117 2006
rect 14977 1971 15068 2001
rect 14977 1937 15000 1971
rect 15034 1937 15068 1971
rect 15102 1937 15117 2001
rect 14977 1929 15117 1937
rect 14977 1902 15068 1929
rect 14977 1868 15000 1902
rect 15034 1868 15068 1902
rect 15102 1868 15117 1929
rect 14977 1857 15117 1868
rect 14977 1833 15068 1857
rect 14977 1799 15000 1833
rect 15034 1799 15068 1833
rect 15102 1799 15117 1857
rect 14977 1785 15117 1799
rect 14977 1764 15068 1785
rect 14977 1730 15000 1764
rect 15034 1730 15068 1764
rect 15102 1730 15117 1785
rect 14977 1713 15117 1730
rect 14977 1695 15068 1713
rect 14977 1661 15000 1695
rect 15034 1661 15068 1695
rect 15102 1661 15117 1713
rect 14977 1641 15117 1661
rect 14977 1626 15068 1641
rect 14977 1592 15000 1626
rect 15034 1592 15068 1626
rect 15102 1592 15117 1641
rect 14977 1569 15117 1592
rect 14977 1557 15068 1569
rect 14977 1523 15000 1557
rect 15034 1523 15068 1557
rect 15102 1523 15117 1569
rect 14977 1497 15117 1523
rect 14977 1488 15068 1497
rect 14977 1454 15000 1488
rect 15034 1454 15068 1488
rect 15102 1454 15117 1497
rect 14977 1425 15117 1454
rect 14977 1419 15068 1425
rect 14977 1385 15000 1419
rect 15034 1385 15068 1419
rect 15102 1385 15117 1425
rect 310 1322 402 1368
rect 14977 1353 15117 1385
rect 14977 1350 15068 1353
rect 14977 1316 15000 1350
rect 15034 1316 15068 1350
rect 15102 1316 15117 1353
rect 7044 1282 14917 1288
rect 14977 1282 15117 1316
rect 68 1281 15117 1282
rect 68 1257 15068 1281
rect 68 1251 7068 1257
rect 3537 1217 3565 1251
rect 3611 1217 3637 1251
rect 3679 1217 3709 1251
rect 3747 1217 3781 1251
rect 3815 1217 3849 1251
rect 3887 1217 3917 1251
rect 3959 1217 3985 1251
rect 4031 1217 4053 1251
rect 4103 1217 4121 1251
rect 4175 1217 4189 1251
rect 4247 1217 4257 1251
rect 4319 1217 4325 1251
rect 4391 1217 4393 1251
rect 4427 1217 4429 1251
rect 4495 1217 4501 1251
rect 4563 1217 4573 1251
rect 4631 1217 4645 1251
rect 4699 1217 4717 1251
rect 4767 1217 4789 1251
rect 4835 1217 4861 1251
rect 4903 1217 4933 1251
rect 4971 1217 5005 1251
rect 5039 1217 5073 1251
rect 5111 1217 5141 1251
rect 5183 1217 5209 1251
rect 5255 1217 5277 1251
rect 5327 1217 5345 1251
rect 5399 1217 5413 1251
rect 5471 1217 5481 1251
rect 5543 1217 5549 1251
rect 5615 1217 5617 1251
rect 5651 1217 5653 1251
rect 5719 1217 5725 1251
rect 5787 1217 5797 1251
rect 5855 1217 5869 1251
rect 5923 1217 5941 1251
rect 5991 1217 6013 1251
rect 6059 1217 6085 1251
rect 6127 1217 6157 1251
rect 6195 1217 6229 1251
rect 6263 1217 6297 1251
rect 6335 1217 6365 1251
rect 6407 1217 6433 1251
rect 6479 1217 6501 1251
rect 6551 1217 6569 1251
rect 6623 1217 6637 1251
rect 6695 1217 6705 1251
rect 6767 1217 6773 1251
rect 6839 1217 6841 1251
rect 6875 1217 6877 1251
rect 6943 1239 7068 1251
rect 6943 1217 6988 1239
rect 7022 1223 7068 1239
rect 7102 1223 7137 1257
rect 7171 1223 7206 1257
rect 7240 1223 7275 1257
rect 7309 1223 7344 1257
rect 7378 1223 7413 1257
rect 7447 1223 7482 1257
rect 7516 1223 7551 1257
rect 7585 1223 7620 1257
rect 7654 1223 7689 1257
rect 7723 1223 7758 1257
rect 7792 1223 7827 1257
rect 7861 1223 7896 1257
rect 7930 1223 7965 1257
rect 7999 1223 8034 1257
rect 8068 1223 8103 1257
rect 8137 1223 8172 1257
rect 8206 1223 8241 1257
rect 8275 1223 8310 1257
rect 8344 1223 8379 1257
rect 8413 1223 8448 1257
rect 8482 1223 8517 1257
rect 8551 1223 8586 1257
rect 8620 1223 8655 1257
rect 8689 1223 8724 1257
rect 8758 1223 8793 1257
rect 8827 1223 8862 1257
rect 8896 1223 8931 1257
rect 8965 1223 9000 1257
rect 9034 1223 9069 1257
rect 9103 1223 9138 1257
rect 9172 1223 9207 1257
rect 9241 1223 9276 1257
rect 9310 1223 9345 1257
rect 9379 1223 9414 1257
rect 9448 1223 9483 1257
rect 9517 1223 9552 1257
rect 9586 1223 9621 1257
rect 9655 1223 9690 1257
rect 9724 1223 9759 1257
rect 7022 1217 9759 1223
rect 14893 1247 15068 1257
rect 15102 1247 15117 1281
rect 14893 1244 15117 1247
rect 14893 1217 14932 1244
rect 14966 1217 15000 1244
rect 7022 1193 7069 1217
rect 6988 1189 7069 1193
rect 7103 1189 7142 1217
rect 7176 1189 7215 1217
rect 7249 1189 7288 1217
rect 7322 1189 7361 1217
rect 7395 1189 7434 1217
rect 7468 1189 7507 1217
rect 7541 1189 7580 1217
rect 7614 1189 7653 1217
rect 7687 1189 7726 1217
rect 7760 1189 7799 1217
rect 7833 1189 7872 1217
rect 7906 1189 7945 1217
rect 7979 1189 8018 1217
rect 8052 1189 8091 1217
rect 8125 1189 8164 1217
rect 8198 1189 8237 1217
rect 8271 1189 8310 1217
rect 8344 1189 8383 1217
rect 8417 1189 8456 1217
rect 8490 1189 8528 1217
rect 8562 1189 8600 1217
rect 8634 1189 8672 1217
rect 8706 1189 8744 1217
rect 8778 1189 8816 1217
rect 8850 1189 8888 1217
rect 8922 1189 8960 1217
rect 8994 1189 9032 1217
rect 9066 1189 9104 1217
rect 6988 1167 7068 1189
rect 7103 1183 7137 1189
rect 7176 1183 7206 1189
rect 7249 1183 7275 1189
rect 7322 1183 7344 1189
rect 7395 1183 7413 1189
rect 7468 1183 7482 1189
rect 7541 1183 7551 1189
rect 7614 1183 7620 1189
rect 7687 1183 7689 1189
rect 7022 1155 7068 1167
rect 7102 1155 7137 1183
rect 7171 1155 7206 1183
rect 7240 1155 7275 1183
rect 7309 1155 7344 1183
rect 7378 1155 7413 1183
rect 7447 1155 7482 1183
rect 7516 1155 7551 1183
rect 7585 1155 7620 1183
rect 7654 1155 7689 1183
rect 7723 1183 7726 1189
rect 7792 1183 7799 1189
rect 7861 1183 7872 1189
rect 7930 1183 7945 1189
rect 7999 1183 8018 1189
rect 8068 1183 8091 1189
rect 8137 1183 8164 1189
rect 8206 1183 8237 1189
rect 7723 1155 7758 1183
rect 7792 1155 7827 1183
rect 7861 1155 7896 1183
rect 7930 1155 7965 1183
rect 7999 1155 8034 1183
rect 8068 1155 8103 1183
rect 8137 1155 8172 1183
rect 8206 1155 8241 1183
rect 8275 1155 8310 1189
rect 8344 1155 8379 1189
rect 8417 1183 8448 1189
rect 8490 1183 8517 1189
rect 8562 1183 8586 1189
rect 8634 1183 8655 1189
rect 8706 1183 8724 1189
rect 8778 1183 8793 1189
rect 8850 1183 8862 1189
rect 8922 1183 8931 1189
rect 8994 1183 9000 1189
rect 9066 1183 9069 1189
rect 8413 1155 8448 1183
rect 8482 1155 8517 1183
rect 8551 1155 8586 1183
rect 8620 1155 8655 1183
rect 8689 1155 8724 1183
rect 8758 1155 8793 1183
rect 8827 1155 8862 1183
rect 8896 1155 8931 1183
rect 8965 1155 9000 1183
rect 9034 1155 9069 1183
rect 9103 1183 9104 1189
rect 9138 1189 9176 1217
rect 9210 1189 9248 1217
rect 9282 1189 9320 1217
rect 9354 1189 9392 1217
rect 9426 1189 9464 1217
rect 9498 1189 9536 1217
rect 9570 1189 9608 1217
rect 9642 1189 9680 1217
rect 9714 1189 9752 1217
rect 9103 1155 9138 1183
rect 9172 1183 9176 1189
rect 9241 1183 9248 1189
rect 9310 1183 9320 1189
rect 9379 1183 9392 1189
rect 9448 1183 9464 1189
rect 9517 1183 9536 1189
rect 9586 1183 9608 1189
rect 9655 1183 9680 1189
rect 9724 1183 9752 1189
rect 14926 1210 14932 1217
rect 14998 1210 15000 1217
rect 15034 1210 15068 1244
rect 15102 1210 15117 1244
rect 14926 1183 14964 1210
rect 14998 1209 15117 1210
rect 14998 1183 15068 1209
rect 9172 1155 9207 1183
rect 9241 1155 9276 1183
rect 9310 1155 9345 1183
rect 9379 1155 9414 1183
rect 9448 1155 9483 1183
rect 9517 1155 9552 1183
rect 9586 1155 9621 1183
rect 9655 1155 9690 1183
rect 9724 1155 9759 1183
rect 7022 1139 9759 1155
rect 14893 1175 15068 1183
rect 15102 1175 15117 1209
rect 14893 1172 15117 1175
rect 14893 1139 14932 1172
rect 14966 1139 15000 1172
rect 7022 1125 7069 1139
rect 6988 1121 7069 1125
rect 7103 1121 7142 1139
rect 7176 1121 7215 1139
rect 7249 1121 7288 1139
rect 7322 1121 7361 1139
rect 7395 1121 7434 1139
rect 7468 1121 7507 1139
rect 7541 1121 7580 1139
rect 7614 1121 7653 1139
rect 7687 1121 7726 1139
rect 7760 1121 7799 1139
rect 7833 1121 7872 1139
rect 7906 1121 7945 1139
rect 7979 1121 8018 1139
rect 8052 1121 8091 1139
rect 8125 1121 8164 1139
rect 8198 1121 8237 1139
rect 8271 1121 8310 1139
rect 8344 1121 8383 1139
rect 8417 1121 8456 1139
rect 8490 1121 8528 1139
rect 8562 1121 8600 1139
rect 8634 1121 8672 1139
rect 8706 1121 8744 1139
rect 8778 1121 8816 1139
rect 8850 1121 8888 1139
rect 8922 1121 8960 1139
rect 8994 1121 9032 1139
rect 9066 1121 9104 1139
rect 6988 1095 7068 1121
rect 7103 1105 7137 1121
rect 7176 1105 7206 1121
rect 7249 1105 7275 1121
rect 7322 1105 7344 1121
rect 7395 1105 7413 1121
rect 7468 1105 7482 1121
rect 7541 1105 7551 1121
rect 7614 1105 7620 1121
rect 7687 1105 7689 1121
rect 3528 1031 3597 1065
rect 3631 1031 3666 1065
rect 3700 1031 3735 1065
rect 3769 1031 3804 1065
rect 3838 1031 3873 1065
rect 3907 1031 3942 1065
rect 3976 1031 4011 1065
rect 4045 1031 4080 1065
rect 4114 1031 4149 1065
rect 4183 1031 4218 1065
rect 4252 1031 4287 1065
rect 4321 1031 4356 1065
rect 4390 1031 4425 1065
rect 4459 1031 4494 1065
rect 4528 1031 4563 1065
rect 4597 1031 4632 1065
rect 4666 1031 4701 1065
rect 4735 1031 4770 1065
rect 4804 1031 4839 1065
rect 4873 1031 4908 1065
rect 4942 1031 4977 1065
rect 5011 1031 5046 1065
rect 5080 1031 5115 1065
rect 5149 1031 5184 1065
rect 5218 1031 5253 1065
rect 5287 1031 5322 1065
rect 5356 1031 5392 1065
rect 5426 1031 5462 1065
rect 5496 1031 5532 1065
rect 5566 1031 5602 1065
rect 5636 1031 5672 1065
rect 5706 1031 5742 1065
rect 5776 1031 5812 1065
rect 5846 1031 5882 1065
rect 5916 1031 5952 1065
rect 5986 1031 6022 1065
rect 6056 1031 6092 1065
rect 6126 1031 6162 1065
rect 6196 1031 6232 1065
rect 6266 1031 6302 1065
rect 6336 1031 6372 1065
rect 6406 1031 6442 1065
rect 6476 1031 6512 1065
rect 6546 1031 6582 1065
rect 6616 1031 6652 1065
rect 6686 1031 6722 1065
rect 6756 1031 6824 1065
rect 3528 966 6824 1031
rect 3528 949 6790 966
rect 3528 943 3722 949
rect 3562 937 3722 943
rect 3562 915 3592 937
rect 3718 915 3722 937
rect 3772 915 3794 949
rect 3840 915 3866 949
rect 3908 915 3938 949
rect 3976 915 4010 949
rect 4044 915 4078 949
rect 4116 915 4146 949
rect 4188 915 4214 949
rect 4260 915 4282 949
rect 4332 915 4350 949
rect 4404 915 4418 949
rect 4476 915 4486 949
rect 4548 915 4554 949
rect 4620 915 4622 949
rect 4656 915 4658 949
rect 4724 915 4730 949
rect 4792 915 4802 949
rect 4860 915 4874 949
rect 4928 915 4946 949
rect 4996 915 5018 949
rect 5064 915 5090 949
rect 5124 915 5252 949
rect 5302 915 5324 949
rect 5370 915 5396 949
rect 5438 915 5468 949
rect 5506 915 5540 949
rect 5574 915 5608 949
rect 5646 915 5676 949
rect 5718 915 5744 949
rect 5790 915 5812 949
rect 5862 915 5880 949
rect 5934 915 5948 949
rect 6006 915 6016 949
rect 6078 915 6084 949
rect 6150 915 6152 949
rect 6186 915 6188 949
rect 6254 915 6260 949
rect 6322 915 6332 949
rect 6390 915 6404 949
rect 6458 915 6476 949
rect 6526 915 6548 949
rect 6594 915 6620 949
rect 6654 938 6790 949
rect 3528 871 3562 909
rect 3528 799 3562 837
rect 3528 727 3562 765
rect 3528 655 3562 693
rect 3528 583 3562 621
rect 3528 511 3562 549
rect 3528 439 3562 477
rect 3528 367 3562 405
rect 3644 885 3678 901
rect 6704 888 6738 904
rect 3644 813 3678 851
rect 5174 865 5208 881
rect 5174 796 5208 831
rect 3644 741 3678 779
rect 3772 759 3794 793
rect 3840 759 3866 793
rect 3908 759 3938 793
rect 3976 759 4010 793
rect 4044 759 4078 793
rect 4116 759 4146 793
rect 4188 759 4214 793
rect 4260 759 4282 793
rect 4332 759 4350 793
rect 4404 759 4418 793
rect 4476 759 4486 793
rect 4548 759 4554 793
rect 4620 759 4622 793
rect 4656 759 4658 793
rect 4724 759 4730 793
rect 4792 759 4802 793
rect 4860 759 4874 793
rect 4928 759 4946 793
rect 4996 759 5018 793
rect 5064 759 5090 793
rect 6704 816 6738 854
rect 5174 727 5208 762
rect 5302 759 5324 793
rect 5370 759 5396 793
rect 5438 759 5468 793
rect 5506 759 5540 793
rect 5574 759 5608 793
rect 5646 759 5676 793
rect 5718 759 5744 793
rect 5790 759 5812 793
rect 5862 759 5880 793
rect 5934 759 5948 793
rect 6006 759 6016 793
rect 6078 759 6084 793
rect 6150 759 6152 793
rect 6186 759 6188 793
rect 6254 759 6260 793
rect 6322 759 6332 793
rect 6390 759 6404 793
rect 6458 759 6476 793
rect 6526 759 6548 793
rect 6594 759 6620 793
rect 6704 744 6738 782
rect 3644 680 3645 707
rect 3679 680 3717 714
rect 5149 693 5174 714
rect 5149 680 5187 693
rect 6654 680 6692 714
rect 6726 680 6738 710
rect 3644 670 3678 680
rect 5174 658 5208 680
rect 3644 599 3678 636
rect 3772 603 3794 637
rect 3840 603 3866 637
rect 3908 603 3938 637
rect 3976 603 4010 637
rect 4044 603 4078 637
rect 4116 603 4146 637
rect 4188 603 4214 637
rect 4260 603 4282 637
rect 4332 603 4350 637
rect 4404 603 4418 637
rect 4476 603 4486 637
rect 4548 603 4554 637
rect 4620 603 4622 637
rect 4656 603 4658 637
rect 4724 603 4730 637
rect 4792 603 4802 637
rect 4860 603 4874 637
rect 4928 603 4946 637
rect 4996 603 5018 637
rect 5064 603 5090 637
rect 6704 672 6738 680
rect 3644 528 3678 565
rect 3644 457 3678 494
rect 5174 590 5208 624
rect 5302 603 5324 637
rect 5370 603 5396 637
rect 5438 603 5468 637
rect 5506 603 5540 637
rect 5574 603 5608 637
rect 5646 603 5676 637
rect 5718 603 5744 637
rect 5790 603 5812 637
rect 5862 603 5880 637
rect 5934 603 5948 637
rect 6006 603 6016 637
rect 6078 603 6084 637
rect 6150 603 6152 637
rect 6186 603 6188 637
rect 6254 603 6260 637
rect 6322 603 6332 637
rect 6390 603 6404 637
rect 6458 603 6476 637
rect 6526 603 6548 637
rect 6594 603 6620 637
rect 5174 522 5208 556
rect 3772 447 3794 481
rect 3840 447 3866 481
rect 3908 447 3938 481
rect 3976 447 4010 481
rect 4044 447 4078 481
rect 4116 447 4146 481
rect 4188 447 4214 481
rect 4260 447 4282 481
rect 4332 447 4350 481
rect 4404 447 4418 481
rect 4476 447 4486 481
rect 4548 447 4554 481
rect 4620 447 4622 481
rect 4656 447 4658 481
rect 4724 447 4730 481
rect 4792 447 4802 481
rect 4860 447 4874 481
rect 4928 447 4946 481
rect 4996 447 5018 481
rect 5064 447 5090 481
rect 5174 454 5208 488
rect 6704 600 6738 638
rect 6704 528 6738 566
rect 3644 386 3678 423
rect 3644 336 3678 352
rect 5302 447 5324 481
rect 5370 447 5396 481
rect 5438 447 5468 481
rect 5506 447 5540 481
rect 5574 447 5608 481
rect 5646 447 5676 481
rect 5718 447 5744 481
rect 5790 447 5812 481
rect 5862 447 5880 481
rect 5934 447 5948 481
rect 6006 447 6016 481
rect 6078 447 6084 481
rect 6150 447 6152 481
rect 6186 447 6188 481
rect 6254 447 6260 481
rect 6322 447 6332 481
rect 6390 447 6404 481
rect 6458 447 6476 481
rect 6526 447 6548 481
rect 6594 447 6620 481
rect 6704 457 6738 494
rect 5174 386 5208 420
rect 5174 336 5208 352
rect 6704 386 6738 423
rect 6704 336 6738 352
rect 6790 869 6824 932
rect 6790 797 6824 811
rect 6790 725 6824 743
rect 6790 653 6824 675
rect 6790 581 6824 607
rect 6790 509 6824 539
rect 6790 437 6824 471
rect 6790 369 6824 403
rect 3528 294 3562 333
rect 3772 291 3794 325
rect 3840 291 3866 325
rect 3908 291 3938 325
rect 3976 291 4010 325
rect 4044 291 4078 325
rect 4116 291 4146 325
rect 4188 291 4214 325
rect 4260 291 4282 325
rect 4332 291 4350 325
rect 4404 291 4418 325
rect 4476 291 4486 325
rect 4548 291 4554 325
rect 4620 291 4622 325
rect 4656 291 4658 325
rect 4724 291 4730 325
rect 4792 291 4802 325
rect 4860 291 4874 325
rect 4928 291 4946 325
rect 4996 291 5018 325
rect 5064 291 5090 325
rect 5302 291 5324 325
rect 5370 291 5396 325
rect 5438 291 5468 325
rect 5506 291 5540 325
rect 5574 291 5608 325
rect 5646 291 5676 325
rect 5718 291 5744 325
rect 5790 291 5812 325
rect 5862 291 5880 325
rect 5934 291 5948 325
rect 6006 291 6016 325
rect 6078 291 6084 325
rect 6150 291 6152 325
rect 6186 291 6188 325
rect 6254 291 6260 325
rect 6322 291 6332 325
rect 6390 291 6404 325
rect 6458 291 6476 325
rect 6526 291 6548 325
rect 6594 291 6620 325
rect 6790 301 6824 331
rect 3528 221 3562 260
rect 6790 233 6824 259
rect 3562 187 3632 209
rect 3528 175 3632 187
rect 3666 175 3700 209
rect 3738 175 3768 209
rect 3810 175 3836 209
rect 3882 175 3904 209
rect 3954 175 3972 209
rect 4026 175 4040 209
rect 4098 175 4108 209
rect 4170 175 4176 209
rect 4242 175 4244 209
rect 4278 175 4280 209
rect 4346 175 4352 209
rect 4414 175 4424 209
rect 4482 175 4496 209
rect 4550 175 4568 209
rect 4618 175 4640 209
rect 4686 175 4712 209
rect 4754 175 4784 209
rect 4822 175 4856 209
rect 4890 175 4924 209
rect 4962 175 4992 209
rect 5034 175 5060 209
rect 5106 175 5128 209
rect 5178 175 5196 209
rect 5250 175 5264 209
rect 5322 175 5332 209
rect 5394 175 5400 209
rect 5466 175 5468 209
rect 5502 175 5504 209
rect 5570 175 5576 209
rect 5638 175 5648 209
rect 5706 175 5720 209
rect 5774 175 5792 209
rect 5842 175 5864 209
rect 5910 175 5936 209
rect 5978 175 6008 209
rect 6046 175 6080 209
rect 6114 175 6148 209
rect 6186 175 6216 209
rect 6258 175 6284 209
rect 6330 175 6352 209
rect 6402 175 6420 209
rect 6474 175 6488 209
rect 6546 175 6556 209
rect 6618 175 6624 209
rect 6690 175 6692 209
rect 6726 187 6790 209
rect 6726 175 6824 187
rect 7022 1087 7068 1095
rect 7102 1087 7137 1105
rect 7171 1087 7206 1105
rect 7240 1087 7275 1105
rect 7309 1087 7344 1105
rect 7378 1087 7413 1105
rect 7447 1087 7482 1105
rect 7516 1087 7551 1105
rect 7585 1087 7620 1105
rect 7654 1087 7689 1105
rect 7723 1105 7726 1121
rect 7792 1105 7799 1121
rect 7861 1105 7872 1121
rect 7930 1105 7945 1121
rect 7999 1105 8018 1121
rect 8068 1105 8091 1121
rect 8137 1105 8164 1121
rect 8206 1105 8237 1121
rect 7723 1087 7758 1105
rect 7792 1087 7827 1105
rect 7861 1087 7896 1105
rect 7930 1087 7965 1105
rect 7999 1087 8034 1105
rect 8068 1087 8103 1105
rect 8137 1087 8172 1105
rect 8206 1087 8241 1105
rect 8275 1087 8310 1121
rect 8344 1087 8379 1121
rect 8417 1105 8448 1121
rect 8490 1105 8517 1121
rect 8562 1105 8586 1121
rect 8634 1105 8655 1121
rect 8706 1105 8724 1121
rect 8778 1105 8793 1121
rect 8850 1105 8862 1121
rect 8922 1105 8931 1121
rect 8994 1105 9000 1121
rect 9066 1105 9069 1121
rect 8413 1087 8448 1105
rect 8482 1087 8517 1105
rect 8551 1087 8586 1105
rect 8620 1087 8655 1105
rect 8689 1087 8724 1105
rect 8758 1087 8793 1105
rect 8827 1087 8862 1105
rect 8896 1087 8931 1105
rect 8965 1087 9000 1105
rect 9034 1087 9069 1105
rect 9103 1105 9104 1121
rect 9138 1121 9176 1139
rect 9210 1121 9248 1139
rect 9282 1121 9320 1139
rect 9354 1121 9392 1139
rect 9426 1121 9464 1139
rect 9498 1121 9536 1139
rect 9570 1121 9608 1139
rect 9642 1121 9680 1139
rect 9714 1121 9752 1139
rect 9103 1087 9138 1105
rect 9172 1105 9176 1121
rect 9241 1105 9248 1121
rect 9310 1105 9320 1121
rect 9379 1105 9392 1121
rect 9448 1105 9464 1121
rect 9517 1105 9536 1121
rect 9586 1105 9608 1121
rect 9655 1105 9680 1121
rect 9724 1105 9752 1121
rect 14926 1138 14932 1139
rect 14998 1138 15000 1139
rect 15034 1138 15068 1172
rect 15102 1138 15117 1172
rect 14926 1105 14964 1138
rect 14998 1137 15117 1138
rect 14998 1105 15068 1137
rect 9172 1087 9207 1105
rect 9241 1087 9276 1105
rect 9310 1087 9345 1105
rect 9379 1087 9414 1105
rect 9448 1087 9483 1105
rect 9517 1087 9552 1105
rect 9586 1087 9621 1105
rect 9655 1087 9690 1105
rect 9724 1087 9759 1105
rect 7022 1061 9759 1087
rect 14893 1103 15068 1105
rect 15102 1103 15117 1137
rect 14893 1100 15117 1103
rect 14893 1066 14932 1100
rect 14966 1066 15000 1100
rect 15034 1066 15068 1100
rect 15102 1066 15117 1100
rect 14893 1065 15117 1066
rect 14893 1061 15068 1065
rect 7022 1057 7069 1061
rect 6988 1053 7069 1057
rect 7103 1053 7142 1061
rect 7176 1053 7215 1061
rect 7249 1053 7288 1061
rect 7322 1053 7361 1061
rect 7395 1053 7434 1061
rect 7468 1053 7507 1061
rect 7541 1053 7580 1061
rect 7614 1053 7653 1061
rect 7687 1053 7726 1061
rect 7760 1053 7799 1061
rect 7833 1053 7872 1061
rect 7906 1053 7945 1061
rect 7979 1053 8018 1061
rect 8052 1053 8091 1061
rect 8125 1053 8164 1061
rect 8198 1053 8237 1061
rect 8271 1053 8310 1061
rect 8344 1053 8383 1061
rect 8417 1053 8456 1061
rect 8490 1053 8528 1061
rect 8562 1053 8600 1061
rect 8634 1053 8672 1061
rect 8706 1053 8744 1061
rect 8778 1053 8816 1061
rect 8850 1053 8888 1061
rect 8922 1053 8960 1061
rect 8994 1053 9032 1061
rect 9066 1053 9104 1061
rect 6988 1023 7068 1053
rect 7103 1027 7137 1053
rect 7176 1027 7206 1053
rect 7249 1027 7275 1053
rect 7322 1027 7344 1053
rect 7395 1027 7413 1053
rect 7468 1027 7482 1053
rect 7541 1027 7551 1053
rect 7614 1027 7620 1053
rect 7687 1027 7689 1053
rect 7022 1019 7068 1023
rect 7102 1019 7137 1027
rect 7171 1019 7206 1027
rect 7240 1019 7275 1027
rect 7309 1019 7344 1027
rect 7378 1019 7413 1027
rect 7447 1019 7482 1027
rect 7516 1019 7551 1027
rect 7585 1019 7620 1027
rect 7654 1019 7689 1027
rect 7723 1027 7726 1053
rect 7792 1027 7799 1053
rect 7861 1027 7872 1053
rect 7930 1027 7945 1053
rect 7999 1027 8018 1053
rect 8068 1027 8091 1053
rect 8137 1027 8164 1053
rect 8206 1027 8237 1053
rect 7723 1019 7758 1027
rect 7792 1019 7827 1027
rect 7861 1019 7896 1027
rect 7930 1019 7965 1027
rect 7999 1019 8034 1027
rect 8068 1019 8103 1027
rect 8137 1019 8172 1027
rect 8206 1019 8241 1027
rect 8275 1019 8310 1053
rect 8344 1019 8379 1053
rect 8417 1027 8448 1053
rect 8490 1027 8517 1053
rect 8562 1027 8586 1053
rect 8634 1027 8655 1053
rect 8706 1027 8724 1053
rect 8778 1027 8793 1053
rect 8850 1027 8862 1053
rect 8922 1027 8931 1053
rect 8994 1027 9000 1053
rect 9066 1027 9069 1053
rect 8413 1019 8448 1027
rect 8482 1019 8517 1027
rect 8551 1019 8586 1027
rect 8620 1019 8655 1027
rect 8689 1019 8724 1027
rect 8758 1019 8793 1027
rect 8827 1019 8862 1027
rect 8896 1019 8931 1027
rect 8965 1019 9000 1027
rect 9034 1019 9069 1027
rect 9103 1027 9104 1053
rect 9138 1053 9176 1061
rect 9210 1053 9248 1061
rect 9282 1053 9320 1061
rect 9354 1053 9392 1061
rect 9426 1053 9464 1061
rect 9498 1053 9536 1061
rect 9570 1053 9608 1061
rect 9642 1053 9680 1061
rect 9714 1053 9752 1061
rect 9103 1019 9138 1027
rect 9172 1027 9176 1053
rect 9241 1027 9248 1053
rect 9310 1027 9320 1053
rect 9379 1027 9392 1053
rect 9448 1027 9464 1053
rect 9517 1027 9536 1053
rect 9586 1027 9608 1053
rect 9655 1027 9680 1053
rect 9724 1027 9752 1053
rect 14926 1028 14964 1061
rect 14998 1031 15068 1061
rect 15102 1031 15117 1065
rect 14998 1028 15117 1031
rect 14926 1027 14932 1028
rect 14998 1027 15000 1028
rect 9172 1019 9207 1027
rect 9241 1019 9276 1027
rect 9310 1019 9345 1027
rect 9379 1019 9414 1027
rect 9448 1019 9483 1027
rect 9517 1019 9552 1027
rect 9586 1019 9621 1027
rect 9655 1019 9690 1027
rect 9724 1019 9759 1027
rect 14893 1019 14932 1027
rect 7022 994 14932 1019
rect 14966 994 15000 1027
rect 15034 994 15068 1028
rect 15102 994 15117 1028
rect 7022 993 15117 994
rect 7022 989 15068 993
rect 6988 988 14576 989
rect 6988 955 7754 988
rect 7022 947 7754 955
rect 7022 917 7067 947
rect 6988 913 7067 917
rect 7101 918 7137 947
rect 7101 913 7104 918
rect 7171 913 7207 947
rect 7241 913 7277 947
rect 7311 913 7347 947
rect 7381 913 7417 947
rect 7451 913 7487 947
rect 7521 913 7557 947
rect 7591 913 7627 947
rect 7661 913 7696 947
rect 7730 913 7754 947
rect 6988 887 7104 913
rect 7022 884 7104 887
rect 7138 884 7754 913
rect 7022 875 7754 884
rect 7022 845 7067 875
rect 6988 841 7067 845
rect 7101 841 7137 875
rect 7171 841 7207 875
rect 7241 841 7277 875
rect 7311 841 7347 875
rect 7381 841 7417 875
rect 7451 841 7487 875
rect 7521 841 7557 875
rect 7591 841 7627 875
rect 7661 841 7696 875
rect 7730 841 7754 875
rect 6988 819 7754 841
rect 7022 803 7754 819
rect 7022 773 7067 803
rect 6988 769 7067 773
rect 7101 769 7137 803
rect 7171 769 7207 803
rect 7241 769 7277 803
rect 7311 769 7347 803
rect 7381 769 7417 803
rect 7451 769 7487 803
rect 7521 769 7557 803
rect 7591 769 7627 803
rect 7661 769 7696 803
rect 7730 769 7754 803
rect 6988 751 7754 769
rect 7022 731 7754 751
rect 7022 701 7067 731
rect 6988 697 7067 701
rect 7101 697 7137 731
rect 7171 697 7207 731
rect 7241 697 7277 731
rect 7311 697 7347 731
rect 7381 697 7417 731
rect 7451 697 7487 731
rect 7521 697 7557 731
rect 7591 697 7627 731
rect 7661 697 7696 731
rect 7730 697 7754 731
rect 6988 683 7754 697
rect 7022 659 7754 683
rect 7022 629 7067 659
rect 6988 625 7067 629
rect 7101 625 7137 659
rect 7171 625 7207 659
rect 7241 625 7277 659
rect 7311 625 7347 659
rect 7381 625 7417 659
rect 7451 625 7487 659
rect 7521 625 7557 659
rect 7591 625 7627 659
rect 7661 625 7696 659
rect 7730 625 7754 659
rect 6988 615 7754 625
rect 7022 587 7754 615
rect 7022 557 7067 587
rect 6988 553 7067 557
rect 7101 553 7137 587
rect 7171 553 7207 587
rect 7241 553 7277 587
rect 7311 553 7347 587
rect 7381 553 7417 587
rect 7451 553 7487 587
rect 7521 553 7557 587
rect 7591 553 7627 587
rect 7661 553 7696 587
rect 7730 553 7754 587
rect 6988 547 7754 553
rect 7022 515 7754 547
rect 7022 485 7067 515
rect 6988 481 7067 485
rect 7101 481 7137 515
rect 7171 481 7207 515
rect 7241 481 7277 515
rect 7311 481 7347 515
rect 7381 481 7417 515
rect 7451 481 7487 515
rect 7521 481 7557 515
rect 7591 481 7627 515
rect 7661 481 7696 515
rect 7730 481 7754 515
rect 6988 479 7754 481
rect 7022 443 7754 479
rect 7022 413 7067 443
rect 6988 411 7067 413
rect 7022 409 7067 411
rect 7101 409 7137 443
rect 7171 409 7207 443
rect 7241 409 7277 443
rect 7311 409 7347 443
rect 7381 409 7417 443
rect 7451 409 7487 443
rect 7521 409 7557 443
rect 7591 409 7627 443
rect 7661 409 7696 443
rect 7730 409 7754 443
rect 7022 377 7754 409
rect 6988 375 7754 377
rect 7022 369 7754 375
rect 9687 955 14576 988
rect 14610 955 14654 989
rect 14688 955 14732 989
rect 14766 955 14810 989
rect 14844 955 14888 989
rect 14922 956 14966 989
rect 14922 955 14932 956
rect 9687 947 11680 955
rect 9687 913 9711 947
rect 9745 913 9781 947
rect 9815 923 9851 947
rect 9885 923 9921 947
rect 9955 923 9991 947
rect 10025 923 10061 947
rect 9830 913 9851 923
rect 9906 913 9921 923
rect 9982 913 9991 923
rect 10058 913 10061 923
rect 10095 923 10131 947
rect 10165 923 10201 947
rect 10235 923 10271 947
rect 10305 923 10341 947
rect 10375 923 10411 947
rect 10445 923 10481 947
rect 10095 913 10100 923
rect 10165 913 10176 923
rect 10235 913 10251 923
rect 10305 913 10326 923
rect 10375 913 10401 923
rect 10445 913 10476 923
rect 10515 913 10551 947
rect 10585 913 10621 947
rect 10655 923 10691 947
rect 10725 923 10761 947
rect 10795 923 10831 947
rect 10865 923 10901 947
rect 10935 923 10971 947
rect 11005 923 11041 947
rect 10660 913 10691 923
rect 10735 913 10761 923
rect 10810 913 10831 923
rect 10885 913 10901 923
rect 10960 913 10971 923
rect 11035 913 11041 923
rect 11075 923 11111 947
rect 11075 913 11076 923
rect 9687 889 9796 913
rect 9830 889 9872 913
rect 9906 889 9948 913
rect 9982 889 10024 913
rect 10058 889 10100 913
rect 10134 889 10176 913
rect 10210 889 10251 913
rect 10285 889 10326 913
rect 10360 889 10401 913
rect 10435 889 10476 913
rect 10510 889 10551 913
rect 10585 889 10626 913
rect 10660 889 10701 913
rect 10735 889 10776 913
rect 10810 889 10851 913
rect 10885 889 10926 913
rect 10960 889 11001 913
rect 11035 889 11076 913
rect 11110 913 11111 923
rect 11145 923 11181 947
rect 11215 923 11251 947
rect 11285 923 11321 947
rect 11145 913 11151 923
rect 11215 913 11226 923
rect 11285 913 11301 923
rect 11355 913 11391 947
rect 11425 913 11460 947
rect 11494 913 11529 947
rect 11563 913 11598 947
rect 11632 921 11680 947
rect 11714 921 11750 955
rect 11784 921 11820 955
rect 11854 921 11890 955
rect 11924 921 11960 955
rect 11994 921 12030 955
rect 12064 921 12099 955
rect 12133 921 12168 955
rect 12202 921 12237 955
rect 12271 921 12306 955
rect 12340 921 12375 955
rect 12409 921 12444 955
rect 12478 921 12513 955
rect 12547 921 12582 955
rect 12616 921 12651 955
rect 12685 921 12720 955
rect 12754 921 12789 955
rect 12823 921 12858 955
rect 12892 921 12927 955
rect 12961 921 12996 955
rect 13030 921 13065 955
rect 13099 921 13134 955
rect 13168 921 13203 955
rect 13237 921 13272 955
rect 13306 921 13341 955
rect 13375 921 13410 955
rect 13444 921 13479 955
rect 13513 921 13548 955
rect 13582 921 13617 955
rect 13651 921 13686 955
rect 13720 921 13755 955
rect 13789 921 13824 955
rect 13858 921 13893 955
rect 13927 921 13962 955
rect 13996 921 14031 955
rect 14065 921 14100 955
rect 14134 921 14169 955
rect 14203 921 14238 955
rect 14272 921 14307 955
rect 14341 921 14376 955
rect 14410 921 14445 955
rect 14479 921 14514 955
rect 14548 921 14583 955
rect 14617 921 14652 955
rect 14686 921 14721 955
rect 14755 921 14790 955
rect 14824 921 14859 955
rect 14893 922 14932 955
rect 15000 959 15068 989
rect 15102 959 15117 993
rect 15000 956 15117 959
rect 14966 922 15000 955
rect 15034 922 15068 956
rect 15102 922 15117 956
rect 14893 921 15117 922
rect 11632 916 15068 921
rect 11632 913 14576 916
rect 11110 889 11151 913
rect 11185 889 11226 913
rect 11260 889 11301 913
rect 11335 889 14576 913
rect 9687 882 14576 889
rect 14610 882 14654 916
rect 14688 882 14732 916
rect 14766 882 14810 916
rect 14844 882 14888 916
rect 14922 884 14966 916
rect 14922 882 14932 884
rect 9687 875 14932 882
rect 9687 841 9711 875
rect 9745 841 9781 875
rect 9815 841 9851 875
rect 9885 841 9921 875
rect 9955 841 9991 875
rect 10025 841 10061 875
rect 10095 841 10131 875
rect 10165 841 10201 875
rect 10235 841 10271 875
rect 10305 841 10341 875
rect 10375 841 10411 875
rect 10445 841 10481 875
rect 10515 841 10551 875
rect 10585 841 10621 875
rect 10655 841 10691 875
rect 10725 841 10761 875
rect 10795 841 10831 875
rect 10865 841 10901 875
rect 10935 841 10971 875
rect 11005 841 11041 875
rect 11075 841 11111 875
rect 11145 841 11181 875
rect 11215 841 11251 875
rect 11285 841 11321 875
rect 11355 841 11391 875
rect 11425 841 11460 875
rect 11494 841 11529 875
rect 11563 841 11598 875
rect 11632 841 11680 875
rect 11714 841 11750 875
rect 11784 841 11820 875
rect 11854 841 11890 875
rect 11924 841 11960 875
rect 11994 841 12030 875
rect 12064 841 12099 875
rect 12133 841 12168 875
rect 12202 841 12237 875
rect 12271 841 12306 875
rect 12340 841 12375 875
rect 12409 841 12444 875
rect 12478 841 12513 875
rect 12547 841 12582 875
rect 12616 841 12651 875
rect 12685 841 12720 875
rect 12754 841 12789 875
rect 12823 841 12858 875
rect 12892 841 12927 875
rect 12961 841 12996 875
rect 13030 841 13065 875
rect 13099 841 13134 875
rect 13168 841 13203 875
rect 13237 841 13272 875
rect 13306 841 13341 875
rect 13375 841 13410 875
rect 13444 841 13479 875
rect 13513 841 13548 875
rect 13582 841 13617 875
rect 13651 841 13686 875
rect 13720 841 13755 875
rect 13789 841 13824 875
rect 13858 841 13893 875
rect 13927 841 13962 875
rect 13996 841 14031 875
rect 14065 841 14100 875
rect 14134 841 14169 875
rect 14203 841 14238 875
rect 14272 841 14307 875
rect 14341 841 14376 875
rect 14410 841 14445 875
rect 14479 841 14514 875
rect 14548 843 14583 875
rect 14548 841 14576 843
rect 14617 841 14652 875
rect 14686 843 14721 875
rect 14755 843 14790 875
rect 14824 843 14859 875
rect 14893 850 14932 875
rect 15000 887 15068 916
rect 15102 887 15117 921
rect 15000 884 15117 887
rect 14966 850 15000 882
rect 15034 850 15068 884
rect 15102 850 15117 884
rect 14893 849 15117 850
rect 14893 843 15068 849
rect 14688 841 14721 843
rect 14766 841 14790 843
rect 14844 841 14859 843
rect 9687 839 14576 841
rect 9687 805 9796 839
rect 9830 805 9872 839
rect 9906 805 9948 839
rect 9982 805 10024 839
rect 10058 805 10100 839
rect 10134 805 10176 839
rect 10210 805 10251 839
rect 10285 805 10326 839
rect 10360 805 10401 839
rect 10435 805 10476 839
rect 10510 805 10551 839
rect 10585 805 10626 839
rect 10660 805 10701 839
rect 10735 805 10776 839
rect 10810 805 10851 839
rect 10885 805 10926 839
rect 10960 805 11001 839
rect 11035 805 11076 839
rect 11110 805 11151 839
rect 11185 805 11226 839
rect 11260 805 11301 839
rect 11335 809 14576 839
rect 14610 809 14654 841
rect 14688 809 14732 841
rect 14766 809 14810 841
rect 14844 809 14888 841
rect 14922 812 14966 843
rect 14922 809 14932 812
rect 11335 805 14932 809
rect 9687 803 14932 805
rect 9687 769 9711 803
rect 9745 769 9781 803
rect 9815 769 9851 803
rect 9885 769 9921 803
rect 9955 769 9991 803
rect 10025 769 10061 803
rect 10095 769 10131 803
rect 10165 769 10201 803
rect 10235 769 10271 803
rect 10305 769 10341 803
rect 10375 769 10411 803
rect 10445 769 10481 803
rect 10515 769 10551 803
rect 10585 769 10621 803
rect 10655 769 10691 803
rect 10725 769 10761 803
rect 10795 769 10831 803
rect 10865 769 10901 803
rect 10935 769 10971 803
rect 11005 769 11041 803
rect 11075 769 11111 803
rect 11145 769 11181 803
rect 11215 769 11251 803
rect 11285 769 11321 803
rect 11355 769 11391 803
rect 11425 769 11460 803
rect 11494 769 11529 803
rect 11563 769 11598 803
rect 11632 795 14932 803
rect 11632 769 11680 795
rect 9687 761 11680 769
rect 11714 761 11750 795
rect 11784 761 11820 795
rect 11854 761 11890 795
rect 11924 761 11960 795
rect 11994 761 12030 795
rect 12064 761 12099 795
rect 12133 761 12168 795
rect 12202 761 12237 795
rect 12271 761 12306 795
rect 12340 761 12375 795
rect 12409 761 12444 795
rect 12478 761 12513 795
rect 12547 761 12582 795
rect 12616 761 12651 795
rect 12685 761 12720 795
rect 12754 761 12789 795
rect 12823 761 12858 795
rect 12892 761 12927 795
rect 12961 761 12996 795
rect 13030 761 13065 795
rect 13099 761 13134 795
rect 13168 761 13203 795
rect 13237 761 13272 795
rect 13306 761 13341 795
rect 13375 761 13410 795
rect 13444 761 13479 795
rect 13513 761 13548 795
rect 13582 761 13617 795
rect 13651 761 13686 795
rect 13720 761 13755 795
rect 13789 761 13824 795
rect 13858 761 13893 795
rect 13927 761 13962 795
rect 13996 761 14031 795
rect 14065 761 14100 795
rect 14134 761 14169 795
rect 14203 761 14238 795
rect 14272 761 14307 795
rect 14341 761 14376 795
rect 14410 761 14445 795
rect 14479 761 14514 795
rect 14548 770 14583 795
rect 14548 761 14576 770
rect 14617 761 14652 795
rect 14686 770 14721 795
rect 14755 770 14790 795
rect 14824 770 14859 795
rect 14893 778 14932 795
rect 15000 815 15068 843
rect 15102 815 15117 849
rect 15000 812 15117 815
rect 14966 778 15000 809
rect 15034 778 15068 812
rect 15102 778 15117 812
rect 14893 777 15117 778
rect 14893 770 15068 777
rect 14688 761 14721 770
rect 14766 761 14790 770
rect 14844 761 14859 770
rect 9687 755 14576 761
rect 9687 731 9796 755
rect 9830 731 9872 755
rect 9906 731 9948 755
rect 9982 731 10024 755
rect 10058 731 10100 755
rect 10134 731 10176 755
rect 10210 731 10251 755
rect 10285 731 10326 755
rect 10360 731 10401 755
rect 10435 731 10476 755
rect 10510 731 10551 755
rect 10585 731 10626 755
rect 10660 731 10701 755
rect 10735 731 10776 755
rect 10810 731 10851 755
rect 10885 731 10926 755
rect 10960 731 11001 755
rect 11035 731 11076 755
rect 9687 697 9711 731
rect 9745 697 9781 731
rect 9830 721 9851 731
rect 9906 721 9921 731
rect 9982 721 9991 731
rect 10058 721 10061 731
rect 9815 697 9851 721
rect 9885 697 9921 721
rect 9955 697 9991 721
rect 10025 697 10061 721
rect 10095 721 10100 731
rect 10165 721 10176 731
rect 10235 721 10251 731
rect 10305 721 10326 731
rect 10375 721 10401 731
rect 10445 721 10476 731
rect 10095 697 10131 721
rect 10165 697 10201 721
rect 10235 697 10271 721
rect 10305 697 10341 721
rect 10375 697 10411 721
rect 10445 697 10481 721
rect 10515 697 10551 731
rect 10585 697 10621 731
rect 10660 721 10691 731
rect 10735 721 10761 731
rect 10810 721 10831 731
rect 10885 721 10901 731
rect 10960 721 10971 731
rect 11035 721 11041 731
rect 10655 697 10691 721
rect 10725 697 10761 721
rect 10795 697 10831 721
rect 10865 697 10901 721
rect 10935 697 10971 721
rect 11005 697 11041 721
rect 11075 721 11076 731
rect 11110 731 11151 755
rect 11185 731 11226 755
rect 11260 731 11301 755
rect 11335 736 14576 755
rect 14610 736 14654 761
rect 14688 736 14732 761
rect 14766 736 14810 761
rect 14844 736 14888 761
rect 14922 740 14966 770
rect 14922 736 14932 740
rect 11335 731 14932 736
rect 11110 721 11111 731
rect 11075 697 11111 721
rect 11145 721 11151 731
rect 11215 721 11226 731
rect 11285 721 11301 731
rect 11145 697 11181 721
rect 11215 697 11251 721
rect 11285 697 11321 721
rect 11355 697 11391 731
rect 11425 697 11460 731
rect 11494 697 11529 731
rect 11563 697 11598 731
rect 11632 728 14932 731
rect 11632 697 11656 728
rect 9687 671 11656 697
rect 9687 659 9796 671
rect 9830 659 9872 671
rect 9906 659 9948 671
rect 9982 659 10024 671
rect 10058 659 10100 671
rect 10134 659 10176 671
rect 10210 659 10251 671
rect 10285 659 10326 671
rect 10360 659 10401 671
rect 10435 659 10476 671
rect 10510 659 10551 671
rect 10585 659 10626 671
rect 10660 659 10701 671
rect 10735 659 10776 671
rect 10810 659 10851 671
rect 10885 659 10926 671
rect 10960 659 11001 671
rect 11035 659 11076 671
rect 9687 625 9711 659
rect 9745 625 9781 659
rect 9830 637 9851 659
rect 9906 637 9921 659
rect 9982 637 9991 659
rect 10058 637 10061 659
rect 9815 625 9851 637
rect 9885 625 9921 637
rect 9955 625 9991 637
rect 10025 625 10061 637
rect 10095 637 10100 659
rect 10165 637 10176 659
rect 10235 637 10251 659
rect 10305 637 10326 659
rect 10375 637 10401 659
rect 10445 637 10476 659
rect 10095 625 10131 637
rect 10165 625 10201 637
rect 10235 625 10271 637
rect 10305 625 10341 637
rect 10375 625 10411 637
rect 10445 625 10481 637
rect 10515 625 10551 659
rect 10585 625 10621 659
rect 10660 637 10691 659
rect 10735 637 10761 659
rect 10810 637 10831 659
rect 10885 637 10901 659
rect 10960 637 10971 659
rect 11035 637 11041 659
rect 10655 625 10691 637
rect 10725 625 10761 637
rect 10795 625 10831 637
rect 10865 625 10901 637
rect 10935 625 10971 637
rect 11005 625 11041 637
rect 11075 637 11076 659
rect 11110 659 11151 671
rect 11185 659 11226 671
rect 11260 659 11301 671
rect 11335 659 11656 671
rect 11110 637 11111 659
rect 11075 625 11111 637
rect 11145 637 11151 659
rect 11215 637 11226 659
rect 11285 637 11301 659
rect 11145 625 11181 637
rect 11215 625 11251 637
rect 11285 625 11321 637
rect 11355 625 11391 659
rect 11425 625 11460 659
rect 11494 625 11529 659
rect 11563 625 11598 659
rect 11632 625 11656 659
rect 9687 587 11656 625
rect 9687 553 9711 587
rect 9745 553 9781 587
rect 9830 553 9851 587
rect 9906 553 9921 587
rect 9982 553 9991 587
rect 10058 553 10061 587
rect 10095 553 10100 587
rect 10165 553 10176 587
rect 10235 553 10251 587
rect 10305 553 10326 587
rect 10375 553 10401 587
rect 10445 553 10476 587
rect 10515 553 10551 587
rect 10585 553 10621 587
rect 10660 553 10691 587
rect 10735 553 10761 587
rect 10810 553 10831 587
rect 10885 553 10901 587
rect 10960 553 10971 587
rect 11035 553 11041 587
rect 11075 553 11076 587
rect 11110 553 11111 587
rect 11145 553 11151 587
rect 11215 553 11226 587
rect 11285 553 11301 587
rect 11355 553 11391 587
rect 11425 553 11460 587
rect 11494 553 11529 587
rect 11563 553 11598 587
rect 11632 553 11656 587
rect 9687 515 11656 553
rect 9687 481 9711 515
rect 9745 481 9781 515
rect 9815 503 9851 515
rect 9885 503 9921 515
rect 9955 503 9991 515
rect 10025 503 10061 515
rect 9830 481 9851 503
rect 9906 481 9921 503
rect 9982 481 9991 503
rect 10058 481 10061 503
rect 10095 503 10131 515
rect 10165 503 10201 515
rect 10235 503 10271 515
rect 10305 503 10341 515
rect 10375 503 10411 515
rect 10445 503 10481 515
rect 10095 481 10100 503
rect 10165 481 10176 503
rect 10235 481 10251 503
rect 10305 481 10326 503
rect 10375 481 10401 503
rect 10445 481 10476 503
rect 10515 481 10551 515
rect 10585 481 10621 515
rect 10655 503 10691 515
rect 10725 503 10761 515
rect 10795 503 10831 515
rect 10865 503 10901 515
rect 10935 503 10971 515
rect 11005 503 11041 515
rect 10660 481 10691 503
rect 10735 481 10761 503
rect 10810 481 10831 503
rect 10885 481 10901 503
rect 10960 481 10971 503
rect 11035 481 11041 503
rect 11075 503 11111 515
rect 11075 481 11076 503
rect 9687 469 9796 481
rect 9830 469 9872 481
rect 9906 469 9948 481
rect 9982 469 10024 481
rect 10058 469 10100 481
rect 10134 469 10176 481
rect 10210 469 10251 481
rect 10285 469 10326 481
rect 10360 469 10401 481
rect 10435 469 10476 481
rect 10510 469 10551 481
rect 10585 469 10626 481
rect 10660 469 10701 481
rect 10735 469 10776 481
rect 10810 469 10851 481
rect 10885 469 10926 481
rect 10960 469 11001 481
rect 11035 469 11076 481
rect 11110 481 11111 503
rect 11145 503 11181 515
rect 11215 503 11251 515
rect 11285 503 11321 515
rect 11145 481 11151 503
rect 11215 481 11226 503
rect 11285 481 11301 503
rect 11355 481 11391 515
rect 11425 481 11460 515
rect 11494 481 11529 515
rect 11563 481 11598 515
rect 11632 481 11656 515
rect 11110 469 11151 481
rect 11185 469 11226 481
rect 11260 469 11301 481
rect 11335 469 11656 481
rect 9687 443 11656 469
rect 9687 409 9711 443
rect 9745 409 9781 443
rect 9815 409 9851 443
rect 9885 409 9921 443
rect 9955 409 9991 443
rect 10025 409 10061 443
rect 10095 409 10131 443
rect 10165 409 10201 443
rect 10235 409 10271 443
rect 10305 409 10341 443
rect 10375 409 10411 443
rect 10445 409 10481 443
rect 10515 409 10551 443
rect 10585 409 10621 443
rect 10655 409 10691 443
rect 10725 409 10761 443
rect 10795 409 10831 443
rect 10865 409 10901 443
rect 10935 409 10971 443
rect 11005 409 11041 443
rect 11075 409 11111 443
rect 11145 409 11181 443
rect 11215 409 11251 443
rect 11285 409 11321 443
rect 11355 409 11391 443
rect 11425 409 11460 443
rect 11494 409 11529 443
rect 11563 409 11598 443
rect 11632 409 11656 443
rect 9687 369 11656 409
rect 14465 706 14932 728
rect 15000 743 15068 770
rect 15102 743 15117 777
rect 15000 740 15117 743
rect 14966 706 15000 736
rect 15034 706 15068 740
rect 15102 706 15117 740
rect 14465 705 15117 706
rect 14465 697 15068 705
rect 14465 695 14576 697
rect 14610 695 14654 697
rect 14688 695 14732 697
rect 14499 661 14543 695
rect 14610 663 14621 695
rect 14688 663 14698 695
rect 14577 661 14621 663
rect 14655 661 14698 663
rect 14766 695 14810 697
rect 14766 663 14775 695
rect 14732 661 14775 663
rect 14809 663 14810 695
rect 14844 695 14888 697
rect 14844 663 14852 695
rect 14809 661 14852 663
rect 14886 663 14888 695
rect 14922 668 14966 697
rect 14922 663 14932 668
rect 14886 661 14932 663
rect 14465 634 14932 661
rect 15000 671 15068 697
rect 15102 671 15117 705
rect 15000 668 15117 671
rect 14966 634 15000 663
rect 15034 634 15068 668
rect 15102 634 15117 668
rect 14465 633 15117 634
rect 14465 623 15068 633
rect 14465 609 14576 623
rect 14610 609 14654 623
rect 14688 609 14732 623
rect 14499 575 14543 609
rect 14610 589 14621 609
rect 14688 589 14698 609
rect 14577 575 14621 589
rect 14655 575 14698 589
rect 14766 609 14810 623
rect 14766 589 14775 609
rect 14732 575 14775 589
rect 14809 589 14810 609
rect 14844 609 14888 623
rect 14844 589 14852 609
rect 14809 575 14852 589
rect 14886 589 14888 609
rect 14922 596 14966 623
rect 14922 589 14932 596
rect 14886 575 14932 589
rect 14465 562 14932 575
rect 15000 599 15068 623
rect 15102 599 15117 633
rect 15000 596 15117 599
rect 14966 562 15000 589
rect 15034 562 15068 596
rect 15102 562 15117 596
rect 14465 561 15117 562
rect 14465 549 15068 561
rect 14465 523 14576 549
rect 14610 523 14654 549
rect 14688 523 14732 549
rect 14499 489 14543 523
rect 14610 515 14621 523
rect 14688 515 14698 523
rect 14577 489 14621 515
rect 14655 489 14698 515
rect 14766 523 14810 549
rect 14766 515 14775 523
rect 14732 489 14775 515
rect 14809 515 14810 523
rect 14844 523 14888 549
rect 14844 515 14852 523
rect 14809 489 14852 515
rect 14886 515 14888 523
rect 14922 524 14966 549
rect 14922 515 14932 524
rect 14886 490 14932 515
rect 15000 527 15068 549
rect 15102 527 15117 561
rect 15000 524 15117 527
rect 14966 490 15000 515
rect 15034 490 15068 524
rect 15102 490 15117 524
rect 14886 489 15117 490
rect 14465 475 15068 489
rect 14465 441 14576 475
rect 14610 441 14654 475
rect 14688 441 14732 475
rect 14766 441 14810 475
rect 14844 441 14888 475
rect 14922 452 14966 475
rect 14922 441 14932 452
rect 14465 437 14932 441
rect 14499 403 14543 437
rect 14577 403 14621 437
rect 14655 403 14698 437
rect 14732 403 14775 437
rect 14809 403 14852 437
rect 14886 418 14932 437
rect 15000 455 15068 475
rect 15102 455 15117 489
rect 15000 452 15117 455
rect 14966 418 15000 441
rect 15034 418 15068 452
rect 15102 418 15117 452
rect 14886 417 15117 418
rect 14886 403 15068 417
rect 14465 390 15068 403
rect 14465 369 14657 390
rect 7022 367 14657 369
rect 14691 367 14735 390
rect 14769 367 14813 390
rect 14847 367 14891 390
rect 14925 380 14969 390
rect 15003 383 15068 390
rect 15102 383 15117 417
rect 15003 380 15117 383
rect 7022 333 7056 367
rect 7090 333 7125 367
rect 7159 333 7194 367
rect 7228 333 7263 367
rect 7297 333 7332 367
rect 7366 333 7401 367
rect 7435 333 7470 367
rect 7504 333 7539 367
rect 7573 333 7608 367
rect 7642 333 7677 367
rect 7711 333 7746 367
rect 7780 333 7815 367
rect 7849 333 7884 367
rect 7918 333 7953 367
rect 7987 333 8022 367
rect 8056 333 8091 367
rect 8125 333 8160 367
rect 8194 333 8229 367
rect 8263 333 8298 367
rect 8332 333 8367 367
rect 8401 333 8436 367
rect 8470 333 8505 367
rect 8539 333 8574 367
rect 8608 333 8643 367
rect 8677 333 8712 367
rect 8746 333 8781 367
rect 8815 333 8850 367
rect 8884 333 8919 367
rect 8953 333 8988 367
rect 9022 333 9057 367
rect 9091 333 9126 367
rect 9160 333 9195 367
rect 9229 333 9264 367
rect 9298 333 9333 367
rect 9367 333 9402 367
rect 9436 333 9471 367
rect 9505 333 9540 367
rect 9574 333 9609 367
rect 9643 333 9678 367
rect 9712 333 9747 367
rect 9781 333 9816 367
rect 9850 333 9885 367
rect 9919 333 9954 367
rect 9988 333 10023 367
rect 10057 333 10092 367
rect 10126 333 10161 367
rect 10195 333 10230 367
rect 10264 333 10299 367
rect 10333 333 10368 367
rect 10402 333 10437 367
rect 10471 333 10506 367
rect 10540 333 10575 367
rect 10609 333 10643 367
rect 10677 333 10711 367
rect 10745 333 10779 367
rect 10813 333 10847 367
rect 10881 333 10915 367
rect 10949 333 10983 367
rect 11017 333 11051 367
rect 11085 333 11119 367
rect 11153 333 11187 367
rect 11221 333 11255 367
rect 11289 333 11323 367
rect 11357 333 11391 367
rect 11425 333 11459 367
rect 11493 333 11527 367
rect 11561 333 11595 367
rect 11629 333 11663 367
rect 11697 333 11731 367
rect 11765 333 11799 367
rect 11833 333 11867 367
rect 11901 333 11935 367
rect 11969 333 12003 367
rect 12037 333 12071 367
rect 12105 333 12139 367
rect 12173 333 12207 367
rect 12241 333 12275 367
rect 12309 333 12343 367
rect 12377 333 12411 367
rect 12445 333 12479 367
rect 12513 333 12547 367
rect 12581 333 12615 367
rect 12649 333 12683 367
rect 12717 333 12751 367
rect 12785 333 12819 367
rect 12853 333 12887 367
rect 12921 333 12955 367
rect 12989 333 13023 367
rect 13057 333 13091 367
rect 13125 333 13159 367
rect 13193 333 13227 367
rect 13261 333 13295 367
rect 13329 333 13363 367
rect 13397 333 13431 367
rect 13465 333 13499 367
rect 13533 333 13567 367
rect 13601 333 13635 367
rect 13669 333 13703 367
rect 13737 333 13771 367
rect 13805 333 13839 367
rect 13873 333 13907 367
rect 13941 333 13975 367
rect 14009 333 14043 367
rect 14077 333 14111 367
rect 14145 333 14179 367
rect 14213 333 14247 367
rect 14281 333 14315 367
rect 14349 333 14383 367
rect 14417 333 14451 367
rect 14485 333 14519 367
rect 14553 333 14587 367
rect 14621 333 14655 367
rect 14691 356 14723 367
rect 14769 356 14791 367
rect 14847 356 14859 367
rect 14925 356 14932 380
rect 14689 333 14723 356
rect 14757 333 14791 356
rect 14825 333 14859 356
rect 14893 346 14932 356
rect 14966 356 14969 380
rect 14966 346 15000 356
rect 15034 346 15068 380
rect 15102 346 15117 380
rect 14893 345 15117 346
rect 14893 333 15068 345
rect 7022 312 15068 333
rect 7022 309 14657 312
rect 6988 303 14657 309
rect 7022 289 14657 303
rect 14691 289 14735 312
rect 14769 289 14813 312
rect 14847 289 14891 312
rect 14925 308 14969 312
rect 15003 311 15068 312
rect 15102 311 15117 345
rect 15003 308 15117 311
rect 7022 255 7056 289
rect 7090 255 7125 289
rect 7159 255 7194 289
rect 7228 255 7263 289
rect 7297 255 7332 289
rect 7366 255 7401 289
rect 7435 255 7470 289
rect 7504 255 7539 289
rect 7573 255 7608 289
rect 7642 255 7677 289
rect 7711 255 7746 289
rect 7780 255 7815 289
rect 7849 255 7884 289
rect 7918 255 7953 289
rect 7987 255 8022 289
rect 8056 255 8091 289
rect 8125 255 8160 289
rect 8194 255 8229 289
rect 8263 255 8298 289
rect 8332 255 8367 289
rect 8401 255 8436 289
rect 8470 255 8505 289
rect 8539 255 8574 289
rect 8608 255 8643 289
rect 8677 255 8712 289
rect 8746 255 8781 289
rect 8815 255 8850 289
rect 8884 255 8919 289
rect 8953 255 8988 289
rect 9022 255 9057 289
rect 9091 255 9126 289
rect 9160 255 9195 289
rect 9229 255 9264 289
rect 9298 255 9333 289
rect 9367 255 9402 289
rect 9436 255 9471 289
rect 9505 255 9540 289
rect 9574 255 9609 289
rect 9643 255 9678 289
rect 9712 255 9747 289
rect 9781 255 9816 289
rect 9850 255 9885 289
rect 9919 255 9954 289
rect 9988 255 10023 289
rect 10057 255 10092 289
rect 10126 255 10161 289
rect 10195 255 10230 289
rect 10264 255 10299 289
rect 10333 255 10368 289
rect 10402 255 10437 289
rect 10471 255 10506 289
rect 10540 255 10575 289
rect 10609 255 10643 289
rect 10677 255 10711 289
rect 10745 255 10779 289
rect 10813 255 10847 289
rect 10881 255 10915 289
rect 10949 255 10983 289
rect 11017 255 11051 289
rect 11085 255 11119 289
rect 11153 255 11187 289
rect 11221 255 11255 289
rect 11289 255 11323 289
rect 11357 255 11391 289
rect 11425 255 11459 289
rect 11493 255 11527 289
rect 11561 255 11595 289
rect 11629 255 11663 289
rect 11697 255 11731 289
rect 11765 255 11799 289
rect 11833 255 11867 289
rect 11901 255 11935 289
rect 11969 255 12003 289
rect 12037 255 12071 289
rect 12105 255 12139 289
rect 12173 255 12207 289
rect 12241 255 12275 289
rect 12309 255 12343 289
rect 12377 255 12411 289
rect 12445 255 12479 289
rect 12513 255 12547 289
rect 12581 255 12615 289
rect 12649 255 12683 289
rect 12717 255 12751 289
rect 12785 255 12819 289
rect 12853 255 12887 289
rect 12921 255 12955 289
rect 12989 255 13023 289
rect 13057 255 13091 289
rect 13125 255 13159 289
rect 13193 255 13227 289
rect 13261 255 13295 289
rect 13329 255 13363 289
rect 13397 255 13431 289
rect 13465 255 13499 289
rect 13533 255 13567 289
rect 13601 255 13635 289
rect 13669 255 13703 289
rect 13737 255 13771 289
rect 13805 255 13839 289
rect 13873 255 13907 289
rect 13941 255 13975 289
rect 14009 255 14043 289
rect 14077 255 14111 289
rect 14145 255 14179 289
rect 14213 255 14247 289
rect 14281 255 14315 289
rect 14349 255 14383 289
rect 14417 255 14451 289
rect 14485 255 14519 289
rect 14553 255 14587 289
rect 14621 255 14655 289
rect 14691 278 14723 289
rect 14769 278 14791 289
rect 14847 278 14859 289
rect 14925 278 14932 308
rect 14689 255 14723 278
rect 14757 255 14791 278
rect 14825 255 14859 278
rect 14893 274 14932 278
rect 14966 278 14969 308
rect 14966 274 15000 278
rect 15034 274 15068 308
rect 15102 274 15117 308
rect 14893 272 15117 274
rect 14893 255 15068 272
rect 7022 241 15068 255
rect 6988 238 15068 241
rect 15102 238 15117 272
rect 6988 236 15117 238
rect 6988 234 14932 236
rect 6988 231 14657 234
rect 7022 211 14657 231
rect 14691 211 14735 234
rect 14769 211 14813 234
rect 14847 211 14891 234
rect 7022 177 7056 211
rect 7090 177 7125 211
rect 7159 177 7194 211
rect 7228 177 7263 211
rect 7297 177 7332 211
rect 7366 177 7401 211
rect 7435 177 7470 211
rect 7504 177 7539 211
rect 7573 177 7608 211
rect 7642 177 7677 211
rect 7711 177 7746 211
rect 7780 177 7815 211
rect 7849 177 7884 211
rect 7918 177 7953 211
rect 7987 177 8022 211
rect 8056 177 8091 211
rect 8125 177 8160 211
rect 8194 177 8229 211
rect 8263 177 8298 211
rect 8332 177 8367 211
rect 8401 177 8436 211
rect 8470 177 8505 211
rect 8539 177 8574 211
rect 8608 177 8643 211
rect 8677 177 8712 211
rect 8746 177 8781 211
rect 8815 177 8850 211
rect 8884 177 8919 211
rect 8953 177 8988 211
rect 9022 177 9057 211
rect 9091 177 9126 211
rect 9160 177 9195 211
rect 9229 177 9264 211
rect 9298 177 9333 211
rect 9367 177 9402 211
rect 9436 177 9471 211
rect 9505 177 9540 211
rect 9574 177 9609 211
rect 9643 177 9678 211
rect 9712 177 9747 211
rect 9781 177 9816 211
rect 9850 177 9885 211
rect 9919 177 9954 211
rect 9988 177 10023 211
rect 10057 177 10092 211
rect 10126 177 10161 211
rect 10195 177 10230 211
rect 10264 177 10299 211
rect 10333 177 10368 211
rect 10402 177 10437 211
rect 10471 177 10506 211
rect 10540 177 10575 211
rect 10609 177 10643 211
rect 10677 177 10711 211
rect 10745 177 10779 211
rect 10813 177 10847 211
rect 10881 177 10915 211
rect 10949 177 10983 211
rect 11017 177 11051 211
rect 11085 177 11119 211
rect 11153 177 11187 211
rect 11221 177 11255 211
rect 11289 177 11323 211
rect 11357 177 11391 211
rect 11425 177 11459 211
rect 11493 177 11527 211
rect 11561 177 11595 211
rect 11629 177 11663 211
rect 11697 177 11731 211
rect 11765 177 11799 211
rect 11833 177 11867 211
rect 11901 177 11935 211
rect 11969 177 12003 211
rect 12037 177 12071 211
rect 12105 177 12139 211
rect 12173 177 12207 211
rect 12241 177 12275 211
rect 12309 177 12343 211
rect 12377 177 12411 211
rect 12445 177 12479 211
rect 12513 177 12547 211
rect 12581 177 12615 211
rect 12649 177 12683 211
rect 12717 177 12751 211
rect 12785 177 12819 211
rect 12853 177 12887 211
rect 12921 177 12955 211
rect 12989 177 13023 211
rect 13057 177 13091 211
rect 13125 177 13159 211
rect 13193 177 13227 211
rect 13261 177 13295 211
rect 13329 177 13363 211
rect 13397 177 13431 211
rect 13465 177 13499 211
rect 13533 177 13567 211
rect 13601 177 13635 211
rect 13669 177 13703 211
rect 13737 177 13771 211
rect 13805 177 13839 211
rect 13873 177 13907 211
rect 13941 177 13975 211
rect 14009 177 14043 211
rect 14077 177 14111 211
rect 14145 177 14179 211
rect 14213 177 14247 211
rect 14281 177 14315 211
rect 14349 177 14383 211
rect 14417 177 14451 211
rect 14485 177 14519 211
rect 14553 177 14587 211
rect 14621 177 14655 211
rect 14691 200 14723 211
rect 14769 200 14791 211
rect 14847 200 14859 211
rect 14925 202 14932 234
rect 14966 234 15000 236
rect 14966 202 14969 234
rect 15034 202 15068 236
rect 15102 202 15117 236
rect 14925 200 14969 202
rect 15003 200 15117 202
rect 14689 177 14723 200
rect 14757 177 14791 200
rect 14825 177 14859 200
rect 14893 199 15117 200
rect 14893 177 15068 199
rect 7022 173 15068 177
rect 6988 165 15068 173
rect 15102 165 15117 199
rect 6988 164 15117 165
rect 6988 159 14932 164
rect 7022 156 14932 159
rect 7022 133 14657 156
rect 14691 133 14735 156
rect 14769 133 14813 156
rect 14847 133 14891 156
rect 7022 105 7056 133
rect 6988 99 7056 105
rect 7090 99 7125 133
rect 7159 99 7194 133
rect 7228 99 7263 133
rect 7297 99 7332 133
rect 7366 99 7401 133
rect 7435 99 7470 133
rect 7504 99 7539 133
rect 7573 99 7608 133
rect 7642 99 7677 133
rect 7711 99 7746 133
rect 7780 99 7815 133
rect 7849 99 7884 133
rect 7918 99 7953 133
rect 7987 99 8022 133
rect 8056 99 8091 133
rect 8125 99 8160 133
rect 8194 99 8229 133
rect 8263 99 8298 133
rect 8332 99 8367 133
rect 8401 99 8436 133
rect 8470 99 8505 133
rect 8539 99 8574 133
rect 8608 99 8643 133
rect 8677 99 8712 133
rect 8746 99 8781 133
rect 8815 99 8850 133
rect 8884 99 8919 133
rect 8953 99 8988 133
rect 9022 99 9057 133
rect 9091 99 9126 133
rect 9160 99 9195 133
rect 9229 99 9264 133
rect 9298 99 9333 133
rect 9367 99 9402 133
rect 9436 99 9471 133
rect 9505 99 9540 133
rect 9574 99 9609 133
rect 9643 99 9678 133
rect 9712 99 9747 133
rect 9781 99 9816 133
rect 9850 99 9885 133
rect 9919 99 9954 133
rect 9988 99 10023 133
rect 10057 99 10092 133
rect 10126 99 10161 133
rect 10195 99 10230 133
rect 10264 99 10299 133
rect 10333 99 10368 133
rect 10402 99 10437 133
rect 10471 99 10506 133
rect 10540 99 10575 133
rect 10609 99 10643 133
rect 10677 99 10711 133
rect 10745 99 10779 133
rect 10813 99 10847 133
rect 10881 99 10915 133
rect 10949 99 10983 133
rect 11017 99 11051 133
rect 11085 99 11119 133
rect 11153 99 11187 133
rect 11221 99 11255 133
rect 11289 99 11323 133
rect 11357 99 11391 133
rect 11425 99 11459 133
rect 11493 99 11527 133
rect 11561 99 11595 133
rect 11629 99 11663 133
rect 11697 99 11731 133
rect 11765 99 11799 133
rect 11833 99 11867 133
rect 11901 99 11935 133
rect 11969 99 12003 133
rect 12037 99 12071 133
rect 12105 99 12139 133
rect 12173 99 12207 133
rect 12241 99 12275 133
rect 12309 99 12343 133
rect 12377 99 12411 133
rect 12445 99 12479 133
rect 12513 99 12547 133
rect 12581 99 12615 133
rect 12649 99 12683 133
rect 12717 99 12751 133
rect 12785 99 12819 133
rect 12853 99 12887 133
rect 12921 99 12955 133
rect 12989 99 13023 133
rect 13057 99 13091 133
rect 13125 99 13159 133
rect 13193 99 13227 133
rect 13261 99 13295 133
rect 13329 99 13363 133
rect 13397 99 13431 133
rect 13465 99 13499 133
rect 13533 99 13567 133
rect 13601 99 13635 133
rect 13669 99 13703 133
rect 13737 99 13771 133
rect 13805 99 13839 133
rect 13873 99 13907 133
rect 13941 99 13975 133
rect 14009 99 14043 133
rect 14077 99 14111 133
rect 14145 99 14179 133
rect 14213 99 14247 133
rect 14281 99 14315 133
rect 14349 99 14383 133
rect 14417 99 14451 133
rect 14485 99 14519 133
rect 14553 99 14587 133
rect 14621 99 14655 133
rect 14691 122 14723 133
rect 14769 122 14791 133
rect 14847 122 14859 133
rect 14925 130 14932 156
rect 14966 156 15000 164
rect 14966 130 14969 156
rect 15034 130 15068 164
rect 15102 130 15117 164
rect 14925 122 14969 130
rect 15003 126 15117 130
rect 15003 122 15068 126
rect 14689 99 14723 122
rect 14757 99 14791 122
rect 14825 99 14859 122
rect 14893 99 15068 122
rect 6988 92 15068 99
rect 15102 92 15117 126
rect 6988 91 15117 92
rect 6988 77 14932 91
rect 6988 55 14657 77
rect 14691 55 14735 77
rect 14769 55 14813 77
rect 14847 55 14891 77
rect 14925 57 14932 77
rect 14966 77 15000 91
rect 14966 57 14969 77
rect 15034 57 15068 91
rect 15102 57 15117 91
rect 3545 1 3578 23
rect 3612 23 3652 35
rect 3686 23 3726 35
rect 3760 23 3800 35
rect 3834 23 3874 35
rect 3908 23 3948 35
rect 3982 23 4022 35
rect 4056 23 4096 35
rect 4130 23 4170 35
rect 4204 23 4244 35
rect 4278 23 4318 35
rect 4352 23 4392 35
rect 4426 23 4466 35
rect 4500 23 4540 35
rect 4574 23 4614 35
rect 4648 23 4688 35
rect 4722 23 4762 35
rect 4796 23 4836 35
rect 4870 23 4910 35
rect 4944 23 4984 35
rect 5018 23 5058 35
rect 5092 23 5132 35
rect 5166 23 5206 35
rect 5240 23 5280 35
rect 5314 23 5354 35
rect 5388 23 5428 35
rect 5462 23 5502 35
rect 3612 1 3632 23
rect 3686 1 3700 23
rect 3760 1 3768 23
rect 3834 1 3836 23
rect 3545 -11 3632 1
rect 3666 -11 3700 1
rect 3734 -11 3768 1
rect 3802 -11 3836 1
rect 3870 1 3874 23
rect 3938 1 3948 23
rect 4006 1 4022 23
rect 4074 1 4096 23
rect 4142 1 4170 23
rect 3870 -11 3904 1
rect 3938 -11 3972 1
rect 4006 -11 4040 1
rect 4074 -11 4108 1
rect 4142 -11 4176 1
rect 4210 -11 4244 23
rect 4278 -11 4312 23
rect 4352 1 4380 23
rect 4426 1 4448 23
rect 4500 1 4516 23
rect 4574 1 4584 23
rect 4648 1 4652 23
rect 4346 -11 4380 1
rect 4414 -11 4448 1
rect 4482 -11 4516 1
rect 4550 -11 4584 1
rect 4618 -11 4652 1
rect 4686 1 4688 23
rect 4754 1 4762 23
rect 4822 1 4836 23
rect 4890 1 4910 23
rect 4958 1 4984 23
rect 5026 1 5058 23
rect 4686 -11 4720 1
rect 4754 -11 4788 1
rect 4822 -11 4856 1
rect 4890 -11 4924 1
rect 4958 -11 4992 1
rect 5026 -11 5060 1
rect 5094 -11 5128 23
rect 5166 1 5196 23
rect 5240 1 5264 23
rect 5314 1 5332 23
rect 5388 1 5400 23
rect 5462 1 5468 23
rect 5162 -11 5196 1
rect 5230 -11 5264 1
rect 5298 -11 5332 1
rect 5366 -11 5400 1
rect 5434 -11 5468 1
rect 5536 23 5576 35
rect 5610 23 5650 35
rect 5684 23 5724 35
rect 5758 23 5798 35
rect 6988 23 7056 55
rect 5502 -11 5536 1
rect 5570 1 5576 23
rect 5638 1 5650 23
rect 5706 1 5724 23
rect 5774 1 5798 23
rect 5570 -11 5604 1
rect 5638 -11 5672 1
rect 5706 -11 5740 1
rect 5774 -11 5808 1
rect 5842 -11 5876 23
rect 5930 -11 5944 23
rect 6002 -11 6012 23
rect 6074 -11 6080 23
rect 6146 -11 6148 23
rect 6182 -11 6184 23
rect 6250 -11 6256 23
rect 6318 -11 6328 23
rect 6386 -11 6400 23
rect 6454 -11 6472 23
rect 6522 -11 6544 23
rect 6590 -11 6616 23
rect 6658 -11 6688 23
rect 6726 -11 6760 23
rect 6794 -11 6828 23
rect 6866 -11 6896 23
rect 6938 -11 6964 23
rect 7010 21 7056 23
rect 7090 21 7125 55
rect 7159 21 7194 55
rect 7228 21 7263 55
rect 7297 21 7332 55
rect 7366 21 7401 55
rect 7435 21 7470 55
rect 7504 21 7539 55
rect 7573 21 7608 55
rect 7642 21 7677 55
rect 7711 21 7746 55
rect 7780 21 7815 55
rect 7849 21 7884 55
rect 7918 21 7953 55
rect 7987 21 8022 55
rect 8056 21 8091 55
rect 8125 21 8160 55
rect 8194 21 8229 55
rect 8263 21 8298 55
rect 8332 21 8367 55
rect 8401 21 8436 55
rect 8470 21 8505 55
rect 8539 21 8574 55
rect 8608 21 8643 55
rect 8677 21 8712 55
rect 8746 21 8781 55
rect 8815 21 8850 55
rect 8884 21 8919 55
rect 8953 21 8988 55
rect 9022 21 9057 55
rect 9091 21 9126 55
rect 9160 21 9195 55
rect 9229 21 9264 55
rect 9298 21 9333 55
rect 9367 21 9402 55
rect 9436 21 9471 55
rect 9505 21 9540 55
rect 9574 21 9609 55
rect 9643 21 9678 55
rect 9712 21 9747 55
rect 9781 21 9816 55
rect 9850 21 9885 55
rect 9919 21 9954 55
rect 9988 21 10023 55
rect 10057 21 10092 55
rect 10126 21 10161 55
rect 10195 21 10230 55
rect 10264 21 10299 55
rect 10333 21 10368 55
rect 10402 21 10437 55
rect 10471 21 10506 55
rect 10540 21 10575 55
rect 10609 21 10643 55
rect 10677 21 10711 55
rect 10745 21 10779 55
rect 10813 21 10847 55
rect 10881 21 10915 55
rect 10949 21 10983 55
rect 11017 21 11051 55
rect 11085 21 11119 55
rect 11153 21 11187 55
rect 11221 21 11255 55
rect 11289 21 11323 55
rect 11357 21 11391 55
rect 11425 21 11459 55
rect 11493 21 11527 55
rect 11561 21 11595 55
rect 11629 21 11663 55
rect 11697 21 11731 55
rect 11765 21 11799 55
rect 11833 21 11867 55
rect 11901 21 11935 55
rect 11969 21 12003 55
rect 12037 21 12071 55
rect 12105 21 12139 55
rect 12173 21 12207 55
rect 12241 21 12275 55
rect 12309 21 12343 55
rect 12377 21 12411 55
rect 12445 21 12479 55
rect 12513 21 12547 55
rect 12581 21 12615 55
rect 12649 21 12683 55
rect 12717 21 12751 55
rect 12785 21 12819 55
rect 12853 21 12887 55
rect 12921 21 12955 55
rect 12989 21 13023 55
rect 13057 21 13091 55
rect 13125 21 13159 55
rect 13193 21 13227 55
rect 13261 21 13295 55
rect 13329 21 13363 55
rect 13397 21 13431 55
rect 13465 21 13499 55
rect 13533 21 13567 55
rect 13601 21 13635 55
rect 13669 21 13703 55
rect 13737 21 13771 55
rect 13805 21 13839 55
rect 13873 21 13907 55
rect 13941 21 13975 55
rect 14009 21 14043 55
rect 14077 21 14111 55
rect 14145 21 14179 55
rect 14213 21 14247 55
rect 14281 21 14315 55
rect 14349 21 14383 55
rect 14417 21 14451 55
rect 14485 21 14519 55
rect 14553 21 14587 55
rect 14621 21 14655 55
rect 14691 43 14723 55
rect 14769 43 14791 55
rect 14847 43 14859 55
rect 14925 43 14969 57
rect 15003 53 15117 57
rect 15003 43 15068 53
rect 14689 21 14723 43
rect 14757 21 14791 43
rect 14825 21 14859 43
rect 14893 21 15068 43
rect 7010 19 15068 21
rect 15102 19 15117 53
rect 7010 -11 7022 19
rect 5884 -9229 5918 -9191
<< viali >>
rect 131 16459 139 16493
rect 139 16459 165 16493
rect 204 16459 210 16493
rect 210 16459 238 16493
rect 277 16459 281 16493
rect 281 16459 311 16493
rect 350 16459 352 16493
rect 352 16459 384 16493
rect 423 16459 444 16493
rect 444 16459 457 16493
rect 496 16459 513 16493
rect 513 16459 530 16493
rect 569 16459 582 16493
rect 582 16459 603 16493
rect 642 16459 651 16493
rect 651 16459 676 16493
rect 715 16459 720 16493
rect 720 16459 749 16493
rect 788 16459 789 16493
rect 789 16459 822 16493
rect 861 16459 892 16493
rect 892 16459 895 16493
rect 934 16459 961 16493
rect 961 16459 968 16493
rect 1007 16459 1030 16493
rect 1030 16459 1041 16493
rect 1079 16459 1099 16493
rect 1099 16459 1113 16493
rect 1151 16459 1168 16493
rect 1168 16459 1185 16493
rect 1223 16459 1237 16493
rect 1237 16459 1257 16493
rect 1295 16459 1306 16493
rect 1306 16459 1329 16493
rect 1367 16459 1375 16493
rect 1375 16459 1401 16493
rect 1439 16459 1444 16493
rect 1444 16459 1473 16493
rect 1511 16459 1513 16493
rect 1513 16459 1545 16493
rect 1583 16459 1617 16493
rect 1655 16459 1686 16493
rect 1686 16459 1689 16493
rect 1727 16459 1755 16493
rect 1755 16459 1761 16493
rect 1799 16459 1824 16493
rect 1824 16459 1833 16493
rect 1871 16459 1893 16493
rect 1893 16459 1905 16493
rect 1943 16459 1962 16493
rect 1962 16459 1977 16493
rect 2015 16459 2031 16493
rect 2031 16459 2049 16493
rect 2087 16459 2100 16493
rect 2100 16459 2121 16493
rect 2159 16459 2169 16493
rect 2169 16459 2193 16493
rect 2231 16459 2238 16493
rect 2238 16459 2265 16493
rect 2303 16459 2307 16493
rect 2307 16459 2337 16493
rect 2375 16459 2376 16493
rect 2376 16459 2409 16493
rect 2447 16459 2479 16493
rect 2479 16459 2481 16493
rect 2519 16459 2548 16493
rect 2548 16459 2553 16493
rect 2591 16459 2617 16493
rect 2617 16459 2625 16493
rect 2663 16459 2686 16493
rect 2686 16459 2697 16493
rect 2735 16459 2755 16493
rect 2755 16459 2769 16493
rect 2807 16459 2824 16493
rect 2824 16459 2841 16493
rect 2879 16459 2893 16493
rect 2893 16459 2913 16493
rect 2951 16459 2962 16493
rect 2962 16459 2985 16493
rect 3023 16459 3030 16493
rect 3030 16459 3057 16493
rect 3095 16459 3098 16493
rect 3098 16459 3129 16493
rect 3167 16459 3200 16493
rect 3200 16459 3201 16493
rect 3239 16459 3268 16493
rect 3268 16459 3273 16493
rect 3311 16459 3336 16493
rect 3336 16459 3345 16493
rect 3383 16459 3404 16493
rect 3404 16459 3417 16493
rect 3455 16459 3472 16493
rect 3472 16459 3489 16493
rect 3527 16459 3540 16493
rect 3540 16459 3561 16493
rect 3599 16459 3608 16493
rect 3608 16459 3633 16493
rect 3671 16459 3676 16493
rect 3676 16459 3705 16493
rect 3743 16459 3744 16493
rect 3744 16459 3777 16493
rect 3815 16459 3846 16493
rect 3846 16459 3849 16493
rect 3887 16459 3914 16493
rect 3914 16459 3921 16493
rect 3959 16459 3982 16493
rect 3982 16459 3993 16493
rect 4031 16459 4050 16493
rect 4050 16459 4065 16493
rect 4103 16459 4118 16493
rect 4118 16459 4137 16493
rect 4175 16459 4186 16493
rect 4186 16459 4209 16493
rect 4247 16459 4254 16493
rect 4254 16459 4281 16493
rect 4319 16459 4322 16493
rect 4322 16459 4353 16493
rect 4391 16459 4424 16493
rect 4424 16459 4425 16493
rect 4463 16459 4492 16493
rect 4492 16459 4497 16493
rect 4535 16459 4560 16493
rect 4560 16459 4569 16493
rect 4607 16459 4628 16493
rect 4628 16459 4641 16493
rect 4679 16459 4696 16493
rect 4696 16459 4713 16493
rect 4751 16459 4764 16493
rect 4764 16459 4785 16493
rect 4823 16459 4832 16493
rect 4832 16459 4857 16493
rect 4895 16459 4900 16493
rect 4900 16459 4929 16493
rect 4967 16459 4968 16493
rect 4968 16459 5001 16493
rect 5039 16459 5070 16493
rect 5070 16459 5073 16493
rect 5111 16459 5138 16493
rect 5138 16459 5145 16493
rect 5183 16459 5206 16493
rect 5206 16459 5217 16493
rect 5255 16459 5274 16493
rect 5274 16459 5289 16493
rect 5327 16459 5342 16493
rect 5342 16459 5361 16493
rect 5399 16459 5410 16493
rect 5410 16459 5433 16493
rect 5471 16459 5478 16493
rect 5478 16459 5505 16493
rect 5543 16459 5546 16493
rect 5546 16459 5577 16493
rect 5615 16459 5648 16493
rect 5648 16459 5649 16493
rect 5687 16459 5716 16493
rect 5716 16459 5721 16493
rect 5759 16459 5784 16493
rect 5784 16459 5793 16493
rect 5831 16459 5852 16493
rect 5852 16459 5865 16493
rect 5903 16459 5920 16493
rect 5920 16459 5937 16493
rect 5975 16459 5988 16493
rect 5988 16459 6009 16493
rect 6047 16459 6056 16493
rect 6056 16459 6081 16493
rect 6119 16459 6124 16493
rect 6124 16459 6153 16493
rect 6191 16459 6192 16493
rect 6192 16459 6225 16493
rect 6263 16459 6294 16493
rect 6294 16459 6297 16493
rect 6335 16459 6362 16493
rect 6362 16459 6369 16493
rect 6407 16459 6430 16493
rect 6430 16459 6441 16493
rect 6479 16459 6498 16493
rect 6498 16459 6513 16493
rect 6551 16459 6566 16493
rect 6566 16459 6585 16493
rect 6623 16459 6634 16493
rect 6634 16459 6657 16493
rect 6695 16459 6702 16493
rect 6702 16459 6729 16493
rect 6767 16459 6770 16493
rect 6770 16459 6801 16493
rect 6839 16459 6872 16493
rect 6872 16459 6873 16493
rect 6911 16459 6940 16493
rect 6940 16459 6945 16493
rect 6983 16459 7008 16493
rect 7008 16459 7017 16493
rect 7055 16459 7076 16493
rect 7076 16459 7089 16493
rect 7127 16459 7144 16493
rect 7144 16459 7161 16493
rect 7199 16459 7212 16493
rect 7212 16459 7233 16493
rect 7271 16459 7280 16493
rect 7280 16459 7305 16493
rect 7343 16459 7348 16493
rect 7348 16459 7377 16493
rect 7415 16459 7416 16493
rect 7416 16459 7449 16493
rect 7487 16459 7518 16493
rect 7518 16459 7521 16493
rect 7559 16459 7586 16493
rect 7586 16459 7593 16493
rect 7631 16459 7654 16493
rect 7654 16459 7665 16493
rect 7703 16459 7722 16493
rect 7722 16459 7737 16493
rect 7775 16459 7790 16493
rect 7790 16459 7809 16493
rect 7847 16459 7858 16493
rect 7858 16459 7881 16493
rect 7919 16459 7926 16493
rect 7926 16459 7953 16493
rect 7991 16459 7994 16493
rect 7994 16459 8025 16493
rect 8063 16459 8096 16493
rect 8096 16459 8097 16493
rect 8135 16459 8164 16493
rect 8164 16459 8169 16493
rect 8207 16459 8232 16493
rect 8232 16459 8241 16493
rect 8279 16459 8300 16493
rect 8300 16459 8313 16493
rect 8351 16459 8368 16493
rect 8368 16459 8385 16493
rect 8423 16459 8436 16493
rect 8436 16459 8457 16493
rect 8495 16459 8504 16493
rect 8504 16459 8529 16493
rect 8567 16459 8572 16493
rect 8572 16459 8601 16493
rect 8639 16459 8640 16493
rect 8640 16459 8673 16493
rect 8711 16459 8742 16493
rect 8742 16459 8745 16493
rect 8783 16459 8810 16493
rect 8810 16459 8817 16493
rect 8855 16459 8878 16493
rect 8878 16459 8889 16493
rect 8927 16459 8946 16493
rect 8946 16459 8961 16493
rect 8999 16459 9014 16493
rect 9014 16459 9033 16493
rect 9071 16459 9082 16493
rect 9082 16459 9105 16493
rect 9143 16459 9150 16493
rect 9150 16459 9177 16493
rect 9215 16459 9218 16493
rect 9218 16459 9249 16493
rect 9287 16459 9320 16493
rect 9320 16459 9321 16493
rect 9359 16459 9388 16493
rect 9388 16459 9393 16493
rect 9431 16459 9456 16493
rect 9456 16459 9465 16493
rect 9503 16459 9524 16493
rect 9524 16459 9537 16493
rect 9575 16459 9592 16493
rect 9592 16459 9609 16493
rect 9647 16459 9660 16493
rect 9660 16459 9681 16493
rect 9719 16459 9728 16493
rect 9728 16459 9753 16493
rect 9791 16459 9796 16493
rect 9796 16459 9825 16493
rect 9863 16459 9864 16493
rect 9864 16459 9897 16493
rect 9935 16459 9966 16493
rect 9966 16459 9969 16493
rect 10007 16459 10034 16493
rect 10034 16459 10041 16493
rect 10079 16459 10102 16493
rect 10102 16459 10113 16493
rect 10151 16459 10170 16493
rect 10170 16459 10185 16493
rect 10223 16459 10238 16493
rect 10238 16459 10257 16493
rect 10295 16459 10306 16493
rect 10306 16459 10329 16493
rect 10367 16459 10374 16493
rect 10374 16459 10401 16493
rect 10439 16459 10442 16493
rect 10442 16459 10473 16493
rect 10511 16459 10544 16493
rect 10544 16459 10545 16493
rect 10583 16459 10612 16493
rect 10612 16459 10617 16493
rect 10655 16459 10680 16493
rect 10680 16459 10689 16493
rect 10727 16459 10748 16493
rect 10748 16459 10761 16493
rect 10799 16459 10816 16493
rect 10816 16459 10833 16493
rect 10871 16459 10884 16493
rect 10884 16459 10905 16493
rect 10943 16459 10952 16493
rect 10952 16459 10977 16493
rect 11015 16459 11020 16493
rect 11020 16459 11049 16493
rect 11087 16459 11088 16493
rect 11088 16459 11121 16493
rect 11159 16459 11190 16493
rect 11190 16459 11193 16493
rect 11231 16459 11258 16493
rect 11258 16459 11265 16493
rect 11303 16459 11326 16493
rect 11326 16459 11337 16493
rect 11375 16459 11394 16493
rect 11394 16459 11409 16493
rect 11447 16459 11462 16493
rect 11462 16459 11481 16493
rect 11519 16459 11530 16493
rect 11530 16459 11553 16493
rect 11591 16459 11598 16493
rect 11598 16459 11625 16493
rect 11663 16459 11666 16493
rect 11666 16459 11697 16493
rect 11735 16459 11768 16493
rect 11768 16459 11769 16493
rect 11807 16459 11836 16493
rect 11836 16459 11841 16493
rect 11879 16459 11904 16493
rect 11904 16459 11913 16493
rect 11951 16459 11972 16493
rect 11972 16459 11985 16493
rect 12023 16459 12040 16493
rect 12040 16459 12057 16493
rect 12095 16459 12108 16493
rect 12108 16459 12129 16493
rect 12167 16459 12176 16493
rect 12176 16459 12201 16493
rect 12239 16459 12244 16493
rect 12244 16459 12273 16493
rect 12311 16459 12312 16493
rect 12312 16459 12345 16493
rect 12383 16459 12414 16493
rect 12414 16459 12417 16493
rect 12455 16459 12482 16493
rect 12482 16459 12489 16493
rect 12527 16459 12550 16493
rect 12550 16459 12561 16493
rect 12599 16459 12618 16493
rect 12618 16459 12633 16493
rect 12671 16459 12686 16493
rect 12686 16459 12705 16493
rect 12743 16459 12754 16493
rect 12754 16459 12777 16493
rect 12815 16459 12822 16493
rect 12822 16459 12849 16493
rect 12887 16459 12890 16493
rect 12890 16459 12921 16493
rect 12959 16459 12992 16493
rect 12992 16459 12993 16493
rect 13031 16459 13060 16493
rect 13060 16459 13065 16493
rect 13103 16459 13128 16493
rect 13128 16459 13137 16493
rect 13175 16459 13196 16493
rect 13196 16459 13209 16493
rect 13247 16459 13264 16493
rect 13264 16459 13281 16493
rect 13319 16459 13332 16493
rect 13332 16459 13353 16493
rect 13391 16459 13400 16493
rect 13400 16459 13425 16493
rect 13463 16459 13468 16493
rect 13468 16459 13497 16493
rect 13535 16459 13536 16493
rect 13536 16459 13569 16493
rect 13607 16459 13638 16493
rect 13638 16459 13641 16493
rect 13679 16459 13706 16493
rect 13706 16459 13713 16493
rect 13751 16459 13774 16493
rect 13774 16459 13785 16493
rect 13823 16459 13842 16493
rect 13842 16459 13857 16493
rect 13895 16459 13910 16493
rect 13910 16459 13929 16493
rect 13967 16459 13978 16493
rect 13978 16459 14001 16493
rect 14039 16459 14046 16493
rect 14046 16459 14073 16493
rect 14111 16459 14114 16493
rect 14114 16459 14145 16493
rect 14183 16459 14216 16493
rect 14216 16459 14217 16493
rect 14255 16459 14284 16493
rect 14284 16459 14289 16493
rect 14327 16459 14352 16493
rect 14352 16459 14361 16493
rect 14399 16469 14420 16493
rect 14420 16469 14433 16493
rect 14471 16469 14492 16493
rect 14492 16469 14505 16493
rect 14543 16469 14564 16493
rect 14564 16469 14577 16493
rect 14615 16469 14636 16493
rect 14636 16469 14649 16493
rect 14687 16469 14708 16493
rect 14708 16469 14721 16493
rect 14759 16469 14780 16493
rect 14780 16469 14793 16493
rect 14831 16469 14852 16493
rect 14852 16469 14865 16493
rect 14903 16469 14924 16493
rect 14924 16469 14937 16493
rect 14399 16459 14433 16469
rect 14471 16459 14505 16469
rect 14543 16459 14577 16469
rect 14615 16459 14649 16469
rect 14687 16459 14721 16469
rect 14759 16459 14793 16469
rect 14831 16459 14865 16469
rect 14903 16459 14937 16469
rect 59 16391 68 16405
rect 68 16391 93 16405
rect 131 16391 139 16405
rect 139 16391 165 16405
rect 59 16371 93 16391
rect 131 16371 165 16391
rect 3882 15969 3914 15980
rect 3914 15969 3916 15980
rect 3955 15969 3982 15980
rect 3982 15969 3989 15980
rect 4028 15969 4050 15980
rect 4050 15969 4062 15980
rect 4101 15969 4118 15980
rect 4118 15969 4135 15980
rect 4174 15969 4186 15980
rect 4186 15969 4208 15980
rect 4247 15969 4254 15980
rect 4254 15969 4281 15980
rect 4320 15969 4322 15980
rect 4322 15969 4354 15980
rect 4393 15969 4424 15980
rect 4424 15969 4427 15980
rect 4466 15969 4492 15980
rect 4492 15969 4500 15980
rect 4539 15969 4560 15980
rect 4560 15969 4573 15980
rect 4612 15969 4628 15980
rect 4628 15969 4646 15980
rect 4685 15969 4696 15980
rect 4696 15969 4719 15980
rect 4758 15969 4764 15980
rect 4764 15969 4792 15980
rect 4831 15969 4832 15980
rect 4832 15969 4865 15980
rect 4904 15969 4934 15980
rect 4934 15969 4938 15980
rect 4977 15969 5002 15980
rect 5002 15969 5011 15980
rect 5050 15969 5070 15980
rect 5070 15969 5084 15980
rect 5123 15969 5138 15980
rect 5138 15969 5157 15980
rect 5196 15969 5206 15980
rect 5206 15969 5230 15980
rect 5269 15969 5274 15980
rect 5274 15969 5303 15980
rect 3882 15946 3916 15969
rect 3955 15946 3989 15969
rect 4028 15946 4062 15969
rect 4101 15946 4135 15969
rect 4174 15946 4208 15969
rect 4247 15946 4281 15969
rect 4320 15946 4354 15969
rect 4393 15946 4427 15969
rect 4466 15946 4500 15969
rect 4539 15946 4573 15969
rect 4612 15946 4646 15969
rect 4685 15946 4719 15969
rect 4758 15946 4792 15969
rect 4831 15946 4865 15969
rect 4904 15946 4938 15969
rect 4977 15946 5011 15969
rect 5050 15946 5084 15969
rect 5123 15946 5157 15969
rect 5196 15946 5230 15969
rect 5269 15946 5303 15969
rect 5342 15946 5376 15980
rect 5415 15969 5444 15980
rect 5444 15969 5449 15980
rect 5488 15969 5512 15980
rect 5512 15969 5522 15980
rect 5561 15969 5580 15980
rect 5580 15969 5595 15980
rect 5634 15969 5648 15980
rect 5648 15969 5668 15980
rect 5707 15969 5716 15980
rect 5716 15969 5741 15980
rect 5780 15969 5784 15980
rect 5784 15969 5814 15980
rect 5853 15969 5886 15980
rect 5886 15969 5887 15980
rect 5926 15969 5954 15980
rect 5954 15969 5960 15980
rect 5999 15969 6022 15980
rect 6022 15969 6033 15980
rect 6072 15969 6090 15980
rect 6090 15969 6106 15980
rect 6145 15969 6158 15980
rect 6158 15969 6179 15980
rect 6218 15969 6226 15980
rect 6226 15969 6252 15980
rect 6291 15969 6294 15980
rect 6294 15969 6325 15980
rect 6364 15969 6396 15980
rect 6396 15969 6398 15980
rect 6437 15969 6464 15980
rect 6464 15969 6471 15980
rect 6510 15969 6532 15980
rect 6532 15969 6544 15980
rect 6583 15969 6600 15980
rect 6600 15969 6617 15980
rect 6656 15969 6668 15980
rect 6668 15969 6690 15980
rect 6729 15969 6736 15980
rect 6736 15969 6763 15980
rect 6802 15969 6804 15980
rect 6804 15969 6836 15980
rect 6875 15969 6906 15980
rect 6906 15969 6909 15980
rect 6948 15969 6974 15980
rect 6974 15969 6982 15980
rect 7021 15969 7042 15980
rect 7042 15969 7055 15980
rect 7094 15969 7110 15980
rect 7110 15969 7128 15980
rect 7167 15969 7178 15980
rect 7178 15969 7201 15980
rect 7240 15969 7246 15980
rect 7246 15969 7274 15980
rect 7313 15969 7314 15980
rect 7314 15969 7347 15980
rect 7386 15969 7416 15980
rect 7416 15969 7420 15980
rect 7459 15969 7484 15980
rect 7484 15969 7493 15980
rect 7532 15969 7552 15980
rect 7552 15969 7566 15980
rect 7605 15969 7620 15980
rect 7620 15969 7639 15980
rect 7678 15969 7688 15980
rect 7688 15969 7712 15980
rect 7751 15969 7756 15980
rect 7756 15969 7785 15980
rect 7824 15969 7858 15980
rect 7897 15969 7926 15980
rect 7926 15969 7931 15980
rect 7970 15969 7994 15980
rect 7994 15969 8004 15980
rect 8043 15969 8062 15980
rect 8062 15969 8077 15980
rect 8116 15969 8130 15980
rect 8130 15969 8150 15980
rect 8189 15969 8198 15980
rect 8198 15969 8223 15980
rect 8262 15969 8266 15980
rect 8266 15969 8296 15980
rect 8335 15969 8368 15980
rect 8368 15969 8369 15980
rect 8408 15969 8436 15980
rect 8436 15969 8442 15980
rect 8481 15969 8504 15980
rect 8504 15969 8515 15980
rect 8554 15969 8572 15980
rect 8572 15969 8588 15980
rect 8627 15969 8640 15980
rect 8640 15969 8661 15980
rect 8699 15969 8708 15980
rect 8708 15969 8733 15980
rect 8771 15969 8776 15980
rect 8776 15969 8805 15980
rect 8843 15969 8844 15980
rect 8844 15969 8877 15980
rect 8915 15969 8946 15980
rect 8946 15969 8949 15980
rect 8987 15969 9014 15980
rect 9014 15969 9021 15980
rect 9059 15969 9082 15980
rect 9082 15969 9093 15980
rect 9131 15969 9150 15980
rect 9150 15969 9165 15980
rect 9203 15969 9218 15980
rect 9218 15969 9237 15980
rect 9275 15969 9286 15980
rect 9286 15969 9309 15980
rect 9347 15969 9354 15980
rect 9354 15969 9381 15980
rect 9419 15969 9422 15980
rect 9422 15969 9453 15980
rect 9491 15969 9524 15980
rect 9524 15969 9525 15980
rect 9563 15969 9592 15980
rect 9592 15969 9597 15980
rect 9635 15969 9660 15980
rect 9660 15969 9669 15980
rect 9707 15969 9728 15980
rect 9728 15969 9741 15980
rect 9779 15969 9796 15980
rect 9796 15969 9813 15980
rect 9851 15969 9864 15980
rect 9864 15969 9885 15980
rect 9923 15969 9932 15980
rect 9932 15969 9957 15980
rect 9995 15969 10000 15980
rect 10000 15969 10029 15980
rect 10067 15969 10068 15980
rect 10068 15969 10101 15980
rect 10139 15969 10170 15980
rect 10170 15969 10173 15980
rect 10211 15969 10238 15980
rect 10238 15969 10245 15980
rect 10283 15969 10306 15980
rect 10306 15969 10317 15980
rect 10355 15969 10374 15980
rect 10374 15969 10389 15980
rect 10427 15969 10442 15980
rect 10442 15969 10461 15980
rect 10499 15969 10510 15980
rect 10510 15969 10533 15980
rect 10571 15969 10578 15980
rect 10578 15969 10605 15980
rect 10643 15969 10646 15980
rect 10646 15969 10677 15980
rect 10715 15969 10748 15980
rect 10748 15969 10749 15980
rect 10787 15969 10816 15980
rect 10816 15969 10821 15980
rect 10859 15969 10884 15980
rect 10884 15969 10893 15980
rect 10931 15969 10952 15980
rect 10952 15969 10965 15980
rect 11003 15969 11020 15980
rect 11020 15969 11037 15980
rect 11075 15969 11088 15980
rect 11088 15969 11109 15980
rect 11147 15969 11156 15980
rect 11156 15969 11181 15980
rect 11219 15969 11224 15980
rect 11224 15969 11253 15980
rect 11291 15969 11292 15980
rect 11292 15969 11325 15980
rect 11363 15969 11394 15980
rect 11394 15969 11397 15980
rect 11435 15969 11462 15980
rect 11462 15969 11469 15980
rect 11507 15969 11530 15980
rect 11530 15969 11541 15980
rect 11579 15969 11598 15980
rect 11598 15969 11613 15980
rect 11651 15969 11666 15980
rect 11666 15969 11685 15980
rect 11723 15969 11734 15980
rect 11734 15969 11757 15980
rect 11795 15969 11802 15980
rect 11802 15969 11829 15980
rect 11867 15969 11870 15980
rect 11870 15969 11901 15980
rect 11939 15969 11972 15980
rect 11972 15969 11973 15980
rect 12011 15969 12040 15980
rect 12040 15969 12045 15980
rect 12083 15969 12108 15980
rect 12108 15969 12117 15980
rect 12155 15969 12176 15980
rect 12176 15969 12189 15980
rect 12227 15969 12244 15980
rect 12244 15969 12261 15980
rect 12299 15969 12312 15980
rect 12312 15969 12333 15980
rect 12371 15969 12380 15980
rect 12380 15969 12405 15980
rect 12443 15969 12448 15980
rect 12448 15969 12477 15980
rect 12515 15969 12516 15980
rect 12516 15969 12549 15980
rect 12587 15969 12618 15980
rect 12618 15969 12621 15980
rect 12659 15969 12686 15980
rect 12686 15969 12693 15980
rect 12731 15969 12754 15980
rect 12754 15969 12765 15980
rect 12803 15969 12822 15980
rect 12822 15969 12837 15980
rect 12875 15969 12890 15980
rect 12890 15969 12909 15980
rect 12947 15969 12958 15980
rect 12958 15969 12981 15980
rect 13019 15969 13026 15980
rect 13026 15969 13053 15980
rect 13091 15969 13094 15980
rect 13094 15969 13125 15980
rect 13163 15969 13196 15980
rect 13196 15969 13197 15980
rect 13235 15969 13264 15980
rect 13264 15969 13269 15980
rect 13307 15969 13332 15980
rect 13332 15969 13341 15980
rect 13379 15969 13400 15980
rect 13400 15969 13413 15980
rect 13451 15969 13468 15980
rect 13468 15969 13485 15980
rect 13523 15969 13536 15980
rect 13536 15969 13557 15980
rect 13595 15969 13604 15980
rect 13604 15969 13629 15980
rect 13667 15969 13672 15980
rect 13672 15969 13701 15980
rect 13739 15969 13740 15980
rect 13740 15969 13773 15980
rect 13811 15969 13842 15980
rect 13842 15969 13845 15980
rect 13883 15969 13910 15980
rect 13910 15969 13917 15980
rect 13955 15969 13978 15980
rect 13978 15969 13989 15980
rect 14027 15969 14046 15980
rect 14046 15969 14061 15980
rect 14099 15969 14114 15980
rect 14114 15969 14133 15980
rect 14171 15969 14182 15980
rect 14182 15969 14205 15980
rect 14243 15969 14250 15980
rect 14250 15969 14277 15980
rect 14315 15969 14318 15980
rect 14318 15969 14349 15980
rect 5415 15946 5449 15969
rect 5488 15946 5522 15969
rect 5561 15946 5595 15969
rect 5634 15946 5668 15969
rect 5707 15946 5741 15969
rect 5780 15946 5814 15969
rect 5853 15946 5887 15969
rect 5926 15946 5960 15969
rect 5999 15946 6033 15969
rect 6072 15946 6106 15969
rect 6145 15946 6179 15969
rect 6218 15946 6252 15969
rect 6291 15946 6325 15969
rect 6364 15946 6398 15969
rect 6437 15946 6471 15969
rect 6510 15946 6544 15969
rect 6583 15946 6617 15969
rect 6656 15946 6690 15969
rect 6729 15946 6763 15969
rect 6802 15946 6836 15969
rect 6875 15946 6909 15969
rect 6948 15946 6982 15969
rect 7021 15946 7055 15969
rect 7094 15946 7128 15969
rect 7167 15946 7201 15969
rect 7240 15946 7274 15969
rect 7313 15946 7347 15969
rect 7386 15946 7420 15969
rect 7459 15946 7493 15969
rect 7532 15946 7566 15969
rect 7605 15946 7639 15969
rect 7678 15946 7712 15969
rect 7751 15946 7785 15969
rect 7824 15946 7858 15969
rect 7897 15946 7931 15969
rect 7970 15946 8004 15969
rect 8043 15946 8077 15969
rect 8116 15946 8150 15969
rect 8189 15946 8223 15969
rect 8262 15946 8296 15969
rect 8335 15946 8369 15969
rect 8408 15946 8442 15969
rect 8481 15946 8515 15969
rect 8554 15946 8588 15969
rect 8627 15946 8661 15969
rect 8699 15946 8733 15969
rect 8771 15946 8805 15969
rect 8843 15946 8877 15969
rect 8915 15946 8949 15969
rect 8987 15946 9021 15969
rect 9059 15946 9093 15969
rect 9131 15946 9165 15969
rect 9203 15946 9237 15969
rect 9275 15946 9309 15969
rect 9347 15946 9381 15969
rect 9419 15946 9453 15969
rect 9491 15946 9525 15969
rect 9563 15946 9597 15969
rect 9635 15946 9669 15969
rect 9707 15946 9741 15969
rect 9779 15946 9813 15969
rect 9851 15946 9885 15969
rect 9923 15946 9957 15969
rect 9995 15946 10029 15969
rect 10067 15946 10101 15969
rect 10139 15946 10173 15969
rect 10211 15946 10245 15969
rect 10283 15946 10317 15969
rect 10355 15946 10389 15969
rect 10427 15946 10461 15969
rect 10499 15946 10533 15969
rect 10571 15946 10605 15969
rect 10643 15946 10677 15969
rect 10715 15946 10749 15969
rect 10787 15946 10821 15969
rect 10859 15946 10893 15969
rect 10931 15946 10965 15969
rect 11003 15946 11037 15969
rect 11075 15946 11109 15969
rect 11147 15946 11181 15969
rect 11219 15946 11253 15969
rect 11291 15946 11325 15969
rect 11363 15946 11397 15969
rect 11435 15946 11469 15969
rect 11507 15946 11541 15969
rect 11579 15946 11613 15969
rect 11651 15946 11685 15969
rect 11723 15946 11757 15969
rect 11795 15946 11829 15969
rect 11867 15946 11901 15969
rect 11939 15946 11973 15969
rect 12011 15946 12045 15969
rect 12083 15946 12117 15969
rect 12155 15946 12189 15969
rect 12227 15946 12261 15969
rect 12299 15946 12333 15969
rect 12371 15946 12405 15969
rect 12443 15946 12477 15969
rect 12515 15946 12549 15969
rect 12587 15946 12621 15969
rect 12659 15946 12693 15969
rect 12731 15946 12765 15969
rect 12803 15946 12837 15969
rect 12875 15946 12909 15969
rect 12947 15946 12981 15969
rect 13019 15946 13053 15969
rect 13091 15946 13125 15969
rect 13163 15946 13197 15969
rect 13235 15946 13269 15969
rect 13307 15946 13341 15969
rect 13379 15946 13413 15969
rect 13451 15946 13485 15969
rect 13523 15946 13557 15969
rect 13595 15946 13629 15969
rect 13667 15946 13701 15969
rect 13739 15946 13773 15969
rect 13811 15946 13845 15969
rect 13883 15946 13917 15969
rect 13955 15946 13989 15969
rect 14027 15946 14061 15969
rect 14099 15946 14133 15969
rect 14171 15946 14205 15969
rect 14243 15946 14277 15969
rect 14315 15946 14349 15969
rect 14387 15951 14421 15980
rect 14459 15951 14493 15980
rect 14531 15951 14565 15980
rect 14603 15951 14637 15980
rect 14675 15951 14709 15980
rect 14747 15951 14781 15980
rect 14819 15951 14853 15980
rect 14891 15951 14925 15980
rect 14387 15946 14420 15951
rect 14420 15946 14421 15951
rect 14459 15946 14492 15951
rect 14492 15946 14493 15951
rect 14531 15946 14564 15951
rect 14564 15946 14565 15951
rect 14603 15946 14636 15951
rect 14636 15946 14637 15951
rect 14675 15946 14708 15951
rect 14708 15946 14709 15951
rect 14747 15946 14780 15951
rect 14780 15946 14781 15951
rect 14819 15946 14852 15951
rect 14852 15946 14853 15951
rect 14891 15946 14924 15951
rect 14924 15946 14925 15951
rect 3882 15899 3914 15906
rect 3914 15899 3916 15906
rect 3955 15899 3982 15906
rect 3982 15899 3989 15906
rect 4028 15899 4050 15906
rect 4050 15899 4062 15906
rect 4101 15899 4118 15906
rect 4118 15899 4135 15906
rect 4174 15899 4186 15906
rect 4186 15899 4208 15906
rect 4247 15899 4254 15906
rect 4254 15899 4281 15906
rect 4320 15899 4322 15906
rect 4322 15899 4354 15906
rect 4393 15899 4424 15906
rect 4424 15899 4427 15906
rect 4466 15899 4492 15906
rect 4492 15899 4500 15906
rect 4539 15899 4560 15906
rect 4560 15899 4573 15906
rect 4612 15899 4628 15906
rect 4628 15899 4646 15906
rect 4685 15899 4696 15906
rect 4696 15899 4719 15906
rect 4758 15899 4764 15906
rect 4764 15899 4792 15906
rect 4831 15899 4832 15906
rect 4832 15899 4865 15906
rect 4904 15899 4934 15906
rect 4934 15899 4938 15906
rect 4977 15899 5002 15906
rect 5002 15899 5011 15906
rect 5050 15899 5070 15906
rect 5070 15899 5084 15906
rect 5123 15899 5138 15906
rect 5138 15899 5157 15906
rect 5196 15899 5206 15906
rect 5206 15899 5230 15906
rect 5269 15899 5274 15906
rect 5274 15899 5303 15906
rect 3882 15872 3916 15899
rect 3955 15872 3989 15899
rect 4028 15872 4062 15899
rect 4101 15872 4135 15899
rect 4174 15872 4208 15899
rect 4247 15872 4281 15899
rect 4320 15872 4354 15899
rect 4393 15872 4427 15899
rect 4466 15872 4500 15899
rect 4539 15872 4573 15899
rect 4612 15872 4646 15899
rect 4685 15872 4719 15899
rect 4758 15872 4792 15899
rect 4831 15872 4865 15899
rect 4904 15872 4938 15899
rect 4977 15872 5011 15899
rect 5050 15872 5084 15899
rect 5123 15872 5157 15899
rect 5196 15872 5230 15899
rect 5269 15872 5303 15899
rect 5342 15872 5376 15906
rect 5415 15899 5444 15906
rect 5444 15899 5449 15906
rect 5488 15899 5512 15906
rect 5512 15899 5522 15906
rect 5561 15899 5580 15906
rect 5580 15899 5595 15906
rect 5634 15899 5648 15906
rect 5648 15899 5668 15906
rect 5707 15899 5716 15906
rect 5716 15899 5741 15906
rect 5780 15899 5784 15906
rect 5784 15899 5814 15906
rect 5853 15899 5886 15906
rect 5886 15899 5887 15906
rect 5926 15899 5954 15906
rect 5954 15899 5960 15906
rect 5999 15899 6022 15906
rect 6022 15899 6033 15906
rect 6072 15899 6090 15906
rect 6090 15899 6106 15906
rect 6145 15899 6158 15906
rect 6158 15899 6179 15906
rect 6218 15899 6226 15906
rect 6226 15899 6252 15906
rect 6291 15899 6294 15906
rect 6294 15899 6325 15906
rect 6364 15899 6396 15906
rect 6396 15899 6398 15906
rect 6437 15899 6464 15906
rect 6464 15899 6471 15906
rect 6510 15899 6532 15906
rect 6532 15899 6544 15906
rect 6583 15899 6600 15906
rect 6600 15899 6617 15906
rect 6656 15899 6668 15906
rect 6668 15899 6690 15906
rect 6729 15899 6736 15906
rect 6736 15899 6763 15906
rect 6802 15899 6804 15906
rect 6804 15899 6836 15906
rect 6875 15899 6906 15906
rect 6906 15899 6909 15906
rect 6948 15899 6974 15906
rect 6974 15899 6982 15906
rect 7021 15899 7042 15906
rect 7042 15899 7055 15906
rect 7094 15899 7110 15906
rect 7110 15899 7128 15906
rect 7167 15899 7178 15906
rect 7178 15899 7201 15906
rect 7240 15899 7246 15906
rect 7246 15899 7274 15906
rect 7313 15899 7314 15906
rect 7314 15899 7347 15906
rect 7386 15899 7416 15906
rect 7416 15899 7420 15906
rect 7459 15899 7484 15906
rect 7484 15899 7493 15906
rect 7532 15899 7552 15906
rect 7552 15899 7566 15906
rect 7605 15899 7620 15906
rect 7620 15899 7639 15906
rect 7678 15899 7688 15906
rect 7688 15899 7712 15906
rect 7751 15899 7756 15906
rect 7756 15899 7785 15906
rect 7824 15899 7858 15906
rect 7897 15899 7926 15906
rect 7926 15899 7931 15906
rect 7970 15899 7994 15906
rect 7994 15899 8004 15906
rect 8043 15899 8062 15906
rect 8062 15899 8077 15906
rect 8116 15899 8130 15906
rect 8130 15899 8150 15906
rect 8189 15899 8198 15906
rect 8198 15899 8223 15906
rect 8262 15899 8266 15906
rect 8266 15899 8296 15906
rect 8335 15899 8368 15906
rect 8368 15899 8369 15906
rect 8408 15899 8436 15906
rect 8436 15899 8442 15906
rect 8481 15899 8504 15906
rect 8504 15899 8515 15906
rect 8554 15899 8572 15906
rect 8572 15899 8588 15906
rect 8627 15899 8640 15906
rect 8640 15899 8661 15906
rect 8699 15899 8708 15906
rect 8708 15899 8733 15906
rect 8771 15899 8776 15906
rect 8776 15899 8805 15906
rect 8843 15899 8844 15906
rect 8844 15899 8877 15906
rect 8915 15899 8946 15906
rect 8946 15899 8949 15906
rect 8987 15899 9014 15906
rect 9014 15899 9021 15906
rect 9059 15899 9082 15906
rect 9082 15899 9093 15906
rect 9131 15899 9150 15906
rect 9150 15899 9165 15906
rect 9203 15899 9218 15906
rect 9218 15899 9237 15906
rect 9275 15899 9286 15906
rect 9286 15899 9309 15906
rect 9347 15899 9354 15906
rect 9354 15899 9381 15906
rect 9419 15899 9422 15906
rect 9422 15899 9453 15906
rect 9491 15899 9524 15906
rect 9524 15899 9525 15906
rect 9563 15899 9592 15906
rect 9592 15899 9597 15906
rect 9635 15899 9660 15906
rect 9660 15899 9669 15906
rect 9707 15899 9728 15906
rect 9728 15899 9741 15906
rect 9779 15899 9796 15906
rect 9796 15899 9813 15906
rect 9851 15899 9864 15906
rect 9864 15899 9885 15906
rect 9923 15899 9932 15906
rect 9932 15899 9957 15906
rect 9995 15899 10000 15906
rect 10000 15899 10029 15906
rect 10067 15899 10068 15906
rect 10068 15899 10101 15906
rect 10139 15899 10170 15906
rect 10170 15899 10173 15906
rect 10211 15899 10238 15906
rect 10238 15899 10245 15906
rect 10283 15899 10306 15906
rect 10306 15899 10317 15906
rect 10355 15899 10374 15906
rect 10374 15899 10389 15906
rect 10427 15899 10442 15906
rect 10442 15899 10461 15906
rect 10499 15899 10510 15906
rect 10510 15899 10533 15906
rect 10571 15899 10578 15906
rect 10578 15899 10605 15906
rect 10643 15899 10646 15906
rect 10646 15899 10677 15906
rect 10715 15899 10748 15906
rect 10748 15899 10749 15906
rect 10787 15899 10816 15906
rect 10816 15899 10821 15906
rect 10859 15899 10884 15906
rect 10884 15899 10893 15906
rect 10931 15899 10952 15906
rect 10952 15899 10965 15906
rect 11003 15899 11020 15906
rect 11020 15899 11037 15906
rect 11075 15899 11088 15906
rect 11088 15899 11109 15906
rect 11147 15899 11156 15906
rect 11156 15899 11181 15906
rect 11219 15899 11224 15906
rect 11224 15899 11253 15906
rect 11291 15899 11292 15906
rect 11292 15899 11325 15906
rect 11363 15899 11394 15906
rect 11394 15899 11397 15906
rect 11435 15899 11462 15906
rect 11462 15899 11469 15906
rect 11507 15899 11530 15906
rect 11530 15899 11541 15906
rect 11579 15899 11598 15906
rect 11598 15899 11613 15906
rect 11651 15899 11666 15906
rect 11666 15899 11685 15906
rect 11723 15899 11734 15906
rect 11734 15899 11757 15906
rect 11795 15899 11802 15906
rect 11802 15899 11829 15906
rect 11867 15899 11870 15906
rect 11870 15899 11901 15906
rect 11939 15899 11972 15906
rect 11972 15899 11973 15906
rect 12011 15899 12040 15906
rect 12040 15899 12045 15906
rect 12083 15899 12108 15906
rect 12108 15899 12117 15906
rect 12155 15899 12176 15906
rect 12176 15899 12189 15906
rect 12227 15899 12244 15906
rect 12244 15899 12261 15906
rect 12299 15899 12312 15906
rect 12312 15899 12333 15906
rect 12371 15899 12380 15906
rect 12380 15899 12405 15906
rect 12443 15899 12448 15906
rect 12448 15899 12477 15906
rect 12515 15899 12516 15906
rect 12516 15899 12549 15906
rect 12587 15899 12618 15906
rect 12618 15899 12621 15906
rect 12659 15899 12686 15906
rect 12686 15899 12693 15906
rect 12731 15899 12754 15906
rect 12754 15899 12765 15906
rect 12803 15899 12822 15906
rect 12822 15899 12837 15906
rect 12875 15899 12890 15906
rect 12890 15899 12909 15906
rect 12947 15899 12958 15906
rect 12958 15899 12981 15906
rect 13019 15899 13026 15906
rect 13026 15899 13053 15906
rect 13091 15899 13094 15906
rect 13094 15899 13125 15906
rect 13163 15899 13196 15906
rect 13196 15899 13197 15906
rect 13235 15899 13264 15906
rect 13264 15899 13269 15906
rect 13307 15899 13332 15906
rect 13332 15899 13341 15906
rect 13379 15899 13400 15906
rect 13400 15899 13413 15906
rect 13451 15899 13468 15906
rect 13468 15899 13485 15906
rect 13523 15899 13536 15906
rect 13536 15899 13557 15906
rect 13595 15899 13604 15906
rect 13604 15899 13629 15906
rect 13667 15899 13672 15906
rect 13672 15899 13701 15906
rect 13739 15899 13740 15906
rect 13740 15899 13773 15906
rect 13811 15899 13842 15906
rect 13842 15899 13845 15906
rect 13883 15899 13910 15906
rect 13910 15899 13917 15906
rect 13955 15899 13978 15906
rect 13978 15899 13989 15906
rect 14027 15899 14046 15906
rect 14046 15899 14061 15906
rect 14099 15899 14114 15906
rect 14114 15899 14133 15906
rect 14171 15899 14182 15906
rect 14182 15899 14205 15906
rect 14243 15899 14250 15906
rect 14250 15899 14277 15906
rect 14315 15899 14318 15906
rect 14318 15899 14349 15906
rect 5415 15872 5449 15899
rect 5488 15872 5522 15899
rect 5561 15872 5595 15899
rect 5634 15872 5668 15899
rect 5707 15872 5741 15899
rect 5780 15872 5814 15899
rect 5853 15872 5887 15899
rect 5926 15872 5960 15899
rect 5999 15872 6033 15899
rect 6072 15872 6106 15899
rect 6145 15872 6179 15899
rect 6218 15872 6252 15899
rect 6291 15872 6325 15899
rect 6364 15872 6398 15899
rect 6437 15872 6471 15899
rect 6510 15872 6544 15899
rect 6583 15872 6617 15899
rect 6656 15872 6690 15899
rect 6729 15872 6763 15899
rect 6802 15872 6836 15899
rect 6875 15872 6909 15899
rect 6948 15872 6982 15899
rect 7021 15872 7055 15899
rect 7094 15872 7128 15899
rect 7167 15872 7201 15899
rect 7240 15872 7274 15899
rect 7313 15872 7347 15899
rect 7386 15872 7420 15899
rect 7459 15872 7493 15899
rect 7532 15872 7566 15899
rect 7605 15872 7639 15899
rect 7678 15872 7712 15899
rect 7751 15872 7785 15899
rect 7824 15872 7858 15899
rect 7897 15872 7931 15899
rect 7970 15872 8004 15899
rect 8043 15872 8077 15899
rect 8116 15872 8150 15899
rect 8189 15872 8223 15899
rect 8262 15872 8296 15899
rect 8335 15872 8369 15899
rect 8408 15872 8442 15899
rect 8481 15872 8515 15899
rect 8554 15872 8588 15899
rect 8627 15872 8661 15899
rect 8699 15872 8733 15899
rect 8771 15872 8805 15899
rect 8843 15872 8877 15899
rect 8915 15872 8949 15899
rect 8987 15872 9021 15899
rect 9059 15872 9093 15899
rect 9131 15872 9165 15899
rect 9203 15872 9237 15899
rect 9275 15872 9309 15899
rect 9347 15872 9381 15899
rect 9419 15872 9453 15899
rect 9491 15872 9525 15899
rect 9563 15872 9597 15899
rect 9635 15872 9669 15899
rect 9707 15872 9741 15899
rect 9779 15872 9813 15899
rect 9851 15872 9885 15899
rect 9923 15872 9957 15899
rect 9995 15872 10029 15899
rect 10067 15872 10101 15899
rect 10139 15872 10173 15899
rect 10211 15872 10245 15899
rect 10283 15872 10317 15899
rect 10355 15872 10389 15899
rect 10427 15872 10461 15899
rect 10499 15872 10533 15899
rect 10571 15872 10605 15899
rect 10643 15872 10677 15899
rect 10715 15872 10749 15899
rect 10787 15872 10821 15899
rect 10859 15872 10893 15899
rect 10931 15872 10965 15899
rect 11003 15872 11037 15899
rect 11075 15872 11109 15899
rect 11147 15872 11181 15899
rect 11219 15872 11253 15899
rect 11291 15872 11325 15899
rect 11363 15872 11397 15899
rect 11435 15872 11469 15899
rect 11507 15872 11541 15899
rect 11579 15872 11613 15899
rect 11651 15872 11685 15899
rect 11723 15872 11757 15899
rect 11795 15872 11829 15899
rect 11867 15872 11901 15899
rect 11939 15872 11973 15899
rect 12011 15872 12045 15899
rect 12083 15872 12117 15899
rect 12155 15872 12189 15899
rect 12227 15872 12261 15899
rect 12299 15872 12333 15899
rect 12371 15872 12405 15899
rect 12443 15872 12477 15899
rect 12515 15872 12549 15899
rect 12587 15872 12621 15899
rect 12659 15872 12693 15899
rect 12731 15872 12765 15899
rect 12803 15872 12837 15899
rect 12875 15872 12909 15899
rect 12947 15872 12981 15899
rect 13019 15872 13053 15899
rect 13091 15872 13125 15899
rect 13163 15872 13197 15899
rect 13235 15872 13269 15899
rect 13307 15872 13341 15899
rect 13379 15872 13413 15899
rect 13451 15872 13485 15899
rect 13523 15872 13557 15899
rect 13595 15872 13629 15899
rect 13667 15872 13701 15899
rect 13739 15872 13773 15899
rect 13811 15872 13845 15899
rect 13883 15872 13917 15899
rect 13955 15872 13989 15899
rect 14027 15872 14061 15899
rect 14099 15872 14133 15899
rect 14171 15872 14205 15899
rect 14243 15872 14277 15899
rect 14315 15872 14349 15899
rect 14387 15882 14421 15906
rect 14459 15882 14493 15906
rect 14531 15882 14565 15906
rect 14603 15882 14637 15906
rect 14675 15882 14709 15906
rect 14747 15882 14781 15906
rect 14819 15882 14853 15906
rect 14891 15882 14925 15906
rect 14387 15872 14420 15882
rect 14420 15872 14421 15882
rect 14459 15872 14492 15882
rect 14492 15872 14493 15882
rect 14531 15872 14564 15882
rect 14564 15872 14565 15882
rect 14603 15872 14636 15882
rect 14636 15872 14637 15882
rect 14675 15872 14708 15882
rect 14708 15872 14709 15882
rect 14747 15872 14780 15882
rect 14780 15872 14781 15882
rect 14819 15872 14852 15882
rect 14852 15872 14853 15882
rect 14891 15872 14924 15882
rect 14924 15872 14925 15882
rect 3882 15829 3914 15832
rect 3914 15829 3916 15832
rect 3955 15829 3982 15832
rect 3982 15829 3989 15832
rect 4028 15829 4050 15832
rect 4050 15829 4062 15832
rect 4101 15829 4118 15832
rect 4118 15829 4135 15832
rect 4174 15829 4186 15832
rect 4186 15829 4208 15832
rect 4247 15829 4254 15832
rect 4254 15829 4281 15832
rect 4320 15829 4322 15832
rect 4322 15829 4354 15832
rect 4393 15829 4424 15832
rect 4424 15829 4427 15832
rect 4466 15829 4492 15832
rect 4492 15829 4500 15832
rect 4539 15829 4560 15832
rect 4560 15829 4573 15832
rect 4612 15829 4628 15832
rect 4628 15829 4646 15832
rect 4685 15829 4696 15832
rect 4696 15829 4719 15832
rect 4758 15829 4764 15832
rect 4764 15829 4792 15832
rect 4831 15829 4832 15832
rect 4832 15829 4865 15832
rect 4904 15829 4934 15832
rect 4934 15829 4938 15832
rect 4977 15829 5002 15832
rect 5002 15829 5011 15832
rect 5050 15829 5070 15832
rect 5070 15829 5084 15832
rect 5123 15829 5138 15832
rect 5138 15829 5157 15832
rect 5196 15829 5206 15832
rect 5206 15829 5230 15832
rect 5269 15829 5274 15832
rect 5274 15829 5303 15832
rect 99 15777 102 15789
rect 102 15777 133 15789
rect 3882 15798 3916 15829
rect 3955 15798 3989 15829
rect 4028 15798 4062 15829
rect 4101 15798 4135 15829
rect 4174 15798 4208 15829
rect 4247 15798 4281 15829
rect 4320 15798 4354 15829
rect 4393 15798 4427 15829
rect 4466 15798 4500 15829
rect 4539 15798 4573 15829
rect 4612 15798 4646 15829
rect 4685 15798 4719 15829
rect 4758 15798 4792 15829
rect 4831 15798 4865 15829
rect 4904 15798 4938 15829
rect 4977 15798 5011 15829
rect 5050 15798 5084 15829
rect 5123 15798 5157 15829
rect 5196 15798 5230 15829
rect 5269 15798 5303 15829
rect 5342 15798 5376 15832
rect 5415 15829 5444 15832
rect 5444 15829 5449 15832
rect 5488 15829 5512 15832
rect 5512 15829 5522 15832
rect 5561 15829 5580 15832
rect 5580 15829 5595 15832
rect 5634 15829 5648 15832
rect 5648 15829 5668 15832
rect 5707 15829 5716 15832
rect 5716 15829 5741 15832
rect 5780 15829 5784 15832
rect 5784 15829 5814 15832
rect 5853 15829 5886 15832
rect 5886 15829 5887 15832
rect 5926 15829 5954 15832
rect 5954 15829 5960 15832
rect 5999 15829 6022 15832
rect 6022 15829 6033 15832
rect 6072 15829 6090 15832
rect 6090 15829 6106 15832
rect 6145 15829 6158 15832
rect 6158 15829 6179 15832
rect 6218 15829 6226 15832
rect 6226 15829 6252 15832
rect 6291 15829 6294 15832
rect 6294 15829 6325 15832
rect 6364 15829 6396 15832
rect 6396 15829 6398 15832
rect 6437 15829 6464 15832
rect 6464 15829 6471 15832
rect 6510 15829 6532 15832
rect 6532 15829 6544 15832
rect 6583 15829 6600 15832
rect 6600 15829 6617 15832
rect 6656 15829 6668 15832
rect 6668 15829 6690 15832
rect 6729 15829 6736 15832
rect 6736 15829 6763 15832
rect 6802 15829 6804 15832
rect 6804 15829 6836 15832
rect 6875 15829 6906 15832
rect 6906 15829 6909 15832
rect 6948 15829 6974 15832
rect 6974 15829 6982 15832
rect 7021 15829 7042 15832
rect 7042 15829 7055 15832
rect 7094 15829 7110 15832
rect 7110 15829 7128 15832
rect 7167 15829 7178 15832
rect 7178 15829 7201 15832
rect 7240 15829 7246 15832
rect 7246 15829 7274 15832
rect 7313 15829 7314 15832
rect 7314 15829 7347 15832
rect 7386 15829 7416 15832
rect 7416 15829 7420 15832
rect 7459 15829 7484 15832
rect 7484 15829 7493 15832
rect 7532 15829 7552 15832
rect 7552 15829 7566 15832
rect 7605 15829 7620 15832
rect 7620 15829 7639 15832
rect 7678 15829 7688 15832
rect 7688 15829 7712 15832
rect 7751 15829 7756 15832
rect 7756 15829 7785 15832
rect 7824 15829 7858 15832
rect 7897 15829 7926 15832
rect 7926 15829 7931 15832
rect 7970 15829 7994 15832
rect 7994 15829 8004 15832
rect 8043 15829 8062 15832
rect 8062 15829 8077 15832
rect 8116 15829 8130 15832
rect 8130 15829 8150 15832
rect 8189 15829 8198 15832
rect 8198 15829 8223 15832
rect 8262 15829 8266 15832
rect 8266 15829 8296 15832
rect 8335 15829 8368 15832
rect 8368 15829 8369 15832
rect 8408 15829 8436 15832
rect 8436 15829 8442 15832
rect 8481 15829 8504 15832
rect 8504 15829 8515 15832
rect 8554 15829 8572 15832
rect 8572 15829 8588 15832
rect 8627 15829 8640 15832
rect 8640 15829 8661 15832
rect 8699 15829 8708 15832
rect 8708 15829 8733 15832
rect 8771 15829 8776 15832
rect 8776 15829 8805 15832
rect 8843 15829 8844 15832
rect 8844 15829 8877 15832
rect 8915 15829 8946 15832
rect 8946 15829 8949 15832
rect 8987 15829 9014 15832
rect 9014 15829 9021 15832
rect 9059 15829 9082 15832
rect 9082 15829 9093 15832
rect 9131 15829 9150 15832
rect 9150 15829 9165 15832
rect 9203 15829 9218 15832
rect 9218 15829 9237 15832
rect 9275 15829 9286 15832
rect 9286 15829 9309 15832
rect 9347 15829 9354 15832
rect 9354 15829 9381 15832
rect 9419 15829 9422 15832
rect 9422 15829 9453 15832
rect 9491 15829 9524 15832
rect 9524 15829 9525 15832
rect 9563 15829 9592 15832
rect 9592 15829 9597 15832
rect 9635 15829 9660 15832
rect 9660 15829 9669 15832
rect 9707 15829 9728 15832
rect 9728 15829 9741 15832
rect 9779 15829 9796 15832
rect 9796 15829 9813 15832
rect 9851 15829 9864 15832
rect 9864 15829 9885 15832
rect 9923 15829 9932 15832
rect 9932 15829 9957 15832
rect 9995 15829 10000 15832
rect 10000 15829 10029 15832
rect 10067 15829 10068 15832
rect 10068 15829 10101 15832
rect 10139 15829 10170 15832
rect 10170 15829 10173 15832
rect 10211 15829 10238 15832
rect 10238 15829 10245 15832
rect 10283 15829 10306 15832
rect 10306 15829 10317 15832
rect 10355 15829 10374 15832
rect 10374 15829 10389 15832
rect 10427 15829 10442 15832
rect 10442 15829 10461 15832
rect 10499 15829 10510 15832
rect 10510 15829 10533 15832
rect 10571 15829 10578 15832
rect 10578 15829 10605 15832
rect 10643 15829 10646 15832
rect 10646 15829 10677 15832
rect 10715 15829 10748 15832
rect 10748 15829 10749 15832
rect 10787 15829 10816 15832
rect 10816 15829 10821 15832
rect 10859 15829 10884 15832
rect 10884 15829 10893 15832
rect 10931 15829 10952 15832
rect 10952 15829 10965 15832
rect 11003 15829 11020 15832
rect 11020 15829 11037 15832
rect 11075 15829 11088 15832
rect 11088 15829 11109 15832
rect 11147 15829 11156 15832
rect 11156 15829 11181 15832
rect 11219 15829 11224 15832
rect 11224 15829 11253 15832
rect 11291 15829 11292 15832
rect 11292 15829 11325 15832
rect 11363 15829 11394 15832
rect 11394 15829 11397 15832
rect 11435 15829 11462 15832
rect 11462 15829 11469 15832
rect 11507 15829 11530 15832
rect 11530 15829 11541 15832
rect 11579 15829 11598 15832
rect 11598 15829 11613 15832
rect 11651 15829 11666 15832
rect 11666 15829 11685 15832
rect 11723 15829 11734 15832
rect 11734 15829 11757 15832
rect 11795 15829 11802 15832
rect 11802 15829 11829 15832
rect 11867 15829 11870 15832
rect 11870 15829 11901 15832
rect 11939 15829 11972 15832
rect 11972 15829 11973 15832
rect 12011 15829 12040 15832
rect 12040 15829 12045 15832
rect 12083 15829 12108 15832
rect 12108 15829 12117 15832
rect 12155 15829 12176 15832
rect 12176 15829 12189 15832
rect 12227 15829 12244 15832
rect 12244 15829 12261 15832
rect 12299 15829 12312 15832
rect 12312 15829 12333 15832
rect 12371 15829 12380 15832
rect 12380 15829 12405 15832
rect 12443 15829 12448 15832
rect 12448 15829 12477 15832
rect 12515 15829 12516 15832
rect 12516 15829 12549 15832
rect 12587 15829 12618 15832
rect 12618 15829 12621 15832
rect 12659 15829 12686 15832
rect 12686 15829 12693 15832
rect 12731 15829 12754 15832
rect 12754 15829 12765 15832
rect 12803 15829 12822 15832
rect 12822 15829 12837 15832
rect 12875 15829 12890 15832
rect 12890 15829 12909 15832
rect 12947 15829 12958 15832
rect 12958 15829 12981 15832
rect 13019 15829 13026 15832
rect 13026 15829 13053 15832
rect 13091 15829 13094 15832
rect 13094 15829 13125 15832
rect 13163 15829 13196 15832
rect 13196 15829 13197 15832
rect 13235 15829 13264 15832
rect 13264 15829 13269 15832
rect 13307 15829 13332 15832
rect 13332 15829 13341 15832
rect 13379 15829 13400 15832
rect 13400 15829 13413 15832
rect 13451 15829 13468 15832
rect 13468 15829 13485 15832
rect 13523 15829 13536 15832
rect 13536 15829 13557 15832
rect 13595 15829 13604 15832
rect 13604 15829 13629 15832
rect 13667 15829 13672 15832
rect 13672 15829 13701 15832
rect 13739 15829 13740 15832
rect 13740 15829 13773 15832
rect 13811 15829 13842 15832
rect 13842 15829 13845 15832
rect 13883 15829 13910 15832
rect 13910 15829 13917 15832
rect 13955 15829 13978 15832
rect 13978 15829 13989 15832
rect 14027 15829 14046 15832
rect 14046 15829 14061 15832
rect 14099 15829 14114 15832
rect 14114 15829 14133 15832
rect 14171 15829 14182 15832
rect 14182 15829 14205 15832
rect 14243 15829 14250 15832
rect 14250 15829 14277 15832
rect 14315 15829 14318 15832
rect 14318 15829 14349 15832
rect 5415 15798 5449 15829
rect 5488 15798 5522 15829
rect 5561 15798 5595 15829
rect 5634 15798 5668 15829
rect 5707 15798 5741 15829
rect 5780 15798 5814 15829
rect 5853 15798 5887 15829
rect 5926 15798 5960 15829
rect 5999 15798 6033 15829
rect 6072 15798 6106 15829
rect 6145 15798 6179 15829
rect 6218 15798 6252 15829
rect 6291 15798 6325 15829
rect 6364 15798 6398 15829
rect 6437 15798 6471 15829
rect 6510 15798 6544 15829
rect 6583 15798 6617 15829
rect 6656 15798 6690 15829
rect 6729 15798 6763 15829
rect 6802 15798 6836 15829
rect 6875 15798 6909 15829
rect 6948 15798 6982 15829
rect 7021 15798 7055 15829
rect 7094 15798 7128 15829
rect 7167 15798 7201 15829
rect 7240 15798 7274 15829
rect 7313 15798 7347 15829
rect 7386 15798 7420 15829
rect 7459 15798 7493 15829
rect 7532 15798 7566 15829
rect 7605 15798 7639 15829
rect 7678 15798 7712 15829
rect 7751 15798 7785 15829
rect 7824 15798 7858 15829
rect 7897 15798 7931 15829
rect 7970 15798 8004 15829
rect 8043 15798 8077 15829
rect 8116 15798 8150 15829
rect 8189 15798 8223 15829
rect 8262 15798 8296 15829
rect 8335 15798 8369 15829
rect 8408 15798 8442 15829
rect 8481 15798 8515 15829
rect 8554 15798 8588 15829
rect 8627 15798 8661 15829
rect 8699 15798 8733 15829
rect 8771 15798 8805 15829
rect 8843 15798 8877 15829
rect 8915 15798 8949 15829
rect 8987 15798 9021 15829
rect 9059 15798 9093 15829
rect 9131 15798 9165 15829
rect 9203 15798 9237 15829
rect 9275 15798 9309 15829
rect 9347 15798 9381 15829
rect 9419 15798 9453 15829
rect 9491 15798 9525 15829
rect 9563 15798 9597 15829
rect 9635 15798 9669 15829
rect 9707 15798 9741 15829
rect 9779 15798 9813 15829
rect 9851 15798 9885 15829
rect 9923 15798 9957 15829
rect 9995 15798 10029 15829
rect 10067 15798 10101 15829
rect 10139 15798 10173 15829
rect 10211 15798 10245 15829
rect 10283 15798 10317 15829
rect 10355 15798 10389 15829
rect 10427 15798 10461 15829
rect 10499 15798 10533 15829
rect 10571 15798 10605 15829
rect 10643 15798 10677 15829
rect 10715 15798 10749 15829
rect 10787 15798 10821 15829
rect 10859 15798 10893 15829
rect 10931 15798 10965 15829
rect 11003 15798 11037 15829
rect 11075 15798 11109 15829
rect 11147 15798 11181 15829
rect 11219 15798 11253 15829
rect 11291 15798 11325 15829
rect 11363 15798 11397 15829
rect 11435 15798 11469 15829
rect 11507 15798 11541 15829
rect 11579 15798 11613 15829
rect 11651 15798 11685 15829
rect 11723 15798 11757 15829
rect 11795 15798 11829 15829
rect 11867 15798 11901 15829
rect 11939 15798 11973 15829
rect 12011 15798 12045 15829
rect 12083 15798 12117 15829
rect 12155 15798 12189 15829
rect 12227 15798 12261 15829
rect 12299 15798 12333 15829
rect 12371 15798 12405 15829
rect 12443 15798 12477 15829
rect 12515 15798 12549 15829
rect 12587 15798 12621 15829
rect 12659 15798 12693 15829
rect 12731 15798 12765 15829
rect 12803 15798 12837 15829
rect 12875 15798 12909 15829
rect 12947 15798 12981 15829
rect 13019 15798 13053 15829
rect 13091 15798 13125 15829
rect 13163 15798 13197 15829
rect 13235 15798 13269 15829
rect 13307 15798 13341 15829
rect 13379 15798 13413 15829
rect 13451 15798 13485 15829
rect 13523 15798 13557 15829
rect 13595 15798 13629 15829
rect 13667 15798 13701 15829
rect 13739 15798 13773 15829
rect 13811 15798 13845 15829
rect 13883 15798 13917 15829
rect 13955 15798 13989 15829
rect 14027 15798 14061 15829
rect 14099 15798 14133 15829
rect 14171 15798 14205 15829
rect 14243 15798 14277 15829
rect 14315 15798 14349 15829
rect 14387 15813 14421 15832
rect 14459 15813 14493 15832
rect 14531 15813 14565 15832
rect 14603 15813 14637 15832
rect 14675 15813 14709 15832
rect 14747 15813 14781 15832
rect 14819 15813 14853 15832
rect 14891 15813 14925 15832
rect 14387 15798 14420 15813
rect 14420 15798 14421 15813
rect 14459 15798 14492 15813
rect 14492 15798 14493 15813
rect 14531 15798 14564 15813
rect 14564 15798 14565 15813
rect 14603 15798 14636 15813
rect 14636 15798 14637 15813
rect 14675 15798 14708 15813
rect 14708 15798 14709 15813
rect 14747 15798 14780 15813
rect 14780 15798 14781 15813
rect 14819 15798 14852 15813
rect 14852 15798 14853 15813
rect 14891 15798 14924 15813
rect 14924 15798 14925 15813
rect 99 15755 133 15777
rect 99 15708 102 15717
rect 102 15708 133 15717
rect 171 15708 173 15717
rect 173 15708 205 15717
rect 3620 15723 3654 15737
rect 3692 15723 3726 15737
rect 3764 15723 3798 15737
rect 3836 15723 3870 15737
rect 3908 15723 3942 15737
rect 3980 15723 4014 15737
rect 4052 15723 4086 15737
rect 4124 15723 4158 15737
rect 4196 15723 4230 15737
rect 4268 15723 4302 15737
rect 4340 15723 4374 15737
rect 4412 15723 4446 15737
rect 4484 15723 4518 15737
rect 4557 15723 4591 15737
rect 4630 15723 4664 15737
rect 4703 15723 4737 15737
rect 4776 15723 4810 15737
rect 4849 15723 4883 15737
rect 4922 15723 4956 15737
rect 4995 15723 5029 15737
rect 5068 15723 5102 15737
rect 5141 15723 5175 15737
rect 5214 15723 5248 15737
rect 5287 15723 5321 15737
rect 5360 15723 5394 15737
rect 99 15683 133 15708
rect 171 15683 205 15708
rect 427 15689 444 15719
rect 444 15689 461 15719
rect 500 15689 513 15719
rect 513 15689 534 15719
rect 573 15689 582 15719
rect 582 15689 607 15719
rect 646 15689 651 15719
rect 651 15689 680 15719
rect 719 15689 720 15719
rect 720 15689 753 15719
rect 792 15689 823 15719
rect 823 15689 826 15719
rect 865 15689 892 15719
rect 892 15689 899 15719
rect 938 15689 961 15719
rect 961 15689 972 15719
rect 1011 15689 1030 15719
rect 1030 15689 1045 15719
rect 1084 15689 1099 15719
rect 1099 15689 1118 15719
rect 1157 15689 1168 15719
rect 1168 15689 1191 15719
rect 1230 15689 1237 15719
rect 1237 15689 1264 15719
rect 1303 15689 1306 15719
rect 1306 15689 1337 15719
rect 427 15685 461 15689
rect 500 15685 534 15689
rect 573 15685 607 15689
rect 646 15685 680 15689
rect 719 15685 753 15689
rect 792 15685 826 15689
rect 865 15685 899 15689
rect 938 15685 972 15689
rect 1011 15685 1045 15689
rect 1084 15685 1118 15689
rect 1157 15685 1191 15689
rect 1230 15685 1264 15689
rect 1303 15685 1337 15689
rect 1376 15685 1410 15719
rect 1449 15689 1479 15719
rect 1479 15689 1483 15719
rect 1521 15689 1548 15719
rect 1548 15689 1555 15719
rect 1593 15689 1617 15719
rect 1617 15689 1627 15719
rect 1665 15689 1686 15719
rect 1686 15689 1699 15719
rect 1737 15689 1755 15719
rect 1755 15689 1771 15719
rect 1809 15689 1824 15719
rect 1824 15689 1843 15719
rect 1881 15689 1893 15719
rect 1893 15689 1915 15719
rect 1953 15689 1962 15719
rect 1962 15689 1987 15719
rect 2025 15689 2031 15719
rect 2031 15689 2059 15719
rect 2097 15689 2100 15719
rect 2100 15689 2131 15719
rect 2169 15689 2203 15719
rect 2241 15689 2272 15719
rect 2272 15689 2275 15719
rect 2313 15689 2341 15719
rect 2341 15689 2347 15719
rect 2385 15689 2410 15719
rect 2410 15689 2419 15719
rect 2457 15689 2479 15719
rect 2479 15689 2491 15719
rect 2529 15689 2548 15719
rect 2548 15689 2563 15719
rect 2601 15689 2617 15719
rect 2617 15689 2635 15719
rect 2673 15689 2686 15719
rect 2686 15689 2707 15719
rect 2745 15689 2755 15719
rect 2755 15689 2779 15719
rect 2817 15689 2824 15719
rect 2824 15689 2851 15719
rect 2889 15689 2893 15719
rect 2893 15689 2923 15719
rect 2961 15689 2962 15719
rect 2962 15689 2995 15719
rect 3033 15689 3064 15719
rect 3064 15689 3067 15719
rect 3105 15689 3132 15719
rect 3132 15689 3139 15719
rect 3177 15689 3200 15719
rect 3200 15689 3211 15719
rect 3249 15689 3268 15719
rect 3268 15689 3283 15719
rect 3321 15689 3336 15719
rect 3336 15689 3355 15719
rect 3393 15689 3404 15719
rect 3404 15689 3427 15719
rect 3465 15689 3472 15719
rect 3472 15689 3499 15719
rect 3537 15689 3540 15719
rect 3540 15689 3571 15719
rect 3620 15703 3642 15723
rect 3642 15703 3654 15723
rect 3692 15703 3710 15723
rect 3710 15703 3726 15723
rect 3764 15703 3778 15723
rect 3778 15703 3798 15723
rect 3836 15703 3846 15723
rect 3846 15703 3870 15723
rect 3908 15703 3914 15723
rect 3914 15703 3942 15723
rect 3980 15703 3982 15723
rect 3982 15703 4014 15723
rect 4052 15703 4084 15723
rect 4084 15703 4086 15723
rect 4124 15703 4152 15723
rect 4152 15703 4158 15723
rect 4196 15703 4220 15723
rect 4220 15703 4230 15723
rect 4268 15703 4288 15723
rect 4288 15703 4302 15723
rect 4340 15703 4356 15723
rect 4356 15703 4374 15723
rect 4412 15703 4424 15723
rect 4424 15703 4446 15723
rect 4484 15703 4492 15723
rect 4492 15703 4518 15723
rect 4557 15703 4560 15723
rect 4560 15703 4591 15723
rect 4630 15703 4662 15723
rect 4662 15703 4664 15723
rect 4703 15703 4730 15723
rect 4730 15703 4737 15723
rect 4776 15703 4798 15723
rect 4798 15703 4810 15723
rect 4849 15703 4866 15723
rect 4866 15703 4883 15723
rect 4922 15703 4934 15723
rect 4934 15703 4956 15723
rect 4995 15703 5002 15723
rect 5002 15703 5029 15723
rect 5068 15703 5070 15723
rect 5070 15703 5102 15723
rect 5141 15703 5172 15723
rect 5172 15703 5175 15723
rect 5214 15703 5240 15723
rect 5240 15703 5248 15723
rect 5287 15703 5308 15723
rect 5308 15703 5321 15723
rect 5360 15703 5376 15723
rect 5376 15703 5394 15723
rect 1449 15685 1483 15689
rect 1521 15685 1555 15689
rect 1593 15685 1627 15689
rect 1665 15685 1699 15689
rect 1737 15685 1771 15689
rect 1809 15685 1843 15689
rect 1881 15685 1915 15689
rect 1953 15685 1987 15689
rect 2025 15685 2059 15689
rect 2097 15685 2131 15689
rect 2169 15685 2203 15689
rect 2241 15685 2275 15689
rect 2313 15685 2347 15689
rect 2385 15685 2419 15689
rect 2457 15685 2491 15689
rect 2529 15685 2563 15689
rect 2601 15685 2635 15689
rect 2673 15685 2707 15689
rect 2745 15685 2779 15689
rect 2817 15685 2851 15689
rect 2889 15685 2923 15689
rect 2961 15685 2995 15689
rect 3033 15685 3067 15689
rect 3105 15685 3139 15689
rect 3177 15685 3211 15689
rect 3249 15685 3283 15689
rect 3321 15685 3355 15689
rect 3393 15685 3427 15689
rect 3465 15685 3499 15689
rect 3537 15685 3571 15689
rect 69 15605 103 15639
rect 153 15605 187 15639
rect 237 15605 271 15639
rect 321 15605 355 15639
rect 405 15605 439 15639
rect 481 15583 515 15616
rect 5396 15613 5430 15647
rect 481 15582 488 15583
rect 488 15582 515 15583
rect 69 15535 103 15562
rect 153 15535 187 15562
rect 237 15535 271 15562
rect 321 15535 355 15562
rect 405 15549 420 15562
rect 420 15549 439 15562
rect 69 15528 102 15535
rect 102 15528 103 15535
rect 153 15528 173 15535
rect 173 15528 187 15535
rect 237 15528 244 15535
rect 244 15528 271 15535
rect 321 15528 352 15535
rect 352 15528 355 15535
rect 405 15528 439 15549
rect 481 15514 515 15541
rect 5396 15535 5430 15569
rect 481 15507 488 15514
rect 488 15507 515 15514
rect 69 15466 103 15485
rect 153 15466 187 15485
rect 237 15466 271 15485
rect 321 15466 355 15485
rect 405 15480 420 15485
rect 420 15480 439 15485
rect 69 15451 102 15466
rect 102 15451 103 15466
rect 153 15451 173 15466
rect 173 15451 187 15466
rect 237 15451 244 15466
rect 244 15451 271 15466
rect 321 15451 352 15466
rect 352 15451 355 15466
rect 405 15451 439 15480
rect 481 15445 515 15466
rect 481 15432 488 15445
rect 488 15432 515 15445
rect 69 15397 103 15408
rect 153 15397 187 15408
rect 237 15397 271 15408
rect 321 15397 355 15408
rect 69 15374 102 15397
rect 102 15374 103 15397
rect 153 15374 173 15397
rect 173 15374 187 15397
rect 237 15374 244 15397
rect 244 15374 271 15397
rect 321 15374 352 15397
rect 352 15374 355 15397
rect 405 15375 439 15408
rect 481 15375 515 15391
rect 405 15374 420 15375
rect 420 15374 439 15375
rect 481 15357 488 15375
rect 488 15357 515 15375
rect 69 15328 103 15331
rect 153 15328 187 15331
rect 237 15328 271 15331
rect 321 15328 355 15331
rect 69 15297 102 15328
rect 102 15297 103 15328
rect 153 15297 173 15328
rect 173 15297 187 15328
rect 237 15297 244 15328
rect 244 15297 271 15328
rect 321 15297 352 15328
rect 352 15297 355 15328
rect 405 15305 439 15331
rect 481 15305 515 15316
rect 405 15297 420 15305
rect 420 15297 439 15305
rect 481 15282 488 15305
rect 488 15282 515 15305
rect 69 15225 102 15254
rect 102 15225 103 15254
rect 153 15225 173 15254
rect 173 15225 187 15254
rect 237 15225 244 15254
rect 244 15225 271 15254
rect 321 15225 352 15254
rect 352 15225 355 15254
rect 405 15235 439 15254
rect 481 15235 515 15241
rect 69 15220 103 15225
rect 153 15220 187 15225
rect 237 15220 271 15225
rect 321 15220 355 15225
rect 405 15220 420 15235
rect 420 15220 439 15235
rect 481 15207 488 15235
rect 488 15207 515 15235
rect 69 15156 102 15177
rect 102 15156 103 15177
rect 153 15156 173 15177
rect 173 15156 187 15177
rect 237 15156 244 15177
rect 244 15156 271 15177
rect 321 15156 352 15177
rect 352 15156 355 15177
rect 405 15165 439 15177
rect 481 15165 515 15166
rect 69 15143 103 15156
rect 153 15143 187 15156
rect 237 15143 271 15156
rect 321 15143 355 15156
rect 405 15143 420 15165
rect 420 15143 439 15165
rect 481 15132 488 15165
rect 488 15132 515 15165
rect 69 15087 102 15100
rect 102 15087 103 15100
rect 153 15087 173 15100
rect 173 15087 187 15100
rect 237 15087 244 15100
rect 244 15087 271 15100
rect 321 15087 352 15100
rect 352 15087 355 15100
rect 405 15095 439 15100
rect 69 15066 103 15087
rect 153 15066 187 15087
rect 237 15066 271 15087
rect 321 15066 355 15087
rect 405 15066 420 15095
rect 420 15066 439 15095
rect 481 15061 488 15091
rect 488 15061 515 15091
rect 481 15057 515 15061
rect 69 15018 102 15022
rect 102 15018 103 15022
rect 153 15018 173 15022
rect 173 15018 187 15022
rect 237 15018 244 15022
rect 244 15018 271 15022
rect 321 15018 352 15022
rect 352 15018 355 15022
rect 69 14988 103 15018
rect 153 14988 187 15018
rect 237 14988 271 15018
rect 321 14988 355 15018
rect 405 14991 420 15022
rect 420 14991 439 15022
rect 481 14991 488 15016
rect 488 14991 515 15016
rect 405 14988 439 14991
rect 481 14982 515 14991
rect 69 14914 103 14944
rect 153 14914 187 14944
rect 237 14914 271 14944
rect 321 14914 355 14944
rect 405 14921 420 14944
rect 420 14921 439 14944
rect 481 14921 488 14941
rect 488 14921 515 14941
rect 69 14910 102 14914
rect 102 14910 103 14914
rect 153 14910 173 14914
rect 173 14910 187 14914
rect 237 14910 244 14914
rect 244 14910 271 14914
rect 321 14910 352 14914
rect 352 14910 355 14914
rect 405 14910 439 14921
rect 481 14907 515 14921
rect 694 15474 728 15508
rect 766 15474 800 15508
rect 838 15474 872 15508
rect 910 15474 944 15508
rect 982 15474 1016 15508
rect 1054 15474 1088 15508
rect 1126 15474 1160 15508
rect 1198 15474 1232 15508
rect 1270 15474 1304 15508
rect 1342 15474 1376 15508
rect 1414 15474 1448 15508
rect 1486 15474 1520 15508
rect 1558 15474 1592 15508
rect 1630 15474 1664 15508
rect 1702 15474 1736 15508
rect 1774 15474 1808 15508
rect 1846 15474 1880 15508
rect 1918 15474 1952 15508
rect 1990 15474 2024 15508
rect 2062 15474 2096 15508
rect 2134 15474 2168 15508
rect 2206 15474 2240 15508
rect 2278 15474 2312 15508
rect 2350 15474 2384 15508
rect 2422 15474 2456 15508
rect 2494 15474 2528 15508
rect 2566 15474 2600 15508
rect 2638 15474 2672 15508
rect 2710 15474 2744 15508
rect 2782 15474 2816 15508
rect 2854 15474 2888 15508
rect 2926 15474 2960 15508
rect 2998 15474 3032 15508
rect 3070 15474 3104 15508
rect 3142 15474 3176 15508
rect 3214 15474 3248 15508
rect 3286 15474 3320 15508
rect 3358 15474 3392 15508
rect 3430 15474 3464 15508
rect 3502 15474 3536 15508
rect 3574 15474 3608 15508
rect 3646 15474 3680 15508
rect 3718 15474 3752 15508
rect 3790 15474 3824 15508
rect 3862 15474 3896 15508
rect 3935 15474 3969 15508
rect 4017 15470 4051 15504
rect 4094 15470 4128 15504
rect 4171 15470 4205 15504
rect 4248 15470 4282 15504
rect 4325 15470 4359 15504
rect 4402 15470 4436 15504
rect 4479 15470 4513 15504
rect 4556 15470 4590 15504
rect 4632 15470 4666 15504
rect 4708 15470 4742 15504
rect 4784 15470 4818 15504
rect 4860 15470 4894 15504
rect 4936 15470 4970 15504
rect 5012 15470 5046 15504
rect 5088 15470 5122 15504
rect 5164 15470 5198 15504
rect 622 15402 656 15436
rect 710 15387 732 15420
rect 732 15387 744 15420
rect 783 15387 801 15420
rect 801 15387 817 15420
rect 856 15387 870 15420
rect 870 15387 890 15420
rect 929 15387 939 15420
rect 939 15387 963 15420
rect 1002 15387 1008 15420
rect 1008 15387 1036 15420
rect 1075 15387 1077 15420
rect 1077 15387 1109 15420
rect 1148 15387 1181 15420
rect 1181 15387 1182 15420
rect 1221 15387 1250 15420
rect 1250 15387 1255 15420
rect 1294 15387 1319 15420
rect 1319 15387 1328 15420
rect 1367 15387 1388 15420
rect 1388 15387 1401 15420
rect 1440 15387 1457 15420
rect 1457 15387 1474 15420
rect 1513 15387 1526 15420
rect 1526 15387 1547 15420
rect 1586 15387 1595 15420
rect 1595 15387 1620 15420
rect 1659 15387 1664 15420
rect 1664 15387 1693 15420
rect 1732 15387 1733 15420
rect 1733 15387 1766 15420
rect 1805 15387 1836 15420
rect 1836 15387 1839 15420
rect 1878 15387 1905 15420
rect 1905 15387 1912 15420
rect 1951 15387 1974 15420
rect 1974 15387 1985 15420
rect 2024 15387 2043 15420
rect 2043 15387 2058 15420
rect 2097 15387 2112 15420
rect 2112 15387 2131 15420
rect 2170 15387 2181 15420
rect 2181 15387 2204 15420
rect 2243 15387 2250 15420
rect 2250 15387 2277 15420
rect 2316 15387 2319 15420
rect 2319 15387 2350 15420
rect 710 15386 744 15387
rect 783 15386 817 15387
rect 856 15386 890 15387
rect 929 15386 963 15387
rect 1002 15386 1036 15387
rect 1075 15386 1109 15387
rect 1148 15386 1182 15387
rect 1221 15386 1255 15387
rect 1294 15386 1328 15387
rect 1367 15386 1401 15387
rect 1440 15386 1474 15387
rect 1513 15386 1547 15387
rect 1586 15386 1620 15387
rect 1659 15386 1693 15387
rect 1732 15386 1766 15387
rect 1805 15386 1839 15387
rect 1878 15386 1912 15387
rect 1951 15386 1985 15387
rect 2024 15386 2058 15387
rect 2097 15386 2131 15387
rect 2170 15386 2204 15387
rect 2243 15386 2277 15387
rect 2316 15386 2350 15387
rect 2389 15386 2423 15420
rect 2462 15387 2492 15420
rect 2492 15387 2496 15420
rect 2535 15387 2561 15420
rect 2561 15387 2569 15420
rect 2608 15387 2630 15420
rect 2630 15387 2642 15420
rect 2681 15387 2699 15420
rect 2699 15387 2715 15420
rect 2754 15387 2768 15420
rect 2768 15387 2788 15420
rect 2827 15387 2837 15420
rect 2837 15387 2861 15420
rect 2900 15387 2906 15420
rect 2906 15387 2934 15420
rect 2973 15387 2975 15420
rect 2975 15387 3007 15420
rect 3047 15387 3078 15420
rect 3078 15387 3081 15420
rect 3121 15387 3147 15420
rect 3147 15387 3155 15420
rect 3195 15387 3216 15420
rect 3216 15387 3229 15420
rect 3269 15387 3285 15420
rect 3285 15387 3303 15420
rect 3343 15387 3354 15420
rect 3354 15387 3377 15420
rect 3417 15387 3423 15420
rect 3423 15387 3451 15420
rect 3491 15387 3492 15420
rect 3492 15387 3525 15420
rect 3565 15387 3596 15420
rect 3596 15387 3599 15420
rect 3639 15387 3665 15420
rect 3665 15387 3673 15420
rect 3713 15387 3734 15420
rect 3734 15387 3747 15420
rect 3787 15387 3803 15420
rect 3803 15387 3821 15420
rect 3861 15387 3872 15420
rect 3872 15387 3895 15420
rect 3935 15387 3941 15420
rect 3941 15387 3969 15420
rect 4211 15387 4217 15391
rect 4217 15387 4245 15391
rect 4287 15387 4320 15391
rect 4320 15387 4321 15391
rect 4363 15387 4389 15391
rect 4389 15387 4397 15391
rect 4439 15387 4458 15391
rect 4458 15387 4473 15391
rect 4515 15387 4527 15391
rect 4527 15387 4549 15391
rect 4591 15387 4596 15391
rect 4596 15387 4625 15391
rect 4667 15387 4700 15391
rect 4700 15387 4701 15391
rect 4743 15387 4769 15391
rect 4769 15387 4777 15391
rect 4819 15387 4838 15391
rect 4838 15387 4853 15391
rect 4894 15387 4907 15391
rect 4907 15387 4928 15391
rect 4969 15387 4976 15391
rect 4976 15387 5003 15391
rect 5044 15387 5045 15391
rect 5045 15387 5078 15391
rect 5228 15410 5262 15444
rect 2462 15386 2496 15387
rect 2535 15386 2569 15387
rect 2608 15386 2642 15387
rect 2681 15386 2715 15387
rect 2754 15386 2788 15387
rect 2827 15386 2861 15387
rect 2900 15386 2934 15387
rect 2973 15386 3007 15387
rect 3047 15386 3081 15387
rect 3121 15386 3155 15387
rect 3195 15386 3229 15387
rect 3269 15386 3303 15387
rect 3343 15386 3377 15387
rect 3417 15386 3451 15387
rect 3491 15386 3525 15387
rect 3565 15386 3599 15387
rect 3639 15386 3673 15387
rect 3713 15386 3747 15387
rect 3787 15386 3821 15387
rect 3861 15386 3895 15387
rect 3935 15386 3969 15387
rect 622 15328 656 15362
rect 4211 15357 4245 15387
rect 4287 15357 4321 15387
rect 4363 15357 4397 15387
rect 4439 15357 4473 15387
rect 4515 15357 4549 15387
rect 4591 15357 4625 15387
rect 4667 15357 4701 15387
rect 4743 15357 4777 15387
rect 4819 15357 4853 15387
rect 4894 15357 4928 15387
rect 4969 15357 5003 15387
rect 5044 15357 5078 15387
rect 5228 15363 5242 15372
rect 5242 15363 5262 15372
rect 710 15303 744 15337
rect 5228 15338 5262 15363
rect 622 15254 656 15288
rect 710 15220 744 15254
rect 622 15180 656 15214
rect 887 15271 896 15305
rect 896 15271 921 15305
rect 959 15271 964 15305
rect 964 15271 993 15305
rect 1031 15271 1032 15305
rect 1032 15271 1065 15305
rect 1103 15271 1134 15305
rect 1134 15271 1137 15305
rect 1175 15271 1202 15305
rect 1202 15271 1209 15305
rect 1247 15271 1270 15305
rect 1270 15271 1281 15305
rect 1319 15271 1338 15305
rect 1338 15271 1353 15305
rect 1391 15271 1406 15305
rect 1406 15271 1425 15305
rect 1463 15271 1474 15305
rect 1474 15271 1497 15305
rect 1535 15271 1542 15305
rect 1542 15271 1569 15305
rect 1607 15271 1610 15305
rect 1610 15271 1641 15305
rect 1679 15271 1712 15305
rect 1712 15271 1713 15305
rect 1751 15271 1785 15305
rect 1823 15271 1857 15305
rect 1895 15271 1929 15305
rect 1967 15271 1996 15305
rect 1996 15271 2001 15305
rect 2039 15271 2064 15305
rect 2064 15271 2073 15305
rect 2111 15271 2132 15305
rect 2132 15271 2145 15305
rect 2183 15271 2200 15305
rect 2200 15271 2217 15305
rect 2256 15271 2268 15305
rect 2268 15271 2290 15305
rect 2329 15271 2336 15305
rect 2336 15271 2363 15305
rect 2402 15271 2404 15305
rect 2404 15271 2436 15305
rect 2483 15271 2506 15305
rect 2506 15271 2517 15305
rect 2555 15271 2574 15305
rect 2574 15271 2589 15305
rect 2627 15271 2642 15305
rect 2642 15271 2661 15305
rect 2699 15271 2710 15305
rect 2710 15271 2733 15305
rect 2771 15271 2778 15305
rect 2778 15271 2805 15305
rect 2843 15271 2846 15305
rect 2846 15271 2877 15305
rect 2915 15271 2949 15305
rect 2987 15271 3021 15305
rect 3059 15271 3083 15305
rect 3083 15271 3093 15305
rect 3131 15271 3151 15305
rect 3151 15271 3165 15305
rect 3204 15271 3219 15305
rect 3219 15271 3238 15305
rect 3277 15271 3287 15305
rect 3287 15271 3311 15305
rect 3350 15271 3355 15305
rect 3355 15271 3384 15305
rect 3423 15271 3457 15305
rect 3496 15271 3525 15305
rect 3525 15271 3530 15305
rect 3569 15271 3593 15305
rect 3593 15271 3603 15305
rect 3642 15271 3661 15305
rect 3661 15271 3676 15305
rect 3715 15271 3729 15305
rect 3729 15271 3749 15305
rect 3788 15271 3797 15305
rect 3797 15271 3822 15305
rect 3861 15271 3865 15305
rect 3865 15271 3895 15305
rect 3934 15271 3967 15305
rect 3967 15271 3968 15305
rect 4007 15271 4041 15305
rect 4080 15271 4114 15305
rect 5228 15284 5262 15300
rect 5228 15266 5242 15284
rect 5242 15266 5262 15284
rect 622 15106 656 15140
rect 710 15137 744 15171
rect 1832 15169 1854 15203
rect 1854 15169 1866 15203
rect 1906 15169 1940 15203
rect 1980 15169 2014 15203
rect 2054 15169 2088 15203
rect 2128 15169 2162 15203
rect 2202 15169 2236 15203
rect 2276 15169 2310 15203
rect 2350 15169 2384 15203
rect 2424 15169 2458 15203
rect 2498 15169 2532 15203
rect 2572 15169 2606 15203
rect 2646 15169 2680 15203
rect 2720 15169 2754 15203
rect 2794 15169 2828 15203
rect 2868 15169 2902 15203
rect 2942 15169 2973 15203
rect 2973 15169 2976 15203
rect 3016 15169 3050 15203
rect 3090 15169 3124 15203
rect 3164 15169 3198 15203
rect 3238 15169 3272 15203
rect 3312 15169 3346 15203
rect 3386 15169 3420 15203
rect 3460 15169 3494 15203
rect 3534 15169 3568 15203
rect 3607 15169 3641 15203
rect 3680 15169 3714 15203
rect 3753 15169 3787 15203
rect 3826 15169 3860 15203
rect 3899 15169 3933 15203
rect 3972 15169 4006 15203
rect 4045 15169 4060 15203
rect 4060 15169 4079 15203
rect 5228 15194 5262 15228
rect 5228 15150 5262 15156
rect 4211 15129 4245 15136
rect 4287 15129 4321 15136
rect 4363 15129 4397 15136
rect 4439 15129 4473 15136
rect 4515 15129 4549 15136
rect 4591 15129 4625 15136
rect 4667 15129 4701 15136
rect 4743 15129 4777 15136
rect 4819 15129 4853 15136
rect 4894 15129 4928 15136
rect 4969 15129 5003 15136
rect 5044 15129 5078 15136
rect 4211 15102 4238 15129
rect 4238 15102 4245 15129
rect 4287 15102 4306 15129
rect 4306 15102 4321 15129
rect 4363 15102 4374 15129
rect 4374 15102 4397 15129
rect 4439 15102 4442 15129
rect 4442 15102 4473 15129
rect 4515 15102 4544 15129
rect 4544 15102 4549 15129
rect 4591 15102 4612 15129
rect 4612 15102 4625 15129
rect 4667 15102 4680 15129
rect 4680 15102 4701 15129
rect 4743 15102 4748 15129
rect 4748 15102 4777 15129
rect 4819 15102 4850 15129
rect 4850 15102 4853 15129
rect 4894 15102 4918 15129
rect 4918 15102 4928 15129
rect 4969 15102 4986 15129
rect 4986 15102 5003 15129
rect 5044 15102 5054 15129
rect 5054 15102 5078 15129
rect 5228 15122 5242 15150
rect 5242 15122 5262 15150
rect 622 15032 656 15066
rect 710 15055 744 15089
rect 2465 15013 2499 15024
rect 2538 15013 2572 15024
rect 2611 15013 2645 15024
rect 2684 15013 2718 15024
rect 2757 15013 2791 15024
rect 2830 15013 2864 15024
rect 2903 15013 2937 15024
rect 2976 15013 3010 15024
rect 3049 15013 3083 15024
rect 3122 15013 3156 15024
rect 3195 15013 3229 15024
rect 3268 15013 3302 15024
rect 3341 15013 3375 15024
rect 3414 15013 3448 15024
rect 3487 15013 3521 15024
rect 3560 15013 3594 15024
rect 3633 15013 3667 15024
rect 3706 15013 3740 15024
rect 3779 15013 3813 15024
rect 3852 15013 3886 15024
rect 3925 15013 3959 15024
rect 3998 15013 4032 15024
rect 4071 15013 4105 15024
rect 4144 15013 4178 15024
rect 4217 15013 4251 15024
rect 4290 15013 4324 15024
rect 4363 15013 4397 15024
rect 4436 15013 4470 15024
rect 4509 15013 4543 15024
rect 4582 15013 4616 15024
rect 4655 15013 4689 15024
rect 4728 15013 4762 15024
rect 4801 15013 4835 15024
rect 622 14958 656 14992
rect 710 14973 744 15007
rect 783 14979 802 15007
rect 802 14979 817 15007
rect 856 14979 871 15007
rect 871 14979 890 15007
rect 929 14979 940 15007
rect 940 14979 963 15007
rect 1002 14979 1009 15007
rect 1009 14979 1036 15007
rect 1075 14979 1078 15007
rect 1078 14979 1109 15007
rect 783 14973 817 14979
rect 856 14973 890 14979
rect 929 14973 963 14979
rect 1002 14973 1036 14979
rect 1075 14973 1109 14979
rect 1148 14973 1182 15007
rect 1221 14979 1251 15007
rect 1251 14979 1255 15007
rect 1294 14979 1320 15007
rect 1320 14979 1328 15007
rect 1367 14979 1389 15007
rect 1389 14979 1401 15007
rect 1440 14979 1458 15007
rect 1458 14979 1474 15007
rect 1513 14979 1527 15007
rect 1527 14979 1547 15007
rect 1586 14979 1596 15007
rect 1596 14979 1620 15007
rect 1659 14979 1665 15007
rect 1665 14979 1693 15007
rect 1732 14979 1734 15007
rect 1734 14979 1766 15007
rect 1805 14979 1837 15007
rect 1837 14979 1839 15007
rect 1878 14979 1906 15007
rect 1906 14979 1912 15007
rect 1950 14979 1975 15007
rect 1975 14979 1984 15007
rect 2022 14979 2044 15007
rect 2044 14979 2056 15007
rect 2094 14979 2113 15007
rect 2113 14979 2128 15007
rect 2166 14979 2182 15007
rect 2182 14979 2200 15007
rect 2238 14979 2251 15007
rect 2251 14979 2272 15007
rect 2310 14979 2320 15007
rect 2320 14979 2344 15007
rect 2465 14990 2493 15013
rect 2493 14990 2499 15013
rect 2538 14990 2562 15013
rect 2562 14990 2572 15013
rect 2611 14990 2631 15013
rect 2631 14990 2645 15013
rect 2684 14990 2700 15013
rect 2700 14990 2718 15013
rect 2757 14990 2769 15013
rect 2769 14990 2791 15013
rect 2830 14990 2838 15013
rect 2838 14990 2864 15013
rect 2903 14990 2907 15013
rect 2907 14990 2937 15013
rect 2976 14990 3010 15013
rect 3049 14990 3079 15013
rect 3079 14990 3083 15013
rect 3122 14990 3148 15013
rect 3148 14990 3156 15013
rect 3195 14990 3217 15013
rect 3217 14990 3229 15013
rect 3268 14990 3286 15013
rect 3286 14990 3302 15013
rect 3341 14990 3355 15013
rect 3355 14990 3375 15013
rect 3414 14990 3424 15013
rect 3424 14990 3448 15013
rect 3487 14990 3493 15013
rect 3493 14990 3521 15013
rect 3560 14990 3562 15013
rect 3562 14990 3594 15013
rect 3633 14990 3666 15013
rect 3666 14990 3667 15013
rect 3706 14990 3735 15013
rect 3735 14990 3740 15013
rect 3779 14990 3804 15013
rect 3804 14990 3813 15013
rect 3852 14990 3873 15013
rect 3873 14990 3886 15013
rect 3925 14990 3942 15013
rect 3942 14990 3959 15013
rect 3998 14990 4011 15013
rect 4011 14990 4032 15013
rect 4071 14990 4080 15013
rect 4080 14990 4105 15013
rect 4144 14990 4149 15013
rect 4149 14990 4178 15013
rect 4217 14990 4218 15013
rect 4218 14990 4251 15013
rect 4290 14990 4321 15013
rect 4321 14990 4324 15013
rect 4363 14990 4390 15013
rect 4390 14990 4397 15013
rect 4436 14990 4459 15013
rect 4459 14990 4470 15013
rect 4509 14990 4528 15013
rect 4528 14990 4543 15013
rect 4582 14990 4597 15013
rect 4597 14990 4616 15013
rect 4655 14990 4666 15013
rect 4666 14990 4689 15013
rect 4728 14990 4735 15013
rect 4735 14990 4762 15013
rect 4801 14990 4804 15013
rect 4804 14990 4835 15013
rect 4874 14990 4908 15024
rect 4947 15013 4981 15024
rect 5020 15013 5054 15024
rect 5094 15013 5128 15024
rect 5168 15013 5202 15024
rect 4947 14990 4977 15013
rect 4977 14990 4981 15013
rect 5020 14990 5046 15013
rect 5046 14990 5054 15013
rect 5094 14990 5115 15013
rect 5115 14990 5128 15013
rect 5168 14990 5184 15013
rect 5184 14990 5202 15013
rect 1221 14973 1255 14979
rect 1294 14973 1328 14979
rect 1367 14973 1401 14979
rect 1440 14973 1474 14979
rect 1513 14973 1547 14979
rect 1586 14973 1620 14979
rect 1659 14973 1693 14979
rect 1732 14973 1766 14979
rect 1805 14973 1839 14979
rect 1878 14973 1912 14979
rect 1950 14973 1984 14979
rect 2022 14973 2056 14979
rect 2094 14973 2128 14979
rect 2166 14973 2200 14979
rect 2238 14973 2272 14979
rect 2310 14973 2344 14979
rect 694 14885 728 14919
rect 768 14885 802 14919
rect 842 14885 876 14919
rect 916 14885 950 14919
rect 990 14885 1024 14919
rect 1064 14885 1098 14919
rect 1138 14885 1172 14919
rect 1212 14885 1246 14919
rect 1286 14885 1320 14919
rect 1360 14885 1394 14919
rect 1434 14885 1468 14919
rect 1507 14885 1541 14919
rect 1580 14885 1614 14919
rect 1653 14885 1687 14919
rect 1726 14885 1760 14919
rect 1799 14885 1833 14919
rect 1872 14885 1906 14919
rect 1945 14885 1979 14919
rect 2018 14885 2052 14919
rect 2091 14885 2125 14919
rect 2164 14885 2198 14919
rect 2237 14885 2271 14919
rect 2310 14885 2344 14919
rect 5396 15457 5430 15491
rect 5396 15379 5430 15413
rect 5396 15301 5430 15335
rect 5396 15223 5430 15257
rect 5396 15145 5430 15179
rect 5396 15067 5430 15101
rect 5396 14989 5430 15023
rect 5396 14911 5430 14945
rect 69 14845 103 14866
rect 153 14845 187 14866
rect 237 14845 271 14866
rect 321 14845 355 14866
rect 405 14851 420 14866
rect 420 14851 439 14866
rect 481 14851 488 14867
rect 488 14851 515 14867
rect 69 14832 102 14845
rect 102 14832 103 14845
rect 153 14832 173 14845
rect 173 14832 187 14845
rect 237 14832 244 14845
rect 244 14832 271 14845
rect 321 14832 352 14845
rect 352 14832 355 14845
rect 405 14832 439 14851
rect 481 14833 515 14851
rect 5396 14833 5430 14867
rect 12860 15441 12894 15464
rect 12934 15441 12968 15464
rect 13008 15441 13042 15464
rect 13082 15441 13116 15464
rect 13156 15441 13190 15464
rect 13230 15441 13264 15464
rect 13304 15441 13338 15464
rect 13378 15441 13412 15464
rect 13452 15441 13486 15464
rect 13526 15441 13560 15464
rect 13600 15441 13634 15464
rect 13674 15441 13708 15464
rect 13748 15441 13782 15464
rect 13822 15441 13856 15464
rect 13896 15441 13930 15464
rect 13970 15441 14004 15464
rect 14044 15441 14078 15464
rect 14118 15441 14152 15464
rect 14191 15441 14225 15464
rect 14264 15441 14298 15464
rect 14337 15441 14371 15464
rect 12860 15430 12869 15441
rect 12869 15430 12894 15441
rect 12934 15430 12938 15441
rect 12938 15430 12968 15441
rect 13008 15430 13041 15441
rect 13041 15430 13042 15441
rect 13082 15430 13110 15441
rect 13110 15430 13116 15441
rect 13156 15430 13179 15441
rect 13179 15430 13190 15441
rect 13230 15430 13248 15441
rect 13248 15430 13264 15441
rect 13304 15430 13317 15441
rect 13317 15430 13338 15441
rect 13378 15430 13386 15441
rect 13386 15430 13412 15441
rect 13452 15430 13455 15441
rect 13455 15430 13486 15441
rect 13526 15430 13559 15441
rect 13559 15430 13560 15441
rect 13600 15430 13628 15441
rect 13628 15430 13634 15441
rect 13674 15430 13697 15441
rect 13697 15430 13708 15441
rect 13748 15430 13766 15441
rect 13766 15430 13782 15441
rect 13822 15430 13835 15441
rect 13835 15430 13856 15441
rect 13896 15430 13904 15441
rect 13904 15430 13930 15441
rect 13970 15430 13973 15441
rect 13973 15430 14004 15441
rect 14044 15430 14076 15441
rect 14076 15430 14078 15441
rect 14118 15430 14145 15441
rect 14145 15430 14152 15441
rect 14191 15430 14214 15441
rect 14214 15430 14225 15441
rect 14264 15430 14283 15441
rect 14283 15430 14298 15441
rect 14337 15430 14352 15441
rect 14352 15430 14371 15441
rect 14410 15434 14420 15464
rect 14420 15434 14444 15464
rect 14483 15434 14492 15464
rect 14492 15434 14517 15464
rect 14556 15434 14564 15464
rect 14564 15434 14590 15464
rect 14629 15434 14636 15464
rect 14636 15434 14663 15464
rect 14702 15434 14708 15464
rect 14708 15434 14736 15464
rect 14775 15434 14780 15464
rect 14780 15434 14809 15464
rect 14848 15434 14852 15464
rect 14852 15434 14882 15464
rect 14410 15430 14444 15434
rect 14483 15430 14517 15434
rect 14556 15430 14590 15434
rect 14629 15430 14663 15434
rect 14702 15430 14736 15434
rect 14775 15430 14809 15434
rect 14848 15430 14882 15434
rect 12860 15371 12894 15382
rect 12934 15371 12968 15382
rect 13008 15371 13042 15382
rect 13082 15371 13116 15382
rect 13156 15371 13190 15382
rect 13230 15371 13264 15382
rect 13304 15371 13338 15382
rect 13378 15371 13412 15382
rect 13452 15371 13486 15382
rect 13526 15371 13560 15382
rect 13600 15371 13634 15382
rect 13674 15371 13708 15382
rect 13748 15371 13782 15382
rect 13822 15371 13856 15382
rect 13896 15371 13930 15382
rect 13970 15371 14004 15382
rect 14044 15371 14078 15382
rect 14118 15371 14152 15382
rect 14191 15371 14225 15382
rect 14264 15371 14298 15382
rect 14337 15371 14371 15382
rect 12860 15348 12869 15371
rect 12869 15348 12894 15371
rect 12934 15348 12938 15371
rect 12938 15348 12968 15371
rect 13008 15348 13041 15371
rect 13041 15348 13042 15371
rect 13082 15348 13110 15371
rect 13110 15348 13116 15371
rect 13156 15348 13179 15371
rect 13179 15348 13190 15371
rect 13230 15348 13248 15371
rect 13248 15348 13264 15371
rect 13304 15348 13317 15371
rect 13317 15348 13338 15371
rect 13378 15348 13386 15371
rect 13386 15348 13412 15371
rect 13452 15348 13455 15371
rect 13455 15348 13486 15371
rect 13526 15348 13559 15371
rect 13559 15348 13560 15371
rect 13600 15348 13628 15371
rect 13628 15348 13634 15371
rect 13674 15348 13697 15371
rect 13697 15348 13708 15371
rect 13748 15348 13766 15371
rect 13766 15348 13782 15371
rect 13822 15348 13835 15371
rect 13835 15348 13856 15371
rect 13896 15348 13904 15371
rect 13904 15348 13930 15371
rect 13970 15348 13973 15371
rect 13973 15348 14004 15371
rect 14044 15348 14076 15371
rect 14076 15348 14078 15371
rect 14118 15348 14145 15371
rect 14145 15348 14152 15371
rect 14191 15348 14214 15371
rect 14214 15348 14225 15371
rect 14264 15348 14283 15371
rect 14283 15348 14298 15371
rect 14337 15348 14352 15371
rect 14352 15348 14371 15371
rect 14410 15365 14420 15382
rect 14420 15365 14444 15382
rect 14483 15365 14492 15382
rect 14492 15365 14517 15382
rect 14556 15365 14564 15382
rect 14564 15365 14590 15382
rect 14629 15365 14636 15382
rect 14636 15365 14663 15382
rect 14702 15365 14708 15382
rect 14708 15365 14736 15382
rect 14775 15365 14780 15382
rect 14780 15365 14809 15382
rect 14848 15365 14852 15382
rect 14852 15365 14882 15382
rect 14410 15348 14444 15365
rect 14483 15348 14517 15365
rect 14556 15348 14590 15365
rect 14629 15348 14663 15365
rect 14702 15348 14736 15365
rect 14775 15348 14809 15365
rect 14848 15348 14882 15365
rect 12860 15267 12869 15300
rect 12869 15267 12894 15300
rect 12934 15267 12938 15300
rect 12938 15267 12968 15300
rect 13008 15267 13041 15300
rect 13041 15267 13042 15300
rect 13082 15267 13110 15300
rect 13110 15267 13116 15300
rect 13156 15267 13179 15300
rect 13179 15267 13190 15300
rect 13230 15267 13248 15300
rect 13248 15267 13264 15300
rect 13304 15267 13317 15300
rect 13317 15267 13338 15300
rect 13378 15267 13386 15300
rect 13386 15267 13412 15300
rect 13452 15267 13455 15300
rect 13455 15267 13486 15300
rect 13526 15267 13559 15300
rect 13559 15267 13560 15300
rect 13600 15267 13628 15300
rect 13628 15267 13634 15300
rect 13674 15267 13697 15300
rect 13697 15267 13708 15300
rect 13748 15267 13766 15300
rect 13766 15267 13782 15300
rect 13822 15267 13835 15300
rect 13835 15267 13856 15300
rect 13896 15267 13904 15300
rect 13904 15267 13930 15300
rect 13970 15267 13973 15300
rect 13973 15267 14004 15300
rect 14044 15267 14076 15300
rect 14076 15267 14078 15300
rect 14118 15267 14145 15300
rect 14145 15267 14152 15300
rect 14191 15267 14214 15300
rect 14214 15267 14225 15300
rect 14264 15267 14283 15300
rect 14283 15267 14298 15300
rect 14337 15267 14352 15300
rect 14352 15267 14371 15300
rect 12860 15266 12894 15267
rect 12934 15266 12968 15267
rect 13008 15266 13042 15267
rect 13082 15266 13116 15267
rect 13156 15266 13190 15267
rect 13230 15266 13264 15267
rect 13304 15266 13338 15267
rect 13378 15266 13412 15267
rect 13452 15266 13486 15267
rect 13526 15266 13560 15267
rect 13600 15266 13634 15267
rect 13674 15266 13708 15267
rect 13748 15266 13782 15267
rect 13822 15266 13856 15267
rect 13896 15266 13930 15267
rect 13970 15266 14004 15267
rect 14044 15266 14078 15267
rect 14118 15266 14152 15267
rect 14191 15266 14225 15267
rect 14264 15266 14298 15267
rect 14337 15266 14371 15267
rect 14410 15296 14420 15300
rect 14420 15296 14444 15300
rect 14483 15296 14492 15300
rect 14492 15296 14517 15300
rect 14556 15296 14564 15300
rect 14564 15296 14590 15300
rect 14629 15296 14636 15300
rect 14636 15296 14663 15300
rect 14702 15296 14708 15300
rect 14708 15296 14736 15300
rect 14775 15296 14780 15300
rect 14780 15296 14809 15300
rect 14848 15296 14852 15300
rect 14852 15296 14882 15300
rect 14410 15266 14444 15296
rect 14483 15266 14517 15296
rect 14556 15266 14590 15296
rect 14629 15266 14663 15296
rect 14702 15266 14736 15296
rect 14775 15266 14809 15296
rect 14848 15266 14882 15296
rect 12860 15197 12869 15218
rect 12869 15197 12894 15218
rect 12934 15197 12938 15218
rect 12938 15197 12968 15218
rect 13008 15197 13041 15218
rect 13041 15197 13042 15218
rect 13082 15197 13110 15218
rect 13110 15197 13116 15218
rect 13156 15197 13179 15218
rect 13179 15197 13190 15218
rect 13230 15197 13248 15218
rect 13248 15197 13264 15218
rect 13304 15197 13317 15218
rect 13317 15197 13338 15218
rect 13378 15197 13386 15218
rect 13386 15197 13412 15218
rect 13452 15197 13455 15218
rect 13455 15197 13486 15218
rect 13526 15197 13559 15218
rect 13559 15197 13560 15218
rect 13600 15197 13628 15218
rect 13628 15197 13634 15218
rect 13674 15197 13697 15218
rect 13697 15197 13708 15218
rect 13748 15197 13766 15218
rect 13766 15197 13782 15218
rect 13822 15197 13835 15218
rect 13835 15197 13856 15218
rect 13896 15197 13904 15218
rect 13904 15197 13930 15218
rect 13970 15197 13973 15218
rect 13973 15197 14004 15218
rect 14044 15197 14076 15218
rect 14076 15197 14078 15218
rect 14118 15197 14145 15218
rect 14145 15197 14152 15218
rect 14191 15197 14214 15218
rect 14214 15197 14225 15218
rect 14264 15197 14283 15218
rect 14283 15197 14298 15218
rect 14337 15197 14352 15218
rect 14352 15197 14371 15218
rect 12860 15184 12894 15197
rect 12934 15184 12968 15197
rect 13008 15184 13042 15197
rect 13082 15184 13116 15197
rect 13156 15184 13190 15197
rect 13230 15184 13264 15197
rect 13304 15184 13338 15197
rect 13378 15184 13412 15197
rect 13452 15184 13486 15197
rect 13526 15184 13560 15197
rect 13600 15184 13634 15197
rect 13674 15184 13708 15197
rect 13748 15184 13782 15197
rect 13822 15184 13856 15197
rect 13896 15184 13930 15197
rect 13970 15184 14004 15197
rect 14044 15184 14078 15197
rect 14118 15184 14152 15197
rect 14191 15184 14225 15197
rect 14264 15184 14298 15197
rect 14337 15184 14371 15197
rect 14410 15192 14444 15218
rect 14483 15192 14517 15218
rect 14556 15192 14590 15218
rect 14629 15192 14663 15218
rect 14702 15192 14736 15218
rect 14775 15192 14809 15218
rect 14848 15192 14882 15218
rect 14410 15184 14420 15192
rect 14420 15184 14444 15192
rect 14483 15184 14492 15192
rect 14492 15184 14517 15192
rect 14556 15184 14564 15192
rect 14564 15184 14590 15192
rect 14629 15184 14636 15192
rect 14636 15184 14663 15192
rect 14702 15184 14708 15192
rect 14708 15184 14736 15192
rect 14775 15184 14780 15192
rect 14780 15184 14809 15192
rect 14848 15184 14852 15192
rect 14852 15184 14882 15192
rect 12860 15127 12869 15136
rect 12869 15127 12894 15136
rect 12934 15127 12938 15136
rect 12938 15127 12968 15136
rect 13008 15127 13041 15136
rect 13041 15127 13042 15136
rect 13082 15127 13110 15136
rect 13110 15127 13116 15136
rect 13156 15127 13179 15136
rect 13179 15127 13190 15136
rect 13230 15127 13248 15136
rect 13248 15127 13264 15136
rect 13304 15127 13317 15136
rect 13317 15127 13338 15136
rect 13378 15127 13386 15136
rect 13386 15127 13412 15136
rect 13452 15127 13455 15136
rect 13455 15127 13486 15136
rect 13526 15127 13559 15136
rect 13559 15127 13560 15136
rect 13600 15127 13628 15136
rect 13628 15127 13634 15136
rect 13674 15127 13697 15136
rect 13697 15127 13708 15136
rect 13748 15127 13766 15136
rect 13766 15127 13782 15136
rect 13822 15127 13835 15136
rect 13835 15127 13856 15136
rect 13896 15127 13904 15136
rect 13904 15127 13930 15136
rect 13970 15127 13973 15136
rect 13973 15127 14004 15136
rect 14044 15127 14076 15136
rect 14076 15127 14078 15136
rect 14118 15127 14145 15136
rect 14145 15127 14152 15136
rect 14191 15127 14214 15136
rect 14214 15127 14225 15136
rect 14264 15127 14283 15136
rect 14283 15127 14298 15136
rect 14337 15127 14352 15136
rect 14352 15127 14371 15136
rect 12860 15102 12894 15127
rect 12934 15102 12968 15127
rect 13008 15102 13042 15127
rect 13082 15102 13116 15127
rect 13156 15102 13190 15127
rect 13230 15102 13264 15127
rect 13304 15102 13338 15127
rect 13378 15102 13412 15127
rect 13452 15102 13486 15127
rect 13526 15102 13560 15127
rect 13600 15102 13634 15127
rect 13674 15102 13708 15127
rect 13748 15102 13782 15127
rect 13822 15102 13856 15127
rect 13896 15102 13930 15127
rect 13970 15102 14004 15127
rect 14044 15102 14078 15127
rect 14118 15102 14152 15127
rect 14191 15102 14225 15127
rect 14264 15102 14298 15127
rect 14337 15102 14371 15127
rect 14410 15123 14444 15136
rect 14483 15123 14517 15136
rect 14556 15123 14590 15136
rect 14629 15123 14663 15136
rect 14702 15123 14736 15136
rect 14775 15123 14809 15136
rect 14848 15123 14882 15136
rect 14410 15102 14420 15123
rect 14420 15102 14444 15123
rect 14483 15102 14492 15123
rect 14492 15102 14517 15123
rect 14556 15102 14564 15123
rect 14564 15102 14590 15123
rect 14629 15102 14636 15123
rect 14636 15102 14663 15123
rect 14702 15102 14708 15123
rect 14708 15102 14736 15123
rect 14775 15102 14780 15123
rect 14780 15102 14809 15123
rect 14848 15102 14852 15123
rect 14852 15102 14882 15123
rect 12860 15021 12894 15054
rect 12934 15021 12968 15054
rect 13008 15021 13042 15054
rect 13082 15021 13116 15054
rect 13156 15021 13190 15054
rect 13230 15021 13264 15054
rect 13304 15021 13338 15054
rect 13378 15021 13412 15054
rect 13452 15021 13486 15054
rect 13526 15021 13560 15054
rect 13600 15021 13634 15054
rect 13674 15021 13708 15054
rect 13748 15021 13782 15054
rect 13822 15021 13856 15054
rect 13896 15021 13930 15054
rect 13970 15021 14004 15054
rect 14044 15021 14078 15054
rect 14118 15021 14152 15054
rect 14191 15021 14225 15054
rect 14264 15021 14298 15054
rect 14337 15021 14371 15054
rect 12860 15020 12869 15021
rect 12869 15020 12894 15021
rect 12934 15020 12938 15021
rect 12938 15020 12968 15021
rect 13008 15020 13041 15021
rect 13041 15020 13042 15021
rect 13082 15020 13110 15021
rect 13110 15020 13116 15021
rect 13156 15020 13179 15021
rect 13179 15020 13190 15021
rect 13230 15020 13248 15021
rect 13248 15020 13264 15021
rect 13304 15020 13317 15021
rect 13317 15020 13338 15021
rect 13378 15020 13386 15021
rect 13386 15020 13412 15021
rect 13452 15020 13455 15021
rect 13455 15020 13486 15021
rect 13526 15020 13559 15021
rect 13559 15020 13560 15021
rect 13600 15020 13628 15021
rect 13628 15020 13634 15021
rect 13674 15020 13697 15021
rect 13697 15020 13708 15021
rect 13748 15020 13766 15021
rect 13766 15020 13782 15021
rect 13822 15020 13835 15021
rect 13835 15020 13856 15021
rect 13896 15020 13904 15021
rect 13904 15020 13930 15021
rect 13970 15020 13973 15021
rect 13973 15020 14004 15021
rect 14044 15020 14076 15021
rect 14076 15020 14078 15021
rect 14118 15020 14145 15021
rect 14145 15020 14152 15021
rect 14191 15020 14214 15021
rect 14214 15020 14225 15021
rect 14264 15020 14283 15021
rect 14283 15020 14298 15021
rect 14337 15020 14352 15021
rect 14352 15020 14371 15021
rect 14410 15020 14420 15054
rect 14420 15020 14444 15054
rect 14483 15020 14492 15054
rect 14492 15020 14517 15054
rect 14556 15020 14564 15054
rect 14564 15020 14590 15054
rect 14629 15020 14636 15054
rect 14636 15020 14663 15054
rect 14702 15020 14708 15054
rect 14708 15020 14736 15054
rect 14775 15020 14780 15054
rect 14780 15020 14809 15054
rect 14848 15020 14852 15054
rect 14852 15020 14882 15054
rect 12860 14951 12894 14972
rect 12934 14951 12968 14972
rect 13008 14951 13042 14972
rect 13082 14951 13116 14972
rect 13156 14951 13190 14972
rect 13230 14951 13264 14972
rect 13304 14951 13338 14972
rect 13378 14951 13412 14972
rect 13452 14951 13486 14972
rect 13526 14951 13560 14972
rect 13600 14951 13634 14972
rect 13674 14951 13708 14972
rect 13748 14951 13782 14972
rect 13822 14951 13856 14972
rect 13896 14951 13930 14972
rect 13970 14951 14004 14972
rect 14044 14951 14078 14972
rect 14118 14951 14152 14972
rect 14191 14951 14225 14972
rect 14264 14951 14298 14972
rect 14337 14951 14371 14972
rect 12860 14938 12869 14951
rect 12869 14938 12894 14951
rect 12934 14938 12938 14951
rect 12938 14938 12968 14951
rect 13008 14938 13041 14951
rect 13041 14938 13042 14951
rect 13082 14938 13110 14951
rect 13110 14938 13116 14951
rect 13156 14938 13179 14951
rect 13179 14938 13190 14951
rect 13230 14938 13248 14951
rect 13248 14938 13264 14951
rect 13304 14938 13317 14951
rect 13317 14938 13338 14951
rect 13378 14938 13386 14951
rect 13386 14938 13412 14951
rect 13452 14938 13455 14951
rect 13455 14938 13486 14951
rect 13526 14938 13559 14951
rect 13559 14938 13560 14951
rect 13600 14938 13628 14951
rect 13628 14938 13634 14951
rect 13674 14938 13697 14951
rect 13697 14938 13708 14951
rect 13748 14938 13766 14951
rect 13766 14938 13782 14951
rect 13822 14938 13835 14951
rect 13835 14938 13856 14951
rect 13896 14938 13904 14951
rect 13904 14938 13930 14951
rect 13970 14938 13973 14951
rect 13973 14938 14004 14951
rect 14044 14938 14076 14951
rect 14076 14938 14078 14951
rect 14118 14938 14145 14951
rect 14145 14938 14152 14951
rect 14191 14938 14214 14951
rect 14214 14938 14225 14951
rect 14264 14938 14283 14951
rect 14283 14938 14298 14951
rect 14337 14938 14352 14951
rect 14352 14938 14371 14951
rect 14410 14951 14420 14972
rect 14420 14951 14444 14972
rect 14483 14951 14492 14972
rect 14492 14951 14517 14972
rect 14556 14951 14564 14972
rect 14564 14951 14590 14972
rect 14629 14951 14636 14972
rect 14636 14951 14663 14972
rect 14702 14951 14708 14972
rect 14708 14951 14736 14972
rect 14775 14951 14780 14972
rect 14780 14951 14809 14972
rect 14848 14951 14852 14972
rect 14852 14951 14882 14972
rect 14410 14938 14444 14951
rect 14483 14938 14517 14951
rect 14556 14938 14590 14951
rect 14629 14938 14663 14951
rect 14702 14938 14736 14951
rect 14775 14938 14809 14951
rect 14848 14938 14882 14951
rect -484 9510 -482 9514
rect -482 9510 -450 9514
rect -411 9510 -378 9514
rect -378 9510 -377 9514
rect -338 9510 -309 9514
rect -309 9510 -304 9514
rect -265 9510 -240 9514
rect -240 9510 -231 9514
rect -192 9510 -171 9514
rect -171 9510 -158 9514
rect -119 9510 -102 9514
rect -102 9510 -85 9514
rect -484 9480 -450 9510
rect -411 9480 -377 9510
rect -338 9480 -304 9510
rect -265 9480 -231 9510
rect -192 9480 -158 9510
rect -119 9480 -85 9510
rect -46 9480 -33 9514
rect -33 9480 -12 9514
rect 27 9480 61 9514
rect 100 9480 134 9514
rect 173 9480 207 9514
rect 246 9480 280 9514
rect 319 9480 353 9514
rect 392 9480 426 9514
rect 465 9480 499 9514
rect 538 9480 572 9514
rect 611 9480 645 9514
rect 684 9480 718 9514
rect 757 9480 791 9514
rect 830 9480 864 9514
rect 903 9480 937 9514
rect 976 9480 1010 9514
rect 1049 9480 1083 9514
rect 1122 9480 1156 9514
rect 1195 9480 1229 9514
rect 1268 9480 1302 9514
rect 1341 9480 1375 9514
rect 1414 9480 1448 9514
rect 1487 9480 1521 9514
rect 1559 9480 1593 9514
rect 1631 9480 1665 9514
rect 1703 9480 1737 9514
rect 1775 9480 1809 9514
rect 1847 9480 1881 9514
rect 1919 9480 1953 9514
rect 1991 9480 2025 9514
rect 2063 9480 2097 9514
rect 2135 9480 2169 9514
rect 2207 9480 2241 9514
rect 2279 9480 2313 9514
rect 2351 9480 2385 9514
rect 2423 9480 2457 9514
rect 2495 9480 2529 9514
rect 2567 9480 2601 9514
rect 2639 9480 2673 9514
rect 2711 9480 2745 9514
rect 2783 9480 2817 9514
rect 2855 9480 2889 9514
rect 2927 9480 2961 9514
rect 2999 9480 3033 9514
rect 3071 9480 3105 9514
rect 3143 9480 3177 9514
rect 3215 9480 3249 9514
rect 3287 9480 3321 9514
rect 3359 9480 3393 9514
rect 3431 9480 3465 9514
rect 3503 9480 3537 9514
rect 3575 9480 3609 9514
rect 3647 9480 3681 9514
rect 3719 9480 3753 9514
rect 3791 9480 3825 9514
rect 3863 9480 3897 9514
rect 3935 9480 3969 9514
rect 4007 9480 4041 9514
rect 4079 9480 4113 9514
rect 4151 9480 4185 9514
rect 4223 9480 4257 9514
rect 4295 9480 4329 9514
rect 4367 9480 4401 9514
rect 4439 9480 4473 9514
rect 4511 9480 4545 9514
rect 4583 9480 4617 9514
rect 4655 9480 4689 9514
rect 4727 9480 4761 9514
rect 4799 9480 4833 9514
rect 4871 9480 4905 9514
rect 4943 9480 4977 9514
rect 5015 9480 5049 9514
rect 5087 9480 5121 9514
rect 5159 9480 5193 9514
rect 5231 9480 5265 9514
rect 5303 9480 5337 9514
rect 5375 9480 5409 9514
rect 5447 9480 5481 9514
rect 5519 9480 5553 9514
rect 5591 9480 5625 9514
rect 5663 9480 5697 9514
rect 5735 9480 5769 9514
rect 5807 9480 5841 9514
rect 5879 9480 5913 9514
rect 5951 9480 5985 9514
rect 6023 9480 6057 9514
rect 6095 9480 6129 9514
rect 6167 9480 6201 9514
rect 6239 9480 6273 9514
rect 6311 9480 6345 9514
rect 6383 9480 6417 9514
rect 6455 9480 6489 9514
rect 6527 9480 6561 9514
rect 6599 9480 6633 9514
rect 6671 9480 6705 9514
rect 6743 9480 6777 9514
rect 6815 9480 6849 9514
rect 6887 9480 6921 9514
rect 6959 9480 6993 9514
rect 7031 9480 7065 9514
rect 7103 9480 7137 9514
rect 7175 9480 7209 9514
rect 7247 9480 7281 9514
rect 7319 9480 7353 9514
rect 7391 9480 7425 9514
rect 7463 9480 7497 9514
rect 7535 9480 7569 9514
rect 7607 9480 7641 9514
rect 7679 9480 7713 9514
rect 7751 9480 7785 9514
rect 7823 9480 7857 9514
rect 7895 9480 7929 9514
rect 7967 9480 8001 9514
rect 8039 9480 8073 9514
rect 8111 9480 8145 9514
rect 8183 9480 8217 9514
rect 8255 9480 8289 9514
rect 8327 9480 8361 9514
rect 8399 9480 8433 9514
rect 8471 9480 8505 9514
rect 8543 9480 8577 9514
rect 8615 9480 8649 9514
rect 8687 9480 8721 9514
rect 8759 9480 8793 9514
rect 8831 9480 8865 9514
rect 8903 9480 8937 9514
rect 8975 9480 9009 9514
rect 9047 9480 9081 9514
rect 9119 9480 9153 9514
rect 9191 9480 9225 9514
rect 9263 9480 9297 9514
rect 9335 9480 9369 9514
rect 9407 9480 9441 9514
rect 9479 9480 9513 9514
rect 9551 9480 9585 9514
rect 9623 9480 9657 9514
rect 9695 9480 9729 9514
rect 9767 9480 9801 9514
rect 9839 9480 9873 9514
rect 9911 9480 9945 9514
rect 9983 9480 10017 9514
rect 10055 9480 10089 9514
rect 10127 9480 10161 9514
rect 10199 9480 10233 9514
rect 10271 9480 10305 9514
rect 10343 9480 10377 9514
rect 10415 9480 10449 9514
rect 10487 9480 10521 9514
rect 10559 9480 10593 9514
rect 10631 9480 10665 9514
rect 10703 9480 10737 9514
rect 10775 9480 10809 9514
rect 10847 9480 10881 9514
rect 10919 9480 10953 9514
rect 10991 9480 11025 9514
rect 11063 9480 11097 9514
rect 11135 9480 11169 9514
rect 11207 9480 11241 9514
rect 11279 9480 11313 9514
rect 11351 9480 11385 9514
rect 11423 9480 11457 9514
rect 11495 9480 11529 9514
rect 11567 9480 11601 9514
rect 11639 9480 11673 9514
rect 11711 9480 11745 9514
rect 11783 9480 11817 9514
rect 11855 9480 11889 9514
rect 11927 9480 11961 9514
rect 11999 9480 12033 9514
rect 12071 9480 12105 9514
rect 12143 9480 12177 9514
rect 12215 9480 12249 9514
rect 12287 9480 12321 9514
rect 12359 9480 12393 9514
rect 12431 9480 12465 9514
rect 12503 9480 12537 9514
rect 12575 9480 12609 9514
rect 12647 9480 12681 9514
rect 12719 9480 12753 9514
rect 12791 9480 12825 9514
rect 12863 9480 12897 9514
rect 12935 9480 12969 9514
rect 13007 9480 13041 9514
rect 13079 9480 13113 9514
rect 13151 9480 13185 9514
rect 13223 9480 13257 9514
rect 13295 9480 13329 9514
rect 13367 9480 13401 9514
rect 13439 9480 13473 9514
rect 13511 9480 13545 9514
rect 13583 9480 13617 9514
rect 13655 9480 13689 9514
rect 13727 9480 13761 9514
rect 13799 9480 13833 9514
rect -484 9408 -450 9428
rect -411 9408 -377 9428
rect -338 9408 -304 9428
rect -265 9408 -231 9428
rect -192 9408 -158 9428
rect -119 9408 -85 9428
rect -484 9394 -482 9408
rect -482 9394 -450 9408
rect -411 9394 -378 9408
rect -378 9394 -377 9408
rect -338 9394 -309 9408
rect -309 9394 -304 9408
rect -265 9394 -240 9408
rect -240 9394 -231 9408
rect -192 9394 -171 9408
rect -171 9394 -158 9408
rect -119 9394 -102 9408
rect -102 9394 -85 9408
rect -46 9394 -33 9428
rect -33 9394 -12 9428
rect 27 9394 61 9428
rect 100 9394 134 9428
rect 173 9394 207 9428
rect 246 9394 280 9428
rect 319 9394 353 9428
rect 392 9394 426 9428
rect 465 9394 499 9428
rect 538 9394 572 9428
rect 611 9394 645 9428
rect 684 9394 718 9428
rect 757 9394 791 9428
rect 830 9394 864 9428
rect 903 9394 937 9428
rect 976 9394 1010 9428
rect 1049 9394 1083 9428
rect 1122 9394 1156 9428
rect 1195 9394 1229 9428
rect 1268 9394 1302 9428
rect 1341 9394 1375 9428
rect 1414 9394 1448 9428
rect 1487 9394 1521 9428
rect 1559 9394 1593 9428
rect 1631 9394 1665 9428
rect 1703 9394 1737 9428
rect 1775 9394 1809 9428
rect 1847 9394 1881 9428
rect 1919 9394 1953 9428
rect 1991 9394 2025 9428
rect 2063 9394 2097 9428
rect 2135 9394 2169 9428
rect 2207 9394 2241 9428
rect 2279 9394 2313 9428
rect 2351 9394 2385 9428
rect 2423 9394 2457 9428
rect 2495 9394 2529 9428
rect 2567 9394 2601 9428
rect 2639 9394 2673 9428
rect 2711 9394 2745 9428
rect 2783 9394 2817 9428
rect 2855 9394 2889 9428
rect 2927 9394 2961 9428
rect 2999 9394 3033 9428
rect 3071 9394 3105 9428
rect 3143 9394 3177 9428
rect 3215 9394 3249 9428
rect 3287 9394 3321 9428
rect 3359 9394 3393 9428
rect 3431 9394 3465 9428
rect 3503 9394 3537 9428
rect 3575 9394 3609 9428
rect 3647 9394 3681 9428
rect 3719 9394 3753 9428
rect 3791 9394 3825 9428
rect 3863 9394 3897 9428
rect 3935 9394 3969 9428
rect 4007 9394 4041 9428
rect 4079 9394 4113 9428
rect 4151 9394 4185 9428
rect 4223 9394 4257 9428
rect 4295 9394 4329 9428
rect 4367 9394 4401 9428
rect 4439 9394 4473 9428
rect 4511 9394 4545 9428
rect 4583 9394 4617 9428
rect 4655 9394 4689 9428
rect 4727 9394 4761 9428
rect 4799 9394 4833 9428
rect 4871 9394 4905 9428
rect 4943 9394 4977 9428
rect 5015 9394 5049 9428
rect 5087 9394 5121 9428
rect 5159 9394 5193 9428
rect 5231 9394 5265 9428
rect 5303 9394 5337 9428
rect 5375 9394 5409 9428
rect 5447 9394 5481 9428
rect 5519 9394 5553 9428
rect 5591 9394 5625 9428
rect 5663 9394 5697 9428
rect 5735 9394 5769 9428
rect 5807 9394 5841 9428
rect 5879 9394 5913 9428
rect 5951 9394 5985 9428
rect 6023 9394 6057 9428
rect 6095 9394 6129 9428
rect 6167 9394 6201 9428
rect 6239 9394 6273 9428
rect 6311 9394 6345 9428
rect 6383 9394 6417 9428
rect 6455 9394 6489 9428
rect 6527 9394 6561 9428
rect 6599 9394 6633 9428
rect 6671 9394 6705 9428
rect 6743 9394 6777 9428
rect 6815 9394 6849 9428
rect 6887 9394 6921 9428
rect 6959 9394 6993 9428
rect 7031 9394 7065 9428
rect 7103 9394 7137 9428
rect 7175 9394 7209 9428
rect 7247 9394 7281 9428
rect 7319 9394 7353 9428
rect 7391 9394 7425 9428
rect 7463 9394 7497 9428
rect 7535 9394 7569 9428
rect 7607 9394 7641 9428
rect 7679 9394 7713 9428
rect 7751 9394 7785 9428
rect 7823 9394 7857 9428
rect 7895 9394 7929 9428
rect 7967 9394 8001 9428
rect 8039 9394 8073 9428
rect 8111 9394 8145 9428
rect 8183 9394 8217 9428
rect 8255 9394 8289 9428
rect 8327 9394 8361 9428
rect 8399 9394 8433 9428
rect 8471 9394 8505 9428
rect 8543 9394 8577 9428
rect 8615 9394 8649 9428
rect 8687 9394 8721 9428
rect 8759 9394 8793 9428
rect 8831 9394 8865 9428
rect 8903 9394 8937 9428
rect 8975 9394 9009 9428
rect 9047 9394 9081 9428
rect 9119 9394 9153 9428
rect 9191 9394 9225 9428
rect 9263 9394 9297 9428
rect 9335 9394 9369 9428
rect 9407 9394 9441 9428
rect 9479 9394 9513 9428
rect 9551 9394 9585 9428
rect 9623 9394 9657 9428
rect 9695 9394 9729 9428
rect 9767 9394 9801 9428
rect 9839 9394 9873 9428
rect 9911 9394 9945 9428
rect 9983 9394 10017 9428
rect 10055 9394 10089 9428
rect 10127 9394 10161 9428
rect 10199 9394 10233 9428
rect 10271 9394 10305 9428
rect 10343 9394 10377 9428
rect 10415 9394 10449 9428
rect 10487 9394 10521 9428
rect 10559 9394 10593 9428
rect 10631 9394 10665 9428
rect 10703 9394 10737 9428
rect 10775 9394 10809 9428
rect 10847 9394 10881 9428
rect 10919 9394 10953 9428
rect 10991 9394 11025 9428
rect 11063 9394 11097 9428
rect 11135 9394 11169 9428
rect 11207 9394 11241 9428
rect 11279 9394 11313 9428
rect 11351 9394 11385 9428
rect 11423 9394 11457 9428
rect 11495 9394 11529 9428
rect 11567 9394 11601 9428
rect 11639 9394 11673 9428
rect 11711 9394 11745 9428
rect 11783 9394 11817 9428
rect 11855 9394 11889 9428
rect 11927 9394 11961 9428
rect 11999 9394 12033 9428
rect 12071 9394 12105 9428
rect 12143 9394 12177 9428
rect 12215 9394 12249 9428
rect 12287 9394 12321 9428
rect 12359 9394 12393 9428
rect 12431 9394 12465 9428
rect 12503 9394 12537 9428
rect 12575 9394 12609 9428
rect 12647 9394 12681 9428
rect 12719 9394 12753 9428
rect 12791 9394 12825 9428
rect 12863 9394 12897 9428
rect 12935 9394 12969 9428
rect 13007 9394 13041 9428
rect 13079 9394 13113 9428
rect 13151 9394 13185 9428
rect 13223 9394 13257 9428
rect 13295 9394 13329 9428
rect 13367 9394 13401 9428
rect 13439 9394 13473 9428
rect 13511 9394 13545 9428
rect 13583 9394 13617 9428
rect 13655 9394 13689 9428
rect 13727 9394 13761 9428
rect 13799 9394 13833 9428
rect -484 9340 -450 9342
rect -411 9340 -377 9342
rect -338 9340 -304 9342
rect -265 9340 -231 9342
rect -192 9340 -158 9342
rect -119 9340 -85 9342
rect -484 9308 -482 9340
rect -482 9308 -450 9340
rect -411 9308 -378 9340
rect -378 9308 -377 9340
rect -338 9308 -309 9340
rect -309 9308 -304 9340
rect -265 9308 -240 9340
rect -240 9308 -231 9340
rect -192 9308 -171 9340
rect -171 9308 -158 9340
rect -119 9308 -102 9340
rect -102 9308 -85 9340
rect -46 9308 -33 9342
rect -33 9308 -12 9342
rect 27 9308 61 9342
rect 100 9308 134 9342
rect 173 9308 207 9342
rect 246 9308 280 9342
rect 319 9308 353 9342
rect 392 9308 426 9342
rect 465 9308 499 9342
rect 538 9308 572 9342
rect 611 9308 645 9342
rect 684 9308 718 9342
rect 757 9308 791 9342
rect 830 9308 864 9342
rect 903 9308 937 9342
rect 976 9308 1010 9342
rect 1049 9308 1083 9342
rect 1122 9308 1156 9342
rect 1195 9308 1229 9342
rect 1268 9308 1302 9342
rect 1341 9308 1375 9342
rect 1414 9308 1448 9342
rect 1487 9308 1521 9342
rect 1559 9308 1593 9342
rect 1631 9308 1665 9342
rect 1703 9308 1737 9342
rect 1775 9308 1809 9342
rect 1847 9308 1881 9342
rect 1919 9308 1953 9342
rect 1991 9308 2025 9342
rect 2063 9308 2097 9342
rect 2135 9308 2169 9342
rect 2207 9308 2241 9342
rect 2279 9308 2313 9342
rect 2351 9308 2385 9342
rect 2423 9308 2457 9342
rect 2495 9308 2529 9342
rect 2567 9308 2601 9342
rect 2639 9308 2673 9342
rect 2711 9308 2745 9342
rect 2783 9308 2817 9342
rect 2855 9308 2889 9342
rect 2927 9308 2961 9342
rect 2999 9308 3033 9342
rect 3071 9308 3105 9342
rect 3143 9308 3177 9342
rect 3215 9308 3249 9342
rect 3287 9308 3321 9342
rect 3359 9308 3393 9342
rect 3431 9308 3465 9342
rect 3503 9308 3537 9342
rect 3575 9308 3609 9342
rect 3647 9308 3681 9342
rect 3719 9308 3753 9342
rect 3791 9308 3825 9342
rect 3863 9308 3897 9342
rect 3935 9308 3969 9342
rect 4007 9308 4041 9342
rect 4079 9308 4113 9342
rect 4151 9308 4185 9342
rect 4223 9308 4257 9342
rect 4295 9308 4329 9342
rect 4367 9308 4401 9342
rect 4439 9308 4473 9342
rect 4511 9308 4545 9342
rect 4583 9308 4617 9342
rect 4655 9308 4689 9342
rect 4727 9308 4761 9342
rect 4799 9308 4833 9342
rect 4871 9308 4905 9342
rect 4943 9308 4977 9342
rect 5015 9308 5049 9342
rect 5087 9308 5121 9342
rect 5159 9308 5193 9342
rect 5231 9308 5265 9342
rect 5303 9308 5337 9342
rect 5375 9308 5409 9342
rect 5447 9308 5481 9342
rect 5519 9308 5553 9342
rect 5591 9308 5625 9342
rect 5663 9308 5697 9342
rect 5735 9308 5769 9342
rect 5807 9308 5841 9342
rect 5879 9308 5913 9342
rect 5951 9308 5985 9342
rect 6023 9308 6057 9342
rect 6095 9308 6129 9342
rect 6167 9308 6201 9342
rect 6239 9308 6273 9342
rect 6311 9308 6345 9342
rect 6383 9308 6417 9342
rect 6455 9308 6489 9342
rect 6527 9308 6561 9342
rect 6599 9308 6633 9342
rect 6671 9308 6705 9342
rect 6743 9308 6777 9342
rect 6815 9308 6849 9342
rect 6887 9308 6921 9342
rect 6959 9308 6993 9342
rect 7031 9308 7065 9342
rect 7103 9308 7137 9342
rect 7175 9308 7209 9342
rect 7247 9308 7281 9342
rect 7319 9308 7353 9342
rect 7391 9308 7425 9342
rect 7463 9308 7497 9342
rect 7535 9308 7569 9342
rect 7607 9308 7641 9342
rect 7679 9308 7713 9342
rect 7751 9308 7785 9342
rect 7823 9308 7857 9342
rect 7895 9308 7929 9342
rect 7967 9308 8001 9342
rect 8039 9308 8073 9342
rect 8111 9308 8145 9342
rect 8183 9308 8217 9342
rect 8255 9308 8289 9342
rect 8327 9308 8361 9342
rect 8399 9308 8433 9342
rect 8471 9308 8505 9342
rect 8543 9308 8577 9342
rect 8615 9308 8649 9342
rect 8687 9308 8721 9342
rect 8759 9308 8793 9342
rect 8831 9308 8865 9342
rect 8903 9308 8937 9342
rect 8975 9308 9009 9342
rect 9047 9308 9081 9342
rect 9119 9308 9153 9342
rect 9191 9308 9225 9342
rect 9263 9308 9297 9342
rect 9335 9308 9369 9342
rect 9407 9308 9441 9342
rect 9479 9308 9513 9342
rect 9551 9308 9585 9342
rect 9623 9308 9657 9342
rect 9695 9308 9729 9342
rect 9767 9308 9801 9342
rect 9839 9308 9873 9342
rect 9911 9308 9945 9342
rect 9983 9308 10017 9342
rect 10055 9308 10089 9342
rect 10127 9308 10161 9342
rect 10199 9308 10233 9342
rect 10271 9308 10305 9342
rect 10343 9308 10377 9342
rect 10415 9308 10449 9342
rect 10487 9308 10521 9342
rect 10559 9308 10593 9342
rect 10631 9308 10665 9342
rect 10703 9308 10737 9342
rect 10775 9308 10809 9342
rect 10847 9308 10881 9342
rect 10919 9308 10953 9342
rect 10991 9308 11025 9342
rect 11063 9308 11097 9342
rect 11135 9308 11169 9342
rect 11207 9308 11241 9342
rect 11279 9308 11313 9342
rect 11351 9308 11385 9342
rect 11423 9308 11457 9342
rect 11495 9308 11529 9342
rect 11567 9308 11601 9342
rect 11639 9308 11673 9342
rect 11711 9308 11745 9342
rect 11783 9308 11817 9342
rect 11855 9308 11889 9342
rect 11927 9308 11961 9342
rect 11999 9308 12033 9342
rect 12071 9308 12105 9342
rect 12143 9308 12177 9342
rect 12215 9308 12249 9342
rect 12287 9308 12321 9342
rect 12359 9308 12393 9342
rect 12431 9308 12465 9342
rect 12503 9308 12537 9342
rect 12575 9308 12609 9342
rect 12647 9308 12681 9342
rect 12719 9308 12753 9342
rect 12791 9308 12825 9342
rect 12863 9308 12897 9342
rect 12935 9308 12969 9342
rect 13007 9308 13041 9342
rect 13079 9308 13113 9342
rect 13151 9308 13185 9342
rect 13223 9308 13257 9342
rect 13295 9308 13329 9342
rect 13367 9308 13401 9342
rect 13439 9308 13473 9342
rect 13511 9308 13545 9342
rect 13583 9308 13617 9342
rect 13655 9308 13689 9342
rect 13727 9308 13761 9342
rect 13799 9308 13833 9342
rect -484 9238 -482 9256
rect -482 9238 -450 9256
rect -411 9238 -378 9256
rect -378 9238 -377 9256
rect -338 9238 -309 9256
rect -309 9238 -304 9256
rect -265 9238 -240 9256
rect -240 9238 -231 9256
rect -192 9238 -171 9256
rect -171 9238 -158 9256
rect -119 9238 -102 9256
rect -102 9238 -85 9256
rect -484 9222 -450 9238
rect -411 9222 -377 9238
rect -338 9222 -304 9238
rect -265 9222 -231 9238
rect -192 9222 -158 9238
rect -119 9222 -85 9238
rect -46 9222 -33 9256
rect -33 9222 -12 9256
rect 27 9222 61 9256
rect 100 9222 134 9256
rect 173 9222 207 9256
rect 246 9222 280 9256
rect 319 9222 353 9256
rect 392 9222 426 9256
rect 465 9222 499 9256
rect 538 9222 572 9256
rect 611 9222 645 9256
rect 684 9222 718 9256
rect 757 9222 791 9256
rect 830 9222 864 9256
rect 903 9222 937 9256
rect 976 9222 1010 9256
rect 1049 9222 1083 9256
rect 1122 9222 1156 9256
rect 1195 9222 1229 9256
rect 1268 9222 1302 9256
rect 1341 9222 1375 9256
rect 1414 9222 1448 9256
rect 1487 9222 1521 9256
rect 1559 9222 1593 9256
rect 1631 9222 1665 9256
rect 1703 9222 1737 9256
rect 1775 9222 1809 9256
rect 1847 9222 1881 9256
rect 1919 9222 1953 9256
rect 1991 9222 2025 9256
rect 2063 9222 2097 9256
rect 2135 9222 2169 9256
rect 2207 9222 2241 9256
rect 2279 9222 2313 9256
rect 2351 9222 2385 9256
rect 2423 9222 2457 9256
rect 2495 9222 2529 9256
rect 2567 9222 2601 9256
rect 2639 9222 2673 9256
rect 2711 9222 2745 9256
rect 2783 9222 2817 9256
rect 2855 9222 2889 9256
rect 2927 9222 2961 9256
rect 2999 9222 3033 9256
rect 3071 9222 3105 9256
rect 3143 9222 3177 9256
rect 3215 9222 3249 9256
rect 3287 9222 3321 9256
rect 3359 9222 3393 9256
rect 3431 9222 3465 9256
rect 3503 9222 3537 9256
rect 3575 9222 3609 9256
rect 3647 9222 3681 9256
rect 3719 9222 3753 9256
rect 3791 9222 3825 9256
rect 3863 9222 3897 9256
rect 3935 9222 3969 9256
rect 4007 9222 4041 9256
rect 4079 9222 4113 9256
rect 4151 9222 4185 9256
rect 4223 9222 4257 9256
rect 4295 9222 4329 9256
rect 4367 9222 4401 9256
rect 4439 9222 4473 9256
rect 4511 9222 4545 9256
rect 4583 9222 4617 9256
rect 4655 9222 4689 9256
rect 4727 9222 4761 9256
rect 4799 9222 4833 9256
rect 4871 9222 4905 9256
rect 4943 9222 4977 9256
rect 5015 9222 5049 9256
rect 5087 9222 5121 9256
rect 5159 9222 5193 9256
rect 5231 9222 5265 9256
rect 5303 9222 5337 9256
rect 5375 9222 5409 9256
rect 5447 9222 5481 9256
rect 5519 9222 5553 9256
rect 5591 9222 5625 9256
rect 5663 9222 5697 9256
rect 5735 9222 5769 9256
rect 5807 9222 5841 9256
rect 5879 9222 5913 9256
rect 5951 9222 5985 9256
rect 6023 9222 6057 9256
rect 6095 9222 6129 9256
rect 6167 9222 6201 9256
rect 6239 9222 6273 9256
rect 6311 9222 6345 9256
rect 6383 9222 6417 9256
rect 6455 9222 6489 9256
rect 6527 9222 6561 9256
rect 6599 9222 6633 9256
rect 6671 9222 6705 9256
rect 6743 9222 6777 9256
rect 6815 9222 6849 9256
rect 6887 9222 6921 9256
rect 6959 9222 6993 9256
rect 7031 9222 7065 9256
rect 7103 9222 7137 9256
rect 7175 9222 7209 9256
rect 7247 9222 7281 9256
rect 7319 9222 7353 9256
rect 7391 9222 7425 9256
rect 7463 9222 7497 9256
rect 7535 9222 7569 9256
rect 7607 9222 7641 9256
rect 7679 9222 7713 9256
rect 7751 9222 7785 9256
rect 7823 9222 7857 9256
rect 7895 9222 7929 9256
rect 7967 9222 8001 9256
rect 8039 9222 8073 9256
rect 8111 9222 8145 9256
rect 8183 9222 8217 9256
rect 8255 9222 8289 9256
rect 8327 9222 8361 9256
rect 8399 9222 8433 9256
rect 8471 9222 8505 9256
rect 8543 9222 8577 9256
rect 8615 9222 8649 9256
rect 8687 9222 8721 9256
rect 8759 9222 8793 9256
rect 8831 9222 8865 9256
rect 8903 9222 8937 9256
rect 8975 9222 9009 9256
rect 9047 9222 9081 9256
rect 9119 9222 9153 9256
rect 9191 9222 9225 9256
rect 9263 9222 9297 9256
rect 9335 9222 9369 9256
rect 9407 9222 9441 9256
rect 9479 9222 9513 9256
rect 9551 9222 9585 9256
rect 9623 9222 9657 9256
rect 9695 9222 9729 9256
rect 9767 9222 9801 9256
rect 9839 9222 9873 9256
rect 9911 9222 9945 9256
rect 9983 9222 10017 9256
rect 10055 9222 10089 9256
rect 10127 9222 10161 9256
rect 10199 9222 10233 9256
rect 10271 9222 10305 9256
rect 10343 9222 10377 9256
rect 10415 9222 10449 9256
rect 10487 9222 10521 9256
rect 10559 9222 10593 9256
rect 10631 9222 10665 9256
rect 10703 9222 10737 9256
rect 10775 9222 10809 9256
rect 10847 9222 10881 9256
rect 10919 9222 10953 9256
rect 10991 9222 11025 9256
rect 11063 9222 11097 9256
rect 11135 9222 11169 9256
rect 11207 9222 11241 9256
rect 11279 9222 11313 9256
rect 11351 9222 11385 9256
rect 11423 9222 11457 9256
rect 11495 9222 11529 9256
rect 11567 9222 11601 9256
rect 11639 9222 11673 9256
rect 11711 9222 11745 9256
rect 11783 9222 11817 9256
rect 11855 9222 11889 9256
rect 11927 9222 11961 9256
rect 11999 9222 12033 9256
rect 12071 9222 12105 9256
rect 12143 9222 12177 9256
rect 12215 9222 12249 9256
rect 12287 9222 12321 9256
rect 12359 9222 12393 9256
rect 12431 9222 12465 9256
rect 12503 9222 12537 9256
rect 12575 9222 12609 9256
rect 12647 9222 12681 9256
rect 12719 9222 12753 9256
rect 12791 9222 12825 9256
rect 12863 9222 12897 9256
rect 12935 9222 12969 9256
rect 13007 9222 13041 9256
rect 13079 9222 13113 9256
rect 13151 9222 13185 9256
rect 13223 9222 13257 9256
rect 13295 9222 13329 9256
rect 13367 9222 13401 9256
rect 13439 9222 13473 9256
rect 13511 9222 13545 9256
rect 13583 9222 13617 9256
rect 13655 9222 13689 9256
rect 13727 9222 13761 9256
rect 13799 9222 13833 9256
rect -484 9136 -450 9170
rect -411 9136 -377 9170
rect -338 9136 -304 9170
rect -265 9136 -231 9170
rect -192 9136 -158 9170
rect -119 9136 -85 9170
rect -46 9136 -33 9170
rect -33 9136 -12 9170
rect 27 9136 61 9170
rect 100 9136 134 9170
rect 173 9136 207 9170
rect 246 9136 280 9170
rect 319 9136 353 9170
rect 392 9136 426 9170
rect 465 9136 499 9170
rect 538 9136 572 9170
rect 611 9136 645 9170
rect 684 9136 718 9170
rect 757 9136 791 9170
rect 830 9136 864 9170
rect 903 9136 937 9170
rect 976 9136 1010 9170
rect 1049 9136 1083 9170
rect 1122 9136 1156 9170
rect 1195 9136 1229 9170
rect 1268 9136 1302 9170
rect 1341 9136 1375 9170
rect 1414 9136 1448 9170
rect 1487 9136 1521 9170
rect 1559 9136 1593 9170
rect 1631 9136 1665 9170
rect 1703 9136 1737 9170
rect 1775 9136 1809 9170
rect 1847 9136 1881 9170
rect 1919 9136 1953 9170
rect 1991 9136 2025 9170
rect 2063 9136 2097 9170
rect 2135 9136 2169 9170
rect 2207 9136 2241 9170
rect 2279 9136 2313 9170
rect 2351 9136 2385 9170
rect 2423 9136 2457 9170
rect 2495 9136 2529 9170
rect 2567 9136 2601 9170
rect 2639 9136 2673 9170
rect 2711 9136 2745 9170
rect 2783 9136 2817 9170
rect 2855 9136 2889 9170
rect 2927 9136 2961 9170
rect 2999 9136 3033 9170
rect 3071 9136 3105 9170
rect 3143 9136 3177 9170
rect 3215 9136 3249 9170
rect 3287 9136 3321 9170
rect 3359 9136 3393 9170
rect 3431 9136 3465 9170
rect 3503 9136 3537 9170
rect 3575 9136 3609 9170
rect 3647 9136 3681 9170
rect 3719 9136 3753 9170
rect 3791 9136 3825 9170
rect 3863 9136 3897 9170
rect 3935 9136 3969 9170
rect 4007 9136 4041 9170
rect 4079 9136 4113 9170
rect 4151 9136 4185 9170
rect 4223 9136 4257 9170
rect 4295 9136 4329 9170
rect 4367 9136 4401 9170
rect 4439 9136 4473 9170
rect 4511 9136 4545 9170
rect 4583 9136 4617 9170
rect 4655 9136 4689 9170
rect 4727 9136 4761 9170
rect 4799 9136 4833 9170
rect 4871 9136 4905 9170
rect 4943 9136 4977 9170
rect 5015 9136 5049 9170
rect 5087 9136 5121 9170
rect 5159 9136 5193 9170
rect 5231 9136 5265 9170
rect 5303 9136 5337 9170
rect 5375 9136 5409 9170
rect 5447 9136 5481 9170
rect 5519 9136 5553 9170
rect 5591 9136 5625 9170
rect 5663 9136 5697 9170
rect 5735 9136 5769 9170
rect 5807 9136 5841 9170
rect 5879 9136 5913 9170
rect 5951 9136 5985 9170
rect 6023 9136 6057 9170
rect 6095 9136 6129 9170
rect 6167 9136 6201 9170
rect 6239 9136 6273 9170
rect 6311 9136 6345 9170
rect 6383 9136 6417 9170
rect 6455 9136 6489 9170
rect 6527 9136 6561 9170
rect 6599 9136 6633 9170
rect 6671 9136 6705 9170
rect 6743 9136 6777 9170
rect 6815 9136 6849 9170
rect 6887 9136 6921 9170
rect 6959 9136 6993 9170
rect 7031 9136 7065 9170
rect 7103 9136 7137 9170
rect 7175 9136 7209 9170
rect 7247 9136 7281 9170
rect 7319 9136 7353 9170
rect 7391 9136 7425 9170
rect 7463 9136 7497 9170
rect 7535 9136 7569 9170
rect 7607 9136 7641 9170
rect 7679 9136 7713 9170
rect 7751 9136 7785 9170
rect 7823 9136 7857 9170
rect 7895 9136 7929 9170
rect 7967 9136 8001 9170
rect 8039 9136 8073 9170
rect 8111 9136 8145 9170
rect 8183 9136 8217 9170
rect 8255 9136 8289 9170
rect 8327 9136 8361 9170
rect 8399 9136 8433 9170
rect 8471 9136 8505 9170
rect 8543 9136 8577 9170
rect 8615 9136 8649 9170
rect 8687 9136 8721 9170
rect 8759 9136 8793 9170
rect 8831 9136 8865 9170
rect 8903 9136 8937 9170
rect 8975 9136 9009 9170
rect 9047 9136 9081 9170
rect 9119 9136 9153 9170
rect 9191 9136 9225 9170
rect 9263 9136 9297 9170
rect 9335 9136 9369 9170
rect 9407 9136 9441 9170
rect 9479 9136 9513 9170
rect 9551 9136 9585 9170
rect 9623 9136 9657 9170
rect 9695 9136 9729 9170
rect 9767 9136 9801 9170
rect 9839 9136 9873 9170
rect 9911 9136 9945 9170
rect 9983 9136 10017 9170
rect 10055 9136 10089 9170
rect 10127 9136 10161 9170
rect 10199 9136 10233 9170
rect 10271 9136 10305 9170
rect 10343 9136 10377 9170
rect 10415 9136 10449 9170
rect 10487 9136 10521 9170
rect 10559 9136 10593 9170
rect 10631 9136 10665 9170
rect 10703 9136 10737 9170
rect 10775 9136 10809 9170
rect 10847 9136 10881 9170
rect 10919 9136 10953 9170
rect 10991 9136 11025 9170
rect 11063 9136 11097 9170
rect 11135 9136 11169 9170
rect 11207 9136 11241 9170
rect 11279 9136 11313 9170
rect 11351 9136 11385 9170
rect 11423 9136 11457 9170
rect 11495 9136 11529 9170
rect 11567 9136 11601 9170
rect 11639 9136 11673 9170
rect 11711 9136 11745 9170
rect 11783 9136 11817 9170
rect 11855 9136 11889 9170
rect 11927 9136 11961 9170
rect 11999 9136 12033 9170
rect 12071 9136 12105 9170
rect 12143 9136 12177 9170
rect 12215 9136 12249 9170
rect 12287 9136 12321 9170
rect 12359 9136 12393 9170
rect 12431 9136 12465 9170
rect 12503 9136 12537 9170
rect 12575 9136 12609 9170
rect 12647 9136 12681 9170
rect 12719 9136 12753 9170
rect 12791 9136 12825 9170
rect 12863 9136 12897 9170
rect 12935 9136 12969 9170
rect 13007 9136 13041 9170
rect 13079 9136 13113 9170
rect 13151 9136 13185 9170
rect 13223 9136 13257 9170
rect 13295 9136 13329 9170
rect 13367 9136 13401 9170
rect 13439 9136 13473 9170
rect 13511 9136 13545 9170
rect 13583 9136 13617 9170
rect 13655 9136 13689 9170
rect 13727 9136 13761 9170
rect 13799 9136 13833 9170
rect 248 8740 278 8753
rect 278 8740 282 8753
rect 322 8740 348 8753
rect 348 8740 356 8753
rect 396 8740 418 8753
rect 418 8740 430 8753
rect 470 8740 488 8753
rect 488 8740 504 8753
rect 544 8740 558 8753
rect 558 8740 578 8753
rect 618 8740 628 8753
rect 628 8740 652 8753
rect 691 8740 698 8753
rect 698 8740 725 8753
rect 764 8740 768 8753
rect 768 8740 798 8753
rect 837 8740 838 8753
rect 838 8740 871 8753
rect 912 8740 942 8760
rect 942 8740 946 8760
rect 984 8740 1012 8760
rect 1012 8740 1018 8760
rect 1056 8740 1082 8760
rect 1082 8740 1090 8760
rect 1128 8740 1152 8760
rect 1152 8740 1162 8760
rect 1200 8740 1222 8760
rect 1222 8740 1234 8760
rect 1272 8740 1292 8760
rect 1292 8740 1306 8760
rect 1344 8740 1362 8760
rect 1362 8740 1378 8760
rect 1416 8740 1432 8760
rect 1432 8740 1450 8760
rect 1488 8740 1501 8760
rect 1501 8740 1522 8760
rect 1560 8740 1570 8760
rect 1570 8740 1594 8760
rect 1632 8740 1639 8760
rect 1639 8740 1666 8760
rect 1704 8740 1708 8760
rect 1708 8740 1738 8760
rect 1776 8740 1777 8760
rect 1777 8740 1810 8760
rect 1849 8740 1881 8760
rect 1881 8740 1883 8760
rect 1922 8740 1950 8760
rect 1950 8740 1956 8760
rect 1995 8740 2019 8760
rect 2019 8740 2029 8760
rect 2068 8740 2088 8760
rect 2088 8740 2102 8760
rect 2141 8740 2157 8760
rect 2157 8740 2175 8760
rect 2227 8740 2260 8753
rect 2260 8740 2261 8753
rect 2306 8740 2329 8753
rect 2329 8740 2340 8753
rect 2385 8740 2398 8753
rect 2398 8740 2419 8753
rect 2464 8740 2467 8753
rect 2467 8740 2498 8753
rect 2543 8740 2571 8753
rect 2571 8740 2577 8753
rect 2621 8740 2640 8753
rect 2640 8740 2655 8753
rect 2699 8740 2709 8753
rect 2709 8740 2733 8753
rect 2777 8740 2778 8753
rect 2778 8740 2811 8753
rect 2855 8740 2881 8753
rect 2881 8740 2889 8753
rect 248 8719 282 8740
rect 322 8719 356 8740
rect 396 8719 430 8740
rect 470 8719 504 8740
rect 544 8719 578 8740
rect 618 8719 652 8740
rect 691 8719 725 8740
rect 764 8719 798 8740
rect 837 8719 871 8740
rect 912 8726 946 8740
rect 984 8726 1018 8740
rect 1056 8726 1090 8740
rect 1128 8726 1162 8740
rect 1200 8726 1234 8740
rect 1272 8726 1306 8740
rect 1344 8726 1378 8740
rect 1416 8726 1450 8740
rect 1488 8726 1522 8740
rect 1560 8726 1594 8740
rect 1632 8726 1666 8740
rect 1704 8726 1738 8740
rect 1776 8726 1810 8740
rect 1849 8726 1883 8740
rect 1922 8726 1956 8740
rect 1995 8726 2029 8740
rect 2068 8726 2102 8740
rect 2141 8726 2175 8740
rect 2227 8719 2261 8740
rect 2306 8719 2340 8740
rect 2385 8719 2419 8740
rect 2464 8719 2498 8740
rect 2543 8719 2577 8740
rect 2621 8719 2655 8740
rect 2699 8719 2733 8740
rect 2777 8719 2811 8740
rect 2855 8719 2889 8740
rect 2933 8736 2967 8753
rect 3011 8736 3036 8753
rect 3036 8736 3045 8753
rect 3477 8736 3479 8760
rect 3479 8736 3511 8760
rect 3550 8736 3581 8760
rect 3581 8736 3584 8760
rect 3623 8736 3649 8760
rect 3649 8736 3657 8760
rect 3696 8736 3717 8760
rect 3717 8736 3730 8760
rect 3769 8736 3785 8760
rect 3785 8736 3803 8760
rect 3842 8736 3853 8760
rect 3853 8736 3876 8760
rect 3915 8736 3921 8760
rect 3921 8736 3949 8760
rect 3988 8736 3989 8760
rect 3989 8736 4022 8760
rect 4061 8736 4091 8760
rect 4091 8736 4095 8760
rect 4134 8736 4159 8760
rect 4159 8736 4168 8760
rect 4207 8736 4227 8760
rect 4227 8736 4241 8760
rect 4280 8736 4295 8760
rect 4295 8736 4314 8760
rect 4353 8736 4363 8760
rect 4363 8736 4387 8760
rect 4426 8736 4431 8760
rect 4431 8736 4460 8760
rect 4499 8736 4533 8760
rect 4572 8736 4601 8760
rect 4601 8736 4606 8760
rect 4645 8736 4669 8760
rect 4669 8736 4679 8760
rect 4718 8736 4737 8760
rect 4737 8736 4752 8760
rect 4791 8736 4805 8760
rect 4805 8736 4825 8760
rect 4864 8736 4873 8760
rect 4873 8736 4898 8760
rect 4937 8736 4941 8760
rect 4941 8736 4971 8760
rect 5010 8736 5043 8760
rect 5043 8736 5044 8760
rect 5083 8736 5111 8760
rect 5111 8736 5117 8760
rect 5156 8736 5179 8760
rect 5179 8736 5190 8760
rect 5229 8736 5247 8760
rect 5247 8736 5263 8760
rect 5302 8736 5315 8760
rect 5315 8736 5336 8760
rect 5375 8736 5383 8760
rect 5383 8736 5409 8760
rect 5448 8736 5451 8760
rect 5451 8736 5482 8760
rect 5521 8736 5553 8760
rect 5553 8736 5555 8760
rect 5594 8736 5621 8760
rect 5621 8736 5628 8760
rect 5667 8736 5689 8760
rect 5689 8736 5701 8760
rect 5740 8736 5757 8760
rect 5757 8736 5774 8760
rect 5813 8736 5825 8760
rect 5825 8736 5847 8760
rect 5886 8736 5893 8760
rect 5893 8736 5920 8760
rect 5959 8736 5961 8760
rect 5961 8736 5993 8760
rect 6032 8736 6063 8760
rect 6063 8736 6066 8760
rect 6105 8736 6131 8760
rect 6131 8736 6139 8760
rect 6178 8736 6199 8760
rect 6199 8736 6212 8760
rect 6251 8736 6267 8760
rect 6267 8736 6285 8760
rect 6324 8736 6335 8760
rect 6335 8736 6358 8760
rect 6397 8736 6403 8760
rect 6403 8736 6431 8760
rect 6470 8736 6471 8760
rect 6471 8736 6504 8760
rect 6543 8736 6573 8760
rect 6573 8736 6577 8760
rect 6616 8736 6641 8760
rect 6641 8736 6650 8760
rect 6689 8736 6709 8760
rect 6709 8736 6723 8760
rect 6762 8736 6777 8760
rect 6777 8736 6796 8760
rect 6835 8736 6845 8760
rect 6845 8736 6869 8760
rect 6908 8736 6913 8760
rect 6913 8736 6942 8760
rect 2933 8719 2967 8736
rect 3011 8719 3045 8736
rect 3477 8726 3511 8736
rect 3550 8726 3584 8736
rect 3623 8726 3657 8736
rect 3696 8726 3730 8736
rect 3769 8726 3803 8736
rect 3842 8726 3876 8736
rect 3915 8726 3949 8736
rect 3988 8726 4022 8736
rect 4061 8726 4095 8736
rect 4134 8726 4168 8736
rect 4207 8726 4241 8736
rect 4280 8726 4314 8736
rect 4353 8726 4387 8736
rect 4426 8726 4460 8736
rect 4499 8726 4533 8736
rect 4572 8726 4606 8736
rect 4645 8726 4679 8736
rect 4718 8726 4752 8736
rect 4791 8726 4825 8736
rect 4864 8726 4898 8736
rect 4937 8726 4971 8736
rect 5010 8726 5044 8736
rect 5083 8726 5117 8736
rect 5156 8726 5190 8736
rect 5229 8726 5263 8736
rect 5302 8726 5336 8736
rect 5375 8726 5409 8736
rect 5448 8726 5482 8736
rect 5521 8726 5555 8736
rect 5594 8726 5628 8736
rect 5667 8726 5701 8736
rect 5740 8726 5774 8736
rect 5813 8726 5847 8736
rect 5886 8726 5920 8736
rect 5959 8726 5993 8736
rect 6032 8726 6066 8736
rect 6105 8726 6139 8736
rect 6178 8726 6212 8736
rect 6251 8726 6285 8736
rect 6324 8726 6358 8736
rect 6397 8726 6431 8736
rect 6470 8726 6504 8736
rect 6543 8726 6577 8736
rect 6616 8726 6650 8736
rect 6689 8726 6723 8736
rect 6762 8726 6796 8736
rect 6835 8726 6869 8736
rect 6908 8726 6942 8736
rect 6981 8726 7015 8760
rect 7054 8736 7083 8760
rect 7083 8736 7088 8760
rect 7127 8736 7151 8760
rect 7151 8736 7161 8760
rect 7200 8736 7219 8760
rect 7219 8736 7234 8760
rect 7273 8736 7287 8760
rect 7287 8736 7307 8760
rect 7346 8736 7355 8760
rect 7355 8736 7380 8760
rect 7419 8736 7423 8760
rect 7423 8736 7453 8760
rect 7492 8736 7525 8760
rect 7525 8736 7526 8760
rect 7565 8736 7593 8760
rect 7593 8736 7599 8760
rect 7638 8736 7661 8760
rect 7661 8736 7672 8760
rect 7711 8736 7729 8760
rect 7729 8736 7745 8760
rect 7784 8736 7797 8760
rect 7797 8736 7818 8760
rect 7857 8736 7865 8760
rect 7865 8736 7891 8760
rect 7930 8736 7933 8760
rect 7933 8736 7964 8760
rect 8003 8736 8035 8760
rect 8035 8736 8037 8760
rect 8075 8736 8103 8760
rect 8103 8736 8109 8760
rect 8147 8736 8171 8760
rect 8171 8736 8181 8760
rect 8219 8736 8239 8760
rect 8239 8736 8253 8760
rect 8291 8736 8307 8760
rect 8307 8736 8325 8760
rect 8363 8739 8393 8760
rect 8393 8739 8397 8760
rect 8435 8739 8462 8760
rect 8462 8739 8469 8760
rect 8507 8739 8531 8760
rect 8531 8739 8541 8760
rect 8579 8739 8600 8760
rect 8600 8739 8613 8760
rect 8651 8739 8669 8760
rect 8669 8739 8685 8760
rect 8723 8739 8738 8760
rect 8738 8739 8757 8760
rect 8795 8739 8807 8760
rect 8807 8739 8829 8760
rect 8867 8739 8876 8760
rect 8876 8739 8901 8760
rect 8939 8739 8945 8760
rect 8945 8739 8973 8760
rect 9011 8739 9014 8760
rect 9014 8739 9045 8760
rect 9083 8739 9117 8760
rect 9155 8739 9186 8760
rect 9186 8739 9189 8760
rect 9227 8739 9254 8760
rect 9254 8739 9261 8760
rect 9299 8739 9322 8760
rect 9322 8739 9333 8760
rect 9371 8739 9390 8760
rect 9390 8739 9405 8760
rect 9443 8739 9458 8760
rect 9458 8739 9477 8760
rect 9515 8739 9526 8760
rect 9526 8739 9549 8760
rect 9587 8739 9594 8760
rect 9594 8739 9621 8760
rect 9659 8739 9662 8760
rect 9662 8739 9693 8760
rect 9731 8739 9764 8760
rect 9764 8739 9765 8760
rect 9803 8739 9832 8760
rect 9832 8739 9837 8760
rect 9875 8739 9900 8760
rect 9900 8739 9909 8760
rect 9947 8739 9968 8760
rect 9968 8739 9981 8760
rect 10019 8739 10036 8760
rect 10036 8739 10053 8760
rect 10091 8739 10104 8760
rect 10104 8739 10125 8760
rect 10163 8739 10172 8760
rect 10172 8739 10197 8760
rect 10235 8739 10240 8760
rect 10240 8739 10269 8760
rect 10307 8739 10308 8760
rect 10308 8739 10341 8760
rect 10379 8739 10410 8760
rect 10410 8739 10413 8760
rect 10451 8739 10478 8760
rect 10478 8739 10485 8760
rect 10523 8739 10546 8760
rect 10546 8739 10557 8760
rect 10595 8739 10614 8760
rect 10614 8739 10629 8760
rect 10667 8739 10682 8760
rect 10682 8739 10701 8760
rect 10739 8739 10750 8760
rect 10750 8739 10773 8760
rect 10811 8739 10818 8760
rect 10818 8739 10845 8760
rect 10883 8739 10886 8760
rect 10886 8739 10917 8760
rect 10955 8739 10988 8760
rect 10988 8739 10989 8760
rect 11027 8739 11056 8760
rect 11056 8739 11061 8760
rect 11099 8739 11124 8760
rect 11124 8739 11133 8760
rect 11171 8739 11192 8760
rect 11192 8739 11205 8760
rect 11243 8739 11260 8760
rect 11260 8739 11277 8760
rect 11315 8739 11328 8760
rect 11328 8739 11349 8760
rect 11387 8739 11396 8760
rect 11396 8739 11421 8760
rect 11459 8739 11464 8760
rect 11464 8739 11493 8760
rect 11531 8739 11532 8760
rect 11532 8739 11565 8760
rect 11603 8739 11634 8760
rect 11634 8739 11637 8760
rect 11675 8739 11702 8760
rect 11702 8739 11709 8760
rect 11747 8739 11770 8760
rect 11770 8739 11781 8760
rect 11819 8739 11838 8760
rect 11838 8739 11853 8760
rect 11891 8739 11906 8760
rect 11906 8739 11925 8760
rect 11963 8739 11974 8760
rect 11974 8739 11997 8760
rect 12035 8739 12042 8760
rect 12042 8739 12069 8760
rect 12107 8739 12110 8760
rect 12110 8739 12141 8760
rect 12179 8739 12212 8760
rect 12212 8739 12213 8760
rect 12251 8739 12280 8760
rect 12280 8739 12285 8760
rect 12323 8739 12348 8760
rect 12348 8739 12357 8760
rect 12395 8739 12416 8760
rect 12416 8739 12429 8760
rect 12467 8739 12484 8760
rect 12484 8739 12501 8760
rect 12539 8739 12552 8760
rect 12552 8739 12573 8760
rect 12611 8739 12620 8760
rect 12620 8739 12645 8760
rect 12683 8739 12688 8760
rect 12688 8739 12717 8760
rect 12755 8739 12756 8760
rect 12756 8739 12789 8760
rect 12827 8739 12858 8760
rect 12858 8739 12861 8760
rect 12899 8739 12926 8760
rect 12926 8739 12933 8760
rect 12971 8739 12994 8760
rect 12994 8739 13005 8760
rect 13043 8739 13062 8760
rect 13062 8739 13077 8760
rect 13115 8739 13130 8760
rect 13130 8739 13149 8760
rect 13187 8739 13198 8760
rect 13198 8739 13221 8760
rect 13259 8739 13266 8760
rect 13266 8739 13293 8760
rect 13331 8739 13334 8760
rect 13334 8739 13365 8760
rect 13403 8739 13436 8760
rect 13436 8739 13437 8760
rect 13475 8739 13504 8760
rect 13504 8739 13509 8760
rect 13547 8739 13572 8760
rect 13572 8739 13581 8760
rect 13619 8739 13640 8760
rect 13640 8739 13653 8760
rect 13691 8739 13708 8760
rect 13708 8739 13725 8760
rect 13763 8739 13776 8760
rect 13776 8739 13797 8760
rect 13835 8739 13844 8760
rect 13844 8739 13869 8760
rect 13907 8739 13912 8760
rect 13912 8739 13941 8760
rect 13979 8739 13980 8760
rect 13980 8739 14013 8760
rect 14051 8739 14082 8760
rect 14082 8739 14085 8760
rect 14123 8739 14150 8760
rect 14150 8739 14157 8760
rect 14195 8739 14218 8760
rect 14218 8739 14229 8760
rect 14267 8739 14286 8760
rect 14286 8739 14301 8760
rect 14339 8739 14354 8760
rect 14354 8739 14373 8760
rect 14411 8739 14422 8760
rect 14422 8739 14445 8760
rect 14483 8739 14490 8760
rect 14490 8739 14517 8760
rect 14555 8739 14558 8760
rect 14558 8739 14589 8760
rect 14627 8739 14660 8760
rect 14660 8739 14661 8760
rect 14699 8739 14728 8760
rect 14728 8739 14733 8760
rect 14771 8739 14796 8760
rect 14796 8739 14805 8760
rect 14843 8739 14864 8760
rect 14864 8739 14877 8760
rect 7054 8726 7088 8736
rect 7127 8726 7161 8736
rect 7200 8726 7234 8736
rect 7273 8726 7307 8736
rect 7346 8726 7380 8736
rect 7419 8726 7453 8736
rect 7492 8726 7526 8736
rect 7565 8726 7599 8736
rect 7638 8726 7672 8736
rect 7711 8726 7745 8736
rect 7784 8726 7818 8736
rect 7857 8726 7891 8736
rect 7930 8726 7964 8736
rect 8003 8726 8037 8736
rect 8075 8726 8109 8736
rect 8147 8726 8181 8736
rect 8219 8726 8253 8736
rect 8291 8726 8325 8736
rect 8363 8726 8397 8739
rect 8435 8726 8469 8739
rect 8507 8726 8541 8739
rect 8579 8726 8613 8739
rect 8651 8726 8685 8739
rect 8723 8726 8757 8739
rect 8795 8726 8829 8739
rect 8867 8726 8901 8739
rect 8939 8726 8973 8739
rect 9011 8726 9045 8739
rect 9083 8726 9117 8739
rect 9155 8726 9189 8739
rect 9227 8726 9261 8739
rect 9299 8726 9333 8739
rect 9371 8726 9405 8739
rect 9443 8726 9477 8739
rect 9515 8726 9549 8739
rect 9587 8726 9621 8739
rect 9659 8726 9693 8739
rect 9731 8726 9765 8739
rect 9803 8726 9837 8739
rect 9875 8726 9909 8739
rect 9947 8726 9981 8739
rect 10019 8726 10053 8739
rect 10091 8726 10125 8739
rect 10163 8726 10197 8739
rect 10235 8726 10269 8739
rect 10307 8726 10341 8739
rect 10379 8726 10413 8739
rect 10451 8726 10485 8739
rect 10523 8726 10557 8739
rect 10595 8726 10629 8739
rect 10667 8726 10701 8739
rect 10739 8726 10773 8739
rect 10811 8726 10845 8739
rect 10883 8726 10917 8739
rect 10955 8726 10989 8739
rect 11027 8726 11061 8739
rect 11099 8726 11133 8739
rect 11171 8726 11205 8739
rect 11243 8726 11277 8739
rect 11315 8726 11349 8739
rect 11387 8726 11421 8739
rect 11459 8726 11493 8739
rect 11531 8726 11565 8739
rect 11603 8726 11637 8739
rect 11675 8726 11709 8739
rect 11747 8726 11781 8739
rect 11819 8726 11853 8739
rect 11891 8726 11925 8739
rect 11963 8726 11997 8739
rect 12035 8726 12069 8739
rect 12107 8726 12141 8739
rect 12179 8726 12213 8739
rect 12251 8726 12285 8739
rect 12323 8726 12357 8739
rect 12395 8726 12429 8739
rect 12467 8726 12501 8739
rect 12539 8726 12573 8739
rect 12611 8726 12645 8739
rect 12683 8726 12717 8739
rect 12755 8726 12789 8739
rect 12827 8726 12861 8739
rect 12899 8726 12933 8739
rect 12971 8726 13005 8739
rect 13043 8726 13077 8739
rect 13115 8726 13149 8739
rect 13187 8726 13221 8739
rect 13259 8726 13293 8739
rect 13331 8726 13365 8739
rect 13403 8726 13437 8739
rect 13475 8726 13509 8739
rect 13547 8726 13581 8739
rect 13619 8726 13653 8739
rect 13691 8726 13725 8739
rect 13763 8726 13797 8739
rect 13835 8726 13869 8739
rect 13907 8726 13941 8739
rect 13979 8726 14013 8739
rect 14051 8726 14085 8739
rect 14123 8726 14157 8739
rect 14195 8726 14229 8739
rect 14267 8726 14301 8739
rect 14339 8726 14373 8739
rect 14411 8726 14445 8739
rect 14483 8726 14517 8739
rect 14555 8726 14589 8739
rect 14627 8726 14661 8739
rect 14699 8726 14733 8739
rect 14771 8726 14805 8739
rect 14843 8726 14877 8739
rect 912 8626 946 8636
rect 984 8626 1018 8636
rect 1056 8626 1090 8636
rect 1128 8626 1162 8636
rect 1200 8626 1234 8636
rect 1272 8626 1306 8636
rect 1344 8626 1378 8636
rect 1416 8626 1450 8636
rect 1488 8626 1522 8636
rect 1560 8626 1594 8636
rect 1632 8626 1666 8636
rect 1704 8626 1738 8636
rect 1776 8626 1810 8636
rect 1849 8626 1883 8636
rect 1922 8626 1956 8636
rect 1995 8626 2029 8636
rect 2068 8626 2102 8636
rect 2141 8626 2175 8636
rect 3477 8630 3511 8636
rect 3550 8630 3584 8636
rect 3623 8630 3657 8636
rect 3696 8630 3730 8636
rect 3769 8630 3803 8636
rect 3842 8630 3876 8636
rect 3915 8630 3949 8636
rect 3988 8630 4022 8636
rect 4061 8630 4095 8636
rect 4134 8630 4168 8636
rect 4207 8630 4241 8636
rect 4280 8630 4314 8636
rect 4353 8630 4387 8636
rect 4426 8630 4460 8636
rect 4499 8630 4533 8636
rect 4572 8630 4606 8636
rect 4645 8630 4679 8636
rect 4718 8630 4752 8636
rect 4791 8630 4825 8636
rect 4864 8630 4898 8636
rect 4937 8630 4971 8636
rect 5010 8630 5044 8636
rect 5083 8630 5117 8636
rect 5156 8630 5190 8636
rect 5229 8630 5263 8636
rect 5302 8630 5336 8636
rect 5375 8630 5409 8636
rect 5448 8630 5482 8636
rect 5521 8630 5555 8636
rect 5594 8630 5628 8636
rect 5667 8630 5701 8636
rect 5740 8630 5774 8636
rect 5813 8630 5847 8636
rect 5886 8630 5920 8636
rect 5959 8630 5993 8636
rect 6032 8630 6066 8636
rect 6105 8630 6139 8636
rect 6178 8630 6212 8636
rect 6251 8630 6285 8636
rect 6324 8630 6358 8636
rect 6397 8630 6431 8636
rect 6470 8630 6504 8636
rect 6543 8630 6577 8636
rect 6616 8630 6650 8636
rect 6689 8630 6723 8636
rect 6762 8630 6796 8636
rect 6835 8630 6869 8636
rect 6908 8630 6942 8636
rect 912 8602 942 8626
rect 942 8602 946 8626
rect 984 8602 1012 8626
rect 1012 8602 1018 8626
rect 1056 8602 1082 8626
rect 1082 8602 1090 8626
rect 1128 8602 1152 8626
rect 1152 8602 1162 8626
rect 1200 8602 1222 8626
rect 1222 8602 1234 8626
rect 1272 8602 1292 8626
rect 1292 8602 1306 8626
rect 1344 8602 1362 8626
rect 1362 8602 1378 8626
rect 1416 8602 1432 8626
rect 1432 8602 1450 8626
rect 1488 8602 1501 8626
rect 1501 8602 1522 8626
rect 1560 8602 1570 8626
rect 1570 8602 1594 8626
rect 1632 8602 1639 8626
rect 1639 8602 1666 8626
rect 1704 8602 1708 8626
rect 1708 8602 1738 8626
rect 1776 8602 1777 8626
rect 1777 8602 1810 8626
rect 1849 8602 1881 8626
rect 1881 8602 1883 8626
rect 1922 8602 1950 8626
rect 1950 8602 1956 8626
rect 1995 8602 2019 8626
rect 2019 8602 2029 8626
rect 2068 8602 2088 8626
rect 2088 8602 2102 8626
rect 2141 8602 2157 8626
rect 2157 8602 2175 8626
rect 3477 8602 3479 8630
rect 3479 8602 3511 8630
rect 3550 8602 3581 8630
rect 3581 8602 3584 8630
rect 3623 8602 3649 8630
rect 3649 8602 3657 8630
rect 3696 8602 3717 8630
rect 3717 8602 3730 8630
rect 3769 8602 3785 8630
rect 3785 8602 3803 8630
rect 3842 8602 3853 8630
rect 3853 8602 3876 8630
rect 3915 8602 3921 8630
rect 3921 8602 3949 8630
rect 3988 8602 3989 8630
rect 3989 8602 4022 8630
rect 4061 8602 4091 8630
rect 4091 8602 4095 8630
rect 4134 8602 4159 8630
rect 4159 8602 4168 8630
rect 4207 8602 4227 8630
rect 4227 8602 4241 8630
rect 4280 8602 4295 8630
rect 4295 8602 4314 8630
rect 4353 8602 4363 8630
rect 4363 8602 4387 8630
rect 4426 8602 4431 8630
rect 4431 8602 4460 8630
rect 4499 8602 4533 8630
rect 4572 8602 4601 8630
rect 4601 8602 4606 8630
rect 4645 8602 4669 8630
rect 4669 8602 4679 8630
rect 4718 8602 4737 8630
rect 4737 8602 4752 8630
rect 4791 8602 4805 8630
rect 4805 8602 4825 8630
rect 4864 8602 4873 8630
rect 4873 8602 4898 8630
rect 4937 8602 4941 8630
rect 4941 8602 4971 8630
rect 5010 8602 5043 8630
rect 5043 8602 5044 8630
rect 5083 8602 5111 8630
rect 5111 8602 5117 8630
rect 5156 8602 5179 8630
rect 5179 8602 5190 8630
rect 5229 8602 5247 8630
rect 5247 8602 5263 8630
rect 5302 8602 5315 8630
rect 5315 8602 5336 8630
rect 5375 8602 5383 8630
rect 5383 8602 5409 8630
rect 5448 8602 5451 8630
rect 5451 8602 5482 8630
rect 5521 8602 5553 8630
rect 5553 8602 5555 8630
rect 5594 8602 5621 8630
rect 5621 8602 5628 8630
rect 5667 8602 5689 8630
rect 5689 8602 5701 8630
rect 5740 8602 5757 8630
rect 5757 8602 5774 8630
rect 5813 8602 5825 8630
rect 5825 8602 5847 8630
rect 5886 8602 5893 8630
rect 5893 8602 5920 8630
rect 5959 8602 5961 8630
rect 5961 8602 5993 8630
rect 6032 8602 6063 8630
rect 6063 8602 6066 8630
rect 6105 8602 6131 8630
rect 6131 8602 6139 8630
rect 6178 8602 6199 8630
rect 6199 8602 6212 8630
rect 6251 8602 6267 8630
rect 6267 8602 6285 8630
rect 6324 8602 6335 8630
rect 6335 8602 6358 8630
rect 6397 8602 6403 8630
rect 6403 8602 6431 8630
rect 6470 8602 6471 8630
rect 6471 8602 6504 8630
rect 6543 8602 6573 8630
rect 6573 8602 6577 8630
rect 6616 8602 6641 8630
rect 6641 8602 6650 8630
rect 6689 8602 6709 8630
rect 6709 8602 6723 8630
rect 6762 8602 6777 8630
rect 6777 8602 6796 8630
rect 6835 8602 6845 8630
rect 6845 8602 6869 8630
rect 6908 8602 6913 8630
rect 6913 8602 6942 8630
rect 6981 8602 7015 8636
rect 7054 8630 7088 8636
rect 7127 8630 7161 8636
rect 7200 8630 7234 8636
rect 7273 8630 7307 8636
rect 7346 8630 7380 8636
rect 7419 8630 7453 8636
rect 7492 8630 7526 8636
rect 7565 8630 7599 8636
rect 7638 8630 7672 8636
rect 7711 8630 7745 8636
rect 7784 8630 7818 8636
rect 7857 8630 7891 8636
rect 7930 8630 7964 8636
rect 8003 8630 8037 8636
rect 8075 8630 8109 8636
rect 8147 8630 8181 8636
rect 8219 8630 8253 8636
rect 8291 8630 8325 8636
rect 7054 8602 7083 8630
rect 7083 8602 7088 8630
rect 7127 8602 7151 8630
rect 7151 8602 7161 8630
rect 7200 8602 7219 8630
rect 7219 8602 7234 8630
rect 7273 8602 7287 8630
rect 7287 8602 7307 8630
rect 7346 8602 7355 8630
rect 7355 8602 7380 8630
rect 7419 8602 7423 8630
rect 7423 8602 7453 8630
rect 7492 8602 7525 8630
rect 7525 8602 7526 8630
rect 7565 8602 7593 8630
rect 7593 8602 7599 8630
rect 7638 8602 7661 8630
rect 7661 8602 7672 8630
rect 7711 8602 7729 8630
rect 7729 8602 7745 8630
rect 7784 8602 7797 8630
rect 7797 8602 7818 8630
rect 7857 8602 7865 8630
rect 7865 8602 7891 8630
rect 7930 8602 7933 8630
rect 7933 8602 7964 8630
rect 8003 8602 8035 8630
rect 8035 8602 8037 8630
rect 8075 8602 8103 8630
rect 8103 8602 8109 8630
rect 8147 8602 8171 8630
rect 8171 8602 8181 8630
rect 8219 8602 8239 8630
rect 8239 8602 8253 8630
rect 8291 8602 8307 8630
rect 8307 8602 8325 8630
rect 8363 8613 8397 8636
rect 8435 8613 8469 8636
rect 8507 8613 8541 8636
rect 8579 8613 8613 8636
rect 8651 8613 8685 8636
rect 8723 8613 8757 8636
rect 8795 8613 8829 8636
rect 8867 8613 8901 8636
rect 8939 8613 8973 8636
rect 9011 8613 9045 8636
rect 9083 8613 9117 8636
rect 9155 8613 9189 8636
rect 9227 8613 9261 8636
rect 9299 8613 9333 8636
rect 9371 8613 9405 8636
rect 9443 8613 9477 8636
rect 9515 8613 9549 8636
rect 9587 8613 9621 8636
rect 9659 8613 9693 8636
rect 9731 8613 9765 8636
rect 9803 8613 9837 8636
rect 9875 8613 9909 8636
rect 9947 8613 9981 8636
rect 10019 8613 10053 8636
rect 10091 8613 10125 8636
rect 10163 8613 10197 8636
rect 10235 8613 10269 8636
rect 10307 8613 10341 8636
rect 10379 8613 10413 8636
rect 10451 8613 10485 8636
rect 10523 8613 10557 8636
rect 10595 8613 10629 8636
rect 10667 8613 10701 8636
rect 10739 8613 10773 8636
rect 10811 8613 10845 8636
rect 10883 8613 10917 8636
rect 10955 8613 10989 8636
rect 11027 8613 11061 8636
rect 11099 8613 11133 8636
rect 11171 8613 11205 8636
rect 11243 8613 11277 8636
rect 11315 8613 11349 8636
rect 11387 8613 11421 8636
rect 11459 8613 11493 8636
rect 11531 8613 11565 8636
rect 11603 8613 11637 8636
rect 11675 8613 11709 8636
rect 11747 8613 11781 8636
rect 11819 8613 11853 8636
rect 11891 8613 11925 8636
rect 11963 8613 11997 8636
rect 12035 8613 12069 8636
rect 12107 8613 12141 8636
rect 12179 8613 12213 8636
rect 12251 8613 12285 8636
rect 12323 8613 12357 8636
rect 12395 8613 12429 8636
rect 12467 8613 12501 8636
rect 12539 8613 12573 8636
rect 12611 8613 12645 8636
rect 12683 8613 12717 8636
rect 12755 8613 12789 8636
rect 12827 8613 12861 8636
rect 12899 8613 12933 8636
rect 12971 8613 13005 8636
rect 13043 8613 13077 8636
rect 13115 8613 13149 8636
rect 13187 8613 13221 8636
rect 13259 8613 13293 8636
rect 13331 8613 13365 8636
rect 13403 8613 13437 8636
rect 13475 8613 13509 8636
rect 13547 8613 13581 8636
rect 13619 8613 13653 8636
rect 13691 8613 13725 8636
rect 13763 8613 13797 8636
rect 13835 8613 13869 8636
rect 13907 8613 13941 8636
rect 13979 8613 14013 8636
rect 14051 8613 14085 8636
rect 14123 8613 14157 8636
rect 14195 8613 14229 8636
rect 14267 8613 14301 8636
rect 14339 8613 14373 8636
rect 14411 8613 14445 8636
rect 14483 8613 14517 8636
rect 14555 8613 14589 8636
rect 14627 8613 14661 8636
rect 14699 8613 14733 8636
rect 14771 8613 14805 8636
rect 14843 8613 14877 8636
rect 8363 8602 8393 8613
rect 8393 8602 8397 8613
rect 8435 8602 8462 8613
rect 8462 8602 8469 8613
rect 8507 8602 8531 8613
rect 8531 8602 8541 8613
rect 8579 8602 8600 8613
rect 8600 8602 8613 8613
rect 8651 8602 8669 8613
rect 8669 8602 8685 8613
rect 8723 8602 8738 8613
rect 8738 8602 8757 8613
rect 8795 8602 8807 8613
rect 8807 8602 8829 8613
rect 8867 8602 8876 8613
rect 8876 8602 8901 8613
rect 8939 8602 8945 8613
rect 8945 8602 8973 8613
rect 9011 8602 9014 8613
rect 9014 8602 9045 8613
rect 9083 8602 9117 8613
rect 9155 8602 9186 8613
rect 9186 8602 9189 8613
rect 9227 8602 9254 8613
rect 9254 8602 9261 8613
rect 9299 8602 9322 8613
rect 9322 8602 9333 8613
rect 9371 8602 9390 8613
rect 9390 8602 9405 8613
rect 9443 8602 9458 8613
rect 9458 8602 9477 8613
rect 9515 8602 9526 8613
rect 9526 8602 9549 8613
rect 9587 8602 9594 8613
rect 9594 8602 9621 8613
rect 9659 8602 9662 8613
rect 9662 8602 9693 8613
rect 9731 8602 9764 8613
rect 9764 8602 9765 8613
rect 9803 8602 9832 8613
rect 9832 8602 9837 8613
rect 9875 8602 9900 8613
rect 9900 8602 9909 8613
rect 9947 8602 9968 8613
rect 9968 8602 9981 8613
rect 10019 8602 10036 8613
rect 10036 8602 10053 8613
rect 10091 8602 10104 8613
rect 10104 8602 10125 8613
rect 10163 8602 10172 8613
rect 10172 8602 10197 8613
rect 10235 8602 10240 8613
rect 10240 8602 10269 8613
rect 10307 8602 10308 8613
rect 10308 8602 10341 8613
rect 10379 8602 10410 8613
rect 10410 8602 10413 8613
rect 10451 8602 10478 8613
rect 10478 8602 10485 8613
rect 10523 8602 10546 8613
rect 10546 8602 10557 8613
rect 10595 8602 10614 8613
rect 10614 8602 10629 8613
rect 10667 8602 10682 8613
rect 10682 8602 10701 8613
rect 10739 8602 10750 8613
rect 10750 8602 10773 8613
rect 10811 8602 10818 8613
rect 10818 8602 10845 8613
rect 10883 8602 10886 8613
rect 10886 8602 10917 8613
rect 10955 8602 10988 8613
rect 10988 8602 10989 8613
rect 11027 8602 11056 8613
rect 11056 8602 11061 8613
rect 11099 8602 11124 8613
rect 11124 8602 11133 8613
rect 11171 8602 11192 8613
rect 11192 8602 11205 8613
rect 11243 8602 11260 8613
rect 11260 8602 11277 8613
rect 11315 8602 11328 8613
rect 11328 8602 11349 8613
rect 11387 8602 11396 8613
rect 11396 8602 11421 8613
rect 11459 8602 11464 8613
rect 11464 8602 11493 8613
rect 11531 8602 11532 8613
rect 11532 8602 11565 8613
rect 11603 8602 11634 8613
rect 11634 8602 11637 8613
rect 11675 8602 11702 8613
rect 11702 8602 11709 8613
rect 11747 8602 11770 8613
rect 11770 8602 11781 8613
rect 11819 8602 11838 8613
rect 11838 8602 11853 8613
rect 11891 8602 11906 8613
rect 11906 8602 11925 8613
rect 11963 8602 11974 8613
rect 11974 8602 11997 8613
rect 12035 8602 12042 8613
rect 12042 8602 12069 8613
rect 12107 8602 12110 8613
rect 12110 8602 12141 8613
rect 12179 8602 12212 8613
rect 12212 8602 12213 8613
rect 12251 8602 12280 8613
rect 12280 8602 12285 8613
rect 12323 8602 12348 8613
rect 12348 8602 12357 8613
rect 12395 8602 12416 8613
rect 12416 8602 12429 8613
rect 12467 8602 12484 8613
rect 12484 8602 12501 8613
rect 12539 8602 12552 8613
rect 12552 8602 12573 8613
rect 12611 8602 12620 8613
rect 12620 8602 12645 8613
rect 12683 8602 12688 8613
rect 12688 8602 12717 8613
rect 12755 8602 12756 8613
rect 12756 8602 12789 8613
rect 12827 8602 12858 8613
rect 12858 8602 12861 8613
rect 12899 8602 12926 8613
rect 12926 8602 12933 8613
rect 12971 8602 12994 8613
rect 12994 8602 13005 8613
rect 13043 8602 13062 8613
rect 13062 8602 13077 8613
rect 13115 8602 13130 8613
rect 13130 8602 13149 8613
rect 13187 8602 13198 8613
rect 13198 8602 13221 8613
rect 13259 8602 13266 8613
rect 13266 8602 13293 8613
rect 13331 8602 13334 8613
rect 13334 8602 13365 8613
rect 13403 8602 13436 8613
rect 13436 8602 13437 8613
rect 13475 8602 13504 8613
rect 13504 8602 13509 8613
rect 13547 8602 13572 8613
rect 13572 8602 13581 8613
rect 13619 8602 13640 8613
rect 13640 8602 13653 8613
rect 13691 8602 13708 8613
rect 13708 8602 13725 8613
rect 13763 8602 13776 8613
rect 13776 8602 13797 8613
rect 13835 8602 13844 8613
rect 13844 8602 13869 8613
rect 13907 8602 13912 8613
rect 13912 8602 13941 8613
rect 13979 8602 13980 8613
rect 13980 8602 14013 8613
rect 14051 8602 14082 8613
rect 14082 8602 14085 8613
rect 14123 8602 14150 8613
rect 14150 8602 14157 8613
rect 14195 8602 14218 8613
rect 14218 8602 14229 8613
rect 14267 8602 14286 8613
rect 14286 8602 14301 8613
rect 14339 8602 14354 8613
rect 14354 8602 14373 8613
rect 14411 8602 14422 8613
rect 14422 8602 14445 8613
rect 14483 8602 14490 8613
rect 14490 8602 14517 8613
rect 14555 8602 14558 8613
rect 14558 8602 14589 8613
rect 14627 8602 14660 8613
rect 14660 8602 14661 8613
rect 14699 8602 14728 8613
rect 14728 8602 14733 8613
rect 14771 8602 14796 8613
rect 14796 8602 14805 8613
rect 14843 8602 14864 8613
rect 14864 8602 14877 8613
rect 13992 8533 14026 8546
rect 14076 8533 14110 8546
rect 13992 8512 14014 8533
rect 14014 8512 14026 8533
rect 14076 8512 14082 8533
rect 14082 8512 14110 8533
rect 14185 8499 14218 8512
rect 14218 8499 14219 8512
rect 14257 8499 14286 8512
rect 14286 8499 14291 8512
rect 14329 8499 14354 8512
rect 14354 8499 14363 8512
rect 14401 8499 14422 8512
rect 14422 8499 14435 8512
rect 14473 8499 14490 8512
rect 14490 8499 14507 8512
rect 14185 8478 14219 8499
rect 14257 8478 14291 8499
rect 14329 8478 14363 8499
rect 14401 8478 14435 8499
rect 14473 8478 14507 8499
rect 13992 8453 14026 8474
rect 14076 8453 14110 8474
rect 14614 8453 14648 8462
rect 14692 8453 14726 8462
rect 14770 8453 14804 8462
rect 14848 8453 14882 8462
rect 13992 8440 14014 8453
rect 14014 8440 14026 8453
rect 14076 8440 14082 8453
rect 14082 8440 14110 8453
rect 14185 8419 14218 8435
rect 14218 8419 14219 8435
rect 14257 8419 14286 8435
rect 14286 8419 14291 8435
rect 14329 8419 14354 8435
rect 14354 8419 14363 8435
rect 14401 8419 14422 8435
rect 14422 8419 14435 8435
rect 14473 8419 14490 8435
rect 14490 8419 14507 8435
rect 14614 8428 14626 8453
rect 14626 8428 14648 8453
rect 14692 8428 14694 8453
rect 14694 8428 14726 8453
rect 14770 8428 14796 8453
rect 14796 8428 14804 8453
rect 14848 8428 14864 8453
rect 14864 8428 14882 8453
rect 14926 8433 14960 8462
rect 15004 8433 15038 8462
rect 14926 8428 14932 8433
rect 14932 8428 14960 8433
rect 14185 8401 14219 8419
rect 14257 8401 14291 8419
rect 14329 8401 14363 8419
rect 14401 8401 14435 8419
rect 14473 8401 14507 8419
rect 248 8321 251 8355
rect 251 8321 282 8355
rect 320 8321 353 8355
rect 353 8321 354 8355
rect 392 8321 421 8355
rect 421 8321 426 8355
rect 2456 8321 2461 8355
rect 2461 8321 2490 8355
rect 2528 8321 2529 8355
rect 2529 8321 2562 8355
rect 2600 8321 2631 8355
rect 2631 8321 2634 8355
rect 13992 8367 14026 8401
rect 14076 8367 14110 8401
rect 15004 8428 15034 8433
rect 15034 8428 15038 8433
rect 14185 8357 14219 8358
rect 14257 8357 14291 8358
rect 14329 8357 14363 8358
rect 14401 8357 14435 8358
rect 14473 8357 14507 8358
rect 14614 8357 14648 8388
rect 14692 8357 14726 8388
rect 14770 8357 14804 8388
rect 14848 8357 14882 8388
rect 14926 8361 14960 8388
rect 15004 8361 15038 8388
rect 14185 8324 14198 8357
rect 14198 8324 14219 8357
rect 14257 8324 14268 8357
rect 14268 8324 14291 8357
rect 14329 8324 14338 8357
rect 14338 8324 14363 8357
rect 14401 8324 14408 8357
rect 14408 8324 14435 8357
rect 14473 8324 14478 8357
rect 14478 8324 14507 8357
rect 14614 8354 14618 8357
rect 14618 8354 14648 8357
rect 14692 8354 14724 8357
rect 14724 8354 14726 8357
rect 14770 8354 14794 8357
rect 14794 8354 14804 8357
rect 14848 8354 14864 8357
rect 14864 8354 14882 8357
rect 14926 8354 14932 8361
rect 14932 8354 14960 8361
rect 15004 8354 15034 8361
rect 15034 8354 15038 8361
rect 14614 8283 14648 8314
rect 14692 8283 14726 8314
rect 14770 8283 14804 8314
rect 14848 8283 14882 8314
rect 14926 8289 14960 8314
rect 15004 8289 15038 8314
rect 8509 8239 8615 8254
rect 8509 7933 8510 8239
rect 8510 7933 8612 8239
rect 8612 7933 8615 8239
rect 8509 7932 8615 7933
rect 9596 8239 9630 8247
rect 9678 8239 9712 8247
rect 9596 8213 9612 8239
rect 9612 8213 9630 8239
rect 9678 8213 9712 8239
rect 9596 8110 9612 8144
rect 9612 8110 9630 8144
rect 9678 8110 9712 8144
rect 9596 8007 9612 8041
rect 9612 8007 9630 8041
rect 9678 8007 9712 8041
rect 10314 8239 10348 8247
rect 10396 8239 10430 8247
rect 10314 8213 10348 8239
rect 10396 8213 10416 8239
rect 10416 8213 10430 8239
rect 10314 8110 10348 8144
rect 10396 8110 10416 8144
rect 10416 8110 10430 8144
rect 10314 8007 10348 8041
rect 10396 8007 10416 8041
rect 10416 8007 10430 8041
rect 10804 8239 10838 8254
rect 10898 8239 10932 8254
rect 10804 8220 10816 8239
rect 10816 8220 10838 8239
rect 10898 8220 10918 8239
rect 10918 8220 10932 8239
rect 10804 8145 10816 8179
rect 10816 8145 10838 8179
rect 10898 8145 10918 8179
rect 10918 8145 10932 8179
rect 10804 8070 10816 8104
rect 10816 8070 10838 8104
rect 10898 8070 10918 8104
rect 10918 8070 10932 8104
rect 10804 7994 10816 8028
rect 10816 7994 10838 8028
rect 10898 7994 10918 8028
rect 10918 7994 10932 8028
rect 10804 7933 10816 7952
rect 10816 7933 10838 7952
rect 10898 7933 10918 7952
rect 10918 7933 10932 7952
rect 10804 7918 10838 7933
rect 10898 7918 10932 7933
rect 14185 8249 14198 8280
rect 14198 8249 14219 8280
rect 14257 8249 14268 8280
rect 14268 8249 14291 8280
rect 14329 8249 14338 8280
rect 14338 8249 14363 8280
rect 14401 8249 14408 8280
rect 14408 8249 14435 8280
rect 14473 8249 14478 8280
rect 14478 8249 14507 8280
rect 14614 8280 14618 8283
rect 14618 8280 14648 8283
rect 14692 8280 14724 8283
rect 14724 8280 14726 8283
rect 14770 8280 14794 8283
rect 14794 8280 14804 8283
rect 14848 8280 14864 8283
rect 14864 8280 14882 8283
rect 14926 8280 14932 8289
rect 14932 8280 14960 8289
rect 15004 8280 15034 8289
rect 15034 8280 15038 8289
rect 14185 8246 14219 8249
rect 14257 8246 14291 8249
rect 14329 8246 14363 8249
rect 14401 8246 14435 8249
rect 14473 8246 14507 8249
rect 14614 8209 14648 8240
rect 14692 8209 14726 8240
rect 14770 8209 14804 8240
rect 14848 8209 14882 8240
rect 14926 8217 14960 8240
rect 15004 8217 15038 8240
rect 14185 8175 14198 8202
rect 14198 8175 14219 8202
rect 14257 8175 14268 8202
rect 14268 8175 14291 8202
rect 14329 8175 14338 8202
rect 14338 8175 14363 8202
rect 14401 8175 14408 8202
rect 14408 8175 14435 8202
rect 14473 8175 14478 8202
rect 14478 8175 14507 8202
rect 14614 8206 14618 8209
rect 14618 8206 14648 8209
rect 14692 8206 14724 8209
rect 14724 8206 14726 8209
rect 14770 8206 14794 8209
rect 14794 8206 14804 8209
rect 14848 8206 14864 8209
rect 14864 8206 14882 8209
rect 14926 8206 14932 8217
rect 14932 8206 14960 8217
rect 15004 8206 15034 8217
rect 15034 8206 15038 8217
rect 14185 8168 14219 8175
rect 14257 8168 14291 8175
rect 14329 8168 14363 8175
rect 14401 8168 14435 8175
rect 14473 8168 14507 8175
rect 14614 8135 14648 8166
rect 14692 8135 14726 8166
rect 14770 8135 14804 8166
rect 14848 8135 14882 8166
rect 14926 8145 14960 8166
rect 15004 8145 15038 8166
rect 14431 8101 14444 8115
rect 14444 8101 14465 8115
rect 14511 8101 14514 8115
rect 14514 8101 14545 8115
rect 14614 8132 14618 8135
rect 14618 8132 14648 8135
rect 14692 8132 14724 8135
rect 14724 8132 14726 8135
rect 14770 8132 14794 8135
rect 14794 8132 14804 8135
rect 14848 8132 14864 8135
rect 14864 8132 14882 8135
rect 14926 8132 14932 8145
rect 14932 8132 14960 8145
rect 15004 8132 15034 8145
rect 15034 8132 15038 8145
rect 14431 8081 14465 8101
rect 14511 8081 14545 8101
rect 14614 8061 14648 8092
rect 14692 8061 14726 8092
rect 14770 8061 14804 8092
rect 14848 8061 14882 8092
rect 14926 8073 14960 8092
rect 15004 8073 15038 8092
rect 14431 8027 14444 8033
rect 14444 8027 14465 8033
rect 14511 8027 14514 8033
rect 14514 8027 14545 8033
rect 14614 8058 14618 8061
rect 14618 8058 14648 8061
rect 14692 8058 14724 8061
rect 14724 8058 14726 8061
rect 14770 8058 14794 8061
rect 14794 8058 14804 8061
rect 14848 8058 14864 8061
rect 14864 8058 14882 8061
rect 14926 8058 14932 8073
rect 14932 8058 14960 8073
rect 15004 8058 15034 8073
rect 15034 8058 15038 8073
rect 14431 7999 14465 8027
rect 14511 7999 14545 8027
rect 14614 7987 14648 8018
rect 14692 7987 14726 8018
rect 14770 7987 14804 8018
rect 14848 7987 14882 8018
rect 14926 8001 14960 8018
rect 15004 8001 15038 8018
rect 14614 7984 14618 7987
rect 14618 7984 14648 7987
rect 14692 7984 14724 7987
rect 14724 7984 14726 7987
rect 14770 7984 14794 7987
rect 14794 7984 14804 7987
rect 14848 7984 14864 7987
rect 14864 7984 14882 7987
rect 14926 7984 14932 8001
rect 14932 7984 14960 8001
rect 15004 7984 15034 8001
rect 15034 7984 15038 8001
rect 14431 7916 14465 7950
rect 14511 7916 14545 7950
rect 14614 7913 14648 7944
rect 14692 7913 14726 7944
rect 14770 7913 14804 7944
rect 14848 7913 14882 7944
rect 14926 7929 14960 7944
rect 15004 7929 15038 7944
rect 14614 7910 14618 7913
rect 14618 7910 14648 7913
rect 14692 7910 14724 7913
rect 14724 7910 14726 7913
rect 14770 7910 14794 7913
rect 14794 7910 14804 7913
rect 14848 7910 14864 7913
rect 14864 7910 14882 7913
rect 14926 7910 14932 7929
rect 14932 7910 14960 7929
rect 15004 7910 15034 7929
rect 15034 7910 15038 7929
rect 14614 7839 14648 7870
rect 14692 7839 14726 7870
rect 14770 7839 14804 7870
rect 14848 7839 14882 7870
rect 14926 7857 14960 7870
rect 15004 7857 15038 7870
rect 14614 7836 14618 7839
rect 14618 7836 14648 7839
rect 14692 7836 14724 7839
rect 14724 7836 14726 7839
rect 14770 7836 14794 7839
rect 14794 7836 14804 7839
rect 14848 7836 14864 7839
rect 14864 7836 14882 7839
rect 14926 7836 14932 7857
rect 14932 7836 14960 7857
rect 15004 7836 15034 7857
rect 15034 7836 15038 7857
rect 14614 7762 14648 7796
rect 14692 7762 14726 7796
rect 14770 7762 14804 7796
rect 14848 7762 14882 7796
rect 14926 7785 14960 7796
rect 15004 7785 15038 7796
rect 14926 7762 14932 7785
rect 14932 7762 14960 7785
rect 15004 7762 15034 7785
rect 15034 7762 15038 7785
rect 14614 7715 14626 7722
rect 14626 7715 14648 7722
rect 14692 7715 14694 7722
rect 14694 7715 14726 7722
rect 14770 7715 14796 7722
rect 14796 7715 14804 7722
rect 14848 7715 14864 7722
rect 14864 7715 14882 7722
rect 14614 7688 14648 7715
rect 14692 7688 14726 7715
rect 14770 7688 14804 7715
rect 14848 7688 14882 7715
rect 14926 7713 14960 7722
rect 15004 7713 15038 7722
rect 14926 7688 14932 7713
rect 14932 7688 14960 7713
rect 15004 7688 15034 7713
rect 15034 7688 15038 7713
rect 14614 7640 14648 7648
rect 14692 7640 14726 7648
rect 14770 7640 14804 7648
rect 14848 7640 14882 7648
rect 14926 7641 14960 7648
rect 15004 7641 15038 7648
rect 14614 7614 14626 7640
rect 14626 7614 14648 7640
rect 14692 7614 14694 7640
rect 14694 7614 14726 7640
rect 14770 7614 14796 7640
rect 14796 7614 14804 7640
rect 14848 7614 14864 7640
rect 14864 7614 14882 7640
rect 14926 7614 14932 7641
rect 14932 7614 14960 7641
rect 15004 7614 15034 7641
rect 15034 7614 15038 7641
rect 14614 7556 14648 7574
rect 14692 7556 14726 7574
rect 14770 7556 14804 7574
rect 14848 7556 14882 7574
rect 14926 7569 14960 7574
rect 15004 7569 15038 7574
rect 14614 7540 14626 7556
rect 14626 7540 14648 7556
rect 14692 7540 14694 7556
rect 14694 7540 14726 7556
rect 14770 7540 14796 7556
rect 14796 7540 14804 7556
rect 14848 7540 14864 7556
rect 14864 7540 14882 7556
rect 14926 7540 14932 7569
rect 14932 7540 14960 7569
rect 15004 7540 15034 7569
rect 15034 7540 15038 7569
rect 14614 7472 14648 7499
rect 14692 7472 14726 7499
rect 14770 7472 14804 7499
rect 14848 7472 14882 7499
rect 14926 7497 14960 7499
rect 15004 7497 15038 7499
rect 14614 7465 14626 7472
rect 14626 7465 14648 7472
rect 14692 7465 14694 7472
rect 14694 7465 14726 7472
rect 14770 7465 14796 7472
rect 14796 7465 14804 7472
rect 14848 7465 14864 7472
rect 14864 7465 14882 7472
rect 14926 7465 14932 7497
rect 14932 7465 14960 7497
rect 15004 7465 15034 7497
rect 15034 7465 15038 7497
rect 14614 7390 14648 7424
rect 14692 7390 14726 7424
rect 14770 7390 14804 7424
rect 14848 7390 14882 7424
rect 14926 7391 14932 7424
rect 14932 7391 14960 7424
rect 15004 7391 15034 7424
rect 15034 7391 15038 7424
rect 14926 7390 14960 7391
rect 15004 7390 15038 7391
rect 57 7354 91 7374
rect 132 7354 166 7374
rect 207 7354 241 7374
rect 282 7354 316 7374
rect 357 7354 391 7374
rect 432 7354 466 7374
rect 507 7354 541 7374
rect 582 7354 616 7374
rect 657 7354 691 7374
rect 732 7354 766 7374
rect 807 7354 841 7374
rect 882 7354 916 7374
rect 957 7354 991 7374
rect 1032 7354 1066 7374
rect 1107 7354 1141 7374
rect 1182 7354 1216 7374
rect 1256 7354 1290 7374
rect 1330 7354 1364 7374
rect 57 7340 68 7354
rect 68 7340 91 7354
rect 132 7340 137 7354
rect 137 7340 166 7354
rect 207 7340 240 7354
rect 240 7340 241 7354
rect 282 7340 309 7354
rect 309 7340 316 7354
rect 357 7340 378 7354
rect 378 7340 391 7354
rect 432 7340 447 7354
rect 447 7340 466 7354
rect 507 7340 516 7354
rect 516 7340 541 7354
rect 582 7340 585 7354
rect 585 7340 616 7354
rect 657 7340 689 7354
rect 689 7340 691 7354
rect 732 7340 758 7354
rect 758 7340 766 7354
rect 807 7340 827 7354
rect 827 7340 841 7354
rect 882 7340 896 7354
rect 896 7340 916 7354
rect 957 7340 965 7354
rect 965 7340 991 7354
rect 1032 7340 1033 7354
rect 1033 7340 1066 7354
rect 1107 7340 1135 7354
rect 1135 7340 1141 7354
rect 1182 7340 1203 7354
rect 1203 7340 1216 7354
rect 1256 7340 1271 7354
rect 1271 7340 1290 7354
rect 1330 7340 1339 7354
rect 1339 7340 1364 7354
rect 57 7282 91 7290
rect 132 7282 166 7290
rect 207 7282 241 7290
rect 282 7282 316 7290
rect 357 7282 391 7290
rect 432 7282 466 7290
rect 507 7282 541 7290
rect 582 7282 616 7290
rect 657 7282 691 7290
rect 732 7282 766 7290
rect 807 7282 841 7290
rect 882 7282 916 7290
rect 957 7282 991 7290
rect 1032 7282 1066 7290
rect 1107 7282 1141 7290
rect 1182 7282 1216 7290
rect 1256 7282 1290 7290
rect 1330 7282 1364 7290
rect 57 7256 68 7282
rect 68 7256 91 7282
rect 132 7256 137 7282
rect 137 7256 166 7282
rect 207 7256 240 7282
rect 240 7256 241 7282
rect 282 7256 309 7282
rect 309 7256 316 7282
rect 357 7256 378 7282
rect 378 7256 391 7282
rect 432 7256 447 7282
rect 447 7256 466 7282
rect 507 7256 516 7282
rect 516 7256 541 7282
rect 582 7256 585 7282
rect 585 7256 616 7282
rect 657 7256 689 7282
rect 689 7256 691 7282
rect 732 7256 758 7282
rect 758 7256 766 7282
rect 807 7256 827 7282
rect 827 7256 841 7282
rect 882 7256 896 7282
rect 896 7256 916 7282
rect 957 7256 965 7282
rect 965 7256 991 7282
rect 1032 7256 1033 7282
rect 1033 7256 1066 7282
rect 1107 7256 1135 7282
rect 1135 7256 1141 7282
rect 1182 7256 1203 7282
rect 1203 7256 1216 7282
rect 1256 7256 1271 7282
rect 1271 7256 1290 7282
rect 1330 7256 1339 7282
rect 1339 7256 1364 7282
rect 1431 7210 1465 7220
rect 1504 7210 1538 7220
rect 1577 7210 1611 7220
rect 1650 7210 1684 7220
rect 1723 7210 1757 7220
rect 1796 7210 1830 7220
rect 1869 7210 1903 7220
rect 1942 7210 1976 7220
rect 2015 7210 2049 7220
rect 2088 7210 2122 7220
rect 2161 7210 2195 7220
rect 2234 7210 2268 7220
rect 2307 7210 2341 7220
rect 2380 7210 2414 7220
rect 2453 7210 2487 7220
rect 2526 7210 2560 7220
rect 2599 7210 2633 7220
rect 2672 7210 2706 7220
rect 57 7176 68 7206
rect 68 7176 91 7206
rect 132 7176 137 7206
rect 137 7176 166 7206
rect 207 7176 240 7206
rect 240 7176 241 7206
rect 282 7176 309 7206
rect 309 7176 316 7206
rect 357 7176 378 7206
rect 378 7176 391 7206
rect 432 7176 447 7206
rect 447 7176 466 7206
rect 507 7176 516 7206
rect 516 7176 541 7206
rect 582 7176 585 7206
rect 585 7176 616 7206
rect 657 7176 689 7206
rect 689 7176 691 7206
rect 732 7176 758 7206
rect 758 7176 766 7206
rect 807 7176 827 7206
rect 827 7176 841 7206
rect 882 7176 896 7206
rect 896 7176 916 7206
rect 957 7176 965 7206
rect 965 7176 991 7206
rect 1032 7176 1033 7206
rect 1033 7176 1066 7206
rect 1107 7176 1135 7206
rect 1135 7176 1141 7206
rect 1182 7176 1203 7206
rect 1203 7176 1216 7206
rect 1256 7176 1271 7206
rect 1271 7176 1290 7206
rect 1330 7176 1339 7206
rect 1339 7176 1364 7206
rect 1431 7186 1441 7210
rect 1441 7186 1465 7210
rect 1504 7186 1509 7210
rect 1509 7186 1538 7210
rect 1577 7186 1611 7210
rect 1650 7186 1679 7210
rect 1679 7186 1684 7210
rect 1723 7186 1747 7210
rect 1747 7186 1757 7210
rect 1796 7186 1815 7210
rect 1815 7186 1830 7210
rect 1869 7186 1883 7210
rect 1883 7186 1903 7210
rect 1942 7186 1951 7210
rect 1951 7186 1976 7210
rect 2015 7186 2019 7210
rect 2019 7186 2049 7210
rect 2088 7186 2121 7210
rect 2121 7186 2122 7210
rect 2161 7186 2189 7210
rect 2189 7186 2195 7210
rect 2234 7186 2257 7210
rect 2257 7186 2268 7210
rect 2307 7186 2325 7210
rect 2325 7186 2341 7210
rect 2380 7186 2393 7210
rect 2393 7186 2414 7210
rect 2453 7186 2461 7210
rect 2461 7186 2487 7210
rect 2526 7186 2529 7210
rect 2529 7186 2560 7210
rect 2599 7186 2631 7210
rect 2631 7186 2633 7210
rect 2672 7186 2699 7210
rect 2699 7186 2706 7210
rect 2745 7186 2779 7220
rect 2818 7186 2852 7220
rect 2891 7186 2925 7220
rect 2964 7186 2998 7220
rect 3037 7186 3071 7220
rect 3110 7186 3144 7220
rect 3183 7186 3217 7220
rect 3256 7186 3290 7220
rect 3329 7186 3363 7220
rect 3402 7186 3436 7220
rect 3475 7186 3509 7220
rect 3548 7186 3582 7220
rect 3621 7186 3655 7220
rect 3694 7186 3728 7220
rect 3767 7186 3801 7220
rect 3840 7186 3874 7220
rect 3913 7186 3947 7220
rect 3986 7186 4020 7220
rect 4059 7186 4093 7220
rect 4132 7186 4166 7220
rect 4205 7186 4239 7220
rect 4278 7186 4312 7220
rect 4351 7186 4385 7220
rect 4424 7186 4458 7220
rect 4497 7186 4531 7220
rect 4570 7186 4604 7220
rect 4643 7186 4677 7220
rect 4716 7186 4750 7220
rect 4789 7186 4823 7220
rect 4862 7186 4896 7220
rect 4935 7186 4969 7220
rect 5008 7186 5042 7220
rect 5081 7186 5115 7220
rect 5154 7186 5188 7220
rect 5227 7186 5261 7220
rect 5300 7186 5334 7220
rect 5373 7186 5407 7220
rect 5446 7186 5480 7220
rect 5519 7186 5553 7220
rect 5592 7186 5626 7220
rect 5665 7186 5699 7220
rect 5738 7186 5772 7220
rect 5811 7186 5845 7220
rect 5884 7186 5918 7220
rect 5957 7186 5991 7220
rect 6030 7186 6064 7220
rect 6103 7186 6137 7220
rect 6176 7186 6210 7220
rect 6249 7186 6283 7220
rect 6322 7186 6356 7220
rect 6395 7186 6429 7220
rect 6468 7186 6502 7220
rect 6540 7186 6574 7220
rect 6612 7186 6646 7220
rect 6684 7186 6718 7220
rect 6756 7186 6790 7220
rect 6828 7186 6862 7220
rect 6900 7186 6934 7220
rect 6972 7186 7006 7220
rect 7044 7186 7078 7220
rect 7116 7186 7150 7220
rect 57 7172 91 7176
rect 132 7172 166 7176
rect 207 7172 241 7176
rect 282 7172 316 7176
rect 357 7172 391 7176
rect 432 7172 466 7176
rect 507 7172 541 7176
rect 582 7172 616 7176
rect 657 7172 691 7176
rect 732 7172 766 7176
rect 807 7172 841 7176
rect 882 7172 916 7176
rect 957 7172 991 7176
rect 1032 7172 1066 7176
rect 1107 7172 1141 7176
rect 1182 7172 1216 7176
rect 1256 7172 1290 7176
rect 1330 7172 1364 7176
rect 57 7104 68 7122
rect 68 7104 91 7122
rect 132 7104 137 7122
rect 137 7104 166 7122
rect 207 7104 240 7122
rect 240 7104 241 7122
rect 282 7104 309 7122
rect 309 7104 316 7122
rect 357 7104 378 7122
rect 378 7104 391 7122
rect 432 7104 447 7122
rect 447 7104 466 7122
rect 507 7104 516 7122
rect 516 7104 541 7122
rect 582 7104 585 7122
rect 585 7104 616 7122
rect 657 7104 689 7122
rect 689 7104 691 7122
rect 732 7104 758 7122
rect 758 7104 766 7122
rect 807 7104 827 7122
rect 827 7104 841 7122
rect 882 7104 896 7122
rect 896 7104 916 7122
rect 957 7104 965 7122
rect 965 7104 991 7122
rect 1032 7104 1033 7122
rect 1033 7104 1066 7122
rect 1107 7104 1135 7122
rect 1135 7104 1141 7122
rect 1182 7104 1203 7122
rect 1203 7104 1216 7122
rect 1256 7104 1271 7122
rect 1271 7104 1290 7122
rect 1330 7104 1339 7122
rect 1339 7104 1364 7122
rect 57 7088 91 7104
rect 132 7088 166 7104
rect 207 7088 241 7104
rect 282 7088 316 7104
rect 357 7088 391 7104
rect 432 7088 466 7104
rect 507 7088 541 7104
rect 582 7088 616 7104
rect 657 7088 691 7104
rect 732 7088 766 7104
rect 807 7088 841 7104
rect 882 7088 916 7104
rect 957 7088 991 7104
rect 1032 7088 1066 7104
rect 1107 7088 1141 7104
rect 1182 7088 1216 7104
rect 1256 7088 1290 7104
rect 1330 7088 1364 7104
rect 57 7032 68 7038
rect 68 7032 91 7038
rect 132 7032 137 7038
rect 137 7032 166 7038
rect 207 7032 240 7038
rect 240 7032 241 7038
rect 282 7032 309 7038
rect 309 7032 316 7038
rect 357 7032 378 7038
rect 378 7032 391 7038
rect 432 7032 447 7038
rect 447 7032 466 7038
rect 507 7032 516 7038
rect 516 7032 541 7038
rect 582 7032 585 7038
rect 585 7032 616 7038
rect 657 7032 689 7038
rect 689 7032 691 7038
rect 732 7032 758 7038
rect 758 7032 766 7038
rect 807 7032 827 7038
rect 827 7032 841 7038
rect 882 7032 896 7038
rect 896 7032 916 7038
rect 957 7032 965 7038
rect 965 7032 991 7038
rect 1032 7032 1033 7038
rect 1033 7032 1066 7038
rect 1107 7032 1135 7038
rect 1135 7032 1141 7038
rect 1182 7032 1203 7038
rect 1203 7032 1216 7038
rect 1256 7032 1271 7038
rect 1271 7032 1290 7038
rect 1330 7032 1339 7038
rect 1339 7032 1364 7038
rect 57 7004 91 7032
rect 132 7004 166 7032
rect 207 7004 241 7032
rect 282 7004 316 7032
rect 357 7004 391 7032
rect 432 7004 466 7032
rect 507 7004 541 7032
rect 582 7004 616 7032
rect 657 7004 691 7032
rect 732 7004 766 7032
rect 807 7004 841 7032
rect 882 7004 916 7032
rect 957 7004 991 7032
rect 1032 7004 1066 7032
rect 1107 7004 1141 7032
rect 1182 7004 1216 7032
rect 1256 7004 1290 7032
rect 1330 7004 1364 7032
rect 14614 7315 14648 7349
rect 14692 7315 14726 7349
rect 14770 7315 14804 7349
rect 14848 7315 14882 7349
rect 14926 7319 14932 7349
rect 14932 7319 14960 7349
rect 15004 7319 15034 7349
rect 15034 7319 15038 7349
rect 14926 7315 14960 7319
rect 15004 7315 15038 7319
rect 14614 7248 14626 7274
rect 14626 7248 14648 7274
rect 14692 7248 14694 7274
rect 14694 7248 14726 7274
rect 14770 7248 14796 7274
rect 14796 7248 14804 7274
rect 14848 7248 14864 7274
rect 14864 7248 14882 7274
rect 14614 7240 14648 7248
rect 14692 7240 14726 7248
rect 14770 7240 14804 7248
rect 14848 7240 14882 7248
rect 14926 7247 14932 7274
rect 14932 7247 14960 7274
rect 15004 7247 15034 7274
rect 15034 7247 15038 7274
rect 14926 7240 14960 7247
rect 15004 7240 15038 7247
rect 14614 7176 14626 7199
rect 14626 7176 14648 7199
rect 14692 7176 14694 7199
rect 14694 7176 14726 7199
rect 14770 7176 14796 7199
rect 14796 7176 14804 7199
rect 14848 7176 14864 7199
rect 14864 7176 14882 7199
rect 14614 7165 14648 7176
rect 14692 7165 14726 7176
rect 14770 7165 14804 7176
rect 14848 7165 14882 7176
rect 14926 7175 14932 7199
rect 14932 7175 14960 7199
rect 15004 7175 15034 7199
rect 15034 7175 15038 7199
rect 14926 7165 14960 7175
rect 15004 7165 15038 7175
rect 14614 7104 14626 7124
rect 14626 7104 14648 7124
rect 14692 7104 14694 7124
rect 14694 7104 14726 7124
rect 14770 7104 14796 7124
rect 14796 7104 14804 7124
rect 14848 7104 14864 7124
rect 14864 7104 14882 7124
rect 14614 7090 14648 7104
rect 14692 7090 14726 7104
rect 14770 7090 14804 7104
rect 14848 7090 14882 7104
rect 14926 7103 14932 7124
rect 14932 7103 14960 7124
rect 15004 7103 15034 7124
rect 15034 7103 15038 7124
rect 14926 7090 14960 7103
rect 15004 7090 15038 7103
rect 15068 6805 15102 6825
rect 15068 6791 15102 6805
rect 15068 6731 15102 6753
rect 15068 6719 15102 6731
rect 15068 6657 15102 6681
rect 15068 6647 15102 6657
rect 15068 6583 15102 6609
rect 15068 6575 15102 6583
rect 15068 6509 15102 6537
rect 15068 6503 15102 6509
rect 68 6434 102 6439
rect 141 6434 175 6439
rect 214 6434 248 6439
rect 287 6434 321 6439
rect 360 6434 394 6439
rect 433 6434 467 6439
rect 506 6434 540 6439
rect 579 6434 613 6439
rect 652 6434 686 6439
rect 725 6434 759 6439
rect 798 6434 832 6439
rect 871 6434 905 6439
rect 944 6434 978 6439
rect 1017 6434 1051 6439
rect 1090 6435 15020 6439
rect 15068 6435 15102 6465
rect 1090 6434 14932 6435
rect 68 6405 102 6434
rect 141 6405 171 6434
rect 171 6405 175 6434
rect 214 6405 240 6434
rect 240 6405 248 6434
rect 287 6405 309 6434
rect 309 6405 321 6434
rect 360 6405 378 6434
rect 378 6405 394 6434
rect 433 6405 447 6434
rect 447 6405 467 6434
rect 506 6405 516 6434
rect 516 6405 540 6434
rect 579 6405 585 6434
rect 585 6405 613 6434
rect 652 6405 654 6434
rect 654 6405 686 6434
rect 725 6405 758 6434
rect 758 6405 759 6434
rect 798 6405 827 6434
rect 827 6405 832 6434
rect 871 6405 896 6434
rect 896 6405 905 6434
rect 944 6405 965 6434
rect 965 6405 978 6434
rect 1017 6405 1034 6434
rect 1034 6405 1051 6434
rect 1090 6400 1103 6434
rect 1103 6400 1137 6434
rect 1137 6400 1172 6434
rect 1172 6400 1206 6434
rect 1206 6400 1241 6434
rect 1241 6400 1275 6434
rect 1275 6400 1310 6434
rect 1310 6400 1344 6434
rect 1344 6400 1379 6434
rect 1379 6400 1413 6434
rect 1413 6400 1448 6434
rect 1448 6400 1482 6434
rect 1482 6400 1517 6434
rect 1517 6400 1551 6434
rect 1551 6400 1586 6434
rect 1586 6400 1620 6434
rect 1620 6400 1655 6434
rect 1655 6400 1689 6434
rect 1689 6400 1724 6434
rect 1724 6400 1758 6434
rect 1758 6400 1793 6434
rect 1793 6400 1827 6434
rect 1827 6400 1862 6434
rect 1862 6400 1896 6434
rect 1896 6400 1931 6434
rect 1931 6400 1965 6434
rect 1965 6400 2000 6434
rect 2000 6400 2034 6434
rect 2034 6400 2069 6434
rect 2069 6400 2103 6434
rect 2103 6400 2138 6434
rect 2138 6400 2172 6434
rect 2172 6400 2207 6434
rect 2207 6400 2241 6434
rect 2241 6400 2276 6434
rect 2276 6400 2310 6434
rect 2310 6400 2345 6434
rect 2345 6400 2379 6434
rect 2379 6400 2414 6434
rect 2414 6400 2448 6434
rect 2448 6400 2483 6434
rect 2483 6400 2517 6434
rect 2517 6400 2551 6434
rect 2551 6400 2585 6434
rect 2585 6400 2619 6434
rect 2619 6400 2653 6434
rect 2653 6400 2687 6434
rect 2687 6400 2721 6434
rect 2721 6400 2755 6434
rect 2755 6400 2789 6434
rect 2789 6400 2823 6434
rect 2823 6400 2857 6434
rect 2857 6400 2891 6434
rect 2891 6400 2925 6434
rect 2925 6400 2959 6434
rect 2959 6400 2993 6434
rect 2993 6400 3027 6434
rect 3027 6400 3061 6434
rect 3061 6400 3095 6434
rect 3095 6400 3129 6434
rect 3129 6400 3163 6434
rect 3163 6400 3197 6434
rect 3197 6400 3231 6434
rect 3231 6400 3265 6434
rect 3265 6400 3299 6434
rect 3299 6400 3333 6434
rect 3333 6400 3367 6434
rect 3367 6400 3401 6434
rect 3401 6400 3435 6434
rect 3435 6400 3469 6434
rect 3469 6400 3503 6434
rect 3503 6400 3537 6434
rect 3537 6400 3571 6434
rect 3571 6400 3605 6434
rect 3605 6400 3639 6434
rect 3639 6400 3673 6434
rect 3673 6400 3707 6434
rect 3707 6400 3741 6434
rect 3741 6400 3775 6434
rect 3775 6400 3809 6434
rect 3809 6400 3843 6434
rect 3843 6400 3877 6434
rect 3877 6400 3911 6434
rect 3911 6400 3945 6434
rect 3945 6400 3979 6434
rect 3979 6400 4013 6434
rect 4013 6400 4047 6434
rect 4047 6400 4081 6434
rect 4081 6400 4115 6434
rect 4115 6400 4149 6434
rect 4149 6400 4183 6434
rect 4183 6400 4217 6434
rect 4217 6400 4251 6434
rect 4251 6400 4285 6434
rect 4285 6400 4319 6434
rect 4319 6400 4353 6434
rect 4353 6400 4387 6434
rect 4387 6400 4421 6434
rect 4421 6400 4455 6434
rect 4455 6400 4489 6434
rect 4489 6400 4523 6434
rect 4523 6400 4557 6434
rect 4557 6400 4591 6434
rect 4591 6400 4625 6434
rect 4625 6400 4659 6434
rect 4659 6400 4693 6434
rect 4693 6400 4727 6434
rect 4727 6400 4761 6434
rect 4761 6400 4795 6434
rect 4795 6400 4829 6434
rect 4829 6400 4863 6434
rect 4863 6400 4897 6434
rect 4897 6400 4931 6434
rect 4931 6400 4965 6434
rect 4965 6400 4999 6434
rect 4999 6400 5033 6434
rect 5033 6400 5067 6434
rect 5067 6400 5101 6434
rect 5101 6400 5135 6434
rect 5135 6400 5169 6434
rect 5169 6400 5203 6434
rect 5203 6400 5237 6434
rect 5237 6400 5271 6434
rect 5271 6400 5305 6434
rect 5305 6400 5339 6434
rect 5339 6400 5373 6434
rect 5373 6400 5407 6434
rect 5407 6400 5441 6434
rect 5441 6400 5475 6434
rect 5475 6400 5509 6434
rect 5509 6400 5543 6434
rect 5543 6400 5577 6434
rect 5577 6400 5611 6434
rect 5611 6400 5645 6434
rect 5645 6400 5679 6434
rect 5679 6400 5713 6434
rect 5713 6400 5747 6434
rect 5747 6400 5781 6434
rect 5781 6400 5815 6434
rect 5815 6400 5849 6434
rect 5849 6400 5883 6434
rect 5883 6400 5917 6434
rect 5917 6400 5951 6434
rect 5951 6400 5985 6434
rect 5985 6400 6019 6434
rect 6019 6400 6053 6434
rect 6053 6400 6087 6434
rect 6087 6400 6121 6434
rect 6121 6400 6155 6434
rect 6155 6400 6189 6434
rect 6189 6400 6223 6434
rect 6223 6400 6257 6434
rect 6257 6400 6291 6434
rect 6291 6400 6325 6434
rect 6325 6400 6359 6434
rect 6359 6400 6393 6434
rect 6393 6400 6427 6434
rect 6427 6400 6461 6434
rect 6461 6400 6495 6434
rect 6495 6400 6529 6434
rect 6529 6400 6563 6434
rect 6563 6400 6597 6434
rect 6597 6400 6631 6434
rect 6631 6400 6665 6434
rect 6665 6400 6699 6434
rect 6699 6400 6733 6434
rect 6733 6400 6767 6434
rect 6767 6400 6801 6434
rect 6801 6400 6835 6434
rect 6835 6400 6869 6434
rect 6869 6400 6903 6434
rect 6903 6400 6937 6434
rect 6937 6400 6971 6434
rect 6971 6400 7005 6434
rect 7005 6400 7039 6434
rect 7039 6400 7073 6434
rect 7073 6400 7107 6434
rect 7107 6400 7141 6434
rect 7141 6400 7175 6434
rect 7175 6400 7209 6434
rect 7209 6400 7243 6434
rect 7243 6400 7277 6434
rect 7277 6400 7311 6434
rect 7311 6400 7345 6434
rect 7345 6400 7379 6434
rect 7379 6400 7413 6434
rect 7413 6400 7447 6434
rect 7447 6400 7481 6434
rect 7481 6400 7515 6434
rect 7515 6400 7549 6434
rect 7549 6400 7583 6434
rect 7583 6400 7617 6434
rect 7617 6400 7651 6434
rect 7651 6400 7685 6434
rect 7685 6400 7719 6434
rect 7719 6400 7753 6434
rect 7753 6400 7787 6434
rect 7787 6400 7821 6434
rect 7821 6400 7855 6434
rect 7855 6400 7889 6434
rect 7889 6400 7923 6434
rect 7923 6400 7957 6434
rect 7957 6400 7991 6434
rect 7991 6400 8025 6434
rect 8025 6400 8059 6434
rect 8059 6400 8093 6434
rect 8093 6400 8127 6434
rect 8127 6400 8161 6434
rect 8161 6400 8195 6434
rect 8195 6400 8229 6434
rect 8229 6400 8263 6434
rect 8263 6400 8297 6434
rect 8297 6400 8331 6434
rect 8331 6400 8365 6434
rect 8365 6400 8399 6434
rect 8399 6400 8433 6434
rect 8433 6400 8467 6434
rect 8467 6400 8501 6434
rect 8501 6400 8535 6434
rect 8535 6400 8569 6434
rect 8569 6400 8603 6434
rect 8603 6400 8637 6434
rect 8637 6400 8671 6434
rect 8671 6400 8705 6434
rect 8705 6400 8739 6434
rect 8739 6400 8773 6434
rect 8773 6400 8807 6434
rect 8807 6400 8841 6434
rect 8841 6400 8875 6434
rect 8875 6400 8909 6434
rect 8909 6400 8943 6434
rect 8943 6400 8977 6434
rect 8977 6400 9011 6434
rect 9011 6400 9045 6434
rect 9045 6400 9079 6434
rect 9079 6400 9113 6434
rect 9113 6400 9147 6434
rect 9147 6400 9181 6434
rect 9181 6400 9215 6434
rect 9215 6400 9249 6434
rect 9249 6400 9283 6434
rect 9283 6400 9317 6434
rect 9317 6400 9351 6434
rect 9351 6400 9385 6434
rect 9385 6400 9419 6434
rect 9419 6400 9453 6434
rect 9453 6400 9487 6434
rect 9487 6400 9521 6434
rect 9521 6400 9555 6434
rect 9555 6400 9589 6434
rect 9589 6400 9623 6434
rect 9623 6400 9657 6434
rect 9657 6400 9691 6434
rect 9691 6400 9725 6434
rect 9725 6400 9759 6434
rect 9759 6400 9793 6434
rect 9793 6400 9827 6434
rect 9827 6400 9861 6434
rect 9861 6400 9895 6434
rect 9895 6400 9929 6434
rect 9929 6400 9963 6434
rect 9963 6400 9997 6434
rect 9997 6400 10031 6434
rect 10031 6400 10065 6434
rect 10065 6400 10099 6434
rect 10099 6400 10133 6434
rect 10133 6400 10167 6434
rect 10167 6400 10201 6434
rect 10201 6400 10235 6434
rect 10235 6400 10269 6434
rect 10269 6400 10303 6434
rect 10303 6400 10337 6434
rect 10337 6400 10371 6434
rect 10371 6400 10405 6434
rect 10405 6400 10439 6434
rect 10439 6400 10473 6434
rect 10473 6400 10507 6434
rect 10507 6400 10541 6434
rect 10541 6400 10575 6434
rect 10575 6400 10609 6434
rect 10609 6400 10643 6434
rect 10643 6400 10677 6434
rect 10677 6400 10711 6434
rect 10711 6400 10745 6434
rect 10745 6400 10779 6434
rect 10779 6400 10813 6434
rect 10813 6400 10847 6434
rect 10847 6400 10881 6434
rect 10881 6400 10915 6434
rect 10915 6400 10949 6434
rect 10949 6400 10983 6434
rect 10983 6400 11017 6434
rect 11017 6400 11051 6434
rect 11051 6400 11085 6434
rect 11085 6400 11119 6434
rect 11119 6400 11153 6434
rect 11153 6400 11187 6434
rect 11187 6400 11221 6434
rect 11221 6400 11255 6434
rect 11255 6400 11289 6434
rect 11289 6400 11323 6434
rect 11323 6400 11357 6434
rect 11357 6400 11391 6434
rect 11391 6400 11425 6434
rect 11425 6400 11459 6434
rect 11459 6400 11493 6434
rect 11493 6400 11527 6434
rect 11527 6400 11561 6434
rect 11561 6400 11595 6434
rect 11595 6400 11629 6434
rect 11629 6400 11663 6434
rect 11663 6400 11697 6434
rect 11697 6400 11731 6434
rect 11731 6400 11765 6434
rect 11765 6400 11799 6434
rect 11799 6400 11833 6434
rect 11833 6400 11867 6434
rect 11867 6400 11901 6434
rect 11901 6400 11935 6434
rect 11935 6400 11969 6434
rect 11969 6400 12003 6434
rect 12003 6400 12037 6434
rect 12037 6400 12071 6434
rect 12071 6400 12105 6434
rect 12105 6400 12139 6434
rect 12139 6400 12173 6434
rect 12173 6400 12207 6434
rect 12207 6400 12241 6434
rect 12241 6400 12275 6434
rect 12275 6400 12309 6434
rect 12309 6400 12343 6434
rect 12343 6400 12377 6434
rect 12377 6400 12411 6434
rect 12411 6400 12445 6434
rect 12445 6400 12479 6434
rect 12479 6400 12513 6434
rect 12513 6400 12547 6434
rect 12547 6400 12581 6434
rect 12581 6400 12615 6434
rect 12615 6400 12649 6434
rect 12649 6400 12683 6434
rect 12683 6400 12717 6434
rect 12717 6400 12751 6434
rect 12751 6400 12785 6434
rect 12785 6400 12819 6434
rect 12819 6400 12853 6434
rect 12853 6400 12887 6434
rect 12887 6400 12921 6434
rect 12921 6400 12955 6434
rect 12955 6400 12989 6434
rect 12989 6400 13023 6434
rect 13023 6400 13057 6434
rect 13057 6400 13091 6434
rect 13091 6400 13125 6434
rect 13125 6400 13159 6434
rect 13159 6400 13193 6434
rect 13193 6400 13227 6434
rect 13227 6400 13261 6434
rect 13261 6400 13295 6434
rect 13295 6400 13329 6434
rect 13329 6400 13363 6434
rect 13363 6400 13397 6434
rect 13397 6400 13431 6434
rect 13431 6400 13465 6434
rect 13465 6400 13499 6434
rect 13499 6400 13533 6434
rect 13533 6400 13567 6434
rect 13567 6400 13601 6434
rect 13601 6400 13635 6434
rect 13635 6400 13669 6434
rect 13669 6400 13703 6434
rect 13703 6400 13737 6434
rect 13737 6400 13771 6434
rect 13771 6400 13805 6434
rect 13805 6400 13839 6434
rect 13839 6400 13873 6434
rect 13873 6400 13907 6434
rect 13907 6400 13941 6434
rect 13941 6400 13975 6434
rect 13975 6400 14009 6434
rect 14009 6400 14043 6434
rect 14043 6400 14077 6434
rect 14077 6400 14111 6434
rect 14111 6400 14145 6434
rect 14145 6400 14179 6434
rect 14179 6400 14213 6434
rect 14213 6400 14247 6434
rect 14247 6400 14281 6434
rect 14281 6400 14315 6434
rect 14315 6400 14349 6434
rect 14349 6400 14383 6434
rect 14383 6400 14417 6434
rect 14417 6400 14451 6434
rect 14451 6400 14485 6434
rect 14485 6400 14519 6434
rect 14519 6400 14553 6434
rect 14553 6400 14587 6434
rect 14587 6400 14621 6434
rect 14621 6400 14655 6434
rect 14655 6400 14689 6434
rect 14689 6400 14723 6434
rect 14723 6400 14757 6434
rect 14757 6400 14791 6434
rect 14791 6400 14825 6434
rect 14825 6400 14859 6434
rect 14859 6400 14893 6434
rect 14893 6401 14932 6434
rect 14932 6401 14966 6435
rect 14966 6401 15000 6435
rect 15000 6401 15020 6435
rect 15068 6431 15102 6435
rect 14893 6400 15020 6401
rect 68 6360 102 6367
rect 141 6360 175 6367
rect 214 6360 248 6367
rect 287 6360 321 6367
rect 360 6360 394 6367
rect 433 6360 467 6367
rect 506 6360 540 6367
rect 579 6360 613 6367
rect 652 6360 686 6367
rect 725 6360 759 6367
rect 798 6360 832 6367
rect 871 6360 905 6367
rect 944 6360 978 6367
rect 1017 6360 1051 6367
rect 1090 6360 15020 6400
rect 15068 6360 15102 6393
rect 68 6333 102 6360
rect 141 6333 171 6360
rect 171 6333 175 6360
rect 214 6333 240 6360
rect 240 6333 248 6360
rect 287 6333 309 6360
rect 309 6333 321 6360
rect 360 6333 378 6360
rect 378 6333 394 6360
rect 433 6333 447 6360
rect 447 6333 467 6360
rect 506 6333 516 6360
rect 516 6333 540 6360
rect 579 6333 585 6360
rect 585 6333 613 6360
rect 652 6333 654 6360
rect 654 6333 686 6360
rect 725 6333 758 6360
rect 758 6333 759 6360
rect 798 6333 827 6360
rect 827 6333 832 6360
rect 871 6333 896 6360
rect 896 6333 905 6360
rect 944 6333 965 6360
rect 965 6333 978 6360
rect 1017 6333 1034 6360
rect 1034 6333 1051 6360
rect 1090 6326 1103 6360
rect 1103 6326 1137 6360
rect 1137 6326 1172 6360
rect 1172 6326 1206 6360
rect 1206 6326 1241 6360
rect 1241 6326 1275 6360
rect 1275 6326 1310 6360
rect 1310 6326 1344 6360
rect 1344 6326 1379 6360
rect 1379 6326 1413 6360
rect 1413 6326 1448 6360
rect 1448 6326 1482 6360
rect 1482 6326 1517 6360
rect 1517 6326 1551 6360
rect 1551 6326 1586 6360
rect 1586 6326 1620 6360
rect 1620 6326 1655 6360
rect 1655 6326 1689 6360
rect 1689 6326 1724 6360
rect 1724 6326 1758 6360
rect 1758 6326 1793 6360
rect 1793 6326 1827 6360
rect 1827 6326 1862 6360
rect 1862 6326 1896 6360
rect 1896 6326 1931 6360
rect 1931 6326 1965 6360
rect 1965 6326 2000 6360
rect 2000 6326 2034 6360
rect 2034 6326 2069 6360
rect 2069 6326 2103 6360
rect 2103 6326 2138 6360
rect 2138 6326 2172 6360
rect 2172 6326 2207 6360
rect 2207 6326 2241 6360
rect 2241 6326 2276 6360
rect 2276 6326 2310 6360
rect 2310 6326 2345 6360
rect 2345 6326 2379 6360
rect 2379 6326 2414 6360
rect 2414 6326 2448 6360
rect 2448 6326 2483 6360
rect 2483 6326 2517 6360
rect 2517 6326 2551 6360
rect 2551 6326 2585 6360
rect 2585 6326 2619 6360
rect 2619 6326 2653 6360
rect 2653 6326 2687 6360
rect 2687 6326 2721 6360
rect 2721 6326 2755 6360
rect 2755 6326 2789 6360
rect 2789 6326 2823 6360
rect 2823 6326 2857 6360
rect 2857 6326 2891 6360
rect 2891 6326 2925 6360
rect 2925 6326 2959 6360
rect 2959 6326 2993 6360
rect 2993 6326 3027 6360
rect 3027 6326 3061 6360
rect 3061 6326 3095 6360
rect 3095 6326 3129 6360
rect 3129 6326 3163 6360
rect 3163 6326 3197 6360
rect 3197 6326 3231 6360
rect 3231 6326 3265 6360
rect 3265 6326 3299 6360
rect 3299 6326 3333 6360
rect 3333 6326 3367 6360
rect 3367 6326 3401 6360
rect 3401 6326 3435 6360
rect 3435 6326 3469 6360
rect 3469 6326 3503 6360
rect 3503 6326 3537 6360
rect 3537 6326 3571 6360
rect 3571 6326 3605 6360
rect 3605 6326 3639 6360
rect 3639 6326 3673 6360
rect 3673 6326 3707 6360
rect 3707 6326 3741 6360
rect 3741 6326 3775 6360
rect 3775 6326 3809 6360
rect 3809 6326 3843 6360
rect 3843 6326 3877 6360
rect 3877 6326 3911 6360
rect 3911 6326 3945 6360
rect 3945 6326 3979 6360
rect 3979 6326 4013 6360
rect 4013 6326 4047 6360
rect 4047 6326 4081 6360
rect 4081 6326 4115 6360
rect 4115 6326 4149 6360
rect 4149 6326 4183 6360
rect 4183 6326 4217 6360
rect 4217 6326 4251 6360
rect 4251 6326 4285 6360
rect 4285 6326 4319 6360
rect 4319 6326 4353 6360
rect 4353 6326 4387 6360
rect 4387 6326 4421 6360
rect 4421 6326 4455 6360
rect 4455 6326 4489 6360
rect 4489 6326 4523 6360
rect 4523 6326 4557 6360
rect 4557 6326 4591 6360
rect 4591 6326 4625 6360
rect 4625 6326 4659 6360
rect 4659 6326 4693 6360
rect 4693 6326 4727 6360
rect 4727 6326 4761 6360
rect 4761 6326 4795 6360
rect 4795 6326 4829 6360
rect 4829 6326 4863 6360
rect 4863 6326 4897 6360
rect 4897 6326 4931 6360
rect 4931 6326 4965 6360
rect 4965 6326 4999 6360
rect 4999 6326 5033 6360
rect 5033 6326 5067 6360
rect 5067 6326 5101 6360
rect 5101 6326 5135 6360
rect 5135 6326 5169 6360
rect 5169 6326 5203 6360
rect 5203 6326 5237 6360
rect 5237 6326 5271 6360
rect 5271 6326 5305 6360
rect 5305 6326 5339 6360
rect 5339 6326 5373 6360
rect 5373 6326 5407 6360
rect 5407 6326 5441 6360
rect 5441 6326 5475 6360
rect 5475 6326 5509 6360
rect 5509 6326 5543 6360
rect 5543 6326 5577 6360
rect 5577 6326 5611 6360
rect 5611 6326 5645 6360
rect 5645 6326 5679 6360
rect 5679 6326 5713 6360
rect 5713 6326 5747 6360
rect 5747 6326 5781 6360
rect 5781 6326 5815 6360
rect 5815 6326 5849 6360
rect 5849 6326 5883 6360
rect 5883 6326 5917 6360
rect 5917 6326 5951 6360
rect 5951 6326 5985 6360
rect 5985 6326 6019 6360
rect 6019 6326 6053 6360
rect 6053 6326 6087 6360
rect 6087 6326 6121 6360
rect 6121 6326 6155 6360
rect 6155 6326 6189 6360
rect 6189 6326 6223 6360
rect 6223 6326 6257 6360
rect 6257 6326 6291 6360
rect 6291 6326 6325 6360
rect 6325 6326 6359 6360
rect 6359 6326 6393 6360
rect 6393 6326 6427 6360
rect 6427 6326 6461 6360
rect 6461 6326 6495 6360
rect 6495 6326 6529 6360
rect 6529 6326 6563 6360
rect 6563 6326 6597 6360
rect 6597 6326 6631 6360
rect 6631 6326 6665 6360
rect 6665 6326 6699 6360
rect 6699 6326 6733 6360
rect 6733 6326 6767 6360
rect 6767 6326 6801 6360
rect 6801 6326 6835 6360
rect 6835 6326 6869 6360
rect 6869 6326 6903 6360
rect 6903 6326 6937 6360
rect 6937 6326 6971 6360
rect 6971 6326 7005 6360
rect 7005 6326 7039 6360
rect 7039 6326 7073 6360
rect 7073 6326 7107 6360
rect 7107 6326 7141 6360
rect 7141 6326 7175 6360
rect 7175 6326 7209 6360
rect 7209 6326 7243 6360
rect 7243 6326 7277 6360
rect 7277 6326 7311 6360
rect 7311 6326 7345 6360
rect 7345 6326 7379 6360
rect 7379 6326 7413 6360
rect 7413 6326 7447 6360
rect 7447 6326 7481 6360
rect 7481 6326 7515 6360
rect 7515 6326 7549 6360
rect 7549 6326 7583 6360
rect 7583 6326 7617 6360
rect 7617 6326 7651 6360
rect 7651 6326 7685 6360
rect 7685 6326 7719 6360
rect 7719 6326 7753 6360
rect 7753 6326 7787 6360
rect 7787 6326 7821 6360
rect 7821 6326 7855 6360
rect 7855 6326 7889 6360
rect 7889 6326 7923 6360
rect 7923 6326 7957 6360
rect 7957 6326 7991 6360
rect 7991 6326 8025 6360
rect 8025 6326 8059 6360
rect 8059 6326 8093 6360
rect 8093 6326 8127 6360
rect 8127 6326 8161 6360
rect 8161 6326 8195 6360
rect 8195 6326 8229 6360
rect 8229 6326 8263 6360
rect 8263 6326 8297 6360
rect 8297 6326 8331 6360
rect 8331 6326 8365 6360
rect 8365 6326 8399 6360
rect 8399 6326 8433 6360
rect 8433 6326 8467 6360
rect 8467 6326 8501 6360
rect 8501 6326 8535 6360
rect 8535 6326 8569 6360
rect 8569 6326 8603 6360
rect 8603 6326 8637 6360
rect 8637 6326 8671 6360
rect 8671 6326 8705 6360
rect 8705 6326 8739 6360
rect 8739 6326 8773 6360
rect 8773 6326 8807 6360
rect 8807 6326 8841 6360
rect 8841 6326 8875 6360
rect 8875 6326 8909 6360
rect 8909 6326 8943 6360
rect 8943 6326 8977 6360
rect 8977 6326 9011 6360
rect 9011 6326 9045 6360
rect 9045 6326 9079 6360
rect 9079 6326 9113 6360
rect 9113 6326 9147 6360
rect 9147 6326 9181 6360
rect 9181 6326 9215 6360
rect 9215 6326 9249 6360
rect 9249 6326 9283 6360
rect 9283 6326 9317 6360
rect 9317 6326 9351 6360
rect 9351 6326 9385 6360
rect 9385 6326 9419 6360
rect 9419 6326 9453 6360
rect 9453 6326 9487 6360
rect 9487 6326 9521 6360
rect 9521 6326 9555 6360
rect 9555 6326 9589 6360
rect 9589 6326 9623 6360
rect 9623 6326 9657 6360
rect 9657 6326 9691 6360
rect 9691 6326 9725 6360
rect 9725 6326 9759 6360
rect 9759 6326 9793 6360
rect 9793 6326 9827 6360
rect 9827 6326 9861 6360
rect 9861 6326 9895 6360
rect 9895 6326 9929 6360
rect 9929 6326 9963 6360
rect 9963 6326 9997 6360
rect 9997 6326 10031 6360
rect 10031 6326 10065 6360
rect 10065 6326 10099 6360
rect 10099 6326 10133 6360
rect 10133 6326 10167 6360
rect 10167 6326 10201 6360
rect 10201 6326 10235 6360
rect 10235 6326 10269 6360
rect 10269 6326 10303 6360
rect 10303 6326 10337 6360
rect 10337 6326 10371 6360
rect 10371 6326 10405 6360
rect 10405 6326 10439 6360
rect 10439 6326 10473 6360
rect 10473 6326 10507 6360
rect 10507 6326 10541 6360
rect 10541 6326 10575 6360
rect 10575 6326 10609 6360
rect 10609 6326 10643 6360
rect 10643 6326 10677 6360
rect 10677 6326 10711 6360
rect 10711 6326 10745 6360
rect 10745 6326 10779 6360
rect 10779 6326 10813 6360
rect 10813 6326 10847 6360
rect 10847 6326 10881 6360
rect 10881 6326 10915 6360
rect 10915 6326 10949 6360
rect 10949 6326 10983 6360
rect 10983 6326 11017 6360
rect 11017 6326 11051 6360
rect 11051 6326 11085 6360
rect 11085 6326 11119 6360
rect 11119 6326 11153 6360
rect 11153 6326 11187 6360
rect 11187 6326 11221 6360
rect 11221 6326 11255 6360
rect 11255 6326 11289 6360
rect 11289 6326 11323 6360
rect 11323 6326 11357 6360
rect 11357 6326 11391 6360
rect 11391 6326 11425 6360
rect 11425 6326 11459 6360
rect 11459 6326 11493 6360
rect 11493 6326 11527 6360
rect 11527 6326 11561 6360
rect 11561 6326 11595 6360
rect 11595 6326 11629 6360
rect 11629 6326 11663 6360
rect 11663 6326 11697 6360
rect 11697 6326 11731 6360
rect 11731 6326 11765 6360
rect 11765 6326 11799 6360
rect 11799 6326 11833 6360
rect 11833 6326 11867 6360
rect 11867 6326 11901 6360
rect 11901 6326 11935 6360
rect 11935 6326 11969 6360
rect 11969 6326 12003 6360
rect 12003 6326 12037 6360
rect 12037 6326 12071 6360
rect 12071 6326 12105 6360
rect 12105 6326 12139 6360
rect 12139 6326 12173 6360
rect 12173 6326 12207 6360
rect 12207 6326 12241 6360
rect 12241 6326 12275 6360
rect 12275 6326 12309 6360
rect 12309 6326 12343 6360
rect 12343 6326 12377 6360
rect 12377 6326 12411 6360
rect 12411 6326 12445 6360
rect 12445 6326 12479 6360
rect 12479 6326 12513 6360
rect 12513 6326 12547 6360
rect 12547 6326 12581 6360
rect 12581 6326 12615 6360
rect 12615 6326 12649 6360
rect 12649 6326 12683 6360
rect 12683 6326 12717 6360
rect 12717 6326 12751 6360
rect 12751 6326 12785 6360
rect 12785 6326 12819 6360
rect 12819 6326 12853 6360
rect 12853 6326 12887 6360
rect 12887 6326 12921 6360
rect 12921 6326 12955 6360
rect 12955 6326 12989 6360
rect 12989 6326 13023 6360
rect 13023 6326 13057 6360
rect 13057 6326 13091 6360
rect 13091 6326 13125 6360
rect 13125 6326 13159 6360
rect 13159 6326 13193 6360
rect 13193 6326 13227 6360
rect 13227 6326 13261 6360
rect 13261 6326 13295 6360
rect 13295 6326 13329 6360
rect 13329 6326 13363 6360
rect 13363 6326 13397 6360
rect 13397 6326 13431 6360
rect 13431 6326 13465 6360
rect 13465 6326 13499 6360
rect 13499 6326 13533 6360
rect 13533 6326 13567 6360
rect 13567 6326 13601 6360
rect 13601 6326 13635 6360
rect 13635 6326 13669 6360
rect 13669 6326 13703 6360
rect 13703 6326 13737 6360
rect 13737 6326 13771 6360
rect 13771 6326 13805 6360
rect 13805 6326 13839 6360
rect 13839 6326 13873 6360
rect 13873 6326 13907 6360
rect 13907 6326 13941 6360
rect 13941 6326 13975 6360
rect 13975 6326 14009 6360
rect 14009 6326 14043 6360
rect 14043 6326 14077 6360
rect 14077 6326 14111 6360
rect 14111 6326 14145 6360
rect 14145 6326 14179 6360
rect 14179 6326 14213 6360
rect 14213 6326 14247 6360
rect 14247 6326 14281 6360
rect 14281 6326 14315 6360
rect 14315 6326 14349 6360
rect 14349 6326 14383 6360
rect 14383 6326 14417 6360
rect 14417 6326 14451 6360
rect 14451 6326 14485 6360
rect 14485 6326 14519 6360
rect 14519 6326 14553 6360
rect 14553 6326 14587 6360
rect 14587 6326 14621 6360
rect 14621 6326 14655 6360
rect 14655 6326 14689 6360
rect 14689 6326 14723 6360
rect 14723 6326 14757 6360
rect 14757 6326 14791 6360
rect 14791 6326 14825 6360
rect 14825 6326 14859 6360
rect 14859 6326 14893 6360
rect 14893 6326 14932 6360
rect 14932 6326 14966 6360
rect 14966 6326 15000 6360
rect 15000 6326 15020 6360
rect 15068 6359 15102 6360
rect 68 6286 102 6295
rect 141 6286 175 6295
rect 214 6286 248 6295
rect 287 6286 321 6295
rect 360 6286 394 6295
rect 433 6286 467 6295
rect 506 6286 540 6295
rect 579 6286 613 6295
rect 652 6286 686 6295
rect 725 6286 759 6295
rect 798 6286 832 6295
rect 871 6286 905 6295
rect 944 6286 978 6295
rect 1017 6286 1051 6295
rect 1090 6286 15020 6326
rect 15068 6287 15102 6321
rect 68 6261 102 6286
rect 141 6261 171 6286
rect 171 6261 175 6286
rect 214 6261 240 6286
rect 240 6261 248 6286
rect 287 6261 309 6286
rect 309 6261 321 6286
rect 360 6261 378 6286
rect 378 6261 394 6286
rect 433 6261 447 6286
rect 447 6261 467 6286
rect 506 6261 516 6286
rect 516 6261 540 6286
rect 579 6261 585 6286
rect 585 6261 613 6286
rect 652 6261 654 6286
rect 654 6261 686 6286
rect 725 6261 758 6286
rect 758 6261 759 6286
rect 798 6261 827 6286
rect 827 6261 832 6286
rect 871 6261 896 6286
rect 896 6261 905 6286
rect 944 6261 965 6286
rect 965 6261 978 6286
rect 1017 6261 1034 6286
rect 1034 6261 1051 6286
rect 1090 6252 1103 6286
rect 1103 6252 1137 6286
rect 1137 6252 1172 6286
rect 1172 6252 1206 6286
rect 1206 6252 1241 6286
rect 1241 6252 1275 6286
rect 1275 6252 1310 6286
rect 1310 6252 1344 6286
rect 1344 6252 1379 6286
rect 1379 6252 1413 6286
rect 1413 6252 1448 6286
rect 1448 6252 1482 6286
rect 1482 6252 1517 6286
rect 1517 6252 1551 6286
rect 1551 6252 1586 6286
rect 1586 6252 1620 6286
rect 1620 6252 1655 6286
rect 1655 6252 1689 6286
rect 1689 6252 1724 6286
rect 1724 6252 1758 6286
rect 1758 6252 1793 6286
rect 1793 6252 1827 6286
rect 1827 6252 1862 6286
rect 1862 6252 1896 6286
rect 1896 6252 1931 6286
rect 1931 6252 1965 6286
rect 1965 6252 2000 6286
rect 2000 6252 2034 6286
rect 2034 6252 2069 6286
rect 2069 6252 2103 6286
rect 2103 6252 2138 6286
rect 2138 6252 2172 6286
rect 2172 6252 2207 6286
rect 2207 6252 2241 6286
rect 2241 6252 2276 6286
rect 2276 6252 2310 6286
rect 2310 6252 2345 6286
rect 2345 6252 2379 6286
rect 2379 6252 2414 6286
rect 2414 6252 2448 6286
rect 2448 6252 2483 6286
rect 2483 6252 2517 6286
rect 2517 6252 2551 6286
rect 2551 6252 2585 6286
rect 2585 6252 2619 6286
rect 2619 6252 2653 6286
rect 2653 6252 2687 6286
rect 2687 6252 2721 6286
rect 2721 6252 2755 6286
rect 2755 6252 2789 6286
rect 2789 6252 2823 6286
rect 2823 6252 2857 6286
rect 2857 6252 2891 6286
rect 2891 6252 2925 6286
rect 2925 6252 2959 6286
rect 2959 6252 2993 6286
rect 2993 6252 3027 6286
rect 3027 6252 3061 6286
rect 3061 6252 3095 6286
rect 3095 6252 3129 6286
rect 3129 6252 3163 6286
rect 3163 6252 3197 6286
rect 3197 6252 3231 6286
rect 3231 6252 3265 6286
rect 3265 6252 3299 6286
rect 3299 6252 3333 6286
rect 3333 6252 3367 6286
rect 3367 6252 3401 6286
rect 3401 6252 3435 6286
rect 3435 6252 3469 6286
rect 3469 6252 3503 6286
rect 3503 6252 3537 6286
rect 3537 6252 3571 6286
rect 3571 6252 3605 6286
rect 3605 6252 3639 6286
rect 3639 6252 3673 6286
rect 3673 6252 3707 6286
rect 3707 6252 3741 6286
rect 3741 6252 3775 6286
rect 3775 6252 3809 6286
rect 3809 6252 3843 6286
rect 3843 6252 3877 6286
rect 3877 6252 3911 6286
rect 3911 6252 3945 6286
rect 3945 6252 3979 6286
rect 3979 6252 4013 6286
rect 4013 6252 4047 6286
rect 4047 6252 4081 6286
rect 4081 6252 4115 6286
rect 4115 6252 4149 6286
rect 4149 6252 4183 6286
rect 4183 6252 4217 6286
rect 4217 6252 4251 6286
rect 4251 6252 4285 6286
rect 4285 6252 4319 6286
rect 4319 6252 4353 6286
rect 4353 6252 4387 6286
rect 4387 6252 4421 6286
rect 4421 6252 4455 6286
rect 4455 6252 4489 6286
rect 4489 6252 4523 6286
rect 4523 6252 4557 6286
rect 4557 6252 4591 6286
rect 4591 6252 4625 6286
rect 4625 6252 4659 6286
rect 4659 6252 4693 6286
rect 4693 6252 4727 6286
rect 4727 6252 4761 6286
rect 4761 6252 4795 6286
rect 4795 6252 4829 6286
rect 4829 6252 4863 6286
rect 4863 6252 4897 6286
rect 4897 6252 4931 6286
rect 4931 6252 4965 6286
rect 4965 6252 4999 6286
rect 4999 6252 5033 6286
rect 5033 6252 5067 6286
rect 5067 6252 5101 6286
rect 5101 6252 5135 6286
rect 5135 6252 5169 6286
rect 5169 6252 5203 6286
rect 5203 6252 5237 6286
rect 5237 6252 5271 6286
rect 5271 6252 5305 6286
rect 5305 6252 5339 6286
rect 5339 6252 5373 6286
rect 5373 6252 5407 6286
rect 5407 6252 5441 6286
rect 5441 6252 5475 6286
rect 5475 6252 5509 6286
rect 5509 6252 5543 6286
rect 5543 6252 5577 6286
rect 5577 6252 5611 6286
rect 5611 6252 5645 6286
rect 5645 6252 5679 6286
rect 5679 6252 5713 6286
rect 5713 6252 5747 6286
rect 5747 6252 5781 6286
rect 5781 6252 5815 6286
rect 5815 6252 5849 6286
rect 5849 6252 5883 6286
rect 5883 6252 5917 6286
rect 5917 6252 5951 6286
rect 5951 6252 5985 6286
rect 5985 6252 6019 6286
rect 6019 6252 6053 6286
rect 6053 6252 6087 6286
rect 6087 6252 6121 6286
rect 6121 6252 6155 6286
rect 6155 6252 6189 6286
rect 6189 6252 6223 6286
rect 6223 6252 6257 6286
rect 6257 6252 6291 6286
rect 6291 6252 6325 6286
rect 6325 6252 6359 6286
rect 6359 6252 6393 6286
rect 6393 6252 6427 6286
rect 6427 6252 6461 6286
rect 6461 6252 6495 6286
rect 6495 6252 6529 6286
rect 6529 6252 6563 6286
rect 6563 6252 6597 6286
rect 6597 6252 6631 6286
rect 6631 6252 6665 6286
rect 6665 6252 6699 6286
rect 6699 6252 6733 6286
rect 6733 6252 6767 6286
rect 6767 6252 6801 6286
rect 6801 6252 6835 6286
rect 6835 6252 6869 6286
rect 6869 6252 6903 6286
rect 6903 6252 6937 6286
rect 6937 6252 6971 6286
rect 6971 6252 7005 6286
rect 7005 6252 7039 6286
rect 7039 6252 7073 6286
rect 7073 6252 7107 6286
rect 7107 6252 7141 6286
rect 7141 6252 7175 6286
rect 7175 6252 7209 6286
rect 7209 6252 7243 6286
rect 7243 6252 7277 6286
rect 7277 6252 7311 6286
rect 7311 6252 7345 6286
rect 7345 6252 7379 6286
rect 7379 6252 7413 6286
rect 7413 6252 7447 6286
rect 7447 6252 7481 6286
rect 7481 6252 7515 6286
rect 7515 6252 7549 6286
rect 7549 6252 7583 6286
rect 7583 6252 7617 6286
rect 7617 6252 7651 6286
rect 7651 6252 7685 6286
rect 7685 6252 7719 6286
rect 7719 6252 7753 6286
rect 7753 6252 7787 6286
rect 7787 6252 7821 6286
rect 7821 6252 7855 6286
rect 7855 6252 7889 6286
rect 7889 6252 7923 6286
rect 7923 6252 7957 6286
rect 7957 6252 7991 6286
rect 7991 6252 8025 6286
rect 8025 6252 8059 6286
rect 8059 6252 8093 6286
rect 8093 6252 8127 6286
rect 8127 6252 8161 6286
rect 8161 6252 8195 6286
rect 8195 6252 8229 6286
rect 8229 6252 8263 6286
rect 8263 6252 8297 6286
rect 8297 6252 8331 6286
rect 8331 6252 8365 6286
rect 8365 6252 8399 6286
rect 8399 6252 8433 6286
rect 8433 6252 8467 6286
rect 8467 6252 8501 6286
rect 8501 6252 8535 6286
rect 8535 6252 8569 6286
rect 8569 6252 8603 6286
rect 8603 6252 8637 6286
rect 8637 6252 8671 6286
rect 8671 6252 8705 6286
rect 8705 6252 8739 6286
rect 8739 6252 8773 6286
rect 8773 6252 8807 6286
rect 8807 6252 8841 6286
rect 8841 6252 8875 6286
rect 8875 6252 8909 6286
rect 8909 6252 8943 6286
rect 8943 6252 8977 6286
rect 8977 6252 9011 6286
rect 9011 6252 9045 6286
rect 9045 6252 9079 6286
rect 9079 6252 9113 6286
rect 9113 6252 9147 6286
rect 9147 6252 9181 6286
rect 9181 6252 9215 6286
rect 9215 6252 9249 6286
rect 9249 6252 9283 6286
rect 9283 6252 9317 6286
rect 9317 6252 9351 6286
rect 9351 6252 9385 6286
rect 9385 6252 9419 6286
rect 9419 6252 9453 6286
rect 9453 6252 9487 6286
rect 9487 6252 9521 6286
rect 9521 6252 9555 6286
rect 9555 6252 9589 6286
rect 9589 6252 9623 6286
rect 9623 6252 9657 6286
rect 9657 6252 9691 6286
rect 9691 6252 9725 6286
rect 9725 6252 9759 6286
rect 9759 6252 9793 6286
rect 9793 6252 9827 6286
rect 9827 6252 9861 6286
rect 9861 6252 9895 6286
rect 9895 6252 9929 6286
rect 9929 6252 9963 6286
rect 9963 6252 9997 6286
rect 9997 6252 10031 6286
rect 10031 6252 10065 6286
rect 10065 6252 10099 6286
rect 10099 6252 10133 6286
rect 10133 6252 10167 6286
rect 10167 6252 10201 6286
rect 10201 6252 10235 6286
rect 10235 6252 10269 6286
rect 10269 6252 10303 6286
rect 10303 6252 10337 6286
rect 10337 6252 10371 6286
rect 10371 6252 10405 6286
rect 10405 6252 10439 6286
rect 10439 6252 10473 6286
rect 10473 6252 10507 6286
rect 10507 6252 10541 6286
rect 10541 6252 10575 6286
rect 10575 6252 10609 6286
rect 10609 6252 10643 6286
rect 10643 6252 10677 6286
rect 10677 6252 10711 6286
rect 10711 6252 10745 6286
rect 10745 6252 10779 6286
rect 10779 6252 10813 6286
rect 10813 6252 10847 6286
rect 10847 6252 10881 6286
rect 10881 6252 10915 6286
rect 10915 6252 10949 6286
rect 10949 6252 10983 6286
rect 10983 6252 11017 6286
rect 11017 6252 11051 6286
rect 11051 6252 11085 6286
rect 11085 6252 11119 6286
rect 11119 6252 11153 6286
rect 11153 6252 11187 6286
rect 11187 6252 11221 6286
rect 11221 6252 11255 6286
rect 11255 6252 11289 6286
rect 11289 6252 11323 6286
rect 11323 6252 11357 6286
rect 11357 6252 11391 6286
rect 11391 6252 11425 6286
rect 11425 6252 11459 6286
rect 11459 6252 11493 6286
rect 11493 6252 11527 6286
rect 11527 6252 11561 6286
rect 11561 6252 11595 6286
rect 11595 6252 11629 6286
rect 11629 6252 11663 6286
rect 11663 6252 11697 6286
rect 11697 6252 11731 6286
rect 11731 6252 11765 6286
rect 11765 6252 11799 6286
rect 11799 6252 11833 6286
rect 11833 6252 11867 6286
rect 11867 6252 11901 6286
rect 11901 6252 11935 6286
rect 11935 6252 11969 6286
rect 11969 6252 12003 6286
rect 12003 6252 12037 6286
rect 12037 6252 12071 6286
rect 12071 6252 12105 6286
rect 12105 6252 12139 6286
rect 12139 6252 12173 6286
rect 12173 6252 12207 6286
rect 12207 6252 12241 6286
rect 12241 6252 12275 6286
rect 12275 6252 12309 6286
rect 12309 6252 12343 6286
rect 12343 6252 12377 6286
rect 12377 6252 12411 6286
rect 12411 6252 12445 6286
rect 12445 6252 12479 6286
rect 12479 6252 12513 6286
rect 12513 6252 12547 6286
rect 12547 6252 12581 6286
rect 12581 6252 12615 6286
rect 12615 6252 12649 6286
rect 12649 6252 12683 6286
rect 12683 6252 12717 6286
rect 12717 6252 12751 6286
rect 12751 6252 12785 6286
rect 12785 6252 12819 6286
rect 12819 6252 12853 6286
rect 12853 6252 12887 6286
rect 12887 6252 12921 6286
rect 12921 6252 12955 6286
rect 12955 6252 12989 6286
rect 12989 6252 13023 6286
rect 13023 6252 13057 6286
rect 13057 6252 13091 6286
rect 13091 6252 13125 6286
rect 13125 6252 13159 6286
rect 13159 6252 13193 6286
rect 13193 6252 13227 6286
rect 13227 6252 13261 6286
rect 13261 6252 13295 6286
rect 13295 6252 13329 6286
rect 13329 6252 13363 6286
rect 13363 6252 13397 6286
rect 13397 6252 13431 6286
rect 13431 6252 13465 6286
rect 13465 6252 13499 6286
rect 13499 6252 13533 6286
rect 13533 6252 13567 6286
rect 13567 6252 13601 6286
rect 13601 6252 13635 6286
rect 13635 6252 13669 6286
rect 13669 6252 13703 6286
rect 13703 6252 13737 6286
rect 13737 6252 13771 6286
rect 13771 6252 13805 6286
rect 13805 6252 13839 6286
rect 13839 6252 13873 6286
rect 13873 6252 13907 6286
rect 13907 6252 13941 6286
rect 13941 6252 13975 6286
rect 13975 6252 14009 6286
rect 14009 6252 14043 6286
rect 14043 6252 14077 6286
rect 14077 6252 14111 6286
rect 14111 6252 14145 6286
rect 14145 6252 14179 6286
rect 14179 6252 14213 6286
rect 14213 6252 14247 6286
rect 14247 6252 14281 6286
rect 14281 6252 14315 6286
rect 14315 6252 14349 6286
rect 14349 6252 14383 6286
rect 14383 6252 14417 6286
rect 14417 6252 14451 6286
rect 14451 6252 14485 6286
rect 14485 6252 14519 6286
rect 14519 6252 14553 6286
rect 14553 6252 14587 6286
rect 14587 6252 14621 6286
rect 14621 6252 14655 6286
rect 14655 6252 14689 6286
rect 14689 6252 14723 6286
rect 14723 6252 14757 6286
rect 14757 6252 14791 6286
rect 14791 6252 14825 6286
rect 14825 6252 14859 6286
rect 14859 6252 14893 6286
rect 14893 6285 15020 6286
rect 14893 6252 14932 6285
rect 1090 6251 14932 6252
rect 14932 6251 14966 6285
rect 14966 6251 15000 6285
rect 15000 6251 15020 6285
rect 68 6212 102 6223
rect 141 6212 175 6223
rect 214 6212 248 6223
rect 287 6212 321 6223
rect 360 6212 394 6223
rect 433 6212 467 6223
rect 506 6212 540 6223
rect 579 6212 613 6223
rect 652 6212 686 6223
rect 725 6212 759 6223
rect 798 6212 832 6223
rect 871 6212 905 6223
rect 944 6212 978 6223
rect 1017 6212 1051 6223
rect 1090 6212 15020 6251
rect 15068 6215 15102 6249
rect 68 6189 102 6212
rect 141 6189 171 6212
rect 171 6189 175 6212
rect 214 6189 240 6212
rect 240 6189 248 6212
rect 287 6189 309 6212
rect 309 6189 321 6212
rect 360 6189 378 6212
rect 378 6189 394 6212
rect 433 6189 447 6212
rect 447 6189 467 6212
rect 506 6189 516 6212
rect 516 6189 540 6212
rect 579 6189 585 6212
rect 585 6189 613 6212
rect 652 6189 654 6212
rect 654 6189 686 6212
rect 725 6189 758 6212
rect 758 6189 759 6212
rect 798 6189 827 6212
rect 827 6189 832 6212
rect 871 6189 896 6212
rect 896 6189 905 6212
rect 944 6189 965 6212
rect 965 6189 978 6212
rect 1017 6189 1034 6212
rect 1034 6189 1051 6212
rect 1090 6178 1103 6212
rect 1103 6178 1137 6212
rect 1137 6178 1172 6212
rect 1172 6178 1206 6212
rect 1206 6178 1241 6212
rect 1241 6178 1275 6212
rect 1275 6178 1310 6212
rect 1310 6178 1344 6212
rect 1344 6178 1379 6212
rect 1379 6178 1413 6212
rect 1413 6178 1448 6212
rect 1448 6178 1482 6212
rect 1482 6178 1517 6212
rect 1517 6178 1551 6212
rect 1551 6178 1586 6212
rect 1586 6178 1620 6212
rect 1620 6178 1655 6212
rect 1655 6178 1689 6212
rect 1689 6178 1724 6212
rect 1724 6178 1758 6212
rect 1758 6178 1793 6212
rect 1793 6178 1827 6212
rect 1827 6178 1862 6212
rect 1862 6178 1896 6212
rect 1896 6178 1931 6212
rect 1931 6178 1965 6212
rect 1965 6178 2000 6212
rect 2000 6178 2034 6212
rect 2034 6178 2069 6212
rect 2069 6178 2103 6212
rect 2103 6178 2138 6212
rect 2138 6178 2172 6212
rect 2172 6178 2207 6212
rect 2207 6178 2241 6212
rect 2241 6178 2276 6212
rect 2276 6178 2310 6212
rect 2310 6178 2345 6212
rect 2345 6178 2379 6212
rect 2379 6178 2414 6212
rect 2414 6178 2448 6212
rect 2448 6178 2483 6212
rect 2483 6178 2517 6212
rect 2517 6178 2551 6212
rect 2551 6178 2585 6212
rect 2585 6178 2619 6212
rect 2619 6178 2653 6212
rect 2653 6178 2687 6212
rect 2687 6178 2721 6212
rect 2721 6178 2755 6212
rect 2755 6178 2789 6212
rect 2789 6178 2823 6212
rect 2823 6178 2857 6212
rect 2857 6178 2891 6212
rect 2891 6178 2925 6212
rect 2925 6178 2959 6212
rect 2959 6178 2993 6212
rect 2993 6178 3027 6212
rect 3027 6178 3061 6212
rect 3061 6178 3095 6212
rect 3095 6178 3129 6212
rect 3129 6178 3163 6212
rect 3163 6178 3197 6212
rect 3197 6178 3231 6212
rect 3231 6178 3265 6212
rect 3265 6178 3299 6212
rect 3299 6178 3333 6212
rect 3333 6178 3367 6212
rect 3367 6178 3401 6212
rect 3401 6178 3435 6212
rect 3435 6178 3469 6212
rect 3469 6178 3503 6212
rect 3503 6178 3537 6212
rect 3537 6178 3571 6212
rect 3571 6178 3605 6212
rect 3605 6178 3639 6212
rect 3639 6178 3673 6212
rect 3673 6178 3707 6212
rect 3707 6178 3741 6212
rect 3741 6178 3775 6212
rect 3775 6178 3809 6212
rect 3809 6178 3843 6212
rect 3843 6178 3877 6212
rect 3877 6178 3911 6212
rect 3911 6178 3945 6212
rect 3945 6178 3979 6212
rect 3979 6178 4013 6212
rect 4013 6178 4047 6212
rect 4047 6178 4081 6212
rect 4081 6178 4115 6212
rect 4115 6178 4149 6212
rect 4149 6178 4183 6212
rect 4183 6178 4217 6212
rect 4217 6178 4251 6212
rect 4251 6178 4285 6212
rect 4285 6178 4319 6212
rect 4319 6178 4353 6212
rect 4353 6178 4387 6212
rect 4387 6178 4421 6212
rect 4421 6178 4455 6212
rect 4455 6178 4489 6212
rect 4489 6178 4523 6212
rect 4523 6178 4557 6212
rect 4557 6178 4591 6212
rect 4591 6178 4625 6212
rect 4625 6178 4659 6212
rect 4659 6178 4693 6212
rect 4693 6178 4727 6212
rect 4727 6178 4761 6212
rect 4761 6178 4795 6212
rect 4795 6178 4829 6212
rect 4829 6178 4863 6212
rect 4863 6178 4897 6212
rect 4897 6178 4931 6212
rect 4931 6178 4965 6212
rect 4965 6178 4999 6212
rect 4999 6178 5033 6212
rect 5033 6178 5067 6212
rect 5067 6178 5101 6212
rect 5101 6178 5135 6212
rect 5135 6178 5169 6212
rect 5169 6178 5203 6212
rect 5203 6178 5237 6212
rect 5237 6178 5271 6212
rect 5271 6178 5305 6212
rect 5305 6178 5339 6212
rect 5339 6178 5373 6212
rect 5373 6178 5407 6212
rect 5407 6178 5441 6212
rect 5441 6178 5475 6212
rect 5475 6178 5509 6212
rect 5509 6178 5543 6212
rect 5543 6178 5577 6212
rect 5577 6178 5611 6212
rect 5611 6178 5645 6212
rect 5645 6178 5679 6212
rect 5679 6178 5713 6212
rect 5713 6178 5747 6212
rect 5747 6178 5781 6212
rect 5781 6178 5815 6212
rect 5815 6178 5849 6212
rect 5849 6178 5883 6212
rect 5883 6178 5917 6212
rect 5917 6178 5951 6212
rect 5951 6178 5985 6212
rect 5985 6178 6019 6212
rect 6019 6178 6053 6212
rect 6053 6178 6087 6212
rect 6087 6178 6121 6212
rect 6121 6178 6155 6212
rect 6155 6178 6189 6212
rect 6189 6178 6223 6212
rect 6223 6178 6257 6212
rect 6257 6178 6291 6212
rect 6291 6178 6325 6212
rect 6325 6178 6359 6212
rect 6359 6178 6393 6212
rect 6393 6178 6427 6212
rect 6427 6178 6461 6212
rect 6461 6178 6495 6212
rect 6495 6178 6529 6212
rect 6529 6178 6563 6212
rect 6563 6178 6597 6212
rect 6597 6178 6631 6212
rect 6631 6178 6665 6212
rect 6665 6178 6699 6212
rect 6699 6178 6733 6212
rect 6733 6178 6767 6212
rect 6767 6178 6801 6212
rect 6801 6178 6835 6212
rect 6835 6178 6869 6212
rect 6869 6178 6903 6212
rect 6903 6178 6937 6212
rect 6937 6178 6971 6212
rect 6971 6178 7005 6212
rect 7005 6178 7039 6212
rect 7039 6178 7073 6212
rect 7073 6178 7107 6212
rect 7107 6178 7141 6212
rect 7141 6178 7175 6212
rect 7175 6178 7209 6212
rect 7209 6178 7243 6212
rect 7243 6178 7277 6212
rect 7277 6178 7311 6212
rect 7311 6178 7345 6212
rect 7345 6178 7379 6212
rect 7379 6178 7413 6212
rect 7413 6178 7447 6212
rect 7447 6178 7481 6212
rect 7481 6178 7515 6212
rect 7515 6178 7549 6212
rect 7549 6178 7583 6212
rect 7583 6178 7617 6212
rect 7617 6178 7651 6212
rect 7651 6178 7685 6212
rect 7685 6178 7719 6212
rect 7719 6178 7753 6212
rect 7753 6178 7787 6212
rect 7787 6178 7821 6212
rect 7821 6178 7855 6212
rect 7855 6178 7889 6212
rect 7889 6178 7923 6212
rect 7923 6178 7957 6212
rect 7957 6178 7991 6212
rect 7991 6178 8025 6212
rect 8025 6178 8059 6212
rect 8059 6178 8093 6212
rect 8093 6178 8127 6212
rect 8127 6178 8161 6212
rect 8161 6178 8195 6212
rect 8195 6178 8229 6212
rect 8229 6178 8263 6212
rect 8263 6178 8297 6212
rect 8297 6178 8331 6212
rect 8331 6178 8365 6212
rect 8365 6178 8399 6212
rect 8399 6178 8433 6212
rect 8433 6178 8467 6212
rect 8467 6178 8501 6212
rect 8501 6178 8535 6212
rect 8535 6178 8569 6212
rect 8569 6178 8603 6212
rect 8603 6178 8637 6212
rect 8637 6178 8671 6212
rect 8671 6178 8705 6212
rect 8705 6178 8739 6212
rect 8739 6178 8773 6212
rect 8773 6178 8807 6212
rect 8807 6178 8841 6212
rect 8841 6178 8875 6212
rect 8875 6178 8909 6212
rect 8909 6178 8943 6212
rect 8943 6178 8977 6212
rect 8977 6178 9011 6212
rect 9011 6178 9045 6212
rect 9045 6178 9079 6212
rect 9079 6178 9113 6212
rect 9113 6178 9147 6212
rect 9147 6178 9181 6212
rect 9181 6178 9215 6212
rect 9215 6178 9249 6212
rect 9249 6178 9283 6212
rect 9283 6178 9317 6212
rect 9317 6178 9351 6212
rect 9351 6178 9385 6212
rect 9385 6178 9419 6212
rect 9419 6178 9453 6212
rect 9453 6178 9487 6212
rect 9487 6178 9521 6212
rect 9521 6178 9555 6212
rect 9555 6178 9589 6212
rect 9589 6178 9623 6212
rect 9623 6178 9657 6212
rect 9657 6178 9691 6212
rect 9691 6178 9725 6212
rect 9725 6178 9759 6212
rect 9759 6178 9793 6212
rect 9793 6178 9827 6212
rect 9827 6178 9861 6212
rect 9861 6178 9895 6212
rect 9895 6178 9929 6212
rect 9929 6178 9963 6212
rect 9963 6178 9997 6212
rect 9997 6178 10031 6212
rect 10031 6178 10065 6212
rect 10065 6178 10099 6212
rect 10099 6178 10133 6212
rect 10133 6178 10167 6212
rect 10167 6178 10201 6212
rect 10201 6178 10235 6212
rect 10235 6178 10269 6212
rect 10269 6178 10303 6212
rect 10303 6178 10337 6212
rect 10337 6178 10371 6212
rect 10371 6178 10405 6212
rect 10405 6178 10439 6212
rect 10439 6178 10473 6212
rect 10473 6178 10507 6212
rect 10507 6178 10541 6212
rect 10541 6178 10575 6212
rect 10575 6178 10609 6212
rect 10609 6178 10643 6212
rect 10643 6178 10677 6212
rect 10677 6178 10711 6212
rect 10711 6178 10745 6212
rect 10745 6178 10779 6212
rect 10779 6178 10813 6212
rect 10813 6178 10847 6212
rect 10847 6178 10881 6212
rect 10881 6178 10915 6212
rect 10915 6178 10949 6212
rect 10949 6178 10983 6212
rect 10983 6178 11017 6212
rect 11017 6178 11051 6212
rect 11051 6178 11085 6212
rect 11085 6178 11119 6212
rect 11119 6178 11153 6212
rect 11153 6178 11187 6212
rect 11187 6178 11221 6212
rect 11221 6178 11255 6212
rect 11255 6178 11289 6212
rect 11289 6178 11323 6212
rect 11323 6178 11357 6212
rect 11357 6178 11391 6212
rect 11391 6178 11425 6212
rect 11425 6178 11459 6212
rect 11459 6178 11493 6212
rect 11493 6178 11527 6212
rect 11527 6178 11561 6212
rect 11561 6178 11595 6212
rect 11595 6178 11629 6212
rect 11629 6178 11663 6212
rect 11663 6178 11697 6212
rect 11697 6178 11731 6212
rect 11731 6178 11765 6212
rect 11765 6178 11799 6212
rect 11799 6178 11833 6212
rect 11833 6178 11867 6212
rect 11867 6178 11901 6212
rect 11901 6178 11935 6212
rect 11935 6178 11969 6212
rect 11969 6178 12003 6212
rect 12003 6178 12037 6212
rect 12037 6178 12071 6212
rect 12071 6178 12105 6212
rect 12105 6178 12139 6212
rect 12139 6178 12173 6212
rect 12173 6178 12207 6212
rect 12207 6178 12241 6212
rect 12241 6178 12275 6212
rect 12275 6178 12309 6212
rect 12309 6178 12343 6212
rect 12343 6178 12377 6212
rect 12377 6178 12411 6212
rect 12411 6178 12445 6212
rect 12445 6178 12479 6212
rect 12479 6178 12513 6212
rect 12513 6178 12547 6212
rect 12547 6178 12581 6212
rect 12581 6178 12615 6212
rect 12615 6178 12649 6212
rect 12649 6178 12683 6212
rect 12683 6178 12717 6212
rect 12717 6178 12751 6212
rect 12751 6178 12785 6212
rect 12785 6178 12819 6212
rect 12819 6178 12853 6212
rect 12853 6178 12887 6212
rect 12887 6178 12921 6212
rect 12921 6178 12955 6212
rect 12955 6178 12989 6212
rect 12989 6178 13023 6212
rect 13023 6178 13057 6212
rect 13057 6178 13091 6212
rect 13091 6178 13125 6212
rect 13125 6178 13159 6212
rect 13159 6178 13193 6212
rect 13193 6178 13227 6212
rect 13227 6178 13261 6212
rect 13261 6178 13295 6212
rect 13295 6178 13329 6212
rect 13329 6178 13363 6212
rect 13363 6178 13397 6212
rect 13397 6178 13431 6212
rect 13431 6178 13465 6212
rect 13465 6178 13499 6212
rect 13499 6178 13533 6212
rect 13533 6178 13567 6212
rect 13567 6178 13601 6212
rect 13601 6178 13635 6212
rect 13635 6178 13669 6212
rect 13669 6178 13703 6212
rect 13703 6178 13737 6212
rect 13737 6178 13771 6212
rect 13771 6178 13805 6212
rect 13805 6178 13839 6212
rect 13839 6178 13873 6212
rect 13873 6178 13907 6212
rect 13907 6178 13941 6212
rect 13941 6178 13975 6212
rect 13975 6178 14009 6212
rect 14009 6178 14043 6212
rect 14043 6178 14077 6212
rect 14077 6178 14111 6212
rect 14111 6178 14145 6212
rect 14145 6178 14179 6212
rect 14179 6178 14213 6212
rect 14213 6178 14247 6212
rect 14247 6178 14281 6212
rect 14281 6178 14315 6212
rect 14315 6178 14349 6212
rect 14349 6178 14383 6212
rect 14383 6178 14417 6212
rect 14417 6178 14451 6212
rect 14451 6178 14485 6212
rect 14485 6178 14519 6212
rect 14519 6178 14553 6212
rect 14553 6178 14587 6212
rect 14587 6178 14621 6212
rect 14621 6178 14655 6212
rect 14655 6178 14689 6212
rect 14689 6178 14723 6212
rect 14723 6178 14757 6212
rect 14757 6178 14791 6212
rect 14791 6178 14825 6212
rect 14825 6178 14859 6212
rect 14859 6178 14893 6212
rect 14893 6210 15020 6212
rect 14893 6178 14932 6210
rect 1090 6176 14932 6178
rect 14932 6176 14966 6210
rect 14966 6176 15000 6210
rect 15000 6176 15020 6210
rect 15068 6176 15102 6177
rect 68 6138 102 6151
rect 141 6138 175 6151
rect 214 6138 248 6151
rect 287 6138 321 6151
rect 360 6138 394 6151
rect 433 6138 467 6151
rect 506 6138 540 6151
rect 579 6138 613 6151
rect 652 6138 686 6151
rect 725 6138 759 6151
rect 798 6138 832 6151
rect 871 6138 905 6151
rect 944 6138 978 6151
rect 1017 6138 1051 6151
rect 1090 6138 15020 6176
rect 15068 6143 15102 6176
rect 68 6117 102 6138
rect 141 6117 171 6138
rect 171 6117 175 6138
rect 214 6117 240 6138
rect 240 6117 248 6138
rect 287 6117 309 6138
rect 309 6117 321 6138
rect 360 6117 378 6138
rect 378 6117 394 6138
rect 433 6117 447 6138
rect 447 6117 467 6138
rect 506 6117 516 6138
rect 516 6117 540 6138
rect 579 6117 585 6138
rect 585 6117 613 6138
rect 652 6117 654 6138
rect 654 6117 686 6138
rect 725 6117 758 6138
rect 758 6117 759 6138
rect 798 6117 827 6138
rect 827 6117 832 6138
rect 871 6117 896 6138
rect 896 6117 905 6138
rect 944 6117 965 6138
rect 965 6117 978 6138
rect 1017 6117 1034 6138
rect 1034 6117 1051 6138
rect 1090 6117 1103 6138
rect 1103 6117 1137 6138
rect 1137 6117 1172 6138
rect 1172 6117 1206 6138
rect 1206 6117 1241 6138
rect 1241 6117 1275 6138
rect 1275 6117 1310 6138
rect 1310 6117 1344 6138
rect 1344 6117 1379 6138
rect 1379 6117 1413 6138
rect 1413 6117 1448 6138
rect 1448 6117 1482 6138
rect 1482 6117 1517 6138
rect 1517 6117 1551 6138
rect 1551 6117 1586 6138
rect 1586 6117 1620 6138
rect 1620 6117 1655 6138
rect 1655 6117 1689 6138
rect 1689 6117 1724 6138
rect 1724 6117 1758 6138
rect 1758 6117 1793 6138
rect 1793 6117 1827 6138
rect 1827 6117 1862 6138
rect 1862 6117 1896 6138
rect 1896 6117 1931 6138
rect 1931 6117 1965 6138
rect 1965 6117 2000 6138
rect 2000 6117 2034 6138
rect 2034 6117 2069 6138
rect 2069 6117 2103 6138
rect 2103 6117 2138 6138
rect 2138 6117 2172 6138
rect 2172 6117 2207 6138
rect 2207 6117 2241 6138
rect 2241 6117 2276 6138
rect 2276 6117 2310 6138
rect 2310 6117 2345 6138
rect 2345 6117 2379 6138
rect 2379 6117 2414 6138
rect 2414 6117 2448 6138
rect 2448 6117 2483 6138
rect 2483 6117 2517 6138
rect 2517 6117 2551 6138
rect 2551 6117 2585 6138
rect 2585 6117 2619 6138
rect 2619 6117 2653 6138
rect 2653 6117 2687 6138
rect 2687 6117 2721 6138
rect 2721 6117 2755 6138
rect 2755 6117 2789 6138
rect 2789 6117 2823 6138
rect 2823 6117 2857 6138
rect 2857 6117 2891 6138
rect 2891 6117 2925 6138
rect 2925 6117 2959 6138
rect 2959 6117 2993 6138
rect 2993 6117 3027 6138
rect 3027 6117 3061 6138
rect 3061 6117 3095 6138
rect 3095 6117 3129 6138
rect 3129 6117 3163 6138
rect 3163 6117 3197 6138
rect 3197 6117 3231 6138
rect 3231 6117 3265 6138
rect 3265 6117 3299 6138
rect 3299 6117 3333 6138
rect 3333 6117 3367 6138
rect 3367 6117 3401 6138
rect 3401 6117 3435 6138
rect 3435 6117 3469 6138
rect 3469 6117 3503 6138
rect 3503 6117 3537 6138
rect 3537 6117 3571 6138
rect 3571 6117 3605 6138
rect 3605 6117 3639 6138
rect 3639 6117 3673 6138
rect 3673 6117 3707 6138
rect 3707 6117 3741 6138
rect 3741 6117 3775 6138
rect 3775 6117 3809 6138
rect 3809 6117 3843 6138
rect 3843 6117 3877 6138
rect 3877 6117 3911 6138
rect 3911 6117 3945 6138
rect 3945 6117 3979 6138
rect 3979 6117 4013 6138
rect 4013 6117 4047 6138
rect 4047 6117 4081 6138
rect 4081 6117 4115 6138
rect 4115 6117 4149 6138
rect 4149 6117 4183 6138
rect 4183 6117 4217 6138
rect 4217 6117 4251 6138
rect 4251 6117 4285 6138
rect 4285 6117 4319 6138
rect 4319 6117 4353 6138
rect 4353 6117 4387 6138
rect 4387 6117 4421 6138
rect 4421 6117 4455 6138
rect 4455 6117 4489 6138
rect 4489 6117 4523 6138
rect 4523 6117 4557 6138
rect 4557 6117 4591 6138
rect 4591 6117 4625 6138
rect 4625 6117 4659 6138
rect 4659 6117 4693 6138
rect 4693 6117 4727 6138
rect 4727 6117 4761 6138
rect 4761 6117 4795 6138
rect 4795 6117 4829 6138
rect 4829 6117 4863 6138
rect 4863 6117 4897 6138
rect 4897 6117 4931 6138
rect 4931 6117 4965 6138
rect 4965 6117 4999 6138
rect 4999 6117 5033 6138
rect 5033 6117 5067 6138
rect 5067 6117 5101 6138
rect 5101 6117 5135 6138
rect 5135 6117 5169 6138
rect 5169 6117 5203 6138
rect 5203 6117 5237 6138
rect 5237 6117 5271 6138
rect 5271 6117 5305 6138
rect 5305 6117 5339 6138
rect 5339 6117 5373 6138
rect 5373 6117 5407 6138
rect 5407 6117 5441 6138
rect 5441 6117 5475 6138
rect 5475 6117 5509 6138
rect 5509 6117 5543 6138
rect 5543 6117 5577 6138
rect 5577 6117 5611 6138
rect 5611 6117 5645 6138
rect 5645 6117 5679 6138
rect 5679 6117 5713 6138
rect 5713 6117 5747 6138
rect 5747 6117 5781 6138
rect 5781 6117 5815 6138
rect 5815 6117 5849 6138
rect 5849 6117 5883 6138
rect 5883 6117 5917 6138
rect 5917 6117 5951 6138
rect 5951 6117 5985 6138
rect 5985 6117 6019 6138
rect 6019 6117 6053 6138
rect 6053 6117 6087 6138
rect 6087 6117 6121 6138
rect 6121 6117 6155 6138
rect 6155 6117 6189 6138
rect 6189 6117 6223 6138
rect 6223 6117 6257 6138
rect 6257 6117 6291 6138
rect 6291 6117 6325 6138
rect 6325 6117 6359 6138
rect 6359 6117 6393 6138
rect 6393 6117 6427 6138
rect 6427 6117 6461 6138
rect 6461 6117 6495 6138
rect 6495 6117 6529 6138
rect 6529 6117 6563 6138
rect 6563 6117 6597 6138
rect 6597 6117 6631 6138
rect 6631 6117 6665 6138
rect 6665 6117 6699 6138
rect 6699 6117 6733 6138
rect 6733 6117 6767 6138
rect 6767 6117 6801 6138
rect 6801 6117 6835 6138
rect 6835 6117 6869 6138
rect 6869 6117 6903 6138
rect 6903 6117 6937 6138
rect 6937 6117 6971 6138
rect 6971 6117 7005 6138
rect 7005 6117 7039 6138
rect 7039 6117 7073 6138
rect 7073 6117 7107 6138
rect 7107 6117 7141 6138
rect 7141 6117 7175 6138
rect 7175 6117 7209 6138
rect 7209 6117 7243 6138
rect 7243 6117 7277 6138
rect 7277 6117 7311 6138
rect 7311 6117 7345 6138
rect 7345 6117 7379 6138
rect 7379 6117 7413 6138
rect 7413 6117 7447 6138
rect 7447 6117 7481 6138
rect 7481 6117 7515 6138
rect 7515 6117 7549 6138
rect 7549 6117 7583 6138
rect 7583 6117 7617 6138
rect 7617 6117 7651 6138
rect 7651 6117 7685 6138
rect 7685 6117 7719 6138
rect 7719 6117 7753 6138
rect 7753 6117 7787 6138
rect 7787 6117 7821 6138
rect 7821 6117 7855 6138
rect 7855 6117 7889 6138
rect 7889 6117 7923 6138
rect 7923 6117 7957 6138
rect 7957 6117 7991 6138
rect 7991 6117 8025 6138
rect 8025 6117 8059 6138
rect 8059 6117 8093 6138
rect 8093 6117 8127 6138
rect 8127 6117 8161 6138
rect 8161 6117 8195 6138
rect 8195 6117 8229 6138
rect 8229 6117 8263 6138
rect 8263 6117 8297 6138
rect 8297 6117 8331 6138
rect 8331 6117 8365 6138
rect 8365 6117 8399 6138
rect 8399 6117 8433 6138
rect 8433 6117 8467 6138
rect 8467 6117 8501 6138
rect 8501 6117 8535 6138
rect 8535 6117 8569 6138
rect 8569 6117 8603 6138
rect 8603 6117 8637 6138
rect 8637 6117 8671 6138
rect 8671 6117 8705 6138
rect 8705 6117 8739 6138
rect 8739 6117 8773 6138
rect 8773 6117 8807 6138
rect 8807 6117 8841 6138
rect 8841 6117 8875 6138
rect 8875 6117 8909 6138
rect 8909 6117 8943 6138
rect 8943 6117 8977 6138
rect 8977 6117 9011 6138
rect 9011 6117 9045 6138
rect 9045 6117 9079 6138
rect 9079 6117 9113 6138
rect 9113 6117 9147 6138
rect 9147 6117 9181 6138
rect 9181 6117 9215 6138
rect 9215 6117 9249 6138
rect 9249 6117 9283 6138
rect 9283 6117 9317 6138
rect 9317 6117 9351 6138
rect 9351 6117 9385 6138
rect 9385 6117 9419 6138
rect 9419 6117 9453 6138
rect 9453 6117 9487 6138
rect 9487 6117 9521 6138
rect 9521 6117 9555 6138
rect 9555 6117 9589 6138
rect 9589 6117 9623 6138
rect 9623 6117 9657 6138
rect 9657 6117 9691 6138
rect 9691 6117 9725 6138
rect 9725 6117 9759 6138
rect 9759 6117 9793 6138
rect 9793 6117 9827 6138
rect 9827 6117 9861 6138
rect 9861 6117 9895 6138
rect 9895 6117 9929 6138
rect 9929 6117 9963 6138
rect 9963 6117 9997 6138
rect 9997 6117 10031 6138
rect 10031 6117 10065 6138
rect 10065 6117 10099 6138
rect 10099 6117 10133 6138
rect 10133 6117 10167 6138
rect 10167 6117 10201 6138
rect 10201 6117 10235 6138
rect 10235 6117 10269 6138
rect 10269 6117 10303 6138
rect 10303 6117 10337 6138
rect 10337 6117 10371 6138
rect 10371 6117 10405 6138
rect 10405 6117 10439 6138
rect 10439 6117 10473 6138
rect 10473 6117 10507 6138
rect 10507 6117 10541 6138
rect 10541 6117 10575 6138
rect 10575 6117 10609 6138
rect 10609 6117 10643 6138
rect 10643 6117 10677 6138
rect 10677 6117 10711 6138
rect 10711 6117 10745 6138
rect 10745 6117 10779 6138
rect 10779 6117 10813 6138
rect 10813 6117 10847 6138
rect 10847 6117 10881 6138
rect 10881 6117 10915 6138
rect 10915 6117 10949 6138
rect 10949 6117 10983 6138
rect 10983 6117 11017 6138
rect 11017 6117 11051 6138
rect 11051 6117 11085 6138
rect 11085 6117 11119 6138
rect 11119 6117 11153 6138
rect 11153 6117 11187 6138
rect 11187 6117 11221 6138
rect 11221 6117 11255 6138
rect 11255 6117 11289 6138
rect 11289 6117 11323 6138
rect 11323 6117 11357 6138
rect 11357 6117 11391 6138
rect 11391 6117 11425 6138
rect 11425 6117 11459 6138
rect 11459 6117 11493 6138
rect 11493 6117 11527 6138
rect 11527 6117 11561 6138
rect 11561 6117 11595 6138
rect 11595 6117 11629 6138
rect 11629 6117 11663 6138
rect 11663 6117 11697 6138
rect 11697 6117 11731 6138
rect 11731 6117 11765 6138
rect 11765 6117 11799 6138
rect 11799 6117 11833 6138
rect 11833 6117 11867 6138
rect 11867 6117 11901 6138
rect 11901 6117 11935 6138
rect 11935 6117 11969 6138
rect 11969 6117 12003 6138
rect 12003 6117 12037 6138
rect 12037 6117 12071 6138
rect 12071 6117 12105 6138
rect 12105 6117 12139 6138
rect 12139 6117 12173 6138
rect 12173 6117 12207 6138
rect 12207 6117 12241 6138
rect 12241 6117 12275 6138
rect 12275 6117 12309 6138
rect 12309 6117 12343 6138
rect 12343 6117 12377 6138
rect 12377 6117 12411 6138
rect 12411 6117 12445 6138
rect 12445 6117 12479 6138
rect 12479 6117 12513 6138
rect 12513 6117 12547 6138
rect 12547 6117 12581 6138
rect 12581 6117 12615 6138
rect 12615 6117 12649 6138
rect 12649 6117 12683 6138
rect 12683 6117 12717 6138
rect 12717 6117 12751 6138
rect 12751 6117 12785 6138
rect 12785 6117 12819 6138
rect 12819 6117 12853 6138
rect 12853 6117 12887 6138
rect 12887 6117 12921 6138
rect 12921 6117 12955 6138
rect 12955 6117 12989 6138
rect 12989 6117 13023 6138
rect 13023 6117 13057 6138
rect 13057 6117 13091 6138
rect 13091 6117 13125 6138
rect 13125 6117 13159 6138
rect 13159 6117 13193 6138
rect 13193 6117 13227 6138
rect 13227 6117 13261 6138
rect 13261 6117 13295 6138
rect 13295 6117 13329 6138
rect 13329 6117 13363 6138
rect 13363 6117 13397 6138
rect 13397 6117 13431 6138
rect 13431 6117 13465 6138
rect 13465 6117 13499 6138
rect 13499 6117 13533 6138
rect 13533 6117 13567 6138
rect 13567 6117 13601 6138
rect 13601 6117 13635 6138
rect 13635 6117 13669 6138
rect 13669 6117 13703 6138
rect 13703 6117 13737 6138
rect 13737 6117 13771 6138
rect 13771 6117 13805 6138
rect 13805 6117 13839 6138
rect 13839 6117 13873 6138
rect 13873 6117 13907 6138
rect 13907 6117 13941 6138
rect 13941 6117 13975 6138
rect 13975 6117 14009 6138
rect 14009 6117 14043 6138
rect 14043 6117 14077 6138
rect 14077 6117 14111 6138
rect 14111 6117 14145 6138
rect 14145 6117 14179 6138
rect 14179 6117 14213 6138
rect 14213 6117 14247 6138
rect 14247 6117 14281 6138
rect 14281 6117 14315 6138
rect 14315 6117 14349 6138
rect 14349 6117 14383 6138
rect 14383 6117 14417 6138
rect 14417 6117 14451 6138
rect 14451 6117 14485 6138
rect 14485 6117 14519 6138
rect 14519 6117 14553 6138
rect 14553 6117 14587 6138
rect 14587 6117 14621 6138
rect 14621 6117 14655 6138
rect 14655 6117 14689 6138
rect 14689 6117 14723 6138
rect 14723 6117 14757 6138
rect 14757 6117 14791 6138
rect 14791 6117 14825 6138
rect 14825 6117 14859 6138
rect 14859 6117 14893 6138
rect 14893 6135 15020 6138
rect 14893 6117 14932 6135
rect 14932 6117 14966 6135
rect 14966 6117 15000 6135
rect 15000 6117 15020 6135
rect 15068 6101 15102 6105
rect 15068 6071 15102 6101
rect 15068 6026 15102 6033
rect 15068 5999 15102 6026
rect 15068 5954 15102 5961
rect 15068 5927 15102 5954
rect 15068 5855 15102 5889
rect 15068 5783 15102 5817
rect 15068 5711 15102 5745
rect 15068 5639 15102 5673
rect 15068 5567 15102 5601
rect 15068 5495 15102 5529
rect 15068 5423 15102 5457
rect 15068 5351 15102 5385
rect 15068 5279 15102 5313
rect 15068 5207 15102 5241
rect 15068 5135 15102 5169
rect 15068 5063 15102 5097
rect 15068 4991 15102 5025
rect 15068 4919 15102 4953
rect 15068 4847 15102 4881
rect 15068 4775 15102 4809
rect 15068 4703 15102 4737
rect 15068 4631 15102 4665
rect 15068 4559 15102 4593
rect 15068 4490 15102 4521
rect 15068 4487 15102 4490
rect 15068 4421 15102 4449
rect 15068 4415 15102 4421
rect 15068 4352 15102 4377
rect 15068 4343 15102 4352
rect 15068 4283 15102 4305
rect 15068 4271 15102 4283
rect 15068 4214 15102 4233
rect 15068 4199 15102 4214
rect 15068 4145 15102 4161
rect 15068 4127 15102 4145
rect 15068 4076 15102 4089
rect 15068 4055 15102 4076
rect 15068 4007 15102 4017
rect 15068 3983 15102 4007
rect 15068 3938 15102 3945
rect 15068 3911 15102 3938
rect 15068 3869 15102 3873
rect 15068 3839 15102 3869
rect 15068 3800 15102 3801
rect 15068 3767 15102 3800
rect 15068 3696 15102 3729
rect 15068 3695 15102 3696
rect 15068 3627 15102 3657
rect 15068 3623 15102 3627
rect 15068 3558 15102 3585
rect 15068 3551 15102 3558
rect 15068 3489 15102 3513
rect 15068 3479 15102 3489
rect 15068 3420 15102 3441
rect 15068 3407 15102 3420
rect 15068 3351 15102 3369
rect 15068 3335 15102 3351
rect 15068 3282 15102 3297
rect 15068 3263 15102 3282
rect 15068 3213 15102 3225
rect 15068 3191 15102 3213
rect 15068 3144 15102 3153
rect 15068 3119 15102 3144
rect 15068 3075 15102 3081
rect 15068 3047 15102 3075
rect 15068 3006 15102 3009
rect 15068 2975 15102 3006
rect 15068 2903 15102 2937
rect 15068 2834 15102 2865
rect 15068 2831 15102 2834
rect 15068 2765 15102 2793
rect 15068 2759 15102 2765
rect 15068 2696 15102 2721
rect 15068 2687 15102 2696
rect 15068 2627 15102 2649
rect 15068 2615 15102 2627
rect 15068 2558 15102 2577
rect 15068 2543 15102 2558
rect 15068 2489 15102 2505
rect 15068 2471 15102 2489
rect 15068 2420 15102 2433
rect 15068 2399 15102 2420
rect 15068 2351 15102 2361
rect 15068 2327 15102 2351
rect 15068 2282 15102 2289
rect 15068 2255 15102 2282
rect 15068 2213 15102 2217
rect 15068 2183 15102 2213
rect 15068 2144 15102 2145
rect 15068 2111 15102 2144
rect 15068 2040 15102 2073
rect 15068 2039 15102 2040
rect 15068 1971 15102 2001
rect 15068 1967 15102 1971
rect 15068 1902 15102 1929
rect 15068 1895 15102 1902
rect 15068 1833 15102 1857
rect 15068 1823 15102 1833
rect 15068 1764 15102 1785
rect 15068 1751 15102 1764
rect 15068 1695 15102 1713
rect 15068 1679 15102 1695
rect 15068 1626 15102 1641
rect 15068 1607 15102 1626
rect 15068 1557 15102 1569
rect 15068 1535 15102 1557
rect 15068 1488 15102 1497
rect 15068 1463 15102 1488
rect 15068 1419 15102 1425
rect 15068 1391 15102 1419
rect 15068 1350 15102 1353
rect 15068 1319 15102 1350
rect 3565 1217 3577 1251
rect 3577 1217 3599 1251
rect 3637 1217 3645 1251
rect 3645 1217 3671 1251
rect 3709 1217 3713 1251
rect 3713 1217 3743 1251
rect 3781 1217 3815 1251
rect 3853 1217 3883 1251
rect 3883 1217 3887 1251
rect 3925 1217 3951 1251
rect 3951 1217 3959 1251
rect 3997 1217 4019 1251
rect 4019 1217 4031 1251
rect 4069 1217 4087 1251
rect 4087 1217 4103 1251
rect 4141 1217 4155 1251
rect 4155 1217 4175 1251
rect 4213 1217 4223 1251
rect 4223 1217 4247 1251
rect 4285 1217 4291 1251
rect 4291 1217 4319 1251
rect 4357 1217 4359 1251
rect 4359 1217 4391 1251
rect 4429 1217 4461 1251
rect 4461 1217 4463 1251
rect 4501 1217 4529 1251
rect 4529 1217 4535 1251
rect 4573 1217 4597 1251
rect 4597 1217 4607 1251
rect 4645 1217 4665 1251
rect 4665 1217 4679 1251
rect 4717 1217 4733 1251
rect 4733 1217 4751 1251
rect 4789 1217 4801 1251
rect 4801 1217 4823 1251
rect 4861 1217 4869 1251
rect 4869 1217 4895 1251
rect 4933 1217 4937 1251
rect 4937 1217 4967 1251
rect 5005 1217 5039 1251
rect 5077 1217 5107 1251
rect 5107 1217 5111 1251
rect 5149 1217 5175 1251
rect 5175 1217 5183 1251
rect 5221 1217 5243 1251
rect 5243 1217 5255 1251
rect 5293 1217 5311 1251
rect 5311 1217 5327 1251
rect 5365 1217 5379 1251
rect 5379 1217 5399 1251
rect 5437 1217 5447 1251
rect 5447 1217 5471 1251
rect 5509 1217 5515 1251
rect 5515 1217 5543 1251
rect 5581 1217 5583 1251
rect 5583 1217 5615 1251
rect 5653 1217 5685 1251
rect 5685 1217 5687 1251
rect 5725 1217 5753 1251
rect 5753 1217 5759 1251
rect 5797 1217 5821 1251
rect 5821 1217 5831 1251
rect 5869 1217 5889 1251
rect 5889 1217 5903 1251
rect 5941 1217 5957 1251
rect 5957 1217 5975 1251
rect 6013 1217 6025 1251
rect 6025 1217 6047 1251
rect 6085 1217 6093 1251
rect 6093 1217 6119 1251
rect 6157 1217 6161 1251
rect 6161 1217 6191 1251
rect 6229 1217 6263 1251
rect 6301 1217 6331 1251
rect 6331 1217 6335 1251
rect 6373 1217 6399 1251
rect 6399 1217 6407 1251
rect 6445 1217 6467 1251
rect 6467 1217 6479 1251
rect 6517 1217 6535 1251
rect 6535 1217 6551 1251
rect 6589 1217 6603 1251
rect 6603 1217 6623 1251
rect 6661 1217 6671 1251
rect 6671 1217 6695 1251
rect 6733 1217 6739 1251
rect 6739 1217 6767 1251
rect 6805 1217 6807 1251
rect 6807 1217 6839 1251
rect 6877 1217 6909 1251
rect 6909 1217 6911 1251
rect 6988 1227 7022 1239
rect 6988 1205 7022 1227
rect 15068 1247 15102 1281
rect 7069 1189 7103 1217
rect 7142 1189 7176 1217
rect 7215 1189 7249 1217
rect 7288 1189 7322 1217
rect 7361 1189 7395 1217
rect 7434 1189 7468 1217
rect 7507 1189 7541 1217
rect 7580 1189 7614 1217
rect 7653 1189 7687 1217
rect 7726 1189 7760 1217
rect 7799 1189 7833 1217
rect 7872 1189 7906 1217
rect 7945 1189 7979 1217
rect 8018 1189 8052 1217
rect 8091 1189 8125 1217
rect 8164 1189 8198 1217
rect 8237 1189 8271 1217
rect 8310 1189 8344 1217
rect 8383 1189 8417 1217
rect 8456 1189 8490 1217
rect 8528 1189 8562 1217
rect 8600 1189 8634 1217
rect 8672 1189 8706 1217
rect 8744 1189 8778 1217
rect 8816 1189 8850 1217
rect 8888 1189 8922 1217
rect 8960 1189 8994 1217
rect 9032 1189 9066 1217
rect 7069 1183 7102 1189
rect 7102 1183 7103 1189
rect 7142 1183 7171 1189
rect 7171 1183 7176 1189
rect 7215 1183 7240 1189
rect 7240 1183 7249 1189
rect 7288 1183 7309 1189
rect 7309 1183 7322 1189
rect 7361 1183 7378 1189
rect 7378 1183 7395 1189
rect 7434 1183 7447 1189
rect 7447 1183 7468 1189
rect 7507 1183 7516 1189
rect 7516 1183 7541 1189
rect 7580 1183 7585 1189
rect 7585 1183 7614 1189
rect 7653 1183 7654 1189
rect 7654 1183 7687 1189
rect 6988 1159 7022 1167
rect 6988 1133 7022 1159
rect 7726 1183 7758 1189
rect 7758 1183 7760 1189
rect 7799 1183 7827 1189
rect 7827 1183 7833 1189
rect 7872 1183 7896 1189
rect 7896 1183 7906 1189
rect 7945 1183 7965 1189
rect 7965 1183 7979 1189
rect 8018 1183 8034 1189
rect 8034 1183 8052 1189
rect 8091 1183 8103 1189
rect 8103 1183 8125 1189
rect 8164 1183 8172 1189
rect 8172 1183 8198 1189
rect 8237 1183 8241 1189
rect 8241 1183 8271 1189
rect 8310 1183 8344 1189
rect 8383 1183 8413 1189
rect 8413 1183 8417 1189
rect 8456 1183 8482 1189
rect 8482 1183 8490 1189
rect 8528 1183 8551 1189
rect 8551 1183 8562 1189
rect 8600 1183 8620 1189
rect 8620 1183 8634 1189
rect 8672 1183 8689 1189
rect 8689 1183 8706 1189
rect 8744 1183 8758 1189
rect 8758 1183 8778 1189
rect 8816 1183 8827 1189
rect 8827 1183 8850 1189
rect 8888 1183 8896 1189
rect 8896 1183 8922 1189
rect 8960 1183 8965 1189
rect 8965 1183 8994 1189
rect 9032 1183 9034 1189
rect 9034 1183 9066 1189
rect 9104 1183 9138 1217
rect 9176 1189 9210 1217
rect 9248 1189 9282 1217
rect 9320 1189 9354 1217
rect 9392 1189 9426 1217
rect 9464 1189 9498 1217
rect 9536 1189 9570 1217
rect 9608 1189 9642 1217
rect 9680 1189 9714 1217
rect 9176 1183 9207 1189
rect 9207 1183 9210 1189
rect 9248 1183 9276 1189
rect 9276 1183 9282 1189
rect 9320 1183 9345 1189
rect 9345 1183 9354 1189
rect 9392 1183 9414 1189
rect 9414 1183 9426 1189
rect 9464 1183 9483 1189
rect 9483 1183 9498 1189
rect 9536 1183 9552 1189
rect 9552 1183 9570 1189
rect 9608 1183 9621 1189
rect 9621 1183 9642 1189
rect 9680 1183 9690 1189
rect 9690 1183 9714 1189
rect 9752 1183 9759 1217
rect 9759 1183 9786 1217
rect 9824 1183 9858 1217
rect 9896 1183 9930 1217
rect 9968 1183 10002 1217
rect 10040 1183 10074 1217
rect 10112 1183 10146 1217
rect 10184 1183 10218 1217
rect 10256 1183 10290 1217
rect 10328 1183 10362 1217
rect 10400 1183 10434 1217
rect 10472 1183 10506 1217
rect 10544 1183 10578 1217
rect 10616 1183 10650 1217
rect 10688 1183 10722 1217
rect 10760 1183 10794 1217
rect 10832 1183 10866 1217
rect 10904 1183 10938 1217
rect 10976 1183 11010 1217
rect 11048 1183 11082 1217
rect 11120 1183 11154 1217
rect 11192 1183 11226 1217
rect 11264 1183 11298 1217
rect 11336 1183 11370 1217
rect 11408 1183 11442 1217
rect 11480 1183 11514 1217
rect 11552 1183 11586 1217
rect 11624 1183 11658 1217
rect 11696 1183 11730 1217
rect 11768 1183 11802 1217
rect 11840 1183 11874 1217
rect 11912 1183 11946 1217
rect 11984 1183 12018 1217
rect 12056 1183 12090 1217
rect 12139 1183 12173 1217
rect 12212 1183 12246 1217
rect 12285 1183 12319 1217
rect 12358 1183 12392 1217
rect 12431 1183 12465 1217
rect 12504 1183 12538 1217
rect 12577 1183 12611 1217
rect 12650 1183 12684 1217
rect 12723 1183 12757 1217
rect 12796 1183 12830 1217
rect 12869 1183 12903 1217
rect 12942 1183 12976 1217
rect 13015 1183 13049 1217
rect 13088 1183 13122 1217
rect 13161 1183 13195 1217
rect 13234 1183 13268 1217
rect 13307 1183 13341 1217
rect 13380 1183 13414 1217
rect 13452 1183 13486 1217
rect 13524 1183 13558 1217
rect 13596 1183 13630 1217
rect 13668 1183 13702 1217
rect 13740 1183 13774 1217
rect 13812 1183 13846 1217
rect 13884 1183 13918 1217
rect 13956 1183 13990 1217
rect 14028 1183 14062 1217
rect 14100 1183 14134 1217
rect 14172 1183 14206 1217
rect 14244 1183 14278 1217
rect 14316 1183 14350 1217
rect 14388 1183 14422 1217
rect 14460 1183 14494 1217
rect 14532 1183 14566 1217
rect 14604 1183 14638 1217
rect 14676 1183 14710 1217
rect 14748 1183 14782 1217
rect 14820 1183 14854 1217
rect 14892 1183 14893 1217
rect 14893 1183 14926 1217
rect 14964 1210 14966 1217
rect 14966 1210 14998 1217
rect 14964 1183 14998 1210
rect 15068 1175 15102 1209
rect 7069 1121 7103 1139
rect 7142 1121 7176 1139
rect 7215 1121 7249 1139
rect 7288 1121 7322 1139
rect 7361 1121 7395 1139
rect 7434 1121 7468 1139
rect 7507 1121 7541 1139
rect 7580 1121 7614 1139
rect 7653 1121 7687 1139
rect 7726 1121 7760 1139
rect 7799 1121 7833 1139
rect 7872 1121 7906 1139
rect 7945 1121 7979 1139
rect 8018 1121 8052 1139
rect 8091 1121 8125 1139
rect 8164 1121 8198 1139
rect 8237 1121 8271 1139
rect 8310 1121 8344 1139
rect 8383 1121 8417 1139
rect 8456 1121 8490 1139
rect 8528 1121 8562 1139
rect 8600 1121 8634 1139
rect 8672 1121 8706 1139
rect 8744 1121 8778 1139
rect 8816 1121 8850 1139
rect 8888 1121 8922 1139
rect 8960 1121 8994 1139
rect 9032 1121 9066 1139
rect 7069 1105 7102 1121
rect 7102 1105 7103 1121
rect 7142 1105 7171 1121
rect 7171 1105 7176 1121
rect 7215 1105 7240 1121
rect 7240 1105 7249 1121
rect 7288 1105 7309 1121
rect 7309 1105 7322 1121
rect 7361 1105 7378 1121
rect 7378 1105 7395 1121
rect 7434 1105 7447 1121
rect 7447 1105 7468 1121
rect 7507 1105 7516 1121
rect 7516 1105 7541 1121
rect 7580 1105 7585 1121
rect 7585 1105 7614 1121
rect 7653 1105 7654 1121
rect 7654 1105 7687 1121
rect 6988 1091 7022 1095
rect 3528 909 3562 943
rect 3722 915 3738 949
rect 3738 915 3756 949
rect 3794 915 3806 949
rect 3806 915 3828 949
rect 3866 915 3874 949
rect 3874 915 3900 949
rect 3938 915 3942 949
rect 3942 915 3972 949
rect 4010 915 4044 949
rect 4082 915 4112 949
rect 4112 915 4116 949
rect 4154 915 4180 949
rect 4180 915 4188 949
rect 4226 915 4248 949
rect 4248 915 4260 949
rect 4298 915 4316 949
rect 4316 915 4332 949
rect 4370 915 4384 949
rect 4384 915 4404 949
rect 4442 915 4452 949
rect 4452 915 4476 949
rect 4514 915 4520 949
rect 4520 915 4548 949
rect 4586 915 4588 949
rect 4588 915 4620 949
rect 4658 915 4690 949
rect 4690 915 4692 949
rect 4730 915 4758 949
rect 4758 915 4764 949
rect 4802 915 4826 949
rect 4826 915 4836 949
rect 4874 915 4894 949
rect 4894 915 4908 949
rect 4946 915 4962 949
rect 4962 915 4980 949
rect 5018 915 5030 949
rect 5030 915 5052 949
rect 5090 915 5124 949
rect 5252 915 5268 949
rect 5268 915 5286 949
rect 5324 915 5336 949
rect 5336 915 5358 949
rect 5396 915 5404 949
rect 5404 915 5430 949
rect 5468 915 5472 949
rect 5472 915 5502 949
rect 5540 915 5574 949
rect 5612 915 5642 949
rect 5642 915 5646 949
rect 5684 915 5710 949
rect 5710 915 5718 949
rect 5756 915 5778 949
rect 5778 915 5790 949
rect 5828 915 5846 949
rect 5846 915 5862 949
rect 5900 915 5914 949
rect 5914 915 5934 949
rect 5972 915 5982 949
rect 5982 915 6006 949
rect 6044 915 6050 949
rect 6050 915 6078 949
rect 6116 915 6118 949
rect 6118 915 6150 949
rect 6188 915 6220 949
rect 6220 915 6222 949
rect 6260 915 6288 949
rect 6288 915 6294 949
rect 6332 915 6356 949
rect 6356 915 6366 949
rect 6404 915 6424 949
rect 6424 915 6438 949
rect 6476 915 6492 949
rect 6492 915 6510 949
rect 6548 915 6560 949
rect 6560 915 6582 949
rect 6620 915 6654 949
rect 3528 837 3562 871
rect 3528 765 3562 799
rect 3528 693 3562 727
rect 3528 621 3562 655
rect 3528 549 3562 583
rect 3528 477 3562 511
rect 3528 405 3562 439
rect 3528 333 3562 367
rect 3722 759 3738 793
rect 3738 759 3756 793
rect 3794 759 3806 793
rect 3806 759 3828 793
rect 3866 759 3874 793
rect 3874 759 3900 793
rect 3938 759 3942 793
rect 3942 759 3972 793
rect 4010 759 4044 793
rect 4082 759 4112 793
rect 4112 759 4116 793
rect 4154 759 4180 793
rect 4180 759 4188 793
rect 4226 759 4248 793
rect 4248 759 4260 793
rect 4298 759 4316 793
rect 4316 759 4332 793
rect 4370 759 4384 793
rect 4384 759 4404 793
rect 4442 759 4452 793
rect 4452 759 4476 793
rect 4514 759 4520 793
rect 4520 759 4548 793
rect 4586 759 4588 793
rect 4588 759 4620 793
rect 4658 759 4690 793
rect 4690 759 4692 793
rect 4730 759 4758 793
rect 4758 759 4764 793
rect 4802 759 4826 793
rect 4826 759 4836 793
rect 4874 759 4894 793
rect 4894 759 4908 793
rect 4946 759 4962 793
rect 4962 759 4980 793
rect 5018 759 5030 793
rect 5030 759 5052 793
rect 5090 759 5124 793
rect 5252 759 5268 793
rect 5268 759 5286 793
rect 5324 759 5336 793
rect 5336 759 5358 793
rect 5396 759 5404 793
rect 5404 759 5430 793
rect 5468 759 5472 793
rect 5472 759 5502 793
rect 5540 759 5574 793
rect 5612 759 5642 793
rect 5642 759 5646 793
rect 5684 759 5710 793
rect 5710 759 5718 793
rect 5756 759 5778 793
rect 5778 759 5790 793
rect 5828 759 5846 793
rect 5846 759 5862 793
rect 5900 759 5914 793
rect 5914 759 5934 793
rect 5972 759 5982 793
rect 5982 759 6006 793
rect 6044 759 6050 793
rect 6050 759 6078 793
rect 6116 759 6118 793
rect 6118 759 6150 793
rect 6188 759 6220 793
rect 6220 759 6222 793
rect 6260 759 6288 793
rect 6288 759 6294 793
rect 6332 759 6356 793
rect 6356 759 6366 793
rect 6404 759 6424 793
rect 6424 759 6438 793
rect 6476 759 6492 793
rect 6492 759 6510 793
rect 6548 759 6560 793
rect 6560 759 6582 793
rect 6620 759 6654 793
rect 3645 707 3678 714
rect 3678 707 3679 714
rect 3645 680 3679 707
rect 3717 680 3751 714
rect 5115 680 5149 714
rect 5187 693 5208 714
rect 5208 693 5221 714
rect 5187 680 5221 693
rect 6620 680 6654 714
rect 6692 710 6704 714
rect 6704 710 6726 714
rect 6692 680 6726 710
rect 3722 603 3738 637
rect 3738 603 3756 637
rect 3794 603 3806 637
rect 3806 603 3828 637
rect 3866 603 3874 637
rect 3874 603 3900 637
rect 3938 603 3942 637
rect 3942 603 3972 637
rect 4010 603 4044 637
rect 4082 603 4112 637
rect 4112 603 4116 637
rect 4154 603 4180 637
rect 4180 603 4188 637
rect 4226 603 4248 637
rect 4248 603 4260 637
rect 4298 603 4316 637
rect 4316 603 4332 637
rect 4370 603 4384 637
rect 4384 603 4404 637
rect 4442 603 4452 637
rect 4452 603 4476 637
rect 4514 603 4520 637
rect 4520 603 4548 637
rect 4586 603 4588 637
rect 4588 603 4620 637
rect 4658 603 4690 637
rect 4690 603 4692 637
rect 4730 603 4758 637
rect 4758 603 4764 637
rect 4802 603 4826 637
rect 4826 603 4836 637
rect 4874 603 4894 637
rect 4894 603 4908 637
rect 4946 603 4962 637
rect 4962 603 4980 637
rect 5018 603 5030 637
rect 5030 603 5052 637
rect 5090 603 5124 637
rect 5252 603 5268 637
rect 5268 603 5286 637
rect 5324 603 5336 637
rect 5336 603 5358 637
rect 5396 603 5404 637
rect 5404 603 5430 637
rect 5468 603 5472 637
rect 5472 603 5502 637
rect 5540 603 5574 637
rect 5612 603 5642 637
rect 5642 603 5646 637
rect 5684 603 5710 637
rect 5710 603 5718 637
rect 5756 603 5778 637
rect 5778 603 5790 637
rect 5828 603 5846 637
rect 5846 603 5862 637
rect 5900 603 5914 637
rect 5914 603 5934 637
rect 5972 603 5982 637
rect 5982 603 6006 637
rect 6044 603 6050 637
rect 6050 603 6078 637
rect 6116 603 6118 637
rect 6118 603 6150 637
rect 6188 603 6220 637
rect 6220 603 6222 637
rect 6260 603 6288 637
rect 6288 603 6294 637
rect 6332 603 6356 637
rect 6356 603 6366 637
rect 6404 603 6424 637
rect 6424 603 6438 637
rect 6476 603 6492 637
rect 6492 603 6510 637
rect 6548 603 6560 637
rect 6560 603 6582 637
rect 6620 603 6654 637
rect 3722 447 3738 481
rect 3738 447 3756 481
rect 3794 447 3806 481
rect 3806 447 3828 481
rect 3866 447 3874 481
rect 3874 447 3900 481
rect 3938 447 3942 481
rect 3942 447 3972 481
rect 4010 447 4044 481
rect 4082 447 4112 481
rect 4112 447 4116 481
rect 4154 447 4180 481
rect 4180 447 4188 481
rect 4226 447 4248 481
rect 4248 447 4260 481
rect 4298 447 4316 481
rect 4316 447 4332 481
rect 4370 447 4384 481
rect 4384 447 4404 481
rect 4442 447 4452 481
rect 4452 447 4476 481
rect 4514 447 4520 481
rect 4520 447 4548 481
rect 4586 447 4588 481
rect 4588 447 4620 481
rect 4658 447 4690 481
rect 4690 447 4692 481
rect 4730 447 4758 481
rect 4758 447 4764 481
rect 4802 447 4826 481
rect 4826 447 4836 481
rect 4874 447 4894 481
rect 4894 447 4908 481
rect 4946 447 4962 481
rect 4962 447 4980 481
rect 5018 447 5030 481
rect 5030 447 5052 481
rect 5090 447 5124 481
rect 5252 447 5268 481
rect 5268 447 5286 481
rect 5324 447 5336 481
rect 5336 447 5358 481
rect 5396 447 5404 481
rect 5404 447 5430 481
rect 5468 447 5472 481
rect 5472 447 5502 481
rect 5540 447 5574 481
rect 5612 447 5642 481
rect 5642 447 5646 481
rect 5684 447 5710 481
rect 5710 447 5718 481
rect 5756 447 5778 481
rect 5778 447 5790 481
rect 5828 447 5846 481
rect 5846 447 5862 481
rect 5900 447 5914 481
rect 5914 447 5934 481
rect 5972 447 5982 481
rect 5982 447 6006 481
rect 6044 447 6050 481
rect 6050 447 6078 481
rect 6116 447 6118 481
rect 6118 447 6150 481
rect 6188 447 6220 481
rect 6220 447 6222 481
rect 6260 447 6288 481
rect 6288 447 6294 481
rect 6332 447 6356 481
rect 6356 447 6366 481
rect 6404 447 6424 481
rect 6424 447 6438 481
rect 6476 447 6492 481
rect 6492 447 6510 481
rect 6548 447 6560 481
rect 6560 447 6582 481
rect 6620 447 6654 481
rect 6790 845 6824 869
rect 6790 835 6824 845
rect 6790 777 6824 797
rect 6790 763 6824 777
rect 6790 709 6824 725
rect 6790 691 6824 709
rect 6790 641 6824 653
rect 6790 619 6824 641
rect 6790 573 6824 581
rect 6790 547 6824 573
rect 6790 505 6824 509
rect 6790 475 6824 505
rect 6790 403 6824 437
rect 6790 335 6824 365
rect 6790 331 6824 335
rect 3528 260 3562 294
rect 3722 291 3738 325
rect 3738 291 3756 325
rect 3794 291 3806 325
rect 3806 291 3828 325
rect 3866 291 3874 325
rect 3874 291 3900 325
rect 3938 291 3942 325
rect 3942 291 3972 325
rect 4010 291 4044 325
rect 4082 291 4112 325
rect 4112 291 4116 325
rect 4154 291 4180 325
rect 4180 291 4188 325
rect 4226 291 4248 325
rect 4248 291 4260 325
rect 4298 291 4316 325
rect 4316 291 4332 325
rect 4370 291 4384 325
rect 4384 291 4404 325
rect 4442 291 4452 325
rect 4452 291 4476 325
rect 4514 291 4520 325
rect 4520 291 4548 325
rect 4586 291 4588 325
rect 4588 291 4620 325
rect 4658 291 4690 325
rect 4690 291 4692 325
rect 4730 291 4758 325
rect 4758 291 4764 325
rect 4802 291 4826 325
rect 4826 291 4836 325
rect 4874 291 4894 325
rect 4894 291 4908 325
rect 4946 291 4962 325
rect 4962 291 4980 325
rect 5018 291 5030 325
rect 5030 291 5052 325
rect 5090 291 5124 325
rect 5252 291 5268 325
rect 5268 291 5286 325
rect 5324 291 5336 325
rect 5336 291 5358 325
rect 5396 291 5404 325
rect 5404 291 5430 325
rect 5468 291 5472 325
rect 5472 291 5502 325
rect 5540 291 5574 325
rect 5612 291 5642 325
rect 5642 291 5646 325
rect 5684 291 5710 325
rect 5710 291 5718 325
rect 5756 291 5778 325
rect 5778 291 5790 325
rect 5828 291 5846 325
rect 5846 291 5862 325
rect 5900 291 5914 325
rect 5914 291 5934 325
rect 5972 291 5982 325
rect 5982 291 6006 325
rect 6044 291 6050 325
rect 6050 291 6078 325
rect 6116 291 6118 325
rect 6118 291 6150 325
rect 6188 291 6220 325
rect 6220 291 6222 325
rect 6260 291 6288 325
rect 6288 291 6294 325
rect 6332 291 6356 325
rect 6356 291 6366 325
rect 6404 291 6424 325
rect 6424 291 6438 325
rect 6476 291 6492 325
rect 6492 291 6510 325
rect 6548 291 6560 325
rect 6560 291 6582 325
rect 6620 291 6654 325
rect 3528 187 3562 221
rect 6790 267 6824 293
rect 6790 259 6824 267
rect 3632 175 3666 209
rect 3704 175 3734 209
rect 3734 175 3738 209
rect 3776 175 3802 209
rect 3802 175 3810 209
rect 3848 175 3870 209
rect 3870 175 3882 209
rect 3920 175 3938 209
rect 3938 175 3954 209
rect 3992 175 4006 209
rect 4006 175 4026 209
rect 4064 175 4074 209
rect 4074 175 4098 209
rect 4136 175 4142 209
rect 4142 175 4170 209
rect 4208 175 4210 209
rect 4210 175 4242 209
rect 4280 175 4312 209
rect 4312 175 4314 209
rect 4352 175 4380 209
rect 4380 175 4386 209
rect 4424 175 4448 209
rect 4448 175 4458 209
rect 4496 175 4516 209
rect 4516 175 4530 209
rect 4568 175 4584 209
rect 4584 175 4602 209
rect 4640 175 4652 209
rect 4652 175 4674 209
rect 4712 175 4720 209
rect 4720 175 4746 209
rect 4784 175 4788 209
rect 4788 175 4818 209
rect 4856 175 4890 209
rect 4928 175 4958 209
rect 4958 175 4962 209
rect 5000 175 5026 209
rect 5026 175 5034 209
rect 5072 175 5094 209
rect 5094 175 5106 209
rect 5144 175 5162 209
rect 5162 175 5178 209
rect 5216 175 5230 209
rect 5230 175 5250 209
rect 5288 175 5298 209
rect 5298 175 5322 209
rect 5360 175 5366 209
rect 5366 175 5394 209
rect 5432 175 5434 209
rect 5434 175 5466 209
rect 5504 175 5536 209
rect 5536 175 5538 209
rect 5576 175 5604 209
rect 5604 175 5610 209
rect 5648 175 5672 209
rect 5672 175 5682 209
rect 5720 175 5740 209
rect 5740 175 5754 209
rect 5792 175 5808 209
rect 5808 175 5826 209
rect 5864 175 5876 209
rect 5876 175 5898 209
rect 5936 175 5944 209
rect 5944 175 5970 209
rect 6008 175 6012 209
rect 6012 175 6042 209
rect 6080 175 6114 209
rect 6152 175 6182 209
rect 6182 175 6186 209
rect 6224 175 6250 209
rect 6250 175 6258 209
rect 6296 175 6318 209
rect 6318 175 6330 209
rect 6368 175 6386 209
rect 6386 175 6402 209
rect 6440 175 6454 209
rect 6454 175 6474 209
rect 6512 175 6522 209
rect 6522 175 6546 209
rect 6584 175 6590 209
rect 6590 175 6618 209
rect 6656 175 6658 209
rect 6658 175 6690 209
rect 6790 199 6824 221
rect 6790 187 6824 199
rect 6988 1061 7022 1091
rect 7726 1105 7758 1121
rect 7758 1105 7760 1121
rect 7799 1105 7827 1121
rect 7827 1105 7833 1121
rect 7872 1105 7896 1121
rect 7896 1105 7906 1121
rect 7945 1105 7965 1121
rect 7965 1105 7979 1121
rect 8018 1105 8034 1121
rect 8034 1105 8052 1121
rect 8091 1105 8103 1121
rect 8103 1105 8125 1121
rect 8164 1105 8172 1121
rect 8172 1105 8198 1121
rect 8237 1105 8241 1121
rect 8241 1105 8271 1121
rect 8310 1105 8344 1121
rect 8383 1105 8413 1121
rect 8413 1105 8417 1121
rect 8456 1105 8482 1121
rect 8482 1105 8490 1121
rect 8528 1105 8551 1121
rect 8551 1105 8562 1121
rect 8600 1105 8620 1121
rect 8620 1105 8634 1121
rect 8672 1105 8689 1121
rect 8689 1105 8706 1121
rect 8744 1105 8758 1121
rect 8758 1105 8778 1121
rect 8816 1105 8827 1121
rect 8827 1105 8850 1121
rect 8888 1105 8896 1121
rect 8896 1105 8922 1121
rect 8960 1105 8965 1121
rect 8965 1105 8994 1121
rect 9032 1105 9034 1121
rect 9034 1105 9066 1121
rect 9104 1105 9138 1139
rect 9176 1121 9210 1139
rect 9248 1121 9282 1139
rect 9320 1121 9354 1139
rect 9392 1121 9426 1139
rect 9464 1121 9498 1139
rect 9536 1121 9570 1139
rect 9608 1121 9642 1139
rect 9680 1121 9714 1139
rect 9176 1105 9207 1121
rect 9207 1105 9210 1121
rect 9248 1105 9276 1121
rect 9276 1105 9282 1121
rect 9320 1105 9345 1121
rect 9345 1105 9354 1121
rect 9392 1105 9414 1121
rect 9414 1105 9426 1121
rect 9464 1105 9483 1121
rect 9483 1105 9498 1121
rect 9536 1105 9552 1121
rect 9552 1105 9570 1121
rect 9608 1105 9621 1121
rect 9621 1105 9642 1121
rect 9680 1105 9690 1121
rect 9690 1105 9714 1121
rect 9752 1105 9759 1139
rect 9759 1105 9786 1139
rect 9824 1105 9858 1139
rect 9896 1105 9930 1139
rect 9968 1105 10002 1139
rect 10040 1105 10074 1139
rect 10112 1105 10146 1139
rect 10184 1105 10218 1139
rect 10256 1105 10290 1139
rect 10328 1105 10362 1139
rect 10400 1105 10434 1139
rect 10472 1105 10506 1139
rect 10544 1105 10578 1139
rect 10616 1105 10650 1139
rect 10688 1105 10722 1139
rect 10760 1105 10794 1139
rect 10832 1105 10866 1139
rect 10904 1105 10938 1139
rect 10976 1105 11010 1139
rect 11048 1105 11082 1139
rect 11120 1105 11154 1139
rect 11192 1105 11226 1139
rect 11264 1105 11298 1139
rect 11336 1105 11370 1139
rect 11408 1105 11442 1139
rect 11480 1105 11514 1139
rect 11552 1105 11586 1139
rect 11624 1105 11658 1139
rect 11696 1105 11730 1139
rect 11768 1105 11802 1139
rect 11840 1105 11874 1139
rect 11912 1105 11946 1139
rect 11984 1105 12018 1139
rect 12056 1105 12090 1139
rect 12139 1105 12173 1139
rect 12212 1105 12246 1139
rect 12285 1105 12319 1139
rect 12358 1105 12392 1139
rect 12431 1105 12465 1139
rect 12504 1105 12538 1139
rect 12577 1105 12611 1139
rect 12650 1105 12684 1139
rect 12723 1105 12757 1139
rect 12796 1105 12830 1139
rect 12869 1105 12903 1139
rect 12942 1105 12976 1139
rect 13015 1105 13049 1139
rect 13088 1105 13122 1139
rect 13161 1105 13195 1139
rect 13234 1105 13268 1139
rect 13307 1105 13341 1139
rect 13380 1105 13414 1139
rect 13452 1105 13486 1139
rect 13524 1105 13558 1139
rect 13596 1105 13630 1139
rect 13668 1105 13702 1139
rect 13740 1105 13774 1139
rect 13812 1105 13846 1139
rect 13884 1105 13918 1139
rect 13956 1105 13990 1139
rect 14028 1105 14062 1139
rect 14100 1105 14134 1139
rect 14172 1105 14206 1139
rect 14244 1105 14278 1139
rect 14316 1105 14350 1139
rect 14388 1105 14422 1139
rect 14460 1105 14494 1139
rect 14532 1105 14566 1139
rect 14604 1105 14638 1139
rect 14676 1105 14710 1139
rect 14748 1105 14782 1139
rect 14820 1105 14854 1139
rect 14892 1105 14893 1139
rect 14893 1105 14926 1139
rect 14964 1138 14966 1139
rect 14966 1138 14998 1139
rect 14964 1105 14998 1138
rect 15068 1103 15102 1137
rect 7069 1053 7103 1061
rect 7142 1053 7176 1061
rect 7215 1053 7249 1061
rect 7288 1053 7322 1061
rect 7361 1053 7395 1061
rect 7434 1053 7468 1061
rect 7507 1053 7541 1061
rect 7580 1053 7614 1061
rect 7653 1053 7687 1061
rect 7726 1053 7760 1061
rect 7799 1053 7833 1061
rect 7872 1053 7906 1061
rect 7945 1053 7979 1061
rect 8018 1053 8052 1061
rect 8091 1053 8125 1061
rect 8164 1053 8198 1061
rect 8237 1053 8271 1061
rect 8310 1053 8344 1061
rect 8383 1053 8417 1061
rect 8456 1053 8490 1061
rect 8528 1053 8562 1061
rect 8600 1053 8634 1061
rect 8672 1053 8706 1061
rect 8744 1053 8778 1061
rect 8816 1053 8850 1061
rect 8888 1053 8922 1061
rect 8960 1053 8994 1061
rect 9032 1053 9066 1061
rect 7069 1027 7102 1053
rect 7102 1027 7103 1053
rect 7142 1027 7171 1053
rect 7171 1027 7176 1053
rect 7215 1027 7240 1053
rect 7240 1027 7249 1053
rect 7288 1027 7309 1053
rect 7309 1027 7322 1053
rect 7361 1027 7378 1053
rect 7378 1027 7395 1053
rect 7434 1027 7447 1053
rect 7447 1027 7468 1053
rect 7507 1027 7516 1053
rect 7516 1027 7541 1053
rect 7580 1027 7585 1053
rect 7585 1027 7614 1053
rect 7653 1027 7654 1053
rect 7654 1027 7687 1053
rect 6988 989 7022 1023
rect 7726 1027 7758 1053
rect 7758 1027 7760 1053
rect 7799 1027 7827 1053
rect 7827 1027 7833 1053
rect 7872 1027 7896 1053
rect 7896 1027 7906 1053
rect 7945 1027 7965 1053
rect 7965 1027 7979 1053
rect 8018 1027 8034 1053
rect 8034 1027 8052 1053
rect 8091 1027 8103 1053
rect 8103 1027 8125 1053
rect 8164 1027 8172 1053
rect 8172 1027 8198 1053
rect 8237 1027 8241 1053
rect 8241 1027 8271 1053
rect 8310 1027 8344 1053
rect 8383 1027 8413 1053
rect 8413 1027 8417 1053
rect 8456 1027 8482 1053
rect 8482 1027 8490 1053
rect 8528 1027 8551 1053
rect 8551 1027 8562 1053
rect 8600 1027 8620 1053
rect 8620 1027 8634 1053
rect 8672 1027 8689 1053
rect 8689 1027 8706 1053
rect 8744 1027 8758 1053
rect 8758 1027 8778 1053
rect 8816 1027 8827 1053
rect 8827 1027 8850 1053
rect 8888 1027 8896 1053
rect 8896 1027 8922 1053
rect 8960 1027 8965 1053
rect 8965 1027 8994 1053
rect 9032 1027 9034 1053
rect 9034 1027 9066 1053
rect 9104 1027 9138 1061
rect 9176 1053 9210 1061
rect 9248 1053 9282 1061
rect 9320 1053 9354 1061
rect 9392 1053 9426 1061
rect 9464 1053 9498 1061
rect 9536 1053 9570 1061
rect 9608 1053 9642 1061
rect 9680 1053 9714 1061
rect 9176 1027 9207 1053
rect 9207 1027 9210 1053
rect 9248 1027 9276 1053
rect 9276 1027 9282 1053
rect 9320 1027 9345 1053
rect 9345 1027 9354 1053
rect 9392 1027 9414 1053
rect 9414 1027 9426 1053
rect 9464 1027 9483 1053
rect 9483 1027 9498 1053
rect 9536 1027 9552 1053
rect 9552 1027 9570 1053
rect 9608 1027 9621 1053
rect 9621 1027 9642 1053
rect 9680 1027 9690 1053
rect 9690 1027 9714 1053
rect 9752 1027 9759 1061
rect 9759 1027 9786 1061
rect 9824 1027 9858 1061
rect 9896 1027 9930 1061
rect 9968 1027 10002 1061
rect 10040 1027 10074 1061
rect 10112 1027 10146 1061
rect 10184 1027 10218 1061
rect 10256 1027 10290 1061
rect 10328 1027 10362 1061
rect 10400 1027 10434 1061
rect 10472 1027 10506 1061
rect 10544 1027 10578 1061
rect 10616 1027 10650 1061
rect 10688 1027 10722 1061
rect 10760 1027 10794 1061
rect 10832 1027 10866 1061
rect 10904 1027 10938 1061
rect 10976 1027 11010 1061
rect 11048 1027 11082 1061
rect 11120 1027 11154 1061
rect 11192 1027 11226 1061
rect 11264 1027 11298 1061
rect 11336 1027 11370 1061
rect 11408 1027 11442 1061
rect 11480 1027 11514 1061
rect 11552 1027 11586 1061
rect 11624 1027 11658 1061
rect 11696 1027 11730 1061
rect 11768 1027 11802 1061
rect 11840 1027 11874 1061
rect 11912 1027 11946 1061
rect 11984 1027 12018 1061
rect 12056 1027 12090 1061
rect 12139 1027 12173 1061
rect 12212 1027 12246 1061
rect 12285 1027 12319 1061
rect 12358 1027 12392 1061
rect 12431 1027 12465 1061
rect 12504 1027 12538 1061
rect 12577 1027 12611 1061
rect 12650 1027 12684 1061
rect 12723 1027 12757 1061
rect 12796 1027 12830 1061
rect 12869 1027 12903 1061
rect 12942 1027 12976 1061
rect 13015 1027 13049 1061
rect 13088 1027 13122 1061
rect 13161 1027 13195 1061
rect 13234 1027 13268 1061
rect 13307 1027 13341 1061
rect 13380 1027 13414 1061
rect 13452 1027 13486 1061
rect 13524 1027 13558 1061
rect 13596 1027 13630 1061
rect 13668 1027 13702 1061
rect 13740 1027 13774 1061
rect 13812 1027 13846 1061
rect 13884 1027 13918 1061
rect 13956 1027 13990 1061
rect 14028 1027 14062 1061
rect 14100 1027 14134 1061
rect 14172 1027 14206 1061
rect 14244 1027 14278 1061
rect 14316 1027 14350 1061
rect 14388 1027 14422 1061
rect 14460 1027 14494 1061
rect 14532 1027 14566 1061
rect 14604 1027 14638 1061
rect 14676 1027 14710 1061
rect 14748 1027 14782 1061
rect 14820 1027 14854 1061
rect 14892 1027 14893 1061
rect 14893 1027 14926 1061
rect 14964 1028 14998 1061
rect 15068 1031 15102 1065
rect 14964 1027 14966 1028
rect 14966 1027 14998 1028
rect 6988 921 7022 951
rect 6988 917 7022 921
rect 7104 913 7137 918
rect 7137 913 7138 918
rect 7104 884 7138 913
rect 6988 853 7022 879
rect 6988 845 7022 853
rect 6988 785 7022 807
rect 6988 773 7022 785
rect 6988 717 7022 735
rect 6988 701 7022 717
rect 6988 649 7022 663
rect 6988 629 7022 649
rect 6988 581 7022 591
rect 6988 557 7022 581
rect 6988 513 7022 519
rect 6988 485 7022 513
rect 6988 445 7022 447
rect 6988 413 7022 445
rect 6988 343 7022 375
rect 14576 955 14610 989
rect 14654 955 14688 989
rect 14732 955 14766 989
rect 14810 955 14844 989
rect 14888 955 14922 989
rect 9796 913 9815 923
rect 9815 913 9830 923
rect 9872 913 9885 923
rect 9885 913 9906 923
rect 9948 913 9955 923
rect 9955 913 9982 923
rect 10024 913 10025 923
rect 10025 913 10058 923
rect 10100 913 10131 923
rect 10131 913 10134 923
rect 10176 913 10201 923
rect 10201 913 10210 923
rect 10251 913 10271 923
rect 10271 913 10285 923
rect 10326 913 10341 923
rect 10341 913 10360 923
rect 10401 913 10411 923
rect 10411 913 10435 923
rect 10476 913 10481 923
rect 10481 913 10510 923
rect 10551 913 10585 923
rect 10626 913 10655 923
rect 10655 913 10660 923
rect 10701 913 10725 923
rect 10725 913 10735 923
rect 10776 913 10795 923
rect 10795 913 10810 923
rect 10851 913 10865 923
rect 10865 913 10885 923
rect 10926 913 10935 923
rect 10935 913 10960 923
rect 11001 913 11005 923
rect 11005 913 11035 923
rect 9796 889 9830 913
rect 9872 889 9906 913
rect 9948 889 9982 913
rect 10024 889 10058 913
rect 10100 889 10134 913
rect 10176 889 10210 913
rect 10251 889 10285 913
rect 10326 889 10360 913
rect 10401 889 10435 913
rect 10476 889 10510 913
rect 10551 889 10585 913
rect 10626 889 10660 913
rect 10701 889 10735 913
rect 10776 889 10810 913
rect 10851 889 10885 913
rect 10926 889 10960 913
rect 11001 889 11035 913
rect 11076 889 11110 923
rect 11151 913 11181 923
rect 11181 913 11185 923
rect 11226 913 11251 923
rect 11251 913 11260 923
rect 11301 913 11321 923
rect 11321 913 11335 923
rect 14966 955 15000 989
rect 15068 959 15102 993
rect 11151 889 11185 913
rect 11226 889 11260 913
rect 11301 889 11335 913
rect 14576 882 14610 916
rect 14654 882 14688 916
rect 14732 882 14766 916
rect 14810 882 14844 916
rect 14888 882 14922 916
rect 14576 841 14583 843
rect 14583 841 14610 843
rect 14966 882 15000 916
rect 15068 887 15102 921
rect 14654 841 14686 843
rect 14686 841 14688 843
rect 14732 841 14755 843
rect 14755 841 14766 843
rect 14810 841 14824 843
rect 14824 841 14844 843
rect 14888 841 14893 843
rect 14893 841 14922 843
rect 9796 805 9830 839
rect 9872 805 9906 839
rect 9948 805 9982 839
rect 10024 805 10058 839
rect 10100 805 10134 839
rect 10176 805 10210 839
rect 10251 805 10285 839
rect 10326 805 10360 839
rect 10401 805 10435 839
rect 10476 805 10510 839
rect 10551 805 10585 839
rect 10626 805 10660 839
rect 10701 805 10735 839
rect 10776 805 10810 839
rect 10851 805 10885 839
rect 10926 805 10960 839
rect 11001 805 11035 839
rect 11076 805 11110 839
rect 11151 805 11185 839
rect 11226 805 11260 839
rect 11301 805 11335 839
rect 14576 809 14610 841
rect 14654 809 14688 841
rect 14732 809 14766 841
rect 14810 809 14844 841
rect 14888 809 14922 841
rect 14576 761 14583 770
rect 14583 761 14610 770
rect 14966 809 15000 843
rect 15068 815 15102 849
rect 14654 761 14686 770
rect 14686 761 14688 770
rect 14732 761 14755 770
rect 14755 761 14766 770
rect 14810 761 14824 770
rect 14824 761 14844 770
rect 14888 761 14893 770
rect 14893 761 14922 770
rect 9796 731 9830 755
rect 9872 731 9906 755
rect 9948 731 9982 755
rect 10024 731 10058 755
rect 10100 731 10134 755
rect 10176 731 10210 755
rect 10251 731 10285 755
rect 10326 731 10360 755
rect 10401 731 10435 755
rect 10476 731 10510 755
rect 10551 731 10585 755
rect 10626 731 10660 755
rect 10701 731 10735 755
rect 10776 731 10810 755
rect 10851 731 10885 755
rect 10926 731 10960 755
rect 11001 731 11035 755
rect 9796 721 9815 731
rect 9815 721 9830 731
rect 9872 721 9885 731
rect 9885 721 9906 731
rect 9948 721 9955 731
rect 9955 721 9982 731
rect 10024 721 10025 731
rect 10025 721 10058 731
rect 10100 721 10131 731
rect 10131 721 10134 731
rect 10176 721 10201 731
rect 10201 721 10210 731
rect 10251 721 10271 731
rect 10271 721 10285 731
rect 10326 721 10341 731
rect 10341 721 10360 731
rect 10401 721 10411 731
rect 10411 721 10435 731
rect 10476 721 10481 731
rect 10481 721 10510 731
rect 10551 721 10585 731
rect 10626 721 10655 731
rect 10655 721 10660 731
rect 10701 721 10725 731
rect 10725 721 10735 731
rect 10776 721 10795 731
rect 10795 721 10810 731
rect 10851 721 10865 731
rect 10865 721 10885 731
rect 10926 721 10935 731
rect 10935 721 10960 731
rect 11001 721 11005 731
rect 11005 721 11035 731
rect 11076 721 11110 755
rect 11151 731 11185 755
rect 11226 731 11260 755
rect 11301 731 11335 755
rect 14576 736 14610 761
rect 14654 736 14688 761
rect 14732 736 14766 761
rect 14810 736 14844 761
rect 14888 736 14922 761
rect 11151 721 11181 731
rect 11181 721 11185 731
rect 11226 721 11251 731
rect 11251 721 11260 731
rect 11301 721 11321 731
rect 11321 721 11335 731
rect 9796 659 9830 671
rect 9872 659 9906 671
rect 9948 659 9982 671
rect 10024 659 10058 671
rect 10100 659 10134 671
rect 10176 659 10210 671
rect 10251 659 10285 671
rect 10326 659 10360 671
rect 10401 659 10435 671
rect 10476 659 10510 671
rect 10551 659 10585 671
rect 10626 659 10660 671
rect 10701 659 10735 671
rect 10776 659 10810 671
rect 10851 659 10885 671
rect 10926 659 10960 671
rect 11001 659 11035 671
rect 9796 637 9815 659
rect 9815 637 9830 659
rect 9872 637 9885 659
rect 9885 637 9906 659
rect 9948 637 9955 659
rect 9955 637 9982 659
rect 10024 637 10025 659
rect 10025 637 10058 659
rect 10100 637 10131 659
rect 10131 637 10134 659
rect 10176 637 10201 659
rect 10201 637 10210 659
rect 10251 637 10271 659
rect 10271 637 10285 659
rect 10326 637 10341 659
rect 10341 637 10360 659
rect 10401 637 10411 659
rect 10411 637 10435 659
rect 10476 637 10481 659
rect 10481 637 10510 659
rect 10551 637 10585 659
rect 10626 637 10655 659
rect 10655 637 10660 659
rect 10701 637 10725 659
rect 10725 637 10735 659
rect 10776 637 10795 659
rect 10795 637 10810 659
rect 10851 637 10865 659
rect 10865 637 10885 659
rect 10926 637 10935 659
rect 10935 637 10960 659
rect 11001 637 11005 659
rect 11005 637 11035 659
rect 11076 637 11110 671
rect 11151 659 11185 671
rect 11226 659 11260 671
rect 11301 659 11335 671
rect 11151 637 11181 659
rect 11181 637 11185 659
rect 11226 637 11251 659
rect 11251 637 11260 659
rect 11301 637 11321 659
rect 11321 637 11335 659
rect 9796 553 9815 587
rect 9815 553 9830 587
rect 9872 553 9885 587
rect 9885 553 9906 587
rect 9948 553 9955 587
rect 9955 553 9982 587
rect 10024 553 10025 587
rect 10025 553 10058 587
rect 10100 553 10131 587
rect 10131 553 10134 587
rect 10176 553 10201 587
rect 10201 553 10210 587
rect 10251 553 10271 587
rect 10271 553 10285 587
rect 10326 553 10341 587
rect 10341 553 10360 587
rect 10401 553 10411 587
rect 10411 553 10435 587
rect 10476 553 10481 587
rect 10481 553 10510 587
rect 10551 553 10585 587
rect 10626 553 10655 587
rect 10655 553 10660 587
rect 10701 553 10725 587
rect 10725 553 10735 587
rect 10776 553 10795 587
rect 10795 553 10810 587
rect 10851 553 10865 587
rect 10865 553 10885 587
rect 10926 553 10935 587
rect 10935 553 10960 587
rect 11001 553 11005 587
rect 11005 553 11035 587
rect 11076 553 11110 587
rect 11151 553 11181 587
rect 11181 553 11185 587
rect 11226 553 11251 587
rect 11251 553 11260 587
rect 11301 553 11321 587
rect 11321 553 11335 587
rect 9796 481 9815 503
rect 9815 481 9830 503
rect 9872 481 9885 503
rect 9885 481 9906 503
rect 9948 481 9955 503
rect 9955 481 9982 503
rect 10024 481 10025 503
rect 10025 481 10058 503
rect 10100 481 10131 503
rect 10131 481 10134 503
rect 10176 481 10201 503
rect 10201 481 10210 503
rect 10251 481 10271 503
rect 10271 481 10285 503
rect 10326 481 10341 503
rect 10341 481 10360 503
rect 10401 481 10411 503
rect 10411 481 10435 503
rect 10476 481 10481 503
rect 10481 481 10510 503
rect 10551 481 10585 503
rect 10626 481 10655 503
rect 10655 481 10660 503
rect 10701 481 10725 503
rect 10725 481 10735 503
rect 10776 481 10795 503
rect 10795 481 10810 503
rect 10851 481 10865 503
rect 10865 481 10885 503
rect 10926 481 10935 503
rect 10935 481 10960 503
rect 11001 481 11005 503
rect 11005 481 11035 503
rect 9796 469 9830 481
rect 9872 469 9906 481
rect 9948 469 9982 481
rect 10024 469 10058 481
rect 10100 469 10134 481
rect 10176 469 10210 481
rect 10251 469 10285 481
rect 10326 469 10360 481
rect 10401 469 10435 481
rect 10476 469 10510 481
rect 10551 469 10585 481
rect 10626 469 10660 481
rect 10701 469 10735 481
rect 10776 469 10810 481
rect 10851 469 10885 481
rect 10926 469 10960 481
rect 11001 469 11035 481
rect 11076 469 11110 503
rect 11151 481 11181 503
rect 11181 481 11185 503
rect 11226 481 11251 503
rect 11251 481 11260 503
rect 11301 481 11321 503
rect 11321 481 11335 503
rect 11151 469 11185 481
rect 11226 469 11260 481
rect 11301 469 11335 481
rect 14966 736 15000 770
rect 15068 743 15102 777
rect 14576 695 14610 697
rect 14654 695 14688 697
rect 14576 663 14577 695
rect 14577 663 14610 695
rect 14654 663 14655 695
rect 14655 663 14688 695
rect 14732 663 14766 697
rect 14810 663 14844 697
rect 14888 663 14922 697
rect 14966 663 15000 697
rect 15068 671 15102 705
rect 14576 609 14610 623
rect 14654 609 14688 623
rect 14576 589 14577 609
rect 14577 589 14610 609
rect 14654 589 14655 609
rect 14655 589 14688 609
rect 14732 589 14766 623
rect 14810 589 14844 623
rect 14888 589 14922 623
rect 14966 589 15000 623
rect 15068 599 15102 633
rect 14576 523 14610 549
rect 14654 523 14688 549
rect 14576 515 14577 523
rect 14577 515 14610 523
rect 14654 515 14655 523
rect 14655 515 14688 523
rect 14732 515 14766 549
rect 14810 515 14844 549
rect 14888 515 14922 549
rect 14966 515 15000 549
rect 15068 527 15102 561
rect 14576 441 14610 475
rect 14654 441 14688 475
rect 14732 441 14766 475
rect 14810 441 14844 475
rect 14888 441 14922 475
rect 14966 441 15000 475
rect 15068 455 15102 489
rect 14657 367 14691 390
rect 14735 367 14769 390
rect 14813 367 14847 390
rect 14891 367 14925 390
rect 14969 380 15003 390
rect 15068 383 15102 417
rect 6988 341 7022 343
rect 14657 356 14689 367
rect 14689 356 14691 367
rect 14735 356 14757 367
rect 14757 356 14769 367
rect 14813 356 14825 367
rect 14825 356 14847 367
rect 14891 356 14893 367
rect 14893 356 14925 367
rect 14969 356 15000 380
rect 15000 356 15003 380
rect 6988 275 7022 303
rect 14657 289 14691 312
rect 14735 289 14769 312
rect 14813 289 14847 312
rect 14891 289 14925 312
rect 14969 308 15003 312
rect 15068 311 15102 345
rect 6988 269 7022 275
rect 14657 278 14689 289
rect 14689 278 14691 289
rect 14735 278 14757 289
rect 14757 278 14769 289
rect 14813 278 14825 289
rect 14825 278 14847 289
rect 14891 278 14893 289
rect 14893 278 14925 289
rect 14969 278 15000 308
rect 15000 278 15003 308
rect 15068 238 15102 272
rect 6988 207 7022 231
rect 14657 211 14691 234
rect 14735 211 14769 234
rect 14813 211 14847 234
rect 14891 211 14925 234
rect 6988 197 7022 207
rect 14657 200 14689 211
rect 14689 200 14691 211
rect 14735 200 14757 211
rect 14757 200 14769 211
rect 14813 200 14825 211
rect 14825 200 14847 211
rect 14891 200 14893 211
rect 14893 200 14925 211
rect 14969 202 15000 234
rect 15000 202 15003 234
rect 14969 200 15003 202
rect 15068 165 15102 199
rect 6988 139 7022 159
rect 6988 125 7022 139
rect 14657 133 14691 156
rect 14735 133 14769 156
rect 14813 133 14847 156
rect 14891 133 14925 156
rect 14657 122 14689 133
rect 14689 122 14691 133
rect 14735 122 14757 133
rect 14757 122 14769 133
rect 14813 122 14825 133
rect 14825 122 14847 133
rect 14891 122 14893 133
rect 14893 122 14925 133
rect 14969 130 15000 156
rect 15000 130 15003 156
rect 14969 122 15003 130
rect 15068 92 15102 126
rect 14657 55 14691 77
rect 14735 55 14769 77
rect 14813 55 14847 77
rect 14891 55 14925 77
rect 14969 57 15000 77
rect 15000 57 15003 77
rect 3578 1 3612 35
rect 3652 23 3686 35
rect 3726 23 3760 35
rect 3800 23 3834 35
rect 3874 23 3908 35
rect 3948 23 3982 35
rect 4022 23 4056 35
rect 4096 23 4130 35
rect 4170 23 4204 35
rect 4244 23 4278 35
rect 4318 23 4352 35
rect 4392 23 4426 35
rect 4466 23 4500 35
rect 4540 23 4574 35
rect 4614 23 4648 35
rect 4688 23 4722 35
rect 4762 23 4796 35
rect 4836 23 4870 35
rect 4910 23 4944 35
rect 4984 23 5018 35
rect 5058 23 5092 35
rect 5132 23 5166 35
rect 5206 23 5240 35
rect 5280 23 5314 35
rect 5354 23 5388 35
rect 5428 23 5462 35
rect 3652 1 3666 23
rect 3666 1 3686 23
rect 3726 1 3734 23
rect 3734 1 3760 23
rect 3800 1 3802 23
rect 3802 1 3834 23
rect 3874 1 3904 23
rect 3904 1 3908 23
rect 3948 1 3972 23
rect 3972 1 3982 23
rect 4022 1 4040 23
rect 4040 1 4056 23
rect 4096 1 4108 23
rect 4108 1 4130 23
rect 4170 1 4176 23
rect 4176 1 4204 23
rect 4244 1 4278 23
rect 4318 1 4346 23
rect 4346 1 4352 23
rect 4392 1 4414 23
rect 4414 1 4426 23
rect 4466 1 4482 23
rect 4482 1 4500 23
rect 4540 1 4550 23
rect 4550 1 4574 23
rect 4614 1 4618 23
rect 4618 1 4648 23
rect 4688 1 4720 23
rect 4720 1 4722 23
rect 4762 1 4788 23
rect 4788 1 4796 23
rect 4836 1 4856 23
rect 4856 1 4870 23
rect 4910 1 4924 23
rect 4924 1 4944 23
rect 4984 1 4992 23
rect 4992 1 5018 23
rect 5058 1 5060 23
rect 5060 1 5092 23
rect 5132 1 5162 23
rect 5162 1 5166 23
rect 5206 1 5230 23
rect 5230 1 5240 23
rect 5280 1 5298 23
rect 5298 1 5314 23
rect 5354 1 5366 23
rect 5366 1 5388 23
rect 5428 1 5434 23
rect 5434 1 5462 23
rect 5502 1 5536 35
rect 5576 23 5610 35
rect 5650 23 5684 35
rect 5724 23 5758 35
rect 5798 23 5832 35
rect 5576 1 5604 23
rect 5604 1 5610 23
rect 5650 1 5672 23
rect 5672 1 5684 23
rect 5724 1 5740 23
rect 5740 1 5758 23
rect 5798 1 5808 23
rect 5808 1 5832 23
rect 5896 -11 5910 23
rect 5910 -11 5930 23
rect 5968 -11 5978 23
rect 5978 -11 6002 23
rect 6040 -11 6046 23
rect 6046 -11 6074 23
rect 6112 -11 6114 23
rect 6114 -11 6146 23
rect 6184 -11 6216 23
rect 6216 -11 6218 23
rect 6256 -11 6284 23
rect 6284 -11 6290 23
rect 6328 -11 6352 23
rect 6352 -11 6362 23
rect 6400 -11 6420 23
rect 6420 -11 6434 23
rect 6472 -11 6488 23
rect 6488 -11 6506 23
rect 6544 -11 6556 23
rect 6556 -11 6578 23
rect 6616 -11 6624 23
rect 6624 -11 6650 23
rect 6688 -11 6692 23
rect 6692 -11 6722 23
rect 6760 -11 6794 23
rect 6832 -11 6862 23
rect 6862 -11 6866 23
rect 6904 -11 6930 23
rect 6930 -11 6938 23
rect 6976 -11 6998 23
rect 6998 -11 7010 23
rect 14657 43 14689 55
rect 14689 43 14691 55
rect 14735 43 14757 55
rect 14757 43 14769 55
rect 14813 43 14825 55
rect 14825 43 14847 55
rect 14891 43 14893 55
rect 14893 43 14925 55
rect 14969 43 15003 57
rect 15068 19 15102 53
rect 5884 -9191 5918 -9157
rect 5884 -9263 5918 -9229
<< metal1 >>
tri 2275 16499 2281 16505 se
rect 2281 16499 2287 16505
tri 38 16493 44 16499 se
rect 44 16493 2287 16499
tri 23 16478 38 16493 se
rect 38 16478 131 16493
rect 57 16459 131 16478
rect 165 16459 204 16493
rect 238 16459 277 16493
rect 311 16459 350 16493
rect 384 16459 423 16493
rect 457 16459 496 16493
rect 530 16459 569 16493
rect 603 16459 642 16493
rect 676 16459 715 16493
rect 749 16459 788 16493
rect 822 16459 861 16493
rect 895 16459 934 16493
rect 968 16459 1007 16493
rect 1041 16459 1079 16493
rect 1113 16459 1151 16493
rect 1185 16459 1223 16493
rect 1257 16459 1295 16493
rect 1329 16459 1367 16493
rect 1401 16459 1439 16493
rect 1473 16459 1511 16493
rect 1545 16459 1583 16493
rect 1617 16459 1655 16493
rect 1689 16459 1727 16493
rect 1761 16459 1799 16493
rect 1833 16459 1871 16493
rect 1905 16459 1943 16493
rect 1977 16459 2015 16493
rect 2049 16459 2087 16493
rect 2121 16459 2159 16493
rect 2193 16459 2231 16493
rect 2265 16459 2287 16493
rect 57 16453 2287 16459
rect 2339 16453 2369 16505
rect 2421 16499 2427 16505
tri 2427 16499 2433 16505 sw
tri 14089 16499 14095 16505 se
rect 14095 16499 14101 16505
rect 2421 16493 14101 16499
rect 2421 16459 2447 16493
rect 2481 16459 2519 16493
rect 2553 16459 2591 16493
rect 2625 16459 2663 16493
rect 2697 16459 2735 16493
rect 2769 16459 2807 16493
rect 2841 16459 2879 16493
rect 2913 16459 2951 16493
rect 2985 16459 3023 16493
rect 3057 16459 3095 16493
rect 3129 16459 3167 16493
rect 3201 16459 3239 16493
rect 3273 16459 3311 16493
rect 3345 16459 3383 16493
rect 3417 16459 3455 16493
rect 3489 16459 3527 16493
rect 3561 16459 3599 16493
rect 3633 16459 3671 16493
rect 3705 16459 3743 16493
rect 3777 16459 3815 16493
rect 3849 16459 3887 16493
rect 3921 16459 3959 16493
rect 3993 16459 4031 16493
rect 4065 16459 4103 16493
rect 4137 16459 4175 16493
rect 4209 16459 4247 16493
rect 4281 16459 4319 16493
rect 4353 16459 4391 16493
rect 4425 16459 4463 16493
rect 4497 16459 4535 16493
rect 4569 16459 4607 16493
rect 4641 16459 4679 16493
rect 4713 16459 4751 16493
rect 4785 16459 4823 16493
rect 4857 16459 4895 16493
rect 4929 16459 4967 16493
rect 5001 16459 5039 16493
rect 5073 16459 5111 16493
rect 5145 16459 5183 16493
rect 5217 16459 5255 16493
rect 5289 16459 5327 16493
rect 5361 16459 5399 16493
rect 5433 16459 5471 16493
rect 5505 16459 5543 16493
rect 5577 16459 5615 16493
rect 5649 16459 5687 16493
rect 5721 16459 5759 16493
rect 5793 16459 5831 16493
rect 5865 16459 5903 16493
rect 5937 16459 5975 16493
rect 6009 16459 6047 16493
rect 6081 16459 6119 16493
rect 6153 16459 6191 16493
rect 6225 16459 6263 16493
rect 6297 16459 6335 16493
rect 6369 16459 6407 16493
rect 6441 16459 6479 16493
rect 6513 16459 6551 16493
rect 6585 16459 6623 16493
rect 6657 16459 6695 16493
rect 6729 16459 6767 16493
rect 6801 16459 6839 16493
rect 6873 16459 6911 16493
rect 6945 16459 6983 16493
rect 7017 16459 7055 16493
rect 7089 16459 7127 16493
rect 7161 16459 7199 16493
rect 7233 16459 7271 16493
rect 7305 16459 7343 16493
rect 7377 16459 7415 16493
rect 7449 16459 7487 16493
rect 7521 16459 7559 16493
rect 7593 16459 7631 16493
rect 7665 16459 7703 16493
rect 7737 16459 7775 16493
rect 7809 16459 7847 16493
rect 7881 16459 7919 16493
rect 7953 16459 7991 16493
rect 8025 16459 8063 16493
rect 8097 16459 8135 16493
rect 8169 16459 8207 16493
rect 8241 16459 8279 16493
rect 8313 16459 8351 16493
rect 8385 16459 8423 16493
rect 8457 16459 8495 16493
rect 8529 16459 8567 16493
rect 8601 16459 8639 16493
rect 8673 16459 8711 16493
rect 8745 16459 8783 16493
rect 8817 16459 8855 16493
rect 8889 16459 8927 16493
rect 8961 16459 8999 16493
rect 9033 16459 9071 16493
rect 9105 16459 9143 16493
rect 9177 16459 9215 16493
rect 9249 16459 9287 16493
rect 9321 16459 9359 16493
rect 9393 16459 9431 16493
rect 9465 16459 9503 16493
rect 9537 16459 9575 16493
rect 9609 16459 9647 16493
rect 9681 16459 9719 16493
rect 9753 16459 9791 16493
rect 9825 16459 9863 16493
rect 9897 16459 9935 16493
rect 9969 16459 10007 16493
rect 10041 16459 10079 16493
rect 10113 16459 10151 16493
rect 10185 16459 10223 16493
rect 10257 16459 10295 16493
rect 10329 16459 10367 16493
rect 10401 16459 10439 16493
rect 10473 16459 10511 16493
rect 10545 16459 10583 16493
rect 10617 16459 10655 16493
rect 10689 16459 10727 16493
rect 10761 16459 10799 16493
rect 10833 16459 10871 16493
rect 10905 16459 10943 16493
rect 10977 16459 11015 16493
rect 11049 16459 11087 16493
rect 11121 16459 11159 16493
rect 11193 16459 11231 16493
rect 11265 16459 11303 16493
rect 11337 16459 11375 16493
rect 11409 16459 11447 16493
rect 11481 16459 11519 16493
rect 11553 16459 11591 16493
rect 11625 16459 11663 16493
rect 11697 16459 11735 16493
rect 11769 16459 11807 16493
rect 11841 16459 11879 16493
rect 11913 16459 11951 16493
rect 11985 16459 12023 16493
rect 12057 16459 12095 16493
rect 12129 16459 12167 16493
rect 12201 16459 12239 16493
rect 12273 16459 12311 16493
rect 12345 16459 12383 16493
rect 12417 16459 12455 16493
rect 12489 16459 12527 16493
rect 12561 16459 12599 16493
rect 12633 16459 12671 16493
rect 12705 16459 12743 16493
rect 12777 16459 12815 16493
rect 12849 16459 12887 16493
rect 12921 16459 12959 16493
rect 12993 16459 13031 16493
rect 13065 16459 13103 16493
rect 13137 16459 13175 16493
rect 13209 16459 13247 16493
rect 13281 16459 13319 16493
rect 13353 16459 13391 16493
rect 13425 16459 13463 16493
rect 13497 16459 13535 16493
rect 13569 16459 13607 16493
rect 13641 16459 13679 16493
rect 13713 16459 13751 16493
rect 13785 16459 13823 16493
rect 13857 16459 13895 16493
rect 13929 16459 13967 16493
rect 14001 16459 14039 16493
rect 14073 16459 14101 16493
rect 2421 16453 14101 16459
rect 14153 16453 14175 16505
rect 14227 16453 14249 16505
rect 14301 16453 14323 16505
rect 14375 16453 14397 16505
rect 14449 16499 14455 16505
tri 14455 16499 14461 16505 sw
rect 14449 16493 14949 16499
rect 14449 16459 14471 16493
rect 14505 16459 14543 16493
rect 14577 16459 14615 16493
rect 14649 16459 14687 16493
rect 14721 16459 14759 16493
rect 14793 16459 14831 16493
rect 14865 16459 14903 16493
rect 14937 16459 14949 16493
rect 14449 16453 14949 16459
rect 57 16424 238 16453
tri 238 16424 267 16453 nw
rect 57 16411 217 16424
rect 47 16405 217 16411
rect 47 16371 59 16405
rect 93 16371 131 16405
rect 165 16403 217 16405
tri 217 16403 238 16424 nw
rect 385 16418 506 16424
rect 165 16371 177 16403
rect 47 16365 177 16371
rect 57 16363 177 16365
tri 177 16363 217 16403 nw
rect 437 16372 506 16418
rect 558 16372 570 16424
rect 622 16372 1938 16424
rect 1990 16372 2002 16424
rect 2054 16372 3468 16424
rect 3520 16372 3532 16424
rect 3584 16372 7754 16424
rect 7806 16372 7818 16424
rect 7870 16372 9456 16424
rect 9508 16372 9520 16424
rect 9572 16372 10936 16424
rect 10988 16372 11000 16424
rect 11052 16372 12279 16424
rect 12331 16372 12343 16424
rect 12395 16372 13713 16424
rect 13765 16372 13777 16424
rect 13829 16372 14946 16424
rect 14998 16372 15010 16424
rect 15062 16372 15068 16424
rect 437 16366 443 16372
rect 57 16325 139 16363
tri 139 16325 177 16363 nw
rect 385 16354 443 16366
rect 57 16296 110 16325
tri 110 16296 139 16325 nw
rect 437 16344 443 16354
tri 443 16344 471 16372 nw
tri 437 16338 443 16344 nw
rect 385 16296 437 16302
rect 57 16292 106 16296
tri 106 16292 110 16296 nw
rect 740 16292 748 16344
rect 800 16292 812 16344
rect 864 16292 1655 16344
rect 1707 16292 1719 16344
rect 1771 16292 3185 16344
rect 3237 16292 3249 16344
rect 3301 16292 3960 16344
rect 4012 16292 4024 16344
rect 4076 16292 4088 16344
rect 4140 16292 4152 16344
rect 4204 16292 4216 16344
rect 4268 16292 7324 16344
rect 7376 16292 7388 16344
rect 7440 16292 9026 16344
rect 9078 16292 9090 16344
rect 9142 16292 10506 16344
rect 10558 16292 10570 16344
rect 10622 16292 11849 16344
rect 11901 16292 11913 16344
rect 11965 16292 13283 16344
rect 13335 16292 13347 16344
rect 13399 16292 14866 16344
rect 14918 16292 14930 16344
rect 14982 16292 14988 16344
rect 57 16279 93 16292
tri 93 16279 106 16292 nw
rect 57 16273 87 16279
tri 87 16273 93 16279 nw
rect 57 16264 78 16273
tri 78 16264 87 16273 nw
tri 57 16243 78 16264 nw
rect 981 16212 989 16264
rect 1041 16212 1053 16264
rect 1105 16212 1351 16264
rect 1403 16212 1415 16264
rect 1467 16212 5738 16264
rect 5790 16212 5827 16264
rect 5879 16212 5916 16264
rect 5968 16212 6005 16264
rect 6057 16212 6894 16264
rect 6946 16212 6958 16264
rect 7010 16212 8596 16264
rect 8648 16212 8660 16264
rect 8712 16212 10076 16264
rect 10128 16212 10140 16264
rect 10192 16212 11419 16264
rect 11471 16212 11483 16264
rect 11535 16212 12853 16264
rect 12905 16212 12917 16264
rect 12969 16212 14786 16264
rect 14838 16212 14850 16264
rect 14902 16212 14908 16264
rect 359 16145 411 16151
rect 2532 16103 2538 16155
rect 2590 16103 2602 16155
rect 2654 16103 14706 16155
rect 14758 16103 14770 16155
rect 14822 16103 14828 16155
rect 359 16081 411 16093
tri 411 16075 439 16103 sw
rect 411 16029 8191 16075
rect 359 16023 8191 16029
rect 8243 16023 8255 16075
rect 8307 16023 9861 16075
rect 9913 16023 9925 16075
rect 9977 16023 9983 16075
rect 10252 16023 10258 16075
rect 10310 16023 10322 16075
rect 10374 16023 14626 16075
rect 14678 16023 14690 16075
rect 14742 16023 14748 16075
rect 278 15989 3616 15995
rect 330 15943 2162 15989
rect 330 15937 339 15943
rect 278 15925 339 15937
rect 330 15906 339 15925
tri 339 15906 376 15943 nw
tri 2128 15909 2162 15943 ne
rect 2214 15943 3616 15989
rect 3668 15943 3680 15995
rect 3732 15943 3738 15995
rect 3870 15985 14937 15986
rect 3870 15980 4439 15985
rect 4491 15980 4506 15985
rect 4558 15980 4573 15985
rect 4625 15980 4640 15985
rect 4692 15980 4707 15985
rect 4759 15980 4774 15985
rect 4826 15980 4841 15985
rect 4893 15980 4908 15985
rect 3870 15946 3882 15980
rect 3916 15946 3955 15980
rect 3989 15946 4028 15980
rect 4062 15946 4101 15980
rect 4135 15946 4174 15980
rect 4208 15946 4247 15980
rect 4281 15946 4320 15980
rect 4354 15946 4393 15980
rect 4427 15946 4439 15980
rect 4500 15946 4506 15980
rect 4826 15946 4831 15980
rect 4893 15946 4904 15980
rect 2162 15925 2214 15937
tri 330 15897 339 15906 nw
rect 278 15867 330 15873
tri 2214 15909 2248 15943 nw
rect 3870 15933 4439 15946
rect 4491 15933 4506 15946
rect 4558 15933 4573 15946
rect 4625 15933 4640 15946
rect 4692 15933 4707 15946
rect 4759 15933 4774 15946
rect 4826 15933 4841 15946
rect 4893 15933 4908 15946
rect 4960 15933 4975 15985
rect 5027 15933 5042 15985
rect 5094 15933 5108 15985
rect 5160 15933 5174 15985
rect 5226 15980 5240 15985
rect 5292 15980 5306 15985
rect 5358 15980 5372 15985
rect 5424 15980 5438 15985
rect 5490 15980 6198 15985
rect 6250 15980 6269 15985
rect 6321 15980 6339 15985
rect 6391 15980 6409 15985
rect 6461 15980 6479 15985
rect 6531 15980 6549 15985
rect 6601 15980 6619 15985
rect 6671 15980 6689 15985
rect 6741 15980 6759 15985
rect 6811 15980 14103 15985
rect 14155 15980 14201 15985
rect 14253 15980 14298 15985
rect 14350 15980 14395 15985
rect 14447 15980 14937 15985
rect 5230 15946 5240 15980
rect 5303 15946 5306 15980
rect 5522 15946 5561 15980
rect 5595 15946 5634 15980
rect 5668 15946 5707 15980
rect 5741 15946 5780 15980
rect 5814 15946 5853 15980
rect 5887 15946 5926 15980
rect 5960 15946 5999 15980
rect 6033 15946 6072 15980
rect 6106 15946 6145 15980
rect 6179 15946 6198 15980
rect 6252 15946 6269 15980
rect 6325 15946 6339 15980
rect 6398 15946 6409 15980
rect 6471 15946 6479 15980
rect 6544 15946 6549 15980
rect 6617 15946 6619 15980
rect 6836 15946 6875 15980
rect 6909 15946 6948 15980
rect 6982 15946 7021 15980
rect 7055 15946 7094 15980
rect 7128 15946 7167 15980
rect 7201 15946 7240 15980
rect 7274 15946 7313 15980
rect 7347 15946 7386 15980
rect 7420 15946 7459 15980
rect 7493 15946 7532 15980
rect 7566 15946 7605 15980
rect 7639 15946 7678 15980
rect 7712 15946 7751 15980
rect 7785 15946 7824 15980
rect 7858 15946 7897 15980
rect 7931 15946 7970 15980
rect 8004 15946 8043 15980
rect 8077 15946 8116 15980
rect 8150 15946 8189 15980
rect 8223 15946 8262 15980
rect 8296 15946 8335 15980
rect 8369 15946 8408 15980
rect 8442 15946 8481 15980
rect 8515 15946 8554 15980
rect 8588 15946 8627 15980
rect 8661 15946 8699 15980
rect 8733 15946 8771 15980
rect 8805 15946 8843 15980
rect 8877 15946 8915 15980
rect 8949 15946 8987 15980
rect 9021 15946 9059 15980
rect 9093 15946 9131 15980
rect 9165 15946 9203 15980
rect 9237 15946 9275 15980
rect 9309 15946 9347 15980
rect 9381 15946 9419 15980
rect 9453 15946 9491 15980
rect 9525 15946 9563 15980
rect 9597 15946 9635 15980
rect 9669 15946 9707 15980
rect 9741 15946 9779 15980
rect 9813 15946 9851 15980
rect 9885 15946 9923 15980
rect 9957 15946 9995 15980
rect 10029 15946 10067 15980
rect 10101 15946 10139 15980
rect 10173 15946 10211 15980
rect 10245 15946 10283 15980
rect 10317 15946 10355 15980
rect 10389 15946 10427 15980
rect 10461 15946 10499 15980
rect 10533 15946 10571 15980
rect 10605 15946 10643 15980
rect 10677 15946 10715 15980
rect 10749 15946 10787 15980
rect 10821 15946 10859 15980
rect 10893 15946 10931 15980
rect 10965 15946 11003 15980
rect 11037 15946 11075 15980
rect 11109 15946 11147 15980
rect 11181 15946 11219 15980
rect 11253 15946 11291 15980
rect 11325 15946 11363 15980
rect 11397 15946 11435 15980
rect 11469 15946 11507 15980
rect 11541 15946 11579 15980
rect 11613 15946 11651 15980
rect 11685 15946 11723 15980
rect 11757 15946 11795 15980
rect 11829 15946 11867 15980
rect 11901 15946 11939 15980
rect 11973 15946 12011 15980
rect 12045 15946 12083 15980
rect 12117 15946 12155 15980
rect 12189 15946 12227 15980
rect 12261 15946 12299 15980
rect 12333 15946 12371 15980
rect 12405 15946 12443 15980
rect 12477 15946 12515 15980
rect 12586 15946 12587 15980
rect 12621 15946 12659 15980
rect 12693 15946 12731 15980
rect 12765 15946 12803 15980
rect 12837 15946 12875 15980
rect 12909 15946 12947 15980
rect 12981 15946 13019 15980
rect 13053 15946 13091 15980
rect 13125 15946 13163 15980
rect 13197 15946 13235 15980
rect 13269 15946 13307 15980
rect 13341 15946 13379 15980
rect 13413 15946 13451 15980
rect 13485 15946 13523 15980
rect 13557 15946 13595 15980
rect 13629 15946 13667 15980
rect 13701 15946 13739 15980
rect 13773 15946 13811 15980
rect 13845 15946 13883 15980
rect 13917 15946 13955 15980
rect 13989 15946 14027 15980
rect 14061 15946 14099 15980
rect 14155 15946 14171 15980
rect 14277 15946 14298 15980
rect 14350 15946 14387 15980
rect 14447 15946 14459 15980
rect 14493 15946 14531 15980
rect 14565 15946 14603 15980
rect 14637 15946 14675 15980
rect 14709 15946 14747 15980
rect 14781 15946 14819 15980
rect 14853 15946 14891 15980
rect 14925 15946 14937 15980
rect 5226 15933 5240 15946
rect 5292 15933 5306 15946
rect 5358 15933 5372 15946
rect 5424 15933 5438 15946
rect 5490 15933 6198 15946
rect 6250 15933 6269 15946
rect 6321 15933 6339 15946
rect 6391 15933 6409 15946
rect 6461 15933 6479 15946
rect 6531 15933 6549 15946
rect 6601 15933 6619 15946
rect 6671 15933 6689 15946
rect 6741 15933 6759 15946
rect 6811 15933 12534 15946
rect 3870 15928 12534 15933
rect 12586 15933 14103 15946
rect 14155 15933 14201 15946
rect 14253 15933 14298 15946
rect 14350 15933 14395 15946
rect 14447 15933 14937 15946
rect 12586 15928 14937 15933
rect 3870 15917 14937 15928
rect 3870 15915 14103 15917
rect 2162 15867 2214 15873
rect 3870 15906 4439 15915
rect 4491 15906 4506 15915
rect 4558 15906 4573 15915
rect 4625 15906 4640 15915
rect 4692 15906 4707 15915
rect 4759 15906 4774 15915
rect 4826 15906 4841 15915
rect 4893 15906 4908 15915
rect 3870 15872 3882 15906
rect 3916 15872 3955 15906
rect 3989 15872 4028 15906
rect 4062 15872 4101 15906
rect 4135 15872 4174 15906
rect 4208 15872 4247 15906
rect 4281 15872 4320 15906
rect 4354 15872 4393 15906
rect 4427 15872 4439 15906
rect 4500 15872 4506 15906
rect 4826 15872 4831 15906
rect 4893 15872 4904 15906
rect 3870 15863 4439 15872
rect 4491 15863 4506 15872
rect 4558 15863 4573 15872
rect 4625 15863 4640 15872
rect 4692 15863 4707 15872
rect 4759 15863 4774 15872
rect 4826 15863 4841 15872
rect 4893 15863 4908 15872
rect 4960 15863 4975 15915
rect 5027 15863 5042 15915
rect 5094 15863 5108 15915
rect 5160 15863 5174 15915
rect 5226 15906 5240 15915
rect 5292 15906 5306 15915
rect 5358 15906 5372 15915
rect 5424 15906 5438 15915
rect 5490 15906 6198 15915
rect 6250 15906 6269 15915
rect 6321 15906 6339 15915
rect 6391 15906 6409 15915
rect 6461 15906 6479 15915
rect 6531 15906 6549 15915
rect 6601 15906 6619 15915
rect 6671 15906 6689 15915
rect 6741 15906 6759 15915
rect 6811 15906 12534 15915
rect 12586 15906 14103 15915
rect 14155 15906 14201 15917
rect 14253 15906 14298 15917
rect 14350 15906 14395 15917
rect 14447 15906 14937 15917
rect 5230 15872 5240 15906
rect 5303 15872 5306 15906
rect 5522 15872 5561 15906
rect 5595 15872 5634 15906
rect 5668 15872 5707 15906
rect 5741 15872 5780 15906
rect 5814 15872 5853 15906
rect 5887 15872 5926 15906
rect 5960 15872 5999 15906
rect 6033 15872 6072 15906
rect 6106 15872 6145 15906
rect 6179 15872 6198 15906
rect 6252 15872 6269 15906
rect 6325 15872 6339 15906
rect 6398 15872 6409 15906
rect 6471 15872 6479 15906
rect 6544 15872 6549 15906
rect 6617 15872 6619 15906
rect 6836 15872 6875 15906
rect 6909 15872 6948 15906
rect 6982 15872 7021 15906
rect 7055 15872 7094 15906
rect 7128 15872 7167 15906
rect 7201 15872 7240 15906
rect 7274 15872 7313 15906
rect 7347 15872 7386 15906
rect 7420 15872 7459 15906
rect 7493 15872 7532 15906
rect 7566 15872 7605 15906
rect 7639 15872 7678 15906
rect 7712 15872 7751 15906
rect 7785 15872 7824 15906
rect 7858 15872 7897 15906
rect 7931 15872 7970 15906
rect 8004 15872 8043 15906
rect 8077 15872 8116 15906
rect 8150 15872 8189 15906
rect 8223 15872 8262 15906
rect 8296 15872 8335 15906
rect 8369 15872 8408 15906
rect 8442 15872 8481 15906
rect 8515 15872 8554 15906
rect 8588 15872 8627 15906
rect 8661 15872 8699 15906
rect 8733 15872 8771 15906
rect 8805 15872 8843 15906
rect 8877 15872 8915 15906
rect 8949 15872 8987 15906
rect 9021 15872 9059 15906
rect 9093 15872 9131 15906
rect 9165 15872 9203 15906
rect 9237 15872 9275 15906
rect 9309 15872 9347 15906
rect 9381 15872 9419 15906
rect 9453 15872 9491 15906
rect 9525 15872 9563 15906
rect 9597 15872 9635 15906
rect 9669 15872 9707 15906
rect 9741 15872 9779 15906
rect 9813 15872 9851 15906
rect 9885 15872 9923 15906
rect 9957 15872 9995 15906
rect 10029 15872 10067 15906
rect 10101 15872 10139 15906
rect 10173 15872 10211 15906
rect 10245 15872 10283 15906
rect 10317 15872 10355 15906
rect 10389 15872 10427 15906
rect 10461 15872 10499 15906
rect 10533 15872 10571 15906
rect 10605 15872 10643 15906
rect 10677 15872 10715 15906
rect 10749 15872 10787 15906
rect 10821 15872 10859 15906
rect 10893 15872 10931 15906
rect 10965 15872 11003 15906
rect 11037 15872 11075 15906
rect 11109 15872 11147 15906
rect 11181 15872 11219 15906
rect 11253 15872 11291 15906
rect 11325 15872 11363 15906
rect 11397 15872 11435 15906
rect 11469 15872 11507 15906
rect 11541 15872 11579 15906
rect 11613 15872 11651 15906
rect 11685 15872 11723 15906
rect 11757 15872 11795 15906
rect 11829 15872 11867 15906
rect 11901 15872 11939 15906
rect 11973 15872 12011 15906
rect 12045 15872 12083 15906
rect 12117 15872 12155 15906
rect 12189 15872 12227 15906
rect 12261 15872 12299 15906
rect 12333 15872 12371 15906
rect 12405 15872 12443 15906
rect 12477 15872 12515 15906
rect 12586 15872 12587 15906
rect 12621 15872 12659 15906
rect 12693 15872 12731 15906
rect 12765 15872 12803 15906
rect 12837 15872 12875 15906
rect 12909 15872 12947 15906
rect 12981 15872 13019 15906
rect 13053 15872 13091 15906
rect 13125 15872 13163 15906
rect 13197 15872 13235 15906
rect 13269 15872 13307 15906
rect 13341 15872 13379 15906
rect 13413 15872 13451 15906
rect 13485 15872 13523 15906
rect 13557 15872 13595 15906
rect 13629 15872 13667 15906
rect 13701 15872 13739 15906
rect 13773 15872 13811 15906
rect 13845 15872 13883 15906
rect 13917 15872 13955 15906
rect 13989 15872 14027 15906
rect 14061 15872 14099 15906
rect 14155 15872 14171 15906
rect 14277 15872 14298 15906
rect 14350 15872 14387 15906
rect 14447 15872 14459 15906
rect 14493 15872 14531 15906
rect 14565 15872 14603 15906
rect 14637 15872 14675 15906
rect 14709 15872 14747 15906
rect 14781 15872 14819 15906
rect 14853 15872 14891 15906
rect 14925 15872 14937 15906
rect 5226 15863 5240 15872
rect 5292 15863 5306 15872
rect 5358 15863 5372 15872
rect 5424 15863 5438 15872
rect 5490 15863 6198 15872
rect 6250 15863 6269 15872
rect 6321 15863 6339 15872
rect 6391 15863 6409 15872
rect 6461 15863 6479 15872
rect 6531 15863 6549 15872
rect 6601 15863 6619 15872
rect 6671 15863 6689 15872
rect 6741 15863 6759 15872
rect 6811 15863 12534 15872
rect 12586 15865 14103 15872
rect 14155 15865 14201 15872
rect 14253 15865 14298 15872
rect 14350 15865 14395 15872
rect 14447 15865 14937 15872
rect 12586 15863 14937 15865
rect 3870 15850 14937 15863
rect 3870 15845 12534 15850
rect 3870 15832 4439 15845
rect 4491 15832 4506 15845
rect 4558 15832 4573 15845
rect 4625 15832 4640 15845
rect 4692 15832 4707 15845
rect 4759 15832 4774 15845
rect 4826 15832 4841 15845
rect 4893 15832 4908 15845
rect 93 15789 139 15801
rect 3870 15798 3882 15832
rect 3916 15798 3955 15832
rect 3989 15798 4028 15832
rect 4062 15798 4101 15832
rect 4135 15798 4174 15832
rect 4208 15798 4247 15832
rect 4281 15798 4320 15832
rect 4354 15798 4393 15832
rect 4427 15798 4439 15832
rect 4500 15798 4506 15832
rect 4826 15798 4831 15832
rect 4893 15798 4904 15832
rect 3870 15793 4439 15798
rect 4491 15793 4506 15798
rect 4558 15793 4573 15798
rect 4625 15793 4640 15798
rect 4692 15793 4707 15798
rect 4759 15793 4774 15798
rect 4826 15793 4841 15798
rect 4893 15793 4908 15798
rect 4960 15793 4975 15845
rect 5027 15793 5042 15845
rect 5094 15793 5108 15845
rect 5160 15793 5174 15845
rect 5226 15832 5240 15845
rect 5292 15832 5306 15845
rect 5358 15832 5372 15845
rect 5424 15832 5438 15845
rect 5490 15832 6198 15845
rect 6250 15832 6269 15845
rect 6321 15832 6339 15845
rect 6391 15832 6409 15845
rect 6461 15832 6479 15845
rect 6531 15832 6549 15845
rect 6601 15832 6619 15845
rect 6671 15832 6689 15845
rect 6741 15832 6759 15845
rect 6811 15832 12534 15845
rect 12586 15849 14937 15850
rect 12586 15832 14103 15849
rect 14155 15832 14201 15849
rect 14253 15832 14298 15849
rect 14350 15832 14395 15849
rect 14447 15832 14937 15849
rect 5230 15798 5240 15832
rect 5303 15798 5306 15832
rect 5522 15798 5561 15832
rect 5595 15798 5634 15832
rect 5668 15798 5707 15832
rect 5741 15798 5780 15832
rect 5814 15798 5853 15832
rect 5887 15798 5926 15832
rect 5960 15798 5999 15832
rect 6033 15798 6072 15832
rect 6106 15798 6145 15832
rect 6179 15798 6198 15832
rect 6252 15798 6269 15832
rect 6325 15798 6339 15832
rect 6398 15798 6409 15832
rect 6471 15798 6479 15832
rect 6544 15798 6549 15832
rect 6617 15798 6619 15832
rect 6836 15798 6875 15832
rect 6909 15798 6948 15832
rect 6982 15798 7021 15832
rect 7055 15798 7094 15832
rect 7128 15798 7167 15832
rect 7201 15798 7240 15832
rect 7274 15798 7313 15832
rect 7347 15798 7386 15832
rect 7420 15798 7459 15832
rect 7493 15798 7532 15832
rect 7566 15798 7605 15832
rect 7639 15798 7678 15832
rect 7712 15798 7751 15832
rect 7785 15798 7824 15832
rect 7858 15798 7897 15832
rect 7931 15798 7970 15832
rect 8004 15798 8043 15832
rect 8077 15798 8116 15832
rect 8150 15798 8189 15832
rect 8223 15798 8262 15832
rect 8296 15798 8335 15832
rect 8369 15798 8408 15832
rect 8442 15798 8481 15832
rect 8515 15798 8554 15832
rect 8588 15798 8627 15832
rect 8661 15798 8699 15832
rect 8733 15798 8771 15832
rect 8805 15798 8843 15832
rect 8877 15798 8915 15832
rect 8949 15798 8987 15832
rect 9021 15798 9059 15832
rect 9093 15798 9131 15832
rect 9165 15798 9203 15832
rect 9237 15798 9275 15832
rect 9309 15798 9347 15832
rect 9381 15798 9419 15832
rect 9453 15798 9491 15832
rect 9525 15798 9563 15832
rect 9597 15798 9635 15832
rect 9669 15798 9707 15832
rect 9741 15798 9779 15832
rect 9813 15798 9851 15832
rect 9885 15798 9923 15832
rect 9957 15798 9995 15832
rect 10029 15798 10067 15832
rect 10101 15798 10139 15832
rect 10173 15798 10211 15832
rect 10245 15798 10283 15832
rect 10317 15798 10355 15832
rect 10389 15798 10427 15832
rect 10461 15798 10499 15832
rect 10533 15798 10571 15832
rect 10605 15798 10643 15832
rect 10677 15798 10715 15832
rect 10749 15798 10787 15832
rect 10821 15798 10859 15832
rect 10893 15798 10931 15832
rect 10965 15798 11003 15832
rect 11037 15798 11075 15832
rect 11109 15798 11147 15832
rect 11181 15798 11219 15832
rect 11253 15798 11291 15832
rect 11325 15798 11363 15832
rect 11397 15798 11435 15832
rect 11469 15798 11507 15832
rect 11541 15798 11579 15832
rect 11613 15798 11651 15832
rect 11685 15798 11723 15832
rect 11757 15798 11795 15832
rect 11829 15798 11867 15832
rect 11901 15798 11939 15832
rect 11973 15798 12011 15832
rect 12045 15798 12083 15832
rect 12117 15798 12155 15832
rect 12189 15798 12227 15832
rect 12261 15798 12299 15832
rect 12333 15798 12371 15832
rect 12405 15798 12443 15832
rect 12477 15798 12515 15832
rect 12586 15798 12587 15832
rect 12621 15798 12659 15832
rect 12693 15798 12731 15832
rect 12765 15798 12803 15832
rect 12837 15798 12875 15832
rect 12909 15798 12947 15832
rect 12981 15798 13019 15832
rect 13053 15798 13091 15832
rect 13125 15798 13163 15832
rect 13197 15798 13235 15832
rect 13269 15798 13307 15832
rect 13341 15798 13379 15832
rect 13413 15798 13451 15832
rect 13485 15798 13523 15832
rect 13557 15798 13595 15832
rect 13629 15798 13667 15832
rect 13701 15798 13739 15832
rect 13773 15798 13811 15832
rect 13845 15798 13883 15832
rect 13917 15798 13955 15832
rect 13989 15798 14027 15832
rect 14061 15798 14099 15832
rect 14155 15798 14171 15832
rect 14277 15798 14298 15832
rect 14350 15798 14387 15832
rect 14447 15798 14459 15832
rect 14493 15798 14531 15832
rect 14565 15798 14603 15832
rect 14637 15798 14675 15832
rect 14709 15798 14747 15832
rect 14781 15798 14819 15832
rect 14853 15798 14891 15832
rect 14925 15798 14937 15832
rect 5226 15793 5240 15798
rect 5292 15793 5306 15798
rect 5358 15793 5372 15798
rect 5424 15793 5438 15798
rect 5490 15793 6198 15798
rect 6250 15793 6269 15798
rect 6321 15793 6339 15798
rect 6391 15793 6409 15798
rect 6461 15793 6479 15798
rect 6531 15793 6549 15798
rect 6601 15793 6619 15798
rect 6671 15793 6689 15798
rect 6741 15793 6759 15798
rect 6811 15797 14103 15798
rect 14155 15797 14201 15798
rect 14253 15797 14298 15798
rect 14350 15797 14395 15798
rect 14447 15797 14937 15798
rect 6811 15793 14937 15797
rect 3870 15792 14937 15793
rect 93 15755 99 15789
rect 133 15755 139 15789
rect 93 15725 139 15755
tri 3574 15737 3580 15743 se
rect 3580 15737 4439 15743
rect 4491 15737 4506 15743
rect 4558 15737 4573 15743
rect 4625 15737 4640 15743
rect 4692 15737 4707 15743
tri 3562 15725 3574 15737 se
rect 3574 15725 3620 15737
rect 56 15719 3620 15725
rect 56 15717 427 15719
rect 56 15683 99 15717
rect 133 15683 171 15717
rect 205 15685 427 15717
rect 461 15685 500 15719
rect 534 15685 573 15719
rect 607 15685 646 15719
rect 680 15685 719 15719
rect 753 15685 792 15719
rect 826 15685 865 15719
rect 899 15685 938 15719
rect 972 15685 1011 15719
rect 1045 15685 1084 15719
rect 1118 15685 1157 15719
rect 1191 15685 1230 15719
rect 1264 15685 1303 15719
rect 1337 15685 1376 15719
rect 1410 15685 1449 15719
rect 1483 15685 1521 15719
rect 1555 15685 1593 15719
rect 1627 15685 1665 15719
rect 1699 15685 1737 15719
rect 1771 15685 1809 15719
rect 1843 15685 1881 15719
rect 1915 15685 1953 15719
rect 1987 15685 2025 15719
rect 2059 15685 2097 15719
rect 2131 15685 2169 15719
rect 2203 15685 2241 15719
rect 2275 15685 2313 15719
rect 2347 15685 2385 15719
rect 2419 15685 2457 15719
rect 2491 15685 2529 15719
rect 2563 15685 2601 15719
rect 2635 15685 2673 15719
rect 2707 15685 2745 15719
rect 2779 15685 2817 15719
rect 2851 15685 2889 15719
rect 2923 15685 2961 15719
rect 2995 15685 3033 15719
rect 3067 15685 3105 15719
rect 3139 15685 3177 15719
rect 3211 15685 3249 15719
rect 3283 15685 3321 15719
rect 3355 15685 3393 15719
rect 3427 15685 3465 15719
rect 3499 15685 3537 15719
rect 3571 15703 3620 15719
rect 3654 15703 3692 15737
rect 3726 15703 3764 15737
rect 3798 15703 3836 15737
rect 3870 15703 3908 15737
rect 3942 15703 3980 15737
rect 4014 15703 4052 15737
rect 4086 15703 4124 15737
rect 4158 15703 4196 15737
rect 4230 15703 4268 15737
rect 4302 15703 4340 15737
rect 4374 15703 4412 15737
rect 4625 15703 4630 15737
rect 4692 15703 4703 15737
rect 3571 15697 4439 15703
rect 3571 15691 3622 15697
tri 3622 15691 3628 15697 nw
tri 4427 15691 4433 15697 ne
rect 4433 15691 4439 15697
rect 4491 15691 4506 15703
rect 4558 15691 4573 15703
rect 4625 15691 4640 15703
rect 4692 15691 4707 15703
rect 4759 15691 4774 15743
rect 4826 15691 4841 15743
rect 4893 15691 4908 15743
rect 4960 15691 4975 15743
rect 5027 15737 5042 15743
rect 5094 15737 5108 15743
rect 5160 15737 5174 15743
rect 5226 15737 5240 15743
rect 5292 15737 5306 15743
rect 5358 15737 5372 15743
rect 5029 15703 5042 15737
rect 5102 15703 5108 15737
rect 5358 15703 5360 15737
rect 5027 15691 5042 15703
rect 5094 15691 5108 15703
rect 5160 15691 5174 15703
rect 5226 15691 5240 15703
rect 5292 15691 5306 15703
rect 5358 15691 5372 15703
rect 5424 15691 5438 15743
rect 5490 15691 5496 15743
tri 5496 15691 5502 15697 nw
tri 6186 15691 6192 15697 ne
rect 6192 15691 6198 15743
rect 6250 15691 6269 15743
rect 6321 15691 6339 15743
rect 6391 15691 6409 15743
rect 6461 15691 6479 15743
rect 6531 15691 6549 15743
rect 6601 15691 6619 15743
rect 6671 15691 6689 15743
rect 6741 15691 6759 15743
rect 6811 15691 6817 15743
rect 12534 15737 12586 15743
tri 6817 15691 6823 15697 nw
rect 3571 15685 3610 15691
rect 205 15683 3610 15685
rect 56 15679 3610 15683
tri 3610 15679 3622 15691 nw
tri 5359 15679 5371 15691 ne
rect 5371 15679 5436 15691
rect 56 15660 650 15679
tri 650 15660 669 15679 nw
tri 5371 15660 5390 15679 ne
rect 56 15647 637 15660
tri 637 15647 650 15660 nw
rect 5390 15647 5436 15679
rect 56 15639 616 15647
rect 56 15605 69 15639
rect 103 15605 153 15639
rect 187 15605 237 15639
rect 271 15605 321 15639
rect 355 15605 405 15639
rect 439 15626 616 15639
tri 616 15626 637 15647 nw
rect 439 15616 603 15626
rect 439 15605 481 15616
rect 56 15582 481 15605
rect 515 15613 603 15616
tri 603 15613 616 15626 nw
rect 5390 15613 5396 15647
rect 5430 15613 5436 15647
rect 515 15582 559 15613
rect 56 15569 559 15582
tri 559 15569 603 15613 nw
rect 5390 15569 5436 15613
rect 56 15562 552 15569
tri 552 15562 559 15569 nw
rect 56 15528 69 15562
rect 103 15528 153 15562
rect 187 15528 237 15562
rect 271 15528 321 15562
rect 355 15528 405 15562
rect 439 15541 530 15562
rect 439 15528 481 15541
rect 56 15507 481 15528
rect 515 15540 530 15541
tri 530 15540 552 15562 nw
rect 515 15535 525 15540
tri 525 15535 530 15540 nw
rect 5390 15535 5396 15569
rect 5430 15535 5436 15569
rect 515 15507 523 15535
tri 523 15533 525 15535 nw
tri 3981 15520 3983 15522 se
rect 3983 15520 5280 15522
tri 3975 15514 3981 15520 se
rect 3981 15514 5280 15520
rect 56 15485 523 15507
rect 56 15451 69 15485
rect 103 15451 153 15485
rect 187 15451 237 15485
rect 271 15451 321 15485
rect 355 15451 405 15485
rect 439 15466 523 15485
rect 439 15451 481 15466
rect 56 15432 481 15451
rect 515 15432 523 15466
rect 56 15408 523 15432
rect 56 15374 69 15408
rect 103 15374 153 15408
rect 187 15374 237 15408
rect 271 15374 321 15408
rect 355 15374 405 15408
rect 439 15391 523 15408
rect 439 15374 481 15391
rect 56 15357 481 15374
rect 515 15357 523 15391
rect 56 15331 523 15357
rect 56 15297 69 15331
rect 103 15297 153 15331
rect 187 15297 237 15331
rect 271 15297 321 15331
rect 355 15297 405 15331
rect 439 15316 523 15331
rect 439 15297 481 15316
rect 56 15282 481 15297
rect 515 15282 523 15316
rect 56 15254 523 15282
rect 56 15220 69 15254
rect 103 15220 153 15254
rect 187 15220 237 15254
rect 271 15220 321 15254
rect 355 15220 405 15254
rect 439 15241 523 15254
rect 439 15220 481 15241
rect 56 15207 481 15220
rect 515 15207 523 15241
rect 56 15177 523 15207
rect 56 15143 69 15177
rect 103 15143 153 15177
rect 187 15143 237 15177
rect 271 15143 321 15177
rect 355 15143 405 15177
rect 439 15166 523 15177
rect 439 15143 481 15166
rect 56 15132 481 15143
rect 515 15132 523 15166
rect 56 15100 523 15132
rect 56 15066 69 15100
rect 103 15066 153 15100
rect 187 15066 237 15100
rect 271 15066 321 15100
rect 355 15066 405 15100
rect 439 15091 523 15100
rect 439 15066 481 15091
rect 56 15057 481 15066
rect 515 15057 523 15091
rect 56 15022 523 15057
rect 56 14988 69 15022
rect 103 14988 153 15022
rect 187 14988 237 15022
rect 271 14988 321 15022
rect 355 14988 405 15022
rect 439 15016 523 15022
rect 439 14988 481 15016
rect 56 14982 481 14988
rect 515 14982 523 15016
rect 56 14944 523 14982
rect 56 14910 69 14944
rect 103 14910 153 14944
rect 187 14910 237 14944
rect 271 14910 321 14944
rect 355 14910 405 14944
rect 439 14941 523 14944
rect 439 14910 481 14941
rect 56 14907 481 14910
rect 515 14925 523 14941
rect 616 15513 5280 15514
rect 616 15508 4591 15513
rect 616 15474 694 15508
rect 728 15474 766 15508
rect 800 15474 838 15508
rect 872 15474 910 15508
rect 944 15474 982 15508
rect 1016 15474 1054 15508
rect 1088 15474 1126 15508
rect 1160 15474 1198 15508
rect 1232 15474 1270 15508
rect 1304 15474 1342 15508
rect 1376 15474 1414 15508
rect 1448 15474 1486 15508
rect 1520 15474 1558 15508
rect 1592 15474 1630 15508
rect 1664 15474 1702 15508
rect 1736 15474 1774 15508
rect 1808 15474 1846 15508
rect 1880 15474 1918 15508
rect 1952 15474 1990 15508
rect 2024 15474 2062 15508
rect 2096 15474 2134 15508
rect 2168 15474 2206 15508
rect 2240 15474 2278 15508
rect 2312 15474 2350 15508
rect 2384 15474 2422 15508
rect 2456 15474 2494 15508
rect 2528 15474 2566 15508
rect 2600 15474 2638 15508
rect 2672 15474 2710 15508
rect 2744 15474 2782 15508
rect 2816 15474 2854 15508
rect 2888 15474 2926 15508
rect 2960 15474 2998 15508
rect 3032 15474 3070 15508
rect 3104 15474 3142 15508
rect 3176 15474 3214 15508
rect 3248 15474 3286 15508
rect 3320 15474 3358 15508
rect 3392 15474 3430 15508
rect 3464 15474 3502 15508
rect 3536 15474 3574 15508
rect 3608 15474 3646 15508
rect 3680 15474 3718 15508
rect 3752 15474 3790 15508
rect 3824 15474 3862 15508
rect 3896 15474 3935 15508
rect 3969 15504 4591 15508
rect 4643 15504 4658 15513
rect 4710 15504 4725 15513
rect 4777 15504 4792 15513
rect 3969 15474 4017 15504
rect 616 15470 4017 15474
rect 4051 15470 4094 15504
rect 4128 15470 4171 15504
rect 4205 15470 4248 15504
rect 4282 15470 4325 15504
rect 4359 15470 4402 15504
rect 4436 15470 4479 15504
rect 4513 15470 4556 15504
rect 4590 15470 4591 15504
rect 4777 15470 4784 15504
rect 616 15461 4591 15470
rect 4643 15461 4658 15470
rect 4710 15461 4725 15470
rect 4777 15461 4792 15470
rect 4844 15461 4859 15513
rect 4911 15461 4926 15513
rect 4978 15461 4993 15513
rect 5045 15504 5059 15513
rect 5111 15504 5280 15513
rect 5046 15470 5059 15504
rect 5122 15470 5164 15504
rect 5198 15470 5280 15504
rect 5045 15461 5059 15470
rect 5111 15461 5280 15470
rect 616 15452 5280 15461
rect 616 15444 4045 15452
tri 4045 15444 4053 15452 nw
tri 5176 15444 5184 15452 ne
rect 5184 15444 5280 15452
rect 616 15436 4019 15444
rect 616 15402 622 15436
rect 656 15420 4019 15436
rect 656 15402 710 15420
rect 616 15386 710 15402
rect 744 15386 783 15420
rect 817 15386 856 15420
rect 890 15386 929 15420
rect 963 15386 1002 15420
rect 1036 15386 1075 15420
rect 1109 15386 1148 15420
rect 1182 15386 1221 15420
rect 1255 15386 1294 15420
rect 1328 15386 1367 15420
rect 1401 15386 1440 15420
rect 1474 15386 1513 15420
rect 1547 15386 1586 15420
rect 1620 15386 1659 15420
rect 1693 15386 1732 15420
rect 1766 15386 1805 15420
rect 1839 15386 1878 15420
rect 1912 15386 1951 15420
rect 1985 15386 2024 15420
rect 2058 15386 2097 15420
rect 2131 15386 2170 15420
rect 2204 15386 2243 15420
rect 2277 15386 2316 15420
rect 2350 15386 2389 15420
rect 2423 15386 2462 15420
rect 2496 15386 2535 15420
rect 2569 15386 2608 15420
rect 2642 15386 2681 15420
rect 2715 15386 2754 15420
rect 2788 15386 2827 15420
rect 2861 15386 2900 15420
rect 2934 15386 2973 15420
rect 3007 15386 3047 15420
rect 3081 15386 3121 15420
rect 3155 15386 3195 15420
rect 3229 15386 3269 15420
rect 3303 15386 3343 15420
rect 3377 15386 3417 15420
rect 3451 15386 3491 15420
rect 3525 15386 3565 15420
rect 3599 15386 3639 15420
rect 3673 15386 3713 15420
rect 3747 15386 3787 15420
rect 3821 15386 3861 15420
rect 3895 15386 3935 15420
rect 3969 15418 4019 15420
tri 4019 15418 4045 15444 nw
tri 5184 15418 5210 15444 ne
rect 3969 15410 4011 15418
tri 4011 15410 4019 15418 nw
rect 5210 15410 5228 15444
rect 5262 15410 5280 15444
rect 3969 15404 4005 15410
tri 4005 15404 4011 15410 nw
rect 3969 15397 3998 15404
tri 3998 15397 4005 15404 nw
rect 3969 15391 3992 15397
tri 3992 15391 3998 15397 nw
rect 4199 15391 5090 15397
rect 3969 15386 3983 15391
rect 616 15382 3983 15386
tri 3983 15382 3992 15391 nw
rect 616 15380 3981 15382
tri 3981 15380 3983 15382 nw
rect 616 15362 834 15380
rect 616 15328 622 15362
rect 656 15357 834 15362
tri 834 15357 857 15380 nw
rect 4199 15357 4211 15391
rect 4245 15357 4287 15391
rect 4321 15357 4363 15391
rect 4397 15357 4439 15391
rect 4473 15357 4515 15391
rect 4549 15357 4591 15391
rect 4625 15381 4667 15391
rect 4701 15381 4743 15391
rect 4777 15381 4819 15391
rect 4853 15381 4894 15391
rect 4928 15381 4969 15391
rect 5003 15381 5044 15391
rect 4654 15357 4667 15381
rect 4739 15357 4743 15381
rect 4853 15357 4856 15381
rect 4928 15357 4940 15381
rect 5003 15357 5024 15381
rect 5078 15357 5090 15391
rect 656 15338 815 15357
tri 815 15338 834 15357 nw
rect 656 15337 812 15338
rect 656 15328 710 15337
rect 616 15303 710 15328
rect 744 15335 812 15337
tri 812 15335 815 15338 nw
rect 744 15311 788 15335
tri 788 15311 812 15335 nw
rect 4199 15329 4602 15357
rect 4654 15329 4687 15357
rect 4739 15329 4772 15357
rect 4824 15329 4856 15357
rect 4908 15329 4940 15357
rect 4992 15329 5024 15357
rect 5076 15329 5090 15357
rect 744 15305 782 15311
tri 782 15305 788 15311 nw
rect 875 15305 1942 15311
rect 1994 15305 2006 15311
rect 2058 15305 3616 15311
rect 3668 15305 3680 15311
rect 3732 15305 4126 15311
rect 744 15303 750 15305
rect 616 15288 750 15303
rect 616 15254 622 15288
rect 656 15254 750 15288
tri 750 15273 782 15305 nw
rect 875 15271 887 15305
rect 921 15271 959 15305
rect 993 15271 1031 15305
rect 1065 15271 1103 15305
rect 1137 15271 1175 15305
rect 1209 15271 1247 15305
rect 1281 15271 1319 15305
rect 1353 15271 1391 15305
rect 1425 15271 1463 15305
rect 1497 15271 1535 15305
rect 1569 15271 1607 15305
rect 1641 15271 1679 15305
rect 1713 15271 1751 15305
rect 1785 15271 1823 15305
rect 1857 15271 1895 15305
rect 1929 15271 1942 15305
rect 2001 15271 2006 15305
rect 2073 15271 2111 15305
rect 2145 15271 2183 15305
rect 2217 15271 2256 15305
rect 2290 15271 2329 15305
rect 2363 15271 2402 15305
rect 2436 15271 2483 15305
rect 2517 15271 2555 15305
rect 2589 15271 2627 15305
rect 2661 15271 2699 15305
rect 2733 15271 2771 15305
rect 2805 15271 2843 15305
rect 2877 15271 2915 15305
rect 2949 15271 2987 15305
rect 3021 15271 3059 15305
rect 3093 15271 3131 15305
rect 3165 15271 3204 15305
rect 3238 15271 3277 15305
rect 3311 15271 3350 15305
rect 3384 15271 3423 15305
rect 3457 15271 3496 15305
rect 3530 15271 3569 15305
rect 3603 15271 3616 15305
rect 3676 15271 3680 15305
rect 3749 15271 3788 15305
rect 3822 15271 3861 15305
rect 3895 15271 3934 15305
rect 3968 15271 4007 15305
rect 4041 15271 4080 15305
rect 4114 15271 4126 15305
rect 875 15265 1942 15271
tri 1930 15259 1936 15265 ne
rect 1936 15259 1942 15265
rect 1994 15259 2006 15271
rect 2058 15265 3616 15271
rect 2058 15259 2064 15265
tri 2064 15259 2070 15265 nw
tri 3604 15259 3610 15265 ne
rect 3610 15259 3616 15265
rect 3668 15259 3680 15271
rect 3732 15265 4126 15271
rect 4199 15265 5090 15329
rect 3732 15259 3738 15265
tri 3738 15259 3744 15265 nw
rect 616 15220 710 15254
rect 744 15220 750 15254
rect 616 15214 750 15220
rect 616 15180 622 15214
rect 656 15180 750 15214
tri 2475 15209 2481 15215 se
rect 2481 15209 2487 15215
rect 616 15171 750 15180
rect 616 15140 710 15171
rect 616 15106 622 15140
rect 656 15137 710 15140
rect 744 15137 750 15171
rect 1820 15203 2487 15209
rect 1820 15169 1832 15203
rect 1866 15169 1906 15203
rect 1940 15169 1980 15203
rect 2014 15169 2054 15203
rect 2088 15169 2128 15203
rect 2162 15169 2202 15203
rect 2236 15169 2276 15203
rect 2310 15169 2350 15203
rect 2384 15169 2424 15203
rect 2458 15169 2487 15203
rect 1820 15163 2487 15169
rect 2539 15163 2551 15215
rect 2603 15209 2609 15215
tri 2609 15209 2615 15215 sw
rect 4199 15213 4602 15265
rect 4654 15213 4687 15265
rect 4739 15213 4772 15265
rect 4824 15213 4856 15265
rect 4908 15213 4940 15265
rect 4992 15213 5024 15265
rect 5076 15213 5090 15265
rect 2603 15203 4091 15209
rect 2606 15169 2646 15203
rect 2680 15169 2720 15203
rect 2754 15169 2794 15203
rect 2828 15169 2868 15203
rect 2902 15169 2942 15203
rect 2976 15169 3016 15203
rect 3050 15169 3090 15203
rect 3124 15169 3164 15203
rect 3198 15169 3238 15203
rect 3272 15169 3312 15203
rect 3346 15169 3386 15203
rect 3420 15169 3460 15203
rect 3494 15169 3534 15203
rect 3568 15169 3607 15203
rect 3641 15169 3680 15203
rect 3714 15169 3753 15203
rect 3787 15169 3826 15203
rect 3860 15169 3899 15203
rect 3933 15169 3972 15203
rect 4006 15169 4045 15203
rect 4079 15169 4091 15203
rect 2603 15163 4091 15169
rect 656 15106 750 15137
rect 4199 15149 5090 15213
rect 4199 15136 4602 15149
rect 4654 15136 4687 15149
rect 4739 15136 4772 15149
rect 4824 15136 4856 15149
rect 4908 15136 4940 15149
rect 4992 15136 5024 15149
rect 5076 15136 5090 15149
rect 616 15102 750 15106
tri 750 15102 768 15120 sw
rect 4199 15102 4211 15136
rect 4245 15102 4287 15136
rect 4321 15102 4363 15136
rect 4397 15102 4439 15136
rect 4473 15102 4515 15136
rect 4549 15102 4591 15136
rect 4654 15102 4667 15136
rect 4739 15102 4743 15136
rect 4853 15102 4856 15136
rect 4928 15102 4940 15136
rect 5003 15102 5024 15136
rect 5078 15102 5090 15136
rect 616 15101 768 15102
tri 768 15101 769 15102 sw
rect 616 15096 769 15101
tri 769 15096 774 15101 sw
rect 4199 15097 4602 15102
rect 4654 15097 4687 15102
rect 4739 15097 4772 15102
rect 4824 15097 4856 15102
rect 4908 15097 4940 15102
rect 4992 15097 5024 15102
rect 5076 15097 5090 15102
rect 4199 15096 5090 15097
rect 5210 15372 5280 15410
rect 5210 15338 5228 15372
rect 5262 15338 5280 15372
rect 5210 15300 5280 15338
rect 5210 15266 5228 15300
rect 5262 15266 5280 15300
rect 5210 15228 5280 15266
rect 5210 15194 5228 15228
rect 5262 15194 5280 15228
rect 5210 15156 5280 15194
rect 5210 15122 5228 15156
rect 5262 15122 5280 15156
rect 616 15089 774 15096
rect 616 15066 710 15089
rect 616 15032 622 15066
rect 656 15055 710 15066
rect 744 15076 774 15089
tri 774 15076 794 15096 sw
rect 744 15067 794 15076
tri 794 15067 803 15076 sw
tri 5201 15067 5210 15076 se
rect 5210 15067 5280 15122
rect 744 15055 803 15067
rect 656 15054 803 15055
tri 803 15054 816 15067 sw
tri 5188 15054 5201 15067 se
rect 5201 15054 5280 15067
rect 656 15042 816 15054
tri 816 15042 828 15054 sw
tri 5176 15042 5188 15054 se
rect 5188 15042 5280 15054
rect 656 15032 828 15042
rect 616 15024 828 15032
tri 828 15024 846 15042 sw
tri 2322 15024 2340 15042 se
rect 2340 15024 5280 15042
rect 616 15013 846 15024
tri 846 15013 857 15024 sw
tri 2311 15013 2322 15024 se
rect 2322 15013 2465 15024
rect 616 15007 2465 15013
rect 616 14992 710 15007
rect 616 14958 622 14992
rect 656 14973 710 14992
rect 744 14973 783 15007
rect 817 14973 856 15007
rect 890 14973 929 15007
rect 963 14973 1002 15007
rect 1036 14973 1075 15007
rect 1109 14973 1148 15007
rect 1182 14973 1221 15007
rect 1255 14973 1294 15007
rect 1328 14973 1367 15007
rect 1401 14973 1440 15007
rect 1474 14973 1513 15007
rect 1547 14973 1586 15007
rect 1620 14973 1659 15007
rect 1693 14973 1732 15007
rect 1766 14973 1805 15007
rect 1839 14973 1878 15007
rect 1912 14973 1950 15007
rect 1984 14973 2022 15007
rect 2056 14973 2094 15007
rect 2128 14973 2166 15007
rect 2200 14973 2238 15007
rect 2272 14973 2310 15007
rect 2344 14990 2465 15007
rect 2499 14990 2538 15024
rect 2572 14990 2611 15024
rect 2645 14990 2684 15024
rect 2718 14990 2757 15024
rect 2791 14990 2830 15024
rect 2864 14990 2903 15024
rect 2937 14990 2976 15024
rect 3010 14990 3049 15024
rect 3083 14990 3122 15024
rect 3156 14990 3195 15024
rect 3229 14990 3268 15024
rect 3302 14990 3341 15024
rect 3375 14990 3414 15024
rect 3448 14990 3487 15024
rect 3521 14990 3560 15024
rect 3594 14990 3633 15024
rect 3667 14990 3706 15024
rect 3740 14990 3779 15024
rect 3813 14990 3852 15024
rect 3886 14990 3925 15024
rect 3959 14990 3998 15024
rect 4032 14990 4071 15024
rect 4105 14990 4144 15024
rect 4178 14990 4217 15024
rect 4251 14990 4290 15024
rect 4324 14990 4363 15024
rect 4397 14990 4436 15024
rect 4470 14990 4509 15024
rect 4543 14990 4582 15024
rect 4616 14990 4655 15024
rect 4689 14990 4728 15024
rect 4762 14990 4801 15024
rect 4835 14990 4874 15024
rect 4908 14990 4947 15024
rect 4981 14990 5020 15024
rect 5054 14990 5094 15024
rect 5128 14990 5168 15024
rect 5202 14990 5280 15024
rect 2344 14973 5280 14990
rect 656 14972 5280 14973
rect 5390 15491 5436 15535
rect 5390 15457 5396 15491
rect 5430 15457 5436 15491
rect 5390 15413 5436 15457
rect 5390 15379 5396 15413
rect 5430 15379 5436 15413
rect 5390 15335 5436 15379
rect 5390 15301 5396 15335
rect 5430 15301 5436 15335
rect 12534 15667 12586 15685
rect 12534 15597 12586 15615
rect 12534 15527 12586 15545
rect 12534 15457 12586 15475
rect 12534 15386 12586 15405
rect 12534 15328 12586 15334
rect 12848 15464 14894 15470
rect 12848 15430 12860 15464
rect 12894 15430 12934 15464
rect 12968 15430 13008 15464
rect 13042 15430 13082 15464
rect 13116 15430 13156 15464
rect 13190 15430 13230 15464
rect 13264 15430 13304 15464
rect 13338 15430 13378 15464
rect 13412 15430 13452 15464
rect 13486 15430 13526 15464
rect 13560 15430 13600 15464
rect 13634 15430 13674 15464
rect 13708 15430 13748 15464
rect 13782 15430 13822 15464
rect 13856 15430 13896 15464
rect 13930 15430 13970 15464
rect 14004 15430 14044 15464
rect 14078 15459 14118 15464
rect 14152 15459 14191 15464
rect 14225 15459 14264 15464
rect 14298 15459 14337 15464
rect 14371 15459 14410 15464
rect 14444 15459 14483 15464
rect 14078 15430 14101 15459
rect 12848 15407 14101 15430
rect 14153 15407 14175 15459
rect 14227 15407 14249 15459
rect 14301 15407 14323 15459
rect 14375 15407 14397 15459
rect 14449 15430 14483 15459
rect 14517 15430 14556 15464
rect 14590 15430 14629 15464
rect 14663 15430 14702 15464
rect 14736 15430 14775 15464
rect 14809 15430 14848 15464
rect 14882 15430 14894 15464
rect 14449 15407 14894 15430
rect 12848 15394 14894 15407
rect 12848 15382 14101 15394
rect 12848 15348 12860 15382
rect 12894 15348 12934 15382
rect 12968 15348 13008 15382
rect 13042 15348 13082 15382
rect 13116 15348 13156 15382
rect 13190 15348 13230 15382
rect 13264 15348 13304 15382
rect 13338 15348 13378 15382
rect 13412 15348 13452 15382
rect 13486 15348 13526 15382
rect 13560 15348 13600 15382
rect 13634 15348 13674 15382
rect 13708 15348 13748 15382
rect 13782 15348 13822 15382
rect 13856 15348 13896 15382
rect 13930 15348 13970 15382
rect 14004 15348 14044 15382
rect 14078 15348 14101 15382
rect 12848 15342 14101 15348
rect 14153 15342 14175 15394
rect 14227 15342 14249 15394
rect 14301 15342 14323 15394
rect 14375 15342 14397 15394
rect 14449 15382 14894 15394
rect 14449 15348 14483 15382
rect 14517 15348 14556 15382
rect 14590 15348 14629 15382
rect 14663 15348 14702 15382
rect 14736 15348 14775 15382
rect 14809 15348 14848 15382
rect 14882 15348 14894 15382
rect 14449 15342 14894 15348
rect 12848 15328 14894 15342
tri 12534 15322 12540 15328 ne
rect 5390 15257 5436 15301
tri 8177 15259 8183 15265 ne
rect 8183 15259 8189 15311
rect 8241 15259 8255 15311
rect 8307 15259 8313 15311
tri 8313 15259 8319 15265 nw
tri 9849 15259 9855 15265 ne
rect 9855 15259 9861 15311
rect 9913 15259 9927 15311
rect 9979 15259 9985 15311
rect 12848 15300 14101 15328
rect 12848 15266 12860 15300
rect 12894 15266 12934 15300
rect 12968 15266 13008 15300
rect 13042 15266 13082 15300
rect 13116 15266 13156 15300
rect 13190 15266 13230 15300
rect 13264 15266 13304 15300
rect 13338 15266 13378 15300
rect 13412 15266 13452 15300
rect 13486 15266 13526 15300
rect 13560 15266 13600 15300
rect 13634 15266 13674 15300
rect 13708 15266 13748 15300
rect 13782 15266 13822 15300
rect 13856 15266 13896 15300
rect 13930 15266 13970 15300
rect 14004 15266 14044 15300
rect 14078 15276 14101 15300
rect 14153 15276 14175 15328
rect 14227 15276 14249 15328
rect 14301 15276 14323 15328
rect 14375 15276 14397 15328
rect 14449 15300 14894 15328
rect 14449 15276 14483 15300
rect 14078 15266 14118 15276
rect 14152 15266 14191 15276
rect 14225 15266 14264 15276
rect 14298 15266 14337 15276
rect 14371 15266 14410 15276
rect 14444 15266 14483 15276
rect 14517 15266 14556 15300
rect 14590 15266 14629 15300
rect 14663 15266 14702 15300
rect 14736 15266 14775 15300
rect 14809 15266 14848 15300
rect 14882 15266 14894 15300
tri 9985 15259 9991 15265 nw
rect 12848 15262 14894 15266
rect 5390 15223 5396 15257
rect 5430 15223 5436 15257
rect 5390 15179 5436 15223
rect 12848 15218 14101 15262
tri 9654 15209 9660 15215 se
rect 5390 15145 5396 15179
rect 5430 15145 5436 15179
rect 9660 15163 9666 15215
rect 9718 15163 9730 15215
rect 9782 15163 9788 15215
tri 9788 15209 9794 15215 sw
rect 12848 15184 12860 15218
rect 12894 15184 12934 15218
rect 12968 15184 13008 15218
rect 13042 15184 13082 15218
rect 13116 15184 13156 15218
rect 13190 15184 13230 15218
rect 13264 15184 13304 15218
rect 13338 15184 13378 15218
rect 13412 15184 13452 15218
rect 13486 15184 13526 15218
rect 13560 15184 13600 15218
rect 13634 15184 13674 15218
rect 13708 15184 13748 15218
rect 13782 15184 13822 15218
rect 13856 15184 13896 15218
rect 13930 15184 13970 15218
rect 14004 15184 14044 15218
rect 14078 15210 14101 15218
rect 14153 15210 14175 15262
rect 14227 15210 14249 15262
rect 14301 15210 14323 15262
rect 14375 15210 14397 15262
rect 14449 15218 14894 15262
rect 14449 15210 14483 15218
rect 14078 15196 14118 15210
rect 14152 15196 14191 15210
rect 14225 15196 14264 15210
rect 14298 15196 14337 15210
rect 14371 15196 14410 15210
rect 14444 15196 14483 15210
rect 14078 15184 14101 15196
rect 5390 15101 5436 15145
rect 5390 15067 5396 15101
rect 5430 15067 5436 15101
rect 5390 15023 5436 15067
rect 5390 14989 5396 15023
rect 5430 14989 5436 15023
rect 656 14958 2491 14972
rect 616 14945 2491 14958
tri 2491 14945 2518 14972 nw
rect 5390 14945 5436 14989
tri 523 14925 530 14932 sw
rect 515 14919 530 14925
tri 530 14919 536 14925 sw
rect 616 14919 2457 14945
rect 515 14907 536 14919
rect 56 14903 536 14907
tri 536 14903 552 14919 sw
rect 56 14885 552 14903
tri 552 14885 570 14903 sw
rect 616 14885 694 14919
rect 728 14885 768 14919
rect 802 14885 842 14919
rect 876 14885 916 14919
rect 950 14885 990 14919
rect 1024 14885 1064 14919
rect 1098 14885 1138 14919
rect 1172 14885 1212 14919
rect 1246 14885 1286 14919
rect 1320 14885 1360 14919
rect 1394 14885 1434 14919
rect 1468 14885 1507 14919
rect 1541 14885 1580 14919
rect 1614 14885 1653 14919
rect 1687 14885 1726 14919
rect 1760 14885 1799 14919
rect 1833 14885 1872 14919
rect 1906 14885 1945 14919
rect 1979 14885 2018 14919
rect 2052 14885 2091 14919
rect 2125 14885 2164 14919
rect 2198 14885 2237 14919
rect 2271 14885 2310 14919
rect 2344 14911 2457 14919
tri 2457 14911 2491 14945 nw
rect 5390 14911 5396 14945
rect 5430 14911 5436 14945
rect 12848 15144 14101 15184
rect 14153 15144 14175 15196
rect 14227 15144 14249 15196
rect 14301 15144 14323 15196
rect 14375 15144 14397 15196
rect 14449 15184 14483 15196
rect 14517 15184 14556 15218
rect 14590 15184 14629 15218
rect 14663 15184 14702 15218
rect 14736 15184 14775 15218
rect 14809 15184 14848 15218
rect 14882 15184 14894 15218
rect 14449 15144 14894 15184
rect 12848 15136 14894 15144
rect 12848 15102 12860 15136
rect 12894 15102 12934 15136
rect 12968 15102 13008 15136
rect 13042 15102 13082 15136
rect 13116 15102 13156 15136
rect 13190 15102 13230 15136
rect 13264 15102 13304 15136
rect 13338 15102 13378 15136
rect 13412 15102 13452 15136
rect 13486 15102 13526 15136
rect 13560 15102 13600 15136
rect 13634 15102 13674 15136
rect 13708 15102 13748 15136
rect 13782 15102 13822 15136
rect 13856 15102 13896 15136
rect 13930 15102 13970 15136
rect 14004 15102 14044 15136
rect 14078 15130 14118 15136
rect 14152 15130 14191 15136
rect 14225 15130 14264 15136
rect 14298 15130 14337 15136
rect 14371 15130 14410 15136
rect 14444 15130 14483 15136
rect 14078 15102 14101 15130
rect 12848 15078 14101 15102
rect 14153 15078 14175 15130
rect 14227 15078 14249 15130
rect 14301 15078 14323 15130
rect 14375 15078 14397 15130
rect 14449 15102 14483 15130
rect 14517 15102 14556 15136
rect 14590 15102 14629 15136
rect 14663 15102 14702 15136
rect 14736 15102 14775 15136
rect 14809 15102 14848 15136
rect 14882 15102 14894 15136
rect 14449 15078 14894 15102
rect 12848 15064 14894 15078
rect 12848 15054 14101 15064
rect 12848 15020 12860 15054
rect 12894 15020 12934 15054
rect 12968 15020 13008 15054
rect 13042 15020 13082 15054
rect 13116 15020 13156 15054
rect 13190 15020 13230 15054
rect 13264 15020 13304 15054
rect 13338 15020 13378 15054
rect 13412 15020 13452 15054
rect 13486 15020 13526 15054
rect 13560 15020 13600 15054
rect 13634 15020 13674 15054
rect 13708 15020 13748 15054
rect 13782 15020 13822 15054
rect 13856 15020 13896 15054
rect 13930 15020 13970 15054
rect 14004 15020 14044 15054
rect 14078 15020 14101 15054
rect 12848 15012 14101 15020
rect 14153 15012 14175 15064
rect 14227 15012 14249 15064
rect 14301 15012 14323 15064
rect 14375 15012 14397 15064
rect 14449 15054 14894 15064
rect 14449 15020 14483 15054
rect 14517 15020 14556 15054
rect 14590 15020 14629 15054
rect 14663 15020 14702 15054
rect 14736 15020 14775 15054
rect 14809 15020 14848 15054
rect 14882 15020 14894 15054
rect 14449 15012 14894 15020
rect 12848 14998 14894 15012
rect 12848 14972 14101 14998
rect 12848 14938 12860 14972
rect 12894 14938 12934 14972
rect 12968 14938 13008 14972
rect 13042 14938 13082 14972
rect 13116 14938 13156 14972
rect 13190 14938 13230 14972
rect 13264 14938 13304 14972
rect 13338 14938 13378 14972
rect 13412 14938 13452 14972
rect 13486 14938 13526 14972
rect 13560 14938 13600 14972
rect 13634 14938 13674 14972
rect 13708 14938 13748 14972
rect 13782 14938 13822 14972
rect 13856 14938 13896 14972
rect 13930 14938 13970 14972
rect 14004 14938 14044 14972
rect 14078 14946 14101 14972
rect 14153 14946 14175 14998
rect 14227 14946 14249 14998
rect 14301 14946 14323 14998
rect 14375 14946 14397 14998
rect 14449 14972 14894 14998
rect 14449 14946 14483 14972
rect 14078 14938 14118 14946
rect 14152 14938 14191 14946
rect 14225 14938 14264 14946
rect 14298 14938 14337 14946
rect 14371 14938 14410 14946
rect 14444 14938 14483 14946
rect 14517 14938 14556 14972
rect 14590 14938 14629 14972
rect 14663 14938 14702 14972
rect 14736 14938 14775 14972
rect 14809 14938 14848 14972
rect 14882 14938 14894 14972
rect 12848 14932 14894 14938
rect 2344 14885 2425 14911
rect 56 14879 570 14885
tri 570 14879 576 14885 sw
rect 616 14879 2425 14885
tri 2425 14879 2457 14911 nw
rect 56 14867 576 14879
tri 576 14867 588 14879 sw
rect 5390 14867 5436 14911
rect 56 14866 481 14867
rect 56 14832 69 14866
rect 103 14832 153 14866
rect 187 14832 237 14866
rect 271 14832 321 14866
rect 355 14832 405 14866
rect 439 14833 481 14866
rect 515 14839 588 14867
tri 588 14839 616 14867 sw
tri 5362 14839 5390 14867 se
rect 5390 14839 5396 14867
rect 515 14836 616 14839
tri 616 14836 619 14839 sw
tri 5359 14836 5362 14839 se
rect 5362 14836 5396 14839
rect 515 14833 619 14836
tri 619 14833 622 14836 sw
tri 5356 14833 5359 14836 se
rect 5359 14833 5396 14836
rect 5430 14833 5436 14867
rect 439 14832 622 14833
rect 56 14830 622 14832
tri 622 14830 625 14833 sw
tri 5353 14830 5356 14833 se
rect 5356 14830 5436 14833
rect 56 14789 625 14830
tri 625 14789 666 14830 sw
tri 5312 14789 5353 14830 se
rect 5353 14789 5436 14830
tri 344 14767 366 14789 se
rect 366 14782 530 14789
tri 530 14782 537 14789 sw
rect 1861 14783 2007 14789
rect 366 14767 726 14782
rect 344 14739 726 14767
rect 526 14681 726 14739
rect 1913 14731 1955 14783
tri 5290 14767 5312 14789 se
rect 5312 14767 5436 14789
rect 5290 14739 5436 14767
rect 14095 14788 14455 14789
rect 1861 14714 2007 14731
rect 1913 14662 1955 14714
rect 1861 14645 2007 14662
rect 1913 14593 1955 14645
rect 1861 14587 2007 14593
rect 14095 14736 14101 14788
rect 14153 14736 14175 14788
rect 14227 14736 14249 14788
rect 14301 14736 14323 14788
rect 14375 14736 14397 14788
rect 14449 14736 14455 14788
rect 14095 14714 14455 14736
rect 14095 14662 14101 14714
rect 14153 14662 14175 14714
rect 14227 14662 14249 14714
rect 14301 14662 14323 14714
rect 14375 14662 14397 14714
rect 14449 14662 14455 14714
rect 14095 14640 14455 14662
rect 14095 14588 14101 14640
rect 14153 14588 14175 14640
rect 14227 14588 14249 14640
rect 14301 14588 14323 14640
rect 14375 14588 14397 14640
rect 14449 14588 14455 14640
rect 14095 14587 14455 14588
rect 870 13850 1790 13857
rect 870 13798 876 13850
rect 928 13798 942 13850
rect 994 13798 1790 13850
rect 870 13786 1790 13798
rect 870 13734 876 13786
rect 928 13734 942 13786
rect 994 13734 1790 13786
rect 870 13727 1790 13734
rect 2220 13805 2226 13857
rect 2278 13805 2292 13857
rect 2344 13805 2350 13857
rect 2220 13779 2350 13805
rect 2220 13727 2226 13779
rect 2278 13727 2292 13779
rect 2344 13727 2350 13779
rect 2782 13850 2912 13857
rect 2782 13798 2788 13850
rect 2840 13798 2854 13850
rect 2906 13798 2912 13850
rect 2782 13786 2912 13798
rect 2782 13734 2788 13786
rect 2840 13734 2854 13786
rect 2906 13734 2912 13786
rect 2782 13727 2912 13734
rect 3342 13727 3842 13857
rect 3895 13850 4274 13857
rect 3895 13798 3901 13850
rect 3953 13798 3980 13850
rect 4032 13798 4059 13850
rect 4111 13798 4138 13850
rect 4190 13798 4216 13850
rect 4268 13798 4274 13850
rect 3895 13786 4274 13798
rect 3895 13734 3901 13786
rect 3953 13734 3980 13786
rect 4032 13734 4059 13786
rect 4111 13734 4138 13786
rect 4190 13734 4216 13786
rect 4268 13734 4274 13786
rect 3895 13727 4274 13734
rect 4334 13727 4766 13857
rect 4771 13727 5763 13857
rect 6188 13851 7180 13857
rect 6188 13799 6194 13851
rect 6246 13799 6259 13851
rect 6311 13799 6324 13851
rect 6376 13799 6389 13851
rect 6441 13799 6453 13851
rect 6505 13799 6517 13851
rect 6569 13799 6581 13851
rect 6633 13799 6645 13851
rect 6697 13799 6709 13851
rect 6761 13799 6773 13851
rect 6825 13799 6837 13851
rect 6889 13799 7180 13851
rect 6188 13779 7180 13799
rect 6188 13727 6194 13779
rect 6246 13727 6259 13779
rect 6311 13727 6324 13779
rect 6376 13727 6389 13779
rect 6441 13727 6453 13779
rect 6505 13727 6517 13779
rect 6569 13727 6581 13779
rect 6633 13727 6645 13779
rect 6697 13727 6709 13779
rect 6761 13727 6773 13779
rect 6825 13727 6837 13779
rect 6889 13727 7180 13779
rect 7742 13805 7748 13857
rect 7800 13805 7814 13857
rect 7866 13805 7872 13857
rect 7742 13779 7872 13805
rect 7742 13727 7748 13779
rect 7800 13727 7814 13779
rect 7866 13727 7872 13779
rect 8317 13853 9287 13857
rect 8317 13801 8680 13853
rect 8732 13801 8745 13853
rect 8797 13801 8809 13853
rect 8861 13801 8873 13853
rect 8925 13801 9287 13853
rect 8317 13779 9287 13801
rect 8317 13727 8680 13779
rect 8732 13727 8745 13779
rect 8797 13727 8809 13779
rect 8861 13727 8873 13779
rect 8925 13727 9287 13779
rect 9854 13821 10835 13857
rect 9854 13769 10305 13821
rect 10357 13769 10371 13821
rect 10423 13769 10437 13821
rect 10489 13769 10503 13821
rect 10555 13769 10568 13821
rect 10620 13769 10633 13821
rect 10685 13769 10698 13821
rect 10750 13769 10763 13821
rect 10815 13769 10835 13821
rect 9854 13727 10835 13769
rect 11278 13820 12270 13857
rect 11278 13768 11716 13820
rect 11768 13768 11781 13820
rect 11833 13768 11846 13820
rect 11898 13768 11911 13820
rect 11963 13768 11976 13820
rect 12028 13768 12041 13820
rect 12093 13768 12106 13820
rect 12158 13768 12270 13820
rect 11278 13727 12270 13768
rect 12832 13805 13138 13857
rect 13190 13805 13205 13857
rect 13257 13805 13272 13857
rect 13324 13805 13339 13857
rect 13391 13805 13406 13857
rect 13458 13805 13473 13857
rect 13525 13805 13540 13857
rect 13592 13805 14124 13857
rect 12832 13779 14124 13805
rect 12832 13727 13138 13779
rect 13190 13727 13205 13779
rect 13257 13727 13272 13779
rect 13324 13727 13339 13779
rect 13391 13727 13406 13779
rect 13458 13727 13473 13779
rect 13525 13727 13540 13779
rect 13592 13727 14124 13779
rect 535 10030 970 10031
rect 535 9978 541 10030
rect 593 9978 616 10030
rect 668 9978 690 10030
rect 742 9978 764 10030
rect 816 9978 838 10030
rect 890 9978 912 10030
rect 964 9978 970 10030
rect 535 9956 970 9978
rect 535 9904 541 9956
rect 593 9904 616 9956
rect 668 9904 690 9956
rect 742 9904 764 9956
rect 816 9904 838 9956
rect 890 9904 912 9956
rect 964 9904 970 9956
rect 535 9882 970 9904
rect 535 9830 541 9882
rect 593 9830 616 9882
rect 668 9830 690 9882
rect 742 9830 764 9882
rect 816 9830 838 9882
rect 890 9830 912 9882
rect 964 9830 970 9882
rect 535 9829 970 9830
tri 13999 9622 14206 9829 ne
rect -496 9514 13845 9521
rect -496 9480 -484 9514
rect -450 9480 -411 9514
rect -377 9480 -338 9514
rect -304 9480 -265 9514
rect -231 9480 -192 9514
rect -158 9480 -119 9514
rect -85 9480 -46 9514
rect -12 9480 27 9514
rect 61 9480 100 9514
rect 134 9480 173 9514
rect 207 9480 246 9514
rect 280 9480 319 9514
rect 353 9480 392 9514
rect 426 9480 465 9514
rect 499 9480 538 9514
rect 572 9480 611 9514
rect 645 9480 684 9514
rect 718 9480 757 9514
rect 791 9480 830 9514
rect 864 9480 903 9514
rect 937 9480 976 9514
rect 1010 9480 1049 9514
rect 1083 9480 1122 9514
rect 1156 9480 1195 9514
rect 1229 9480 1268 9514
rect 1302 9480 1341 9514
rect 1375 9480 1414 9514
rect 1448 9480 1487 9514
rect 1521 9480 1559 9514
rect 1593 9480 1631 9514
rect 1665 9480 1703 9514
rect 1737 9480 1775 9514
rect 1809 9480 1847 9514
rect 1881 9480 1919 9514
rect 1953 9480 1991 9514
rect 2025 9480 2063 9514
rect 2097 9480 2135 9514
rect 2169 9480 2207 9514
rect 2241 9480 2279 9514
rect 2313 9480 2351 9514
rect 2385 9480 2423 9514
rect 2457 9480 2495 9514
rect 2529 9480 2567 9514
rect 2601 9480 2639 9514
rect 2673 9480 2711 9514
rect 2745 9480 2783 9514
rect 2817 9480 2855 9514
rect 2889 9480 2927 9514
rect 2961 9480 2999 9514
rect 3033 9480 3071 9514
rect 3105 9480 3143 9514
rect 3177 9480 3215 9514
rect 3249 9480 3287 9514
rect 3321 9480 3359 9514
rect 3393 9480 3431 9514
rect 3465 9480 3503 9514
rect 3537 9480 3575 9514
rect 3609 9480 3647 9514
rect 3681 9480 3719 9514
rect 3753 9480 3791 9514
rect 3825 9480 3863 9514
rect 3897 9480 3935 9514
rect 3969 9480 4007 9514
rect 4041 9480 4079 9514
rect 4113 9480 4151 9514
rect 4185 9480 4223 9514
rect 4257 9480 4295 9514
rect 4329 9480 4367 9514
rect 4401 9480 4439 9514
rect 4473 9480 4511 9514
rect 4545 9480 4583 9514
rect 4617 9480 4655 9514
rect 4689 9480 4727 9514
rect 4761 9480 4799 9514
rect 4833 9480 4871 9514
rect 4905 9480 4943 9514
rect 4977 9480 5015 9514
rect 5049 9480 5087 9514
rect 5121 9480 5159 9514
rect 5193 9480 5231 9514
rect 5265 9480 5303 9514
rect 5337 9480 5375 9514
rect 5409 9480 5447 9514
rect 5481 9480 5519 9514
rect 5553 9480 5591 9514
rect 5625 9480 5663 9514
rect 5697 9480 5735 9514
rect 5769 9480 5807 9514
rect 5841 9480 5879 9514
rect 5913 9480 5951 9514
rect 5985 9480 6023 9514
rect 6057 9480 6095 9514
rect 6129 9480 6167 9514
rect 6201 9480 6239 9514
rect 6273 9480 6311 9514
rect 6345 9480 6383 9514
rect 6417 9480 6455 9514
rect 6489 9480 6527 9514
rect 6561 9480 6599 9514
rect 6633 9480 6671 9514
rect 6705 9480 6743 9514
rect 6777 9480 6815 9514
rect 6849 9480 6887 9514
rect 6921 9480 6959 9514
rect 6993 9480 7031 9514
rect 7065 9480 7103 9514
rect 7137 9480 7175 9514
rect 7209 9480 7247 9514
rect 7281 9480 7319 9514
rect 7353 9480 7391 9514
rect 7425 9480 7463 9514
rect 7497 9480 7535 9514
rect 7569 9480 7607 9514
rect 7641 9480 7679 9514
rect 7713 9480 7751 9514
rect 7785 9480 7823 9514
rect 7857 9480 7895 9514
rect 7929 9480 7967 9514
rect 8001 9480 8039 9514
rect 8073 9480 8111 9514
rect 8145 9480 8183 9514
rect 8217 9480 8255 9514
rect 8289 9480 8327 9514
rect 8361 9480 8399 9514
rect 8433 9480 8471 9514
rect 8505 9480 8543 9514
rect 8577 9480 8615 9514
rect 8649 9480 8687 9514
rect 8721 9480 8759 9514
rect 8793 9480 8831 9514
rect 8865 9480 8903 9514
rect 8937 9480 8975 9514
rect 9009 9480 9047 9514
rect 9081 9480 9119 9514
rect 9153 9480 9191 9514
rect 9225 9480 9263 9514
rect 9297 9480 9335 9514
rect 9369 9480 9407 9514
rect 9441 9480 9479 9514
rect 9513 9480 9551 9514
rect 9585 9480 9623 9514
rect 9657 9480 9695 9514
rect 9729 9480 9767 9514
rect 9801 9480 9839 9514
rect 9873 9480 9911 9514
rect 9945 9480 9983 9514
rect 10017 9480 10055 9514
rect 10089 9480 10127 9514
rect 10161 9480 10199 9514
rect 10233 9480 10271 9514
rect 10305 9480 10343 9514
rect 10377 9480 10415 9514
rect 10449 9480 10487 9514
rect 10521 9480 10559 9514
rect 10593 9480 10631 9514
rect 10665 9480 10703 9514
rect 10737 9480 10775 9514
rect 10809 9480 10847 9514
rect 10881 9480 10919 9514
rect 10953 9480 10991 9514
rect 11025 9480 11063 9514
rect 11097 9480 11135 9514
rect 11169 9480 11207 9514
rect 11241 9480 11279 9514
rect 11313 9480 11351 9514
rect 11385 9480 11423 9514
rect 11457 9480 11495 9514
rect 11529 9480 11567 9514
rect 11601 9480 11639 9514
rect 11673 9480 11711 9514
rect 11745 9480 11783 9514
rect 11817 9480 11855 9514
rect 11889 9480 11927 9514
rect 11961 9480 11999 9514
rect 12033 9480 12071 9514
rect 12105 9480 12143 9514
rect 12177 9480 12215 9514
rect 12249 9480 12287 9514
rect 12321 9480 12359 9514
rect 12393 9480 12431 9514
rect 12465 9480 12503 9514
rect 12537 9480 12575 9514
rect 12609 9480 12647 9514
rect 12681 9480 12719 9514
rect 12753 9480 12791 9514
rect 12825 9480 12863 9514
rect 12897 9480 12935 9514
rect 12969 9480 13007 9514
rect 13041 9480 13079 9514
rect 13113 9480 13151 9514
rect 13185 9480 13223 9514
rect 13257 9480 13295 9514
rect 13329 9480 13367 9514
rect 13401 9480 13439 9514
rect 13473 9480 13511 9514
rect 13545 9480 13583 9514
rect 13617 9480 13655 9514
rect 13689 9480 13727 9514
rect 13761 9480 13799 9514
rect 13833 9480 13845 9514
rect -496 9428 13845 9480
rect -496 9394 -484 9428
rect -450 9394 -411 9428
rect -377 9394 -338 9428
rect -304 9394 -265 9428
rect -231 9394 -192 9428
rect -158 9394 -119 9428
rect -85 9394 -46 9428
rect -12 9394 27 9428
rect 61 9394 100 9428
rect 134 9394 173 9428
rect 207 9394 246 9428
rect 280 9394 319 9428
rect 353 9394 392 9428
rect 426 9394 465 9428
rect 499 9394 538 9428
rect 572 9394 611 9428
rect 645 9394 684 9428
rect 718 9394 757 9428
rect 791 9394 830 9428
rect 864 9394 903 9428
rect 937 9394 976 9428
rect 1010 9394 1049 9428
rect 1083 9394 1122 9428
rect 1156 9394 1195 9428
rect 1229 9394 1268 9428
rect 1302 9394 1341 9428
rect 1375 9394 1414 9428
rect 1448 9394 1487 9428
rect 1521 9394 1559 9428
rect 1593 9394 1631 9428
rect 1665 9394 1703 9428
rect 1737 9394 1775 9428
rect 1809 9394 1847 9428
rect 1881 9394 1919 9428
rect 1953 9394 1991 9428
rect 2025 9394 2063 9428
rect 2097 9394 2135 9428
rect 2169 9394 2207 9428
rect 2241 9394 2279 9428
rect 2313 9394 2351 9428
rect 2385 9394 2423 9428
rect 2457 9394 2495 9428
rect 2529 9394 2567 9428
rect 2601 9394 2639 9428
rect 2673 9394 2711 9428
rect 2745 9394 2783 9428
rect 2817 9394 2855 9428
rect 2889 9394 2927 9428
rect 2961 9394 2999 9428
rect 3033 9394 3071 9428
rect 3105 9394 3143 9428
rect 3177 9394 3215 9428
rect 3249 9394 3287 9428
rect 3321 9394 3359 9428
rect 3393 9394 3431 9428
rect 3465 9394 3503 9428
rect 3537 9394 3575 9428
rect 3609 9394 3647 9428
rect 3681 9394 3719 9428
rect 3753 9394 3791 9428
rect 3825 9394 3863 9428
rect 3897 9394 3935 9428
rect 3969 9394 4007 9428
rect 4041 9394 4079 9428
rect 4113 9394 4151 9428
rect 4185 9394 4223 9428
rect 4257 9394 4295 9428
rect 4329 9394 4367 9428
rect 4401 9394 4439 9428
rect 4473 9394 4511 9428
rect 4545 9394 4583 9428
rect 4617 9394 4655 9428
rect 4689 9394 4727 9428
rect 4761 9394 4799 9428
rect 4833 9394 4871 9428
rect 4905 9394 4943 9428
rect 4977 9394 5015 9428
rect 5049 9394 5087 9428
rect 5121 9394 5159 9428
rect 5193 9394 5231 9428
rect 5265 9394 5303 9428
rect 5337 9394 5375 9428
rect 5409 9394 5447 9428
rect 5481 9394 5519 9428
rect 5553 9394 5591 9428
rect 5625 9394 5663 9428
rect 5697 9394 5735 9428
rect 5769 9394 5807 9428
rect 5841 9394 5879 9428
rect 5913 9394 5951 9428
rect 5985 9394 6023 9428
rect 6057 9394 6095 9428
rect 6129 9394 6167 9428
rect 6201 9394 6239 9428
rect 6273 9394 6311 9428
rect 6345 9394 6383 9428
rect 6417 9394 6455 9428
rect 6489 9394 6527 9428
rect 6561 9394 6599 9428
rect 6633 9394 6671 9428
rect 6705 9394 6743 9428
rect 6777 9394 6815 9428
rect 6849 9394 6887 9428
rect 6921 9394 6959 9428
rect 6993 9394 7031 9428
rect 7065 9394 7103 9428
rect 7137 9394 7175 9428
rect 7209 9394 7247 9428
rect 7281 9394 7319 9428
rect 7353 9394 7391 9428
rect 7425 9394 7463 9428
rect 7497 9394 7535 9428
rect 7569 9394 7607 9428
rect 7641 9394 7679 9428
rect 7713 9394 7751 9428
rect 7785 9394 7823 9428
rect 7857 9394 7895 9428
rect 7929 9394 7967 9428
rect 8001 9394 8039 9428
rect 8073 9394 8111 9428
rect 8145 9394 8183 9428
rect 8217 9394 8255 9428
rect 8289 9394 8327 9428
rect 8361 9394 8399 9428
rect 8433 9394 8471 9428
rect 8505 9394 8543 9428
rect 8577 9394 8615 9428
rect 8649 9394 8687 9428
rect 8721 9394 8759 9428
rect 8793 9394 8831 9428
rect 8865 9394 8903 9428
rect 8937 9394 8975 9428
rect 9009 9394 9047 9428
rect 9081 9394 9119 9428
rect 9153 9394 9191 9428
rect 9225 9394 9263 9428
rect 9297 9394 9335 9428
rect 9369 9394 9407 9428
rect 9441 9394 9479 9428
rect 9513 9394 9551 9428
rect 9585 9394 9623 9428
rect 9657 9394 9695 9428
rect 9729 9394 9767 9428
rect 9801 9394 9839 9428
rect 9873 9394 9911 9428
rect 9945 9394 9983 9428
rect 10017 9394 10055 9428
rect 10089 9394 10127 9428
rect 10161 9394 10199 9428
rect 10233 9394 10271 9428
rect 10305 9394 10343 9428
rect 10377 9394 10415 9428
rect 10449 9394 10487 9428
rect 10521 9394 10559 9428
rect 10593 9394 10631 9428
rect 10665 9394 10703 9428
rect 10737 9394 10775 9428
rect 10809 9394 10847 9428
rect 10881 9394 10919 9428
rect 10953 9394 10991 9428
rect 11025 9394 11063 9428
rect 11097 9394 11135 9428
rect 11169 9394 11207 9428
rect 11241 9394 11279 9428
rect 11313 9394 11351 9428
rect 11385 9394 11423 9428
rect 11457 9394 11495 9428
rect 11529 9394 11567 9428
rect 11601 9394 11639 9428
rect 11673 9394 11711 9428
rect 11745 9394 11783 9428
rect 11817 9394 11855 9428
rect 11889 9394 11927 9428
rect 11961 9394 11999 9428
rect 12033 9394 12071 9428
rect 12105 9394 12143 9428
rect 12177 9394 12215 9428
rect 12249 9394 12287 9428
rect 12321 9394 12359 9428
rect 12393 9394 12431 9428
rect 12465 9394 12503 9428
rect 12537 9394 12575 9428
rect 12609 9394 12647 9428
rect 12681 9394 12719 9428
rect 12753 9394 12791 9428
rect 12825 9394 12863 9428
rect 12897 9394 12935 9428
rect 12969 9394 13007 9428
rect 13041 9394 13079 9428
rect 13113 9394 13151 9428
rect 13185 9394 13223 9428
rect 13257 9394 13295 9428
rect 13329 9394 13367 9428
rect 13401 9394 13439 9428
rect 13473 9394 13511 9428
rect 13545 9394 13583 9428
rect 13617 9394 13655 9428
rect 13689 9394 13727 9428
rect 13761 9394 13799 9428
rect 13833 9394 13845 9428
rect -496 9359 13845 9394
rect -496 9342 12258 9359
rect 12310 9342 12335 9359
rect 12387 9342 12412 9359
rect 12464 9342 12488 9359
rect -496 9308 -484 9342
rect -450 9308 -411 9342
rect -377 9308 -338 9342
rect -304 9308 -265 9342
rect -231 9308 -192 9342
rect -158 9308 -119 9342
rect -85 9308 -46 9342
rect -12 9308 27 9342
rect 61 9308 100 9342
rect 134 9308 173 9342
rect 207 9308 246 9342
rect 280 9308 319 9342
rect 353 9308 392 9342
rect 426 9308 465 9342
rect 499 9308 538 9342
rect 572 9308 611 9342
rect 645 9308 684 9342
rect 718 9308 757 9342
rect 791 9308 830 9342
rect 864 9308 903 9342
rect 937 9308 976 9342
rect 1010 9308 1049 9342
rect 1083 9308 1122 9342
rect 1156 9308 1195 9342
rect 1229 9308 1268 9342
rect 1302 9308 1341 9342
rect 1375 9308 1414 9342
rect 1448 9308 1487 9342
rect 1521 9308 1559 9342
rect 1593 9308 1631 9342
rect 1665 9308 1703 9342
rect 1737 9308 1775 9342
rect 1809 9308 1847 9342
rect 1881 9308 1919 9342
rect 1953 9308 1991 9342
rect 2025 9308 2063 9342
rect 2097 9308 2135 9342
rect 2169 9308 2207 9342
rect 2241 9308 2279 9342
rect 2313 9308 2351 9342
rect 2385 9308 2423 9342
rect 2457 9308 2495 9342
rect 2529 9308 2567 9342
rect 2601 9308 2639 9342
rect 2673 9308 2711 9342
rect 2745 9308 2783 9342
rect 2817 9308 2855 9342
rect 2889 9308 2927 9342
rect 2961 9308 2999 9342
rect 3033 9308 3071 9342
rect 3105 9308 3143 9342
rect 3177 9308 3215 9342
rect 3249 9308 3287 9342
rect 3321 9308 3359 9342
rect 3393 9308 3431 9342
rect 3465 9308 3503 9342
rect 3537 9308 3575 9342
rect 3609 9308 3647 9342
rect 3681 9308 3719 9342
rect 3753 9308 3791 9342
rect 3825 9308 3863 9342
rect 3897 9308 3935 9342
rect 3969 9308 4007 9342
rect 4041 9308 4079 9342
rect 4113 9308 4151 9342
rect 4185 9308 4223 9342
rect 4257 9308 4295 9342
rect 4329 9308 4367 9342
rect 4401 9308 4439 9342
rect 4473 9308 4511 9342
rect 4545 9308 4583 9342
rect 4617 9308 4655 9342
rect 4689 9308 4727 9342
rect 4761 9308 4799 9342
rect 4833 9308 4871 9342
rect 4905 9308 4943 9342
rect 4977 9308 5015 9342
rect 5049 9308 5087 9342
rect 5121 9308 5159 9342
rect 5193 9308 5231 9342
rect 5265 9308 5303 9342
rect 5337 9308 5375 9342
rect 5409 9308 5447 9342
rect 5481 9308 5519 9342
rect 5553 9308 5591 9342
rect 5625 9308 5663 9342
rect 5697 9308 5735 9342
rect 5769 9308 5807 9342
rect 5841 9308 5879 9342
rect 5913 9308 5951 9342
rect 5985 9308 6023 9342
rect 6057 9308 6095 9342
rect 6129 9308 6167 9342
rect 6201 9308 6239 9342
rect 6273 9308 6311 9342
rect 6345 9308 6383 9342
rect 6417 9308 6455 9342
rect 6489 9308 6527 9342
rect 6561 9308 6599 9342
rect 6633 9308 6671 9342
rect 6705 9308 6743 9342
rect 6777 9308 6815 9342
rect 6849 9308 6887 9342
rect 6921 9308 6959 9342
rect 6993 9308 7031 9342
rect 7065 9308 7103 9342
rect 7137 9308 7175 9342
rect 7209 9308 7247 9342
rect 7281 9308 7319 9342
rect 7353 9308 7391 9342
rect 7425 9308 7463 9342
rect 7497 9308 7535 9342
rect 7569 9308 7607 9342
rect 7641 9308 7679 9342
rect 7713 9308 7751 9342
rect 7785 9308 7823 9342
rect 7857 9308 7895 9342
rect 7929 9308 7967 9342
rect 8001 9308 8039 9342
rect 8073 9308 8111 9342
rect 8145 9308 8183 9342
rect 8217 9308 8255 9342
rect 8289 9308 8327 9342
rect 8361 9308 8399 9342
rect 8433 9308 8471 9342
rect 8505 9308 8543 9342
rect 8577 9308 8615 9342
rect 8649 9308 8687 9342
rect 8721 9308 8759 9342
rect 8793 9308 8831 9342
rect 8865 9308 8903 9342
rect 8937 9308 8975 9342
rect 9009 9308 9047 9342
rect 9081 9308 9119 9342
rect 9153 9308 9191 9342
rect 9225 9308 9263 9342
rect 9297 9308 9335 9342
rect 9369 9308 9407 9342
rect 9441 9308 9479 9342
rect 9513 9308 9551 9342
rect 9585 9308 9623 9342
rect 9657 9308 9695 9342
rect 9729 9308 9767 9342
rect 9801 9308 9839 9342
rect 9873 9308 9911 9342
rect 9945 9308 9983 9342
rect 10017 9308 10055 9342
rect 10089 9308 10127 9342
rect 10161 9308 10199 9342
rect 10233 9308 10271 9342
rect 10305 9308 10343 9342
rect 10377 9308 10415 9342
rect 10449 9308 10487 9342
rect 10521 9308 10559 9342
rect 10593 9308 10631 9342
rect 10665 9308 10703 9342
rect 10737 9308 10775 9342
rect 10809 9308 10847 9342
rect 10881 9308 10919 9342
rect 10953 9308 10991 9342
rect 11025 9308 11063 9342
rect 11097 9308 11135 9342
rect 11169 9308 11207 9342
rect 11241 9308 11279 9342
rect 11313 9308 11351 9342
rect 11385 9308 11423 9342
rect 11457 9308 11495 9342
rect 11529 9308 11567 9342
rect 11601 9308 11639 9342
rect 11673 9308 11711 9342
rect 11745 9308 11783 9342
rect 11817 9308 11855 9342
rect 11889 9308 11927 9342
rect 11961 9308 11999 9342
rect 12033 9308 12071 9342
rect 12105 9308 12143 9342
rect 12177 9308 12215 9342
rect 12249 9308 12258 9342
rect 12321 9308 12335 9342
rect 12393 9308 12412 9342
rect 12465 9308 12488 9342
rect -496 9307 12258 9308
rect 12310 9307 12335 9308
rect 12387 9307 12412 9308
rect 12464 9307 12488 9308
rect 12540 9307 12564 9359
rect 12616 9342 13845 9359
rect 12616 9308 12647 9342
rect 12681 9308 12719 9342
rect 12753 9308 12791 9342
rect 12825 9308 12863 9342
rect 12897 9308 12935 9342
rect 12969 9308 13007 9342
rect 13041 9308 13079 9342
rect 13113 9308 13151 9342
rect 13185 9308 13223 9342
rect 13257 9308 13295 9342
rect 13329 9308 13367 9342
rect 13401 9308 13439 9342
rect 13473 9308 13511 9342
rect 13545 9308 13583 9342
rect 13617 9308 13655 9342
rect 13689 9308 13727 9342
rect 13761 9308 13799 9342
rect 13833 9308 13845 9342
rect 12616 9307 13845 9308
rect -496 9271 13845 9307
rect -496 9256 12258 9271
rect 12310 9256 12335 9271
rect 12387 9256 12412 9271
rect 12464 9256 12488 9271
rect -496 9222 -484 9256
rect -450 9222 -411 9256
rect -377 9222 -338 9256
rect -304 9222 -265 9256
rect -231 9222 -192 9256
rect -158 9222 -119 9256
rect -85 9222 -46 9256
rect -12 9222 27 9256
rect 61 9222 100 9256
rect 134 9222 173 9256
rect 207 9222 246 9256
rect 280 9222 319 9256
rect 353 9222 392 9256
rect 426 9222 465 9256
rect 499 9222 538 9256
rect 572 9222 611 9256
rect 645 9222 684 9256
rect 718 9222 757 9256
rect 791 9222 830 9256
rect 864 9222 903 9256
rect 937 9222 976 9256
rect 1010 9222 1049 9256
rect 1083 9222 1122 9256
rect 1156 9222 1195 9256
rect 1229 9222 1268 9256
rect 1302 9222 1341 9256
rect 1375 9222 1414 9256
rect 1448 9222 1487 9256
rect 1521 9222 1559 9256
rect 1593 9222 1631 9256
rect 1665 9222 1703 9256
rect 1737 9222 1775 9256
rect 1809 9222 1847 9256
rect 1881 9222 1919 9256
rect 1953 9222 1991 9256
rect 2025 9222 2063 9256
rect 2097 9222 2135 9256
rect 2169 9222 2207 9256
rect 2241 9222 2279 9256
rect 2313 9222 2351 9256
rect 2385 9222 2423 9256
rect 2457 9222 2495 9256
rect 2529 9222 2567 9256
rect 2601 9222 2639 9256
rect 2673 9222 2711 9256
rect 2745 9222 2783 9256
rect 2817 9222 2855 9256
rect 2889 9222 2927 9256
rect 2961 9222 2999 9256
rect 3033 9222 3071 9256
rect 3105 9222 3143 9256
rect 3177 9222 3215 9256
rect 3249 9222 3287 9256
rect 3321 9222 3359 9256
rect 3393 9222 3431 9256
rect 3465 9222 3503 9256
rect 3537 9222 3575 9256
rect 3609 9222 3647 9256
rect 3681 9222 3719 9256
rect 3753 9222 3791 9256
rect 3825 9222 3863 9256
rect 3897 9222 3935 9256
rect 3969 9222 4007 9256
rect 4041 9222 4079 9256
rect 4113 9222 4151 9256
rect 4185 9222 4223 9256
rect 4257 9222 4295 9256
rect 4329 9222 4367 9256
rect 4401 9222 4439 9256
rect 4473 9222 4511 9256
rect 4545 9222 4583 9256
rect 4617 9222 4655 9256
rect 4689 9222 4727 9256
rect 4761 9222 4799 9256
rect 4833 9222 4871 9256
rect 4905 9222 4943 9256
rect 4977 9222 5015 9256
rect 5049 9222 5087 9256
rect 5121 9222 5159 9256
rect 5193 9222 5231 9256
rect 5265 9222 5303 9256
rect 5337 9222 5375 9256
rect 5409 9222 5447 9256
rect 5481 9222 5519 9256
rect 5553 9222 5591 9256
rect 5625 9222 5663 9256
rect 5697 9222 5735 9256
rect 5769 9222 5807 9256
rect 5841 9222 5879 9256
rect 5913 9222 5951 9256
rect 5985 9222 6023 9256
rect 6057 9222 6095 9256
rect 6129 9222 6167 9256
rect 6201 9222 6239 9256
rect 6273 9222 6311 9256
rect 6345 9222 6383 9256
rect 6417 9222 6455 9256
rect 6489 9222 6527 9256
rect 6561 9222 6599 9256
rect 6633 9222 6671 9256
rect 6705 9222 6743 9256
rect 6777 9222 6815 9256
rect 6849 9222 6887 9256
rect 6921 9222 6959 9256
rect 6993 9222 7031 9256
rect 7065 9222 7103 9256
rect 7137 9222 7175 9256
rect 7209 9222 7247 9256
rect 7281 9222 7319 9256
rect 7353 9222 7391 9256
rect 7425 9222 7463 9256
rect 7497 9222 7535 9256
rect 7569 9222 7607 9256
rect 7641 9222 7679 9256
rect 7713 9222 7751 9256
rect 7785 9222 7823 9256
rect 7857 9222 7895 9256
rect 7929 9222 7967 9256
rect 8001 9222 8039 9256
rect 8073 9222 8111 9256
rect 8145 9222 8183 9256
rect 8217 9222 8255 9256
rect 8289 9222 8327 9256
rect 8361 9222 8399 9256
rect 8433 9222 8471 9256
rect 8505 9222 8543 9256
rect 8577 9222 8615 9256
rect 8649 9222 8687 9256
rect 8721 9222 8759 9256
rect 8793 9222 8831 9256
rect 8865 9222 8903 9256
rect 8937 9222 8975 9256
rect 9009 9222 9047 9256
rect 9081 9222 9119 9256
rect 9153 9222 9191 9256
rect 9225 9222 9263 9256
rect 9297 9222 9335 9256
rect 9369 9222 9407 9256
rect 9441 9222 9479 9256
rect 9513 9222 9551 9256
rect 9585 9222 9623 9256
rect 9657 9222 9695 9256
rect 9729 9222 9767 9256
rect 9801 9222 9839 9256
rect 9873 9222 9911 9256
rect 9945 9222 9983 9256
rect 10017 9222 10055 9256
rect 10089 9222 10127 9256
rect 10161 9222 10199 9256
rect 10233 9222 10271 9256
rect 10305 9222 10343 9256
rect 10377 9222 10415 9256
rect 10449 9222 10487 9256
rect 10521 9222 10559 9256
rect 10593 9222 10631 9256
rect 10665 9222 10703 9256
rect 10737 9222 10775 9256
rect 10809 9222 10847 9256
rect 10881 9222 10919 9256
rect 10953 9222 10991 9256
rect 11025 9222 11063 9256
rect 11097 9222 11135 9256
rect 11169 9222 11207 9256
rect 11241 9222 11279 9256
rect 11313 9222 11351 9256
rect 11385 9222 11423 9256
rect 11457 9222 11495 9256
rect 11529 9222 11567 9256
rect 11601 9222 11639 9256
rect 11673 9222 11711 9256
rect 11745 9222 11783 9256
rect 11817 9222 11855 9256
rect 11889 9222 11927 9256
rect 11961 9222 11999 9256
rect 12033 9222 12071 9256
rect 12105 9222 12143 9256
rect 12177 9222 12215 9256
rect 12249 9222 12258 9256
rect 12321 9222 12335 9256
rect 12393 9222 12412 9256
rect 12465 9222 12488 9256
rect -496 9219 12258 9222
rect 12310 9219 12335 9222
rect 12387 9219 12412 9222
rect 12464 9219 12488 9222
rect 12540 9219 12564 9271
rect 12616 9256 13845 9271
rect 12616 9222 12647 9256
rect 12681 9222 12719 9256
rect 12753 9222 12791 9256
rect 12825 9222 12863 9256
rect 12897 9222 12935 9256
rect 12969 9222 13007 9256
rect 13041 9222 13079 9256
rect 13113 9222 13151 9256
rect 13185 9222 13223 9256
rect 13257 9222 13295 9256
rect 13329 9222 13367 9256
rect 13401 9222 13439 9256
rect 13473 9222 13511 9256
rect 13545 9222 13583 9256
rect 13617 9222 13655 9256
rect 13689 9222 13727 9256
rect 13761 9222 13799 9256
rect 13833 9222 13845 9256
rect 12616 9219 13845 9222
rect -496 9183 13845 9219
rect -496 9170 12258 9183
rect 12310 9170 12335 9183
rect 12387 9170 12412 9183
rect 12464 9170 12488 9183
rect -496 9136 -484 9170
rect -450 9136 -411 9170
rect -377 9136 -338 9170
rect -304 9136 -265 9170
rect -231 9136 -192 9170
rect -158 9136 -119 9170
rect -85 9136 -46 9170
rect -12 9136 27 9170
rect 61 9136 100 9170
rect 134 9136 173 9170
rect 207 9136 246 9170
rect 280 9136 319 9170
rect 353 9136 392 9170
rect 426 9136 465 9170
rect 499 9136 538 9170
rect 572 9136 611 9170
rect 645 9136 684 9170
rect 718 9136 757 9170
rect 791 9136 830 9170
rect 864 9136 903 9170
rect 937 9136 976 9170
rect 1010 9136 1049 9170
rect 1083 9136 1122 9170
rect 1156 9136 1195 9170
rect 1229 9136 1268 9170
rect 1302 9136 1341 9170
rect 1375 9136 1414 9170
rect 1448 9136 1487 9170
rect 1521 9136 1559 9170
rect 1593 9136 1631 9170
rect 1665 9136 1703 9170
rect 1737 9136 1775 9170
rect 1809 9136 1847 9170
rect 1881 9136 1919 9170
rect 1953 9136 1991 9170
rect 2025 9136 2063 9170
rect 2097 9136 2135 9170
rect 2169 9136 2207 9170
rect 2241 9136 2279 9170
rect 2313 9136 2351 9170
rect 2385 9136 2423 9170
rect 2457 9136 2495 9170
rect 2529 9136 2567 9170
rect 2601 9136 2639 9170
rect 2673 9136 2711 9170
rect 2745 9136 2783 9170
rect 2817 9136 2855 9170
rect 2889 9136 2927 9170
rect 2961 9136 2999 9170
rect 3033 9136 3071 9170
rect 3105 9136 3143 9170
rect 3177 9136 3215 9170
rect 3249 9136 3287 9170
rect 3321 9136 3359 9170
rect 3393 9136 3431 9170
rect 3465 9136 3503 9170
rect 3537 9136 3575 9170
rect 3609 9136 3647 9170
rect 3681 9136 3719 9170
rect 3753 9136 3791 9170
rect 3825 9136 3863 9170
rect 3897 9136 3935 9170
rect 3969 9136 4007 9170
rect 4041 9136 4079 9170
rect 4113 9136 4151 9170
rect 4185 9136 4223 9170
rect 4257 9136 4295 9170
rect 4329 9136 4367 9170
rect 4401 9136 4439 9170
rect 4473 9136 4511 9170
rect 4545 9136 4583 9170
rect 4617 9136 4655 9170
rect 4689 9136 4727 9170
rect 4761 9136 4799 9170
rect 4833 9136 4871 9170
rect 4905 9136 4943 9170
rect 4977 9136 5015 9170
rect 5049 9136 5087 9170
rect 5121 9136 5159 9170
rect 5193 9136 5231 9170
rect 5265 9136 5303 9170
rect 5337 9136 5375 9170
rect 5409 9136 5447 9170
rect 5481 9136 5519 9170
rect 5553 9136 5591 9170
rect 5625 9136 5663 9170
rect 5697 9136 5735 9170
rect 5769 9136 5807 9170
rect 5841 9136 5879 9170
rect 5913 9136 5951 9170
rect 5985 9136 6023 9170
rect 6057 9136 6095 9170
rect 6129 9136 6167 9170
rect 6201 9136 6239 9170
rect 6273 9136 6311 9170
rect 6345 9136 6383 9170
rect 6417 9136 6455 9170
rect 6489 9136 6527 9170
rect 6561 9136 6599 9170
rect 6633 9136 6671 9170
rect 6705 9136 6743 9170
rect 6777 9136 6815 9170
rect 6849 9136 6887 9170
rect 6921 9136 6959 9170
rect 6993 9136 7031 9170
rect 7065 9136 7103 9170
rect 7137 9136 7175 9170
rect 7209 9136 7247 9170
rect 7281 9136 7319 9170
rect 7353 9136 7391 9170
rect 7425 9136 7463 9170
rect 7497 9136 7535 9170
rect 7569 9136 7607 9170
rect 7641 9136 7679 9170
rect 7713 9136 7751 9170
rect 7785 9136 7823 9170
rect 7857 9136 7895 9170
rect 7929 9136 7967 9170
rect 8001 9136 8039 9170
rect 8073 9136 8111 9170
rect 8145 9136 8183 9170
rect 8217 9136 8255 9170
rect 8289 9136 8327 9170
rect 8361 9136 8399 9170
rect 8433 9136 8471 9170
rect 8505 9136 8543 9170
rect 8577 9136 8615 9170
rect 8649 9136 8687 9170
rect 8721 9136 8759 9170
rect 8793 9136 8831 9170
rect 8865 9136 8903 9170
rect 8937 9136 8975 9170
rect 9009 9136 9047 9170
rect 9081 9136 9119 9170
rect 9153 9136 9191 9170
rect 9225 9136 9263 9170
rect 9297 9136 9335 9170
rect 9369 9136 9407 9170
rect 9441 9136 9479 9170
rect 9513 9136 9551 9170
rect 9585 9136 9623 9170
rect 9657 9136 9695 9170
rect 9729 9136 9767 9170
rect 9801 9136 9839 9170
rect 9873 9136 9911 9170
rect 9945 9136 9983 9170
rect 10017 9136 10055 9170
rect 10089 9136 10127 9170
rect 10161 9136 10199 9170
rect 10233 9136 10271 9170
rect 10305 9136 10343 9170
rect 10377 9136 10415 9170
rect 10449 9136 10487 9170
rect 10521 9136 10559 9170
rect 10593 9136 10631 9170
rect 10665 9136 10703 9170
rect 10737 9136 10775 9170
rect 10809 9136 10847 9170
rect 10881 9136 10919 9170
rect 10953 9136 10991 9170
rect 11025 9136 11063 9170
rect 11097 9136 11135 9170
rect 11169 9136 11207 9170
rect 11241 9136 11279 9170
rect 11313 9136 11351 9170
rect 11385 9136 11423 9170
rect 11457 9136 11495 9170
rect 11529 9136 11567 9170
rect 11601 9136 11639 9170
rect 11673 9136 11711 9170
rect 11745 9136 11783 9170
rect 11817 9136 11855 9170
rect 11889 9136 11927 9170
rect 11961 9136 11999 9170
rect 12033 9136 12071 9170
rect 12105 9136 12143 9170
rect 12177 9136 12215 9170
rect 12249 9136 12258 9170
rect 12321 9136 12335 9170
rect 12393 9136 12412 9170
rect 12465 9136 12488 9170
rect -496 9131 12258 9136
rect 12310 9131 12335 9136
rect 12387 9131 12412 9136
rect 12464 9131 12488 9136
rect 12540 9131 12564 9183
rect 12616 9170 13845 9183
rect 12616 9136 12647 9170
rect 12681 9136 12719 9170
rect 12753 9136 12791 9170
rect 12825 9136 12863 9170
rect 12897 9136 12935 9170
rect 12969 9136 13007 9170
rect 13041 9136 13079 9170
rect 13113 9136 13151 9170
rect 13185 9136 13223 9170
rect 13257 9136 13295 9170
rect 13329 9136 13367 9170
rect 13401 9136 13439 9170
rect 13473 9136 13511 9170
rect 13545 9136 13583 9170
rect 13617 9136 13655 9170
rect 13689 9136 13727 9170
rect 13761 9136 13799 9170
rect 13833 9136 13845 9170
rect 12616 9131 13845 9136
rect -496 9129 13845 9131
rect 14206 9460 15114 9829
rect 14206 9408 14240 9460
rect 14292 9408 14312 9460
rect 14364 9408 14384 9460
rect 14436 9408 14456 9460
rect 14508 9408 14528 9460
rect 14580 9408 14600 9460
rect 14652 9408 15114 9460
rect 14206 9395 15114 9408
rect 14206 9343 14240 9395
rect 14292 9343 14312 9395
rect 14364 9343 14384 9395
rect 14436 9343 14456 9395
rect 14508 9343 14528 9395
rect 14580 9343 14600 9395
rect 14652 9343 15114 9395
rect 14206 9330 15114 9343
rect 14206 9278 14240 9330
rect 14292 9278 14312 9330
rect 14364 9278 14384 9330
rect 14436 9278 14456 9330
rect 14508 9278 14528 9330
rect 14580 9278 14600 9330
rect 14652 9278 15114 9330
rect 14206 9265 15114 9278
rect 14206 9213 14240 9265
rect 14292 9213 14312 9265
rect 14364 9213 14384 9265
rect 14436 9213 14456 9265
rect 14508 9213 14528 9265
rect 14580 9213 14600 9265
rect 14652 9213 15114 9265
rect 14206 9200 15114 9213
rect 14206 9148 14240 9200
rect 14292 9148 14312 9200
rect 14364 9148 14384 9200
rect 14436 9148 14456 9200
rect 14508 9148 14528 9200
rect 14580 9148 14600 9200
rect 14652 9148 15114 9200
rect 14206 9135 15114 9148
rect 14206 9083 14240 9135
rect 14292 9083 14312 9135
rect 14364 9083 14384 9135
rect 14436 9083 14456 9135
rect 14508 9083 14528 9135
rect 14580 9083 14600 9135
rect 14652 9083 15114 9135
rect 14206 9070 15114 9083
rect 14206 9018 14240 9070
rect 14292 9018 14312 9070
rect 14364 9018 14384 9070
rect 14436 9018 14456 9070
rect 14508 9018 14528 9070
rect 14580 9018 14600 9070
rect 14652 9018 15114 9070
rect 14206 9005 15114 9018
tri 14031 8828 14206 9003 se
rect 14206 8953 14240 9005
rect 14292 8953 14312 9005
rect 14364 8953 14384 9005
rect 14436 8953 14456 9005
rect 14508 8953 14528 9005
rect 14580 8953 14600 9005
rect 14652 8953 15114 9005
rect 14206 8940 15114 8953
rect 14206 8888 14240 8940
rect 14292 8888 14312 8940
rect 14364 8888 14384 8940
rect 14436 8888 14456 8940
rect 14508 8888 14528 8940
rect 14580 8888 14600 8940
rect 14652 8888 15114 8940
rect 14206 8875 15114 8888
rect 14206 8828 14240 8875
rect 56 8827 14240 8828
rect 56 8775 541 8827
rect 593 8775 616 8827
rect 668 8775 690 8827
rect 742 8775 764 8827
rect 816 8775 838 8827
rect 890 8775 912 8827
rect 964 8823 14240 8827
rect 14292 8823 14312 8875
rect 14364 8823 14384 8875
rect 14436 8823 14456 8875
rect 14508 8823 14528 8875
rect 14580 8823 14600 8875
rect 14652 8823 15114 8875
rect 964 8810 15114 8823
rect 964 8775 14240 8810
rect 56 8760 14240 8775
rect 14292 8760 14312 8810
rect 14364 8760 14384 8810
rect 14436 8760 14456 8810
rect 14508 8760 14528 8810
rect 14580 8760 14600 8810
rect 14652 8760 15114 8810
rect 56 8753 912 8760
rect 56 8719 248 8753
rect 282 8719 322 8753
rect 356 8719 396 8753
rect 430 8719 470 8753
rect 504 8751 544 8753
rect 578 8751 618 8753
rect 652 8751 691 8753
rect 725 8751 764 8753
rect 798 8751 837 8753
rect 871 8751 912 8753
rect 946 8751 984 8760
rect 504 8719 541 8751
rect 56 8699 541 8719
rect 593 8699 616 8751
rect 668 8699 690 8751
rect 742 8699 764 8751
rect 816 8719 837 8751
rect 816 8699 838 8719
rect 890 8699 912 8751
rect 964 8726 984 8751
rect 1018 8726 1056 8760
rect 1090 8726 1128 8760
rect 1162 8726 1200 8760
rect 1234 8726 1272 8760
rect 1306 8726 1344 8760
rect 1378 8726 1416 8760
rect 1450 8726 1488 8760
rect 1522 8726 1560 8760
rect 1594 8726 1632 8760
rect 1666 8726 1704 8760
rect 1738 8726 1776 8760
rect 1810 8726 1849 8760
rect 1883 8726 1922 8760
rect 1956 8726 1995 8760
rect 2029 8726 2068 8760
rect 2102 8726 2141 8760
rect 2175 8753 3477 8760
rect 2175 8726 2227 8753
rect 964 8719 2227 8726
rect 2261 8719 2306 8753
rect 2340 8719 2385 8753
rect 2419 8719 2464 8753
rect 2498 8719 2543 8753
rect 2577 8719 2621 8753
rect 2655 8719 2699 8753
rect 2733 8719 2777 8753
rect 2811 8719 2855 8753
rect 2889 8719 2933 8753
rect 2967 8719 3011 8753
rect 3045 8726 3477 8753
rect 3511 8726 3550 8760
rect 3584 8726 3623 8760
rect 3657 8726 3696 8760
rect 3730 8726 3769 8760
rect 3803 8726 3842 8760
rect 3876 8726 3915 8760
rect 3949 8726 3988 8760
rect 4022 8726 4061 8760
rect 4095 8726 4134 8760
rect 4168 8726 4207 8760
rect 4241 8726 4280 8760
rect 4314 8726 4353 8760
rect 4387 8726 4426 8760
rect 4460 8726 4499 8760
rect 4533 8726 4572 8760
rect 4606 8726 4645 8760
rect 4679 8726 4718 8760
rect 4752 8726 4791 8760
rect 4825 8726 4864 8760
rect 4898 8726 4937 8760
rect 4971 8726 5010 8760
rect 5044 8726 5083 8760
rect 5117 8726 5156 8760
rect 5190 8726 5229 8760
rect 5263 8726 5302 8760
rect 5336 8726 5375 8760
rect 5409 8726 5448 8760
rect 5482 8726 5521 8760
rect 5555 8726 5594 8760
rect 5628 8726 5667 8760
rect 5701 8726 5740 8760
rect 5774 8726 5813 8760
rect 5847 8726 5886 8760
rect 5920 8726 5959 8760
rect 5993 8726 6032 8760
rect 6066 8726 6105 8760
rect 6139 8726 6178 8760
rect 6212 8726 6251 8760
rect 6285 8726 6324 8760
rect 6358 8726 6397 8760
rect 6431 8726 6470 8760
rect 6504 8726 6543 8760
rect 6577 8726 6616 8760
rect 6650 8726 6689 8760
rect 6723 8726 6762 8760
rect 6796 8726 6835 8760
rect 6869 8726 6908 8760
rect 6942 8726 6981 8760
rect 7015 8726 7054 8760
rect 7088 8726 7127 8760
rect 7161 8726 7200 8760
rect 7234 8726 7273 8760
rect 7307 8726 7346 8760
rect 7380 8726 7419 8760
rect 7453 8726 7492 8760
rect 7526 8726 7565 8760
rect 7599 8726 7638 8760
rect 7672 8726 7711 8760
rect 7745 8726 7784 8760
rect 7818 8726 7857 8760
rect 7891 8726 7930 8760
rect 7964 8726 8003 8760
rect 8037 8726 8075 8760
rect 8109 8726 8147 8760
rect 8181 8726 8219 8760
rect 8253 8726 8291 8760
rect 8325 8726 8363 8760
rect 8397 8726 8435 8760
rect 8469 8726 8507 8760
rect 8541 8726 8579 8760
rect 8613 8726 8651 8760
rect 8685 8726 8723 8760
rect 8757 8726 8795 8760
rect 8829 8726 8867 8760
rect 8901 8726 8939 8760
rect 8973 8726 9011 8760
rect 9045 8726 9083 8760
rect 9117 8726 9155 8760
rect 9189 8726 9227 8760
rect 9261 8726 9299 8760
rect 9333 8726 9371 8760
rect 9405 8726 9443 8760
rect 9477 8726 9515 8760
rect 9549 8726 9587 8760
rect 9621 8726 9659 8760
rect 9693 8726 9731 8760
rect 9765 8726 9803 8760
rect 9837 8726 9875 8760
rect 9909 8726 9947 8760
rect 9981 8726 10019 8760
rect 10053 8726 10091 8760
rect 10125 8726 10163 8760
rect 10197 8726 10235 8760
rect 10269 8726 10307 8760
rect 10341 8726 10379 8760
rect 10413 8726 10451 8760
rect 10485 8726 10523 8760
rect 10557 8726 10595 8760
rect 10629 8726 10667 8760
rect 10701 8726 10739 8760
rect 10773 8726 10811 8760
rect 10845 8726 10883 8760
rect 10917 8726 10955 8760
rect 10989 8726 11027 8760
rect 11061 8726 11099 8760
rect 11133 8726 11171 8760
rect 11205 8726 11243 8760
rect 11277 8726 11315 8760
rect 11349 8726 11387 8760
rect 11421 8726 11459 8760
rect 11493 8726 11531 8760
rect 11565 8726 11603 8760
rect 11637 8726 11675 8760
rect 11709 8726 11747 8760
rect 11781 8726 11819 8760
rect 11853 8726 11891 8760
rect 11925 8726 11963 8760
rect 11997 8726 12035 8760
rect 12069 8726 12107 8760
rect 12141 8726 12179 8760
rect 12213 8726 12251 8760
rect 12285 8726 12323 8760
rect 12357 8726 12395 8760
rect 12429 8726 12467 8760
rect 12501 8726 12539 8760
rect 12573 8726 12611 8760
rect 12645 8726 12683 8760
rect 12717 8726 12755 8760
rect 12789 8726 12827 8760
rect 12861 8726 12899 8760
rect 12933 8726 12971 8760
rect 13005 8726 13043 8760
rect 13077 8726 13115 8760
rect 13149 8726 13187 8760
rect 13221 8726 13259 8760
rect 13293 8726 13331 8760
rect 13365 8726 13403 8760
rect 13437 8726 13475 8760
rect 13509 8726 13547 8760
rect 13581 8726 13619 8760
rect 13653 8726 13691 8760
rect 13725 8726 13763 8760
rect 13797 8726 13835 8760
rect 13869 8726 13907 8760
rect 13941 8726 13979 8760
rect 14013 8726 14051 8760
rect 14085 8726 14123 8760
rect 14157 8726 14195 8760
rect 14229 8758 14240 8760
rect 14301 8758 14312 8760
rect 14373 8758 14384 8760
rect 14445 8758 14456 8760
rect 14517 8758 14528 8760
rect 14589 8758 14600 8760
rect 14229 8745 14267 8758
rect 14301 8745 14339 8758
rect 14373 8745 14411 8758
rect 14445 8745 14483 8758
rect 14517 8745 14555 8758
rect 14589 8745 14627 8758
rect 14229 8726 14240 8745
rect 14301 8726 14312 8745
rect 14373 8726 14384 8745
rect 14445 8726 14456 8745
rect 14517 8726 14528 8745
rect 14589 8726 14600 8745
rect 14661 8726 14699 8760
rect 14733 8726 14771 8760
rect 14805 8726 14843 8760
rect 14877 8726 15114 8760
rect 3045 8719 14240 8726
rect 964 8713 14240 8719
rect 964 8699 2306 8713
tri 2306 8699 2320 8713 nw
tri 3344 8699 3358 8713 ne
rect 3358 8699 14240 8713
tri 728 8693 734 8699 ne
rect 734 8693 2243 8699
tri 734 8636 791 8693 ne
rect 791 8670 2243 8693
rect 791 8636 842 8670
tri 791 8602 825 8636 ne
rect 825 8618 842 8636
rect 894 8618 912 8670
rect 964 8636 2243 8670
tri 2243 8636 2306 8699 nw
tri 3358 8636 3421 8699 ne
rect 3421 8693 14240 8699
rect 14292 8693 14312 8726
rect 14364 8693 14384 8726
rect 14436 8693 14456 8726
rect 14508 8693 14528 8726
rect 14580 8693 14600 8726
rect 14652 8693 15114 8726
rect 3421 8680 15114 8693
rect 3421 8636 14240 8680
rect 14292 8636 14312 8680
rect 14364 8636 14384 8680
rect 14436 8636 14456 8680
rect 14508 8636 14528 8680
rect 14580 8636 14600 8680
rect 14652 8636 15114 8680
rect 964 8618 984 8636
rect 825 8602 912 8618
rect 946 8602 984 8618
rect 1018 8602 1056 8636
rect 1090 8602 1128 8636
rect 1162 8602 1200 8636
rect 1234 8602 1272 8636
rect 1306 8602 1344 8636
rect 1378 8602 1416 8636
rect 1450 8602 1488 8636
rect 1522 8602 1560 8636
rect 1594 8602 1632 8636
rect 1666 8602 1704 8636
rect 1738 8602 1776 8636
rect 1810 8602 1849 8636
rect 1883 8602 1922 8636
rect 1956 8602 1995 8636
rect 2029 8602 2068 8636
rect 2102 8602 2141 8636
rect 2175 8602 2209 8636
tri 2209 8602 2243 8636 nw
tri 3421 8602 3455 8636 ne
rect 3455 8602 3477 8636
rect 3511 8602 3550 8636
rect 3584 8602 3623 8636
rect 3657 8602 3696 8636
rect 3730 8602 3769 8636
rect 3803 8602 3842 8636
rect 3876 8602 3915 8636
rect 3949 8602 3988 8636
rect 4022 8602 4061 8636
rect 4095 8602 4134 8636
rect 4168 8602 4207 8636
rect 4241 8602 4280 8636
rect 4314 8602 4353 8636
rect 4387 8602 4426 8636
rect 4460 8602 4499 8636
rect 4533 8602 4572 8636
rect 4606 8602 4645 8636
rect 4679 8602 4718 8636
rect 4752 8602 4791 8636
rect 4825 8602 4864 8636
rect 4898 8602 4937 8636
rect 4971 8602 5010 8636
rect 5044 8602 5083 8636
rect 5117 8602 5156 8636
rect 5190 8602 5229 8636
rect 5263 8602 5302 8636
rect 5336 8602 5375 8636
rect 5409 8602 5448 8636
rect 5482 8602 5521 8636
rect 5555 8602 5594 8636
rect 5628 8602 5667 8636
rect 5701 8602 5740 8636
rect 5774 8602 5813 8636
rect 5847 8602 5886 8636
rect 5920 8602 5959 8636
rect 5993 8602 6032 8636
rect 6066 8602 6105 8636
rect 6139 8602 6178 8636
rect 6212 8602 6251 8636
rect 6285 8602 6324 8636
rect 6358 8602 6397 8636
rect 6431 8602 6470 8636
rect 6504 8602 6543 8636
rect 6577 8602 6616 8636
rect 6650 8602 6689 8636
rect 6723 8602 6762 8636
rect 6796 8602 6835 8636
rect 6869 8602 6908 8636
rect 6942 8602 6981 8636
rect 7015 8602 7054 8636
rect 7088 8602 7127 8636
rect 7161 8602 7200 8636
rect 7234 8602 7273 8636
rect 7307 8602 7346 8636
rect 7380 8602 7419 8636
rect 7453 8602 7492 8636
rect 7526 8602 7565 8636
rect 7599 8602 7638 8636
rect 7672 8602 7711 8636
rect 7745 8602 7784 8636
rect 7818 8602 7857 8636
rect 7891 8602 7930 8636
rect 7964 8602 8003 8636
rect 8037 8602 8075 8636
rect 8109 8602 8147 8636
rect 8181 8602 8219 8636
rect 8253 8602 8291 8636
rect 8325 8602 8363 8636
rect 8397 8602 8435 8636
rect 8469 8602 8507 8636
rect 8541 8602 8579 8636
rect 8613 8602 8651 8636
rect 8685 8602 8723 8636
rect 8757 8602 8795 8636
rect 8829 8602 8867 8636
rect 8901 8602 8939 8636
rect 8973 8602 9011 8636
rect 9045 8602 9083 8636
rect 9117 8602 9155 8636
rect 9189 8602 9227 8636
rect 9261 8602 9299 8636
rect 9333 8602 9371 8636
rect 9405 8602 9443 8636
rect 9477 8602 9515 8636
rect 9549 8602 9587 8636
rect 9621 8602 9659 8636
rect 9693 8602 9731 8636
rect 9765 8602 9803 8636
rect 9837 8602 9875 8636
rect 9909 8602 9947 8636
rect 9981 8602 10019 8636
rect 10053 8602 10091 8636
rect 10125 8602 10163 8636
rect 10197 8602 10235 8636
rect 10269 8602 10307 8636
rect 10341 8602 10379 8636
rect 10413 8602 10451 8636
rect 10485 8602 10523 8636
rect 10557 8602 10595 8636
rect 10629 8602 10667 8636
rect 10701 8602 10739 8636
rect 10773 8602 10811 8636
rect 10845 8602 10883 8636
rect 10917 8602 10955 8636
rect 10989 8602 11027 8636
rect 11061 8602 11099 8636
rect 11133 8602 11171 8636
rect 11205 8602 11243 8636
rect 11277 8602 11315 8636
rect 11349 8602 11387 8636
rect 11421 8602 11459 8636
rect 11493 8602 11531 8636
rect 11565 8602 11603 8636
rect 11637 8602 11675 8636
rect 11709 8602 11747 8636
rect 11781 8602 11819 8636
rect 11853 8602 11891 8636
rect 11925 8602 11963 8636
rect 11997 8602 12035 8636
rect 12069 8602 12107 8636
rect 12141 8602 12179 8636
rect 12213 8602 12251 8636
rect 12285 8602 12323 8636
rect 12357 8602 12395 8636
rect 12429 8602 12467 8636
rect 12501 8602 12539 8636
rect 12573 8602 12611 8636
rect 12645 8602 12683 8636
rect 12717 8602 12755 8636
rect 12789 8602 12827 8636
rect 12861 8602 12899 8636
rect 12933 8602 12971 8636
rect 13005 8602 13043 8636
rect 13077 8602 13115 8636
rect 13149 8602 13187 8636
rect 13221 8602 13259 8636
rect 13293 8602 13331 8636
rect 13365 8602 13403 8636
rect 13437 8602 13475 8636
rect 13509 8602 13547 8636
rect 13581 8602 13619 8636
rect 13653 8602 13691 8636
rect 13725 8602 13763 8636
rect 13797 8602 13835 8636
rect 13869 8602 13907 8636
rect 13941 8602 13979 8636
rect 14013 8602 14051 8636
rect 14085 8602 14123 8636
rect 14157 8602 14195 8636
rect 14229 8628 14240 8636
rect 14301 8628 14312 8636
rect 14373 8628 14384 8636
rect 14445 8628 14456 8636
rect 14517 8628 14528 8636
rect 14589 8628 14600 8636
rect 14229 8615 14267 8628
rect 14301 8615 14339 8628
rect 14373 8615 14411 8628
rect 14445 8615 14483 8628
rect 14517 8615 14555 8628
rect 14589 8615 14627 8628
rect 14229 8602 14240 8615
rect 14301 8602 14312 8615
rect 14373 8602 14384 8615
rect 14445 8602 14456 8615
rect 14517 8602 14528 8615
rect 14589 8602 14600 8615
rect 14661 8602 14699 8636
rect 14733 8602 14771 8636
rect 14805 8602 14843 8636
rect 14877 8602 15114 8636
tri 825 8595 832 8602 ne
rect 832 8595 2194 8602
tri 832 8587 840 8595 ne
rect 840 8587 2194 8595
tri 2194 8587 2209 8602 nw
tri 3455 8596 3461 8602 ne
rect 3461 8596 14240 8602
tri 3461 8587 3470 8596 ne
rect 3470 8587 14240 8596
tri 13739 8558 13768 8587 ne
rect 13768 8563 14240 8587
rect 14292 8563 14312 8602
rect 14364 8563 14384 8602
rect 14436 8563 14456 8602
rect 14508 8563 14528 8602
rect 14580 8563 14600 8602
rect 14652 8563 15114 8602
rect 13768 8558 15114 8563
tri 13768 8546 13780 8558 ne
rect 13780 8550 15114 8558
rect 13780 8546 14240 8550
tri 13780 8512 13814 8546 ne
rect 13814 8512 13992 8546
rect 14026 8512 14076 8546
rect 14110 8512 14240 8546
tri 13814 8478 13848 8512 ne
rect 13848 8478 14185 8512
rect 14219 8498 14240 8512
rect 14292 8498 14312 8550
rect 14364 8498 14384 8550
rect 14436 8498 14456 8550
rect 14508 8498 14528 8550
rect 14580 8498 14600 8550
rect 14652 8498 15114 8550
rect 14219 8485 14257 8498
rect 14291 8485 14329 8498
rect 14363 8485 14401 8498
rect 14435 8485 14473 8498
rect 14507 8485 15114 8498
rect 14219 8478 14240 8485
tri 13848 8474 13852 8478 ne
rect 13852 8474 14240 8478
tri 13852 8440 13886 8474 ne
rect 13886 8440 13992 8474
rect 14026 8440 14076 8474
rect 14110 8440 14240 8474
tri 13886 8435 13891 8440 ne
rect 13891 8435 14240 8440
tri 13891 8401 13925 8435 ne
rect 13925 8401 14185 8435
rect 14219 8433 14240 8435
rect 14292 8433 14312 8485
rect 14364 8433 14384 8485
rect 14436 8433 14456 8485
rect 14508 8433 14528 8485
rect 14580 8433 14600 8485
rect 14652 8462 15114 8485
rect 14652 8433 14692 8462
rect 14219 8420 14257 8433
rect 14291 8420 14329 8433
rect 14363 8420 14401 8433
rect 14435 8420 14473 8433
rect 14507 8428 14614 8433
rect 14648 8428 14692 8433
rect 14726 8428 14770 8462
rect 14804 8428 14848 8462
rect 14882 8428 14926 8462
rect 14960 8428 15004 8462
rect 15038 8428 15114 8462
rect 14507 8420 15114 8428
rect 14219 8401 14240 8420
tri 13925 8398 13928 8401 ne
rect 13928 8398 13992 8401
tri 402 8361 406 8365 se
rect 406 8361 458 8365
rect 235 8359 458 8361
rect 235 8355 406 8359
rect 235 8321 248 8355
rect 282 8321 320 8355
rect 354 8321 392 8355
rect 235 8315 406 8321
tri 372 8314 373 8315 ne
rect 373 8314 406 8315
tri 373 8287 400 8314 ne
rect 400 8307 406 8314
rect 400 8295 458 8307
rect 400 8287 406 8295
tri 400 8281 406 8287 ne
rect 2444 8355 2647 8398
tri 13928 8367 13959 8398 ne
rect 13959 8367 13992 8398
rect 14026 8367 14076 8401
rect 14110 8368 14240 8401
rect 14292 8368 14312 8420
rect 14364 8368 14384 8420
rect 14436 8368 14456 8420
rect 14508 8368 14528 8420
rect 14580 8368 14600 8420
rect 14652 8388 15114 8420
rect 14652 8368 14692 8388
rect 14110 8367 14614 8368
tri 13959 8358 13968 8367 ne
rect 13968 8358 14614 8367
tri 13968 8355 13971 8358 ne
rect 13971 8355 14185 8358
rect 2444 8321 2456 8355
rect 2490 8321 2528 8355
rect 2562 8321 2600 8355
rect 2634 8321 2647 8355
tri 13971 8324 14002 8355 ne
rect 14002 8324 14185 8355
rect 14219 8354 14257 8358
rect 14291 8354 14329 8358
rect 14363 8354 14401 8358
rect 14435 8354 14473 8358
rect 14507 8354 14614 8358
rect 14648 8354 14692 8368
rect 14726 8354 14770 8388
rect 14804 8354 14848 8388
rect 14882 8354 14926 8388
rect 14960 8354 15004 8388
rect 15038 8354 15114 8388
rect 14219 8324 14240 8354
rect 2444 8268 2647 8321
tri 14002 8314 14012 8324 ne
rect 14012 8314 14240 8324
tri 14012 8287 14039 8314 ne
rect 14039 8302 14240 8314
rect 14292 8302 14312 8354
rect 14364 8302 14384 8354
rect 14436 8302 14456 8354
rect 14508 8302 14528 8354
rect 14580 8302 14600 8354
rect 14652 8314 15114 8354
rect 14652 8302 14692 8314
rect 14039 8288 14614 8302
rect 14648 8288 14692 8302
rect 14039 8287 14240 8288
rect 10798 8281 11156 8287
tri 7008 8254 7014 8260 se
rect 7014 8254 8627 8260
rect 406 8235 458 8243
tri 6989 8235 7008 8254 se
rect 7008 8235 8509 8254
tri 6686 7932 6989 8235 se
rect 6989 7932 8509 8235
rect 8615 7932 8627 8254
rect 9590 8247 9881 8259
rect 9883 8258 10183 8259
rect 9590 8213 9596 8247
rect 9630 8213 9678 8247
rect 9712 8213 9881 8247
rect 9590 8144 9881 8213
rect 9590 8110 9596 8144
rect 9630 8110 9678 8144
rect 9712 8110 9881 8144
rect 9590 8041 9881 8110
rect 9590 8007 9596 8041
rect 9630 8007 9678 8041
rect 9712 8007 9881 8041
rect 9590 7995 9881 8007
rect 9882 7996 10184 8258
rect 10185 8247 10436 8259
rect 10185 8213 10314 8247
rect 10348 8213 10396 8247
rect 10430 8213 10436 8247
rect 10185 8144 10436 8213
rect 10185 8110 10314 8144
rect 10348 8110 10396 8144
rect 10430 8110 10436 8144
rect 10185 8041 10436 8110
rect 10185 8007 10314 8041
rect 10348 8007 10396 8041
rect 10430 8007 10436 8041
rect 9883 7995 10183 7996
rect 10185 7995 10436 8007
rect 10798 8229 10800 8281
rect 10852 8229 10876 8281
rect 10928 8254 10952 8281
rect 10932 8229 10952 8254
rect 11004 8229 11028 8281
rect 11080 8229 11104 8281
rect 10798 8220 10804 8229
rect 10838 8220 10898 8229
rect 10932 8220 11156 8229
rect 10798 8214 11156 8220
rect 10798 8162 10800 8214
rect 10852 8162 10876 8214
rect 10928 8179 10952 8214
rect 10932 8162 10952 8179
rect 11004 8162 11028 8214
rect 11080 8162 11104 8214
rect 10798 8147 10804 8162
rect 10838 8147 10898 8162
rect 10932 8147 11156 8162
rect 10798 8095 10800 8147
rect 10852 8095 10876 8147
rect 10932 8145 10952 8147
rect 10928 8104 10952 8145
rect 10932 8095 10952 8104
rect 11004 8095 11028 8147
rect 11080 8095 11104 8147
rect 10798 8079 10804 8095
rect 10838 8079 10898 8095
rect 10932 8079 11156 8095
rect 10798 8027 10800 8079
rect 10852 8027 10876 8079
rect 10932 8070 10952 8079
rect 10928 8028 10952 8070
rect 10932 8027 10952 8028
rect 11004 8027 11028 8079
rect 11080 8027 11104 8079
rect 10798 8011 10804 8027
rect 10838 8011 10898 8027
rect 10932 8011 11156 8027
tri 6672 7918 6686 7932 se
rect 6686 7926 8627 7932
rect 10798 7959 10800 8011
rect 10852 7959 10876 8011
rect 10932 7994 10952 8011
rect 10928 7959 10952 7994
rect 11004 7959 11028 8011
rect 11080 7959 11104 8011
rect 10798 7952 11156 7959
rect 10798 7943 10804 7952
rect 10838 7943 10898 7952
rect 10932 7943 11156 7952
rect 6686 7918 7144 7926
tri 7144 7918 7152 7926 nw
tri 6670 7916 6672 7918 se
rect 6672 7916 7142 7918
tri 7142 7916 7144 7918 nw
tri 6664 7910 6670 7916 se
rect 6670 7910 7136 7916
tri 7136 7910 7142 7916 nw
tri 6660 7906 6664 7910 se
rect 6664 7906 7132 7910
tri 7132 7906 7136 7910 nw
tri 6624 7870 6660 7906 se
rect 6660 7870 7096 7906
tri 7096 7870 7132 7906 nw
rect 10798 7891 10800 7943
rect 10852 7891 10876 7943
rect 10932 7918 10952 7943
rect 10928 7891 10952 7918
rect 11004 7891 11028 7943
rect 11080 7891 11104 7943
rect 10798 7885 11156 7891
rect 12252 8281 12622 8287
rect 12252 8229 12255 8281
rect 12307 8229 12333 8281
rect 12385 8229 12411 8281
rect 12463 8229 12489 8281
rect 12541 8229 12567 8281
rect 12619 8229 12622 8281
tri 14039 8280 14046 8287 ne
rect 14046 8280 14240 8287
tri 14046 8257 14069 8280 ne
rect 14069 8257 14185 8280
rect 12252 8210 12622 8229
rect 12252 8158 12255 8210
rect 12307 8158 12333 8210
rect 12385 8158 12411 8210
rect 12463 8158 12489 8210
rect 12541 8158 12567 8210
rect 12619 8158 12622 8210
rect 12252 8139 12622 8158
rect 12252 8087 12255 8139
rect 12307 8087 12333 8139
rect 12385 8087 12411 8139
rect 12463 8087 12489 8139
rect 12541 8087 12567 8139
rect 12619 8087 12622 8139
rect 12252 8068 12622 8087
rect 12252 8016 12255 8068
rect 12307 8016 12333 8068
rect 12385 8016 12411 8068
rect 12463 8016 12489 8068
rect 12541 8016 12567 8068
rect 12619 8033 12622 8068
tri 12622 8033 12645 8056 sw
rect 12619 8016 12645 8033
rect 12252 7999 12645 8016
tri 12645 7999 12679 8033 sw
rect 12252 7997 12679 7999
rect 12252 7945 12255 7997
rect 12307 7945 12333 7997
rect 12385 7945 12411 7997
rect 12463 7945 12489 7997
rect 12541 7945 12567 7997
rect 12619 7984 12679 7997
tri 12679 7984 12694 7999 sw
rect 12619 7950 12694 7984
tri 12694 7950 12728 7984 sw
rect 12619 7945 12728 7950
rect 12252 7925 12728 7945
rect 12252 7873 12255 7925
rect 12307 7873 12333 7925
rect 12385 7873 12411 7925
rect 12463 7873 12489 7925
rect 12541 7873 12567 7925
rect 12619 7916 12728 7925
tri 12728 7916 12762 7950 sw
rect 13310 7924 13365 8257
tri 14069 8246 14080 8257 ne
rect 14080 8246 14185 8257
rect 14219 8246 14240 8280
tri 14080 8240 14086 8246 ne
rect 14086 8240 14240 8246
tri 14086 8206 14120 8240 ne
rect 14120 8236 14240 8240
rect 14292 8236 14312 8288
rect 14364 8236 14384 8288
rect 14436 8236 14456 8288
rect 14508 8236 14528 8288
rect 14580 8236 14600 8288
rect 14652 8280 14692 8288
rect 14726 8280 14770 8314
rect 14804 8280 14848 8314
rect 14882 8280 14926 8314
rect 14960 8280 15004 8314
rect 15038 8280 15114 8314
rect 14652 8240 15114 8280
rect 14652 8236 14692 8240
rect 14120 8222 14614 8236
rect 14648 8222 14692 8236
rect 14120 8206 14240 8222
tri 14120 8202 14124 8206 ne
rect 14124 8202 14240 8206
tri 14124 8168 14158 8202 ne
rect 14158 8168 14185 8202
rect 14219 8170 14240 8202
rect 14292 8170 14312 8222
rect 14364 8170 14384 8222
rect 14436 8170 14456 8222
rect 14508 8170 14528 8222
rect 14580 8170 14600 8222
rect 14652 8206 14692 8222
rect 14726 8206 14770 8240
rect 14804 8206 14848 8240
rect 14882 8206 14926 8240
rect 14960 8206 15004 8240
rect 15038 8206 15114 8240
rect 14652 8170 15114 8206
rect 14219 8168 14257 8170
rect 14291 8168 14329 8170
rect 14363 8168 14401 8170
rect 14435 8168 14473 8170
rect 14507 8168 15114 8170
tri 14158 8166 14160 8168 ne
rect 14160 8166 15114 8168
tri 14160 8156 14170 8166 ne
rect 14170 8156 14614 8166
rect 14648 8156 14692 8166
tri 14170 8132 14194 8156 ne
rect 14194 8132 14240 8156
tri 14194 8115 14211 8132 ne
rect 14211 8115 14240 8132
tri 14211 8098 14228 8115 ne
rect 14228 8104 14240 8115
rect 14292 8104 14312 8156
rect 14364 8104 14384 8156
rect 14436 8115 14456 8156
rect 14508 8115 14528 8156
rect 14508 8104 14511 8115
rect 14580 8104 14600 8156
rect 14652 8132 14692 8156
rect 14726 8132 14770 8166
rect 14804 8132 14848 8166
rect 14882 8132 14926 8166
rect 14960 8132 15004 8166
rect 15038 8132 15114 8166
rect 14652 8104 15114 8132
rect 14228 8098 14431 8104
tri 14228 8081 14245 8098 ne
rect 14245 8081 14431 8098
rect 14465 8081 14511 8104
rect 14545 8092 15114 8104
rect 14545 8081 14614 8092
tri 14245 8058 14268 8081 ne
rect 14268 8058 14614 8081
rect 14648 8058 14692 8092
rect 14726 8058 14770 8092
rect 14804 8058 14848 8092
rect 14882 8058 14926 8092
rect 14960 8058 15004 8092
rect 15038 8058 15114 8092
tri 14268 8056 14270 8058 ne
rect 14270 8056 15114 8058
tri 14270 8033 14293 8056 ne
rect 14293 8033 15114 8056
tri 14293 7999 14327 8033 ne
rect 14327 7999 14431 8033
rect 14465 7999 14511 8033
rect 14545 8018 15114 8033
rect 14545 7999 14614 8018
tri 14327 7984 14342 7999 ne
rect 14342 7984 14614 7999
rect 14648 7984 14692 8018
rect 14726 7984 14770 8018
rect 14804 7984 14848 8018
rect 14882 7984 14926 8018
rect 14960 7984 15004 8018
rect 15038 7984 15114 8018
tri 14342 7950 14376 7984 ne
rect 14376 7950 15114 7984
tri 14376 7924 14402 7950 ne
rect 14402 7924 14431 7950
tri 14402 7916 14410 7924 ne
rect 14410 7916 14431 7924
rect 14465 7916 14511 7950
rect 14545 7944 15114 7950
rect 14545 7916 14614 7944
rect 12619 7910 12762 7916
tri 12762 7910 12768 7916 sw
tri 14410 7910 14416 7916 ne
rect 14416 7910 14614 7916
rect 14648 7910 14692 7944
rect 14726 7910 14770 7944
rect 14804 7910 14848 7944
rect 14882 7910 14926 7944
rect 14960 7910 15004 7944
rect 15038 7910 15114 7944
rect 12619 7904 12768 7910
tri 12768 7904 12774 7910 sw
tri 14416 7904 14422 7910 ne
rect 14422 7904 15114 7910
rect 12619 7885 12774 7904
tri 12774 7885 12793 7904 sw
tri 14422 7885 14441 7904 ne
rect 14441 7885 15114 7904
rect 12619 7873 12793 7885
rect 12252 7870 12793 7873
tri 12793 7870 12808 7885 sw
tri 14441 7870 14456 7885 ne
rect 14456 7870 15114 7885
tri 6611 7857 6624 7870 se
rect 6624 7857 7083 7870
tri 7083 7857 7096 7870 nw
rect 12252 7867 12808 7870
tri 12808 7867 12811 7870 sw
tri 14456 7867 14459 7870 ne
rect 14459 7867 14614 7870
tri 12563 7857 12573 7867 ne
rect 12573 7857 12811 7867
tri 12811 7857 12821 7867 sw
tri 14459 7857 14469 7867 ne
rect 14469 7857 14614 7867
rect 278 7851 7062 7857
rect 330 7836 7062 7851
tri 7062 7836 7083 7857 nw
tri 12573 7836 12594 7857 ne
rect 12594 7836 12821 7857
tri 12821 7836 12842 7857 sw
tri 14469 7836 14490 7857 ne
rect 14490 7836 14614 7857
rect 14648 7836 14692 7870
rect 14726 7836 14770 7870
rect 14804 7836 14848 7870
rect 14882 7836 14926 7870
rect 14960 7836 15004 7870
rect 15038 7836 15114 7870
rect 330 7799 7022 7836
rect 278 7796 7022 7799
tri 7022 7796 7062 7836 nw
tri 12594 7796 12634 7836 ne
rect 12634 7796 12842 7836
tri 12842 7796 12882 7836 sw
tri 14490 7796 14530 7836 ne
rect 14530 7796 15114 7836
rect 278 7785 6988 7796
rect 330 7762 6988 7785
tri 6988 7762 7022 7796 nw
tri 12634 7785 12645 7796 ne
rect 12645 7785 12882 7796
tri 12882 7785 12893 7796 sw
tri 14530 7785 14541 7796 ne
rect 14541 7785 14614 7796
tri 12645 7762 12668 7785 ne
rect 12668 7762 12893 7785
tri 12893 7762 12916 7785 sw
tri 14541 7762 14564 7785 ne
rect 14564 7762 14614 7785
rect 14648 7762 14692 7796
rect 14726 7762 14770 7796
rect 14804 7762 14848 7796
rect 14882 7762 14926 7796
rect 14960 7762 15004 7796
rect 15038 7762 15114 7796
rect 330 7733 6948 7762
rect 278 7722 6948 7733
tri 6948 7722 6988 7762 nw
tri 12668 7722 12708 7762 ne
rect 12708 7722 12916 7762
tri 12916 7722 12956 7762 sw
tri 14564 7722 14604 7762 ne
rect 14604 7722 15114 7762
rect 278 7718 6914 7722
rect 330 7688 6914 7718
tri 6914 7688 6948 7722 nw
tri 12708 7688 12742 7722 ne
rect 12742 7718 12956 7722
tri 12956 7718 12960 7722 sw
tri 14604 7718 14608 7722 ne
rect 12742 7688 12960 7718
tri 12960 7688 12990 7718 sw
rect 14608 7688 14614 7722
rect 14648 7688 14692 7722
rect 14726 7688 14770 7722
rect 14804 7688 14848 7722
rect 14882 7688 14926 7722
rect 14960 7688 15004 7722
rect 15038 7688 15114 7722
rect 330 7666 6874 7688
rect 278 7651 6874 7666
tri 25 7614 27 7616 sw
rect 25 7574 27 7614
tri 27 7574 67 7614 sw
rect 330 7648 6874 7651
tri 6874 7648 6914 7688 nw
tri 12742 7648 12782 7688 ne
rect 12782 7648 12990 7688
tri 12990 7648 13030 7688 sw
rect 14608 7648 15114 7688
rect 330 7614 6840 7648
tri 6840 7614 6874 7648 nw
tri 12782 7614 12816 7648 ne
rect 12816 7614 13030 7648
tri 13030 7614 13064 7648 sw
rect 14608 7614 14614 7648
rect 14648 7614 14692 7648
rect 14726 7614 14770 7648
rect 14804 7614 14848 7648
rect 14882 7614 14926 7648
rect 14960 7614 15004 7648
rect 15038 7614 15114 7648
rect 330 7599 6800 7614
rect 278 7584 6800 7599
rect 25 7540 67 7574
tri 67 7540 101 7574 sw
rect 25 7526 101 7540
tri 101 7526 115 7540 sw
rect 330 7574 6800 7584
tri 6800 7574 6840 7614 nw
tri 12816 7574 12856 7614 ne
rect 12856 7574 13064 7614
tri 13064 7574 13104 7614 sw
rect 14608 7574 15114 7614
rect 330 7561 6787 7574
tri 6787 7561 6800 7574 nw
tri 12856 7561 12869 7574 ne
rect 12869 7561 13104 7574
tri 13104 7561 13117 7574 sw
rect 330 7540 6766 7561
tri 6766 7540 6787 7561 nw
rect 330 7532 6752 7540
rect 278 7526 6752 7532
tri 6752 7526 6766 7540 nw
rect 25 7499 115 7526
tri 115 7499 142 7526 sw
rect 11129 7509 11135 7561
rect 11187 7509 11208 7561
rect 11260 7509 11280 7561
rect 11332 7509 11338 7561
tri 12869 7540 12890 7561 ne
rect 12890 7540 13117 7561
tri 13117 7540 13138 7561 sw
rect 14608 7540 14614 7574
rect 14648 7540 14692 7574
rect 14726 7540 14770 7574
rect 14804 7540 14848 7574
rect 14882 7540 14926 7574
rect 14960 7540 15004 7574
rect 15038 7540 15114 7574
tri 12890 7537 12893 7540 ne
rect 25 7465 142 7499
tri 142 7465 176 7499 sw
rect 11129 7481 11338 7509
rect 25 7429 176 7465
tri 176 7429 212 7465 sw
rect 11129 7429 11135 7481
rect 11187 7429 11208 7481
rect 11260 7429 11280 7481
rect 11332 7429 11338 7481
rect 12893 7499 13138 7540
tri 13138 7499 13179 7540 sw
rect 14608 7499 15114 7540
rect 12893 7465 13179 7499
tri 13179 7465 13213 7499 sw
rect 14608 7465 14614 7499
rect 14648 7465 14692 7499
rect 14726 7465 14770 7499
rect 14804 7465 14848 7499
rect 14882 7465 14926 7499
rect 14960 7465 15004 7499
rect 15038 7465 15114 7499
rect 12893 7435 13213 7465
tri 13213 7435 13243 7465 sw
rect 25 7424 212 7429
tri 212 7424 217 7429 sw
rect 25 7390 217 7424
tri 217 7390 251 7424 sw
rect 25 7381 251 7390
tri 251 7381 260 7390 sw
rect 25 7374 1405 7381
rect 25 7340 57 7374
rect 91 7340 132 7374
rect 166 7340 207 7374
rect 241 7340 282 7374
rect 316 7340 357 7374
rect 391 7340 432 7374
rect 466 7340 507 7374
rect 541 7340 582 7374
rect 616 7340 657 7374
rect 691 7340 732 7374
rect 766 7340 807 7374
rect 841 7340 882 7374
rect 916 7340 957 7374
rect 991 7340 1032 7374
rect 1066 7340 1107 7374
rect 1141 7340 1182 7374
rect 1216 7340 1256 7374
rect 1290 7340 1330 7374
rect 1364 7349 1405 7374
tri 1405 7349 1437 7381 sw
rect 1364 7340 1437 7349
rect 25 7315 1437 7340
tri 1437 7315 1471 7349 sw
rect 25 7290 1471 7315
rect 25 7256 57 7290
rect 91 7256 132 7290
rect 166 7256 207 7290
rect 241 7256 282 7290
rect 316 7256 357 7290
rect 391 7256 432 7290
rect 466 7256 507 7290
rect 541 7256 582 7290
rect 616 7256 657 7290
rect 691 7256 732 7290
rect 766 7256 807 7290
rect 841 7256 882 7290
rect 916 7256 957 7290
rect 991 7256 1032 7290
rect 1066 7256 1107 7290
rect 1141 7256 1182 7290
rect 1216 7256 1256 7290
rect 1290 7256 1330 7290
rect 1364 7274 1471 7290
tri 1471 7274 1512 7315 sw
rect 1364 7256 1512 7274
rect 25 7240 1512 7256
tri 1512 7240 1546 7274 sw
rect 25 7226 1546 7240
tri 1546 7226 1560 7240 sw
rect 25 7220 7162 7226
rect 25 7206 1431 7220
rect 25 7172 57 7206
rect 91 7172 132 7206
rect 166 7172 207 7206
rect 241 7172 282 7206
rect 316 7172 357 7206
rect 391 7172 432 7206
rect 466 7172 507 7206
rect 541 7172 582 7206
rect 616 7172 657 7206
rect 691 7172 732 7206
rect 766 7172 807 7206
rect 841 7172 882 7206
rect 916 7172 957 7206
rect 991 7172 1032 7206
rect 1066 7172 1107 7206
rect 1141 7172 1182 7206
rect 1216 7172 1256 7206
rect 1290 7172 1330 7206
rect 1364 7186 1431 7206
rect 1465 7186 1504 7220
rect 1538 7186 1577 7220
rect 1611 7186 1650 7220
rect 1684 7186 1723 7220
rect 1757 7186 1796 7220
rect 1830 7186 1869 7220
rect 1903 7186 1942 7220
rect 1976 7186 2015 7220
rect 2049 7186 2088 7220
rect 2122 7186 2161 7220
rect 2195 7186 2234 7220
rect 2268 7186 2307 7220
rect 2341 7186 2380 7220
rect 2414 7186 2453 7220
rect 2487 7186 2526 7220
rect 2560 7186 2599 7220
rect 2633 7186 2672 7220
rect 2706 7186 2745 7220
rect 2779 7186 2818 7220
rect 2852 7186 2891 7220
rect 2925 7186 2964 7220
rect 2998 7186 3037 7220
rect 3071 7186 3110 7220
rect 3144 7186 3183 7220
rect 3217 7186 3256 7220
rect 3290 7186 3329 7220
rect 3363 7186 3402 7220
rect 3436 7186 3475 7220
rect 3509 7186 3548 7220
rect 3582 7186 3621 7220
rect 3655 7186 3694 7220
rect 3728 7186 3767 7220
rect 3801 7186 3840 7220
rect 3874 7186 3913 7220
rect 3947 7186 3986 7220
rect 4020 7186 4059 7220
rect 4093 7186 4132 7220
rect 4166 7186 4205 7220
rect 4239 7186 4278 7220
rect 4312 7186 4351 7220
rect 4385 7186 4424 7220
rect 4458 7186 4497 7220
rect 4531 7186 4570 7220
rect 4604 7186 4643 7220
rect 4677 7186 4716 7220
rect 4750 7186 4789 7220
rect 4823 7186 4862 7220
rect 4896 7186 4935 7220
rect 4969 7186 5008 7220
rect 5042 7186 5081 7220
rect 5115 7186 5154 7220
rect 5188 7186 5227 7220
rect 5261 7186 5300 7220
rect 5334 7186 5373 7220
rect 5407 7186 5446 7220
rect 5480 7186 5519 7220
rect 5553 7186 5592 7220
rect 5626 7186 5665 7220
rect 5699 7186 5738 7220
rect 5772 7186 5811 7220
rect 5845 7186 5884 7220
rect 5918 7186 5957 7220
rect 5991 7186 6030 7220
rect 6064 7186 6103 7220
rect 6137 7186 6176 7220
rect 6210 7186 6249 7220
rect 6283 7186 6322 7220
rect 6356 7186 6395 7220
rect 6429 7186 6468 7220
rect 6502 7186 6540 7220
rect 6574 7186 6612 7220
rect 6646 7186 6684 7220
rect 6718 7186 6756 7220
rect 6790 7186 6828 7220
rect 6862 7186 6900 7220
rect 6934 7186 6972 7220
rect 7006 7186 7044 7220
rect 7078 7186 7116 7220
rect 7150 7186 7162 7220
rect 1364 7180 7162 7186
rect 1364 7172 1564 7180
rect 25 7165 1564 7172
tri 1564 7165 1579 7180 nw
rect 25 7125 1524 7165
tri 1524 7125 1564 7165 nw
rect 25 7124 1523 7125
tri 1523 7124 1524 7125 nw
tri 7474 7124 7475 7125 se
rect 7475 7124 7873 7125
rect 25 7122 1489 7124
rect 25 7088 57 7122
rect 91 7088 132 7122
rect 166 7088 207 7122
rect 241 7088 282 7122
rect 316 7088 357 7122
rect 391 7088 432 7122
rect 466 7088 507 7122
rect 541 7088 582 7122
rect 616 7088 657 7122
rect 691 7088 732 7122
rect 766 7088 807 7122
rect 841 7088 882 7122
rect 916 7088 957 7122
rect 991 7088 1032 7122
rect 1066 7088 1107 7122
rect 1141 7088 1182 7122
rect 1216 7088 1256 7122
rect 1290 7088 1330 7122
rect 1364 7090 1489 7122
tri 1489 7090 1523 7124 nw
tri 7440 7090 7474 7124 se
rect 7474 7090 7873 7124
rect 1364 7088 1396 7090
rect 25 7038 1396 7088
rect 25 7004 57 7038
rect 91 7004 132 7038
rect 166 7004 207 7038
rect 241 7004 282 7038
rect 316 7004 357 7038
rect 391 7004 432 7038
rect 466 7004 507 7038
rect 541 7004 582 7038
rect 616 7004 657 7038
rect 691 7004 732 7038
rect 766 7004 807 7038
rect 841 7004 882 7038
rect 916 7004 957 7038
rect 991 7004 1032 7038
rect 1066 7004 1107 7038
rect 1141 7004 1182 7038
rect 1216 7004 1256 7038
rect 1290 7004 1330 7038
rect 1364 7004 1396 7038
rect 25 6997 1396 7004
tri 1396 6997 1489 7090 nw
tri 7347 6997 7440 7090 se
rect 7440 6997 7873 7090
tri 7291 6941 7347 6997 se
rect 7347 6995 7873 6997
rect 7347 6941 7475 6995
tri 7475 6941 7529 6995 nw
tri 7230 6880 7291 6941 se
rect 7291 6880 7414 6941
tri 7414 6880 7475 6941 nw
rect 338 6874 7359 6880
rect 390 6825 7359 6874
tri 7359 6825 7414 6880 nw
rect 390 6822 7325 6825
rect 338 6808 7325 6822
rect 390 6791 7325 6808
tri 7325 6791 7359 6825 nw
rect 390 6756 7287 6791
rect 338 6753 7287 6756
tri 7287 6753 7325 6791 nw
rect 338 6750 7284 6753
tri 7284 6750 7287 6753 nw
tri 12882 6647 12893 6658 se
rect 12893 6647 13243 7435
rect 14608 7424 15114 7465
rect 14608 7390 14614 7424
rect 14648 7390 14692 7424
rect 14726 7390 14770 7424
rect 14804 7390 14848 7424
rect 14882 7390 14926 7424
rect 14960 7390 15004 7424
rect 15038 7390 15114 7424
rect 14608 7349 15114 7390
rect 14608 7315 14614 7349
rect 14648 7315 14692 7349
rect 14726 7315 14770 7349
rect 14804 7315 14848 7349
rect 14882 7315 14926 7349
rect 14960 7315 15004 7349
rect 15038 7315 15114 7349
rect 14608 7274 15114 7315
rect 14608 7240 14614 7274
rect 14648 7240 14692 7274
rect 14726 7240 14770 7274
rect 14804 7240 14848 7274
rect 14882 7240 14926 7274
rect 14960 7240 15004 7274
rect 15038 7240 15114 7274
rect 14608 7199 15114 7240
rect 14608 7165 14614 7199
rect 14648 7165 14692 7199
rect 14726 7165 14770 7199
rect 14804 7165 14848 7199
rect 14882 7165 14926 7199
rect 14960 7165 15004 7199
rect 15038 7165 15114 7199
rect 14608 7124 15114 7165
rect 14608 7090 14614 7124
rect 14648 7090 14692 7124
rect 14726 7090 14770 7124
rect 14804 7090 14848 7124
rect 14882 7090 14926 7124
rect 14960 7090 15004 7124
rect 15038 7090 15114 7124
rect 14608 7053 15114 7090
rect 15062 6825 15108 6837
rect 15062 6791 15068 6825
rect 15102 6791 15108 6825
rect 15062 6753 15108 6791
rect 15062 6719 15068 6753
rect 15102 6719 15108 6753
rect 15062 6681 15108 6719
tri 13243 6647 13254 6658 sw
rect 15062 6647 15068 6681
rect 15102 6647 15108 6681
tri 12844 6609 12882 6647 se
rect 12882 6609 13254 6647
tri 13254 6609 13292 6647 sw
rect 15062 6609 15108 6647
tri 12810 6575 12844 6609 se
rect 12844 6575 13292 6609
tri 13292 6575 13326 6609 sw
rect 15062 6575 15068 6609
rect 15102 6575 15108 6609
tri 12772 6537 12810 6575 se
rect 12810 6537 13326 6575
tri 13326 6537 13364 6575 sw
rect 15062 6537 15108 6575
tri 12738 6503 12772 6537 se
rect 12772 6503 13364 6537
tri 13364 6503 13398 6537 sw
rect 15062 6503 15068 6537
rect 15102 6503 15108 6537
tri 12700 6465 12738 6503 se
rect 12738 6465 13398 6503
tri 13398 6465 13436 6503 sw
rect 15062 6465 15108 6503
tri 12685 6450 12700 6465 se
rect 12700 6450 13436 6465
tri 13436 6450 13451 6465 sw
rect 15062 6450 15068 6465
rect 56 6439 15068 6450
rect 56 6405 68 6439
rect 102 6405 141 6439
rect 175 6405 214 6439
rect 248 6405 287 6439
rect 321 6405 360 6439
rect 394 6405 433 6439
rect 467 6405 506 6439
rect 540 6405 579 6439
rect 613 6405 652 6439
rect 686 6405 725 6439
rect 759 6405 798 6439
rect 832 6405 871 6439
rect 905 6405 944 6439
rect 978 6405 1017 6439
rect 1051 6405 1090 6439
rect 56 6367 1090 6405
rect 56 6333 68 6367
rect 102 6333 141 6367
rect 175 6333 214 6367
rect 248 6333 287 6367
rect 321 6333 360 6367
rect 394 6333 433 6367
rect 467 6333 506 6367
rect 540 6333 579 6367
rect 613 6333 652 6367
rect 686 6333 725 6367
rect 759 6333 798 6367
rect 832 6333 871 6367
rect 905 6333 944 6367
rect 978 6333 1017 6367
rect 1051 6333 1090 6367
rect 56 6295 1090 6333
rect 56 6261 68 6295
rect 102 6261 141 6295
rect 175 6261 214 6295
rect 248 6261 287 6295
rect 321 6261 360 6295
rect 394 6261 433 6295
rect 467 6261 506 6295
rect 540 6261 579 6295
rect 613 6261 652 6295
rect 686 6261 725 6295
rect 759 6261 798 6295
rect 832 6261 871 6295
rect 905 6261 944 6295
rect 978 6261 1017 6295
rect 1051 6261 1090 6295
rect 56 6223 1090 6261
rect 56 6189 68 6223
rect 102 6189 141 6223
rect 175 6189 214 6223
rect 248 6189 287 6223
rect 321 6189 360 6223
rect 394 6189 433 6223
rect 467 6189 506 6223
rect 540 6189 579 6223
rect 613 6189 652 6223
rect 686 6189 725 6223
rect 759 6189 798 6223
rect 832 6189 871 6223
rect 905 6189 944 6223
rect 978 6189 1017 6223
rect 1051 6189 1090 6223
rect 56 6151 1090 6189
rect 56 6117 68 6151
rect 102 6117 141 6151
rect 175 6117 214 6151
rect 248 6117 287 6151
rect 321 6117 360 6151
rect 394 6117 433 6151
rect 467 6117 506 6151
rect 540 6117 579 6151
rect 613 6117 652 6151
rect 686 6117 725 6151
rect 759 6117 798 6151
rect 832 6117 871 6151
rect 905 6117 944 6151
rect 978 6117 1017 6151
rect 1051 6117 1090 6151
rect 15020 6431 15068 6439
rect 15102 6450 15108 6465
rect 15102 6431 15114 6450
rect 15020 6393 15114 6431
rect 15020 6359 15068 6393
rect 15102 6359 15114 6393
rect 15020 6321 15114 6359
rect 15020 6287 15068 6321
rect 15102 6287 15114 6321
rect 15020 6249 15114 6287
rect 15020 6215 15068 6249
rect 15102 6215 15114 6249
rect 15020 6177 15114 6215
rect 15020 6143 15068 6177
rect 15102 6143 15114 6177
rect 15020 6117 15114 6143
rect 56 6105 15114 6117
rect 56 6086 15068 6105
rect 14974 6071 15068 6086
rect 15102 6071 15114 6105
rect 14974 6033 15114 6071
rect 14974 5999 15068 6033
rect 15102 5999 15114 6033
rect 14974 5961 15114 5999
rect 14974 5927 15068 5961
rect 15102 5927 15114 5961
rect 14974 5889 15114 5927
rect 14974 5855 15068 5889
rect 15102 5855 15114 5889
rect 14974 5817 15114 5855
rect 14974 5783 15068 5817
rect 15102 5783 15114 5817
rect 14974 5745 15114 5783
rect 14974 5711 15068 5745
rect 15102 5711 15114 5745
rect 14974 5673 15114 5711
rect 14974 5639 15068 5673
rect 15102 5639 15114 5673
rect 14974 5601 15114 5639
rect 510 5568 809 5586
rect 510 5516 516 5568
rect 568 5516 634 5568
rect 686 5516 751 5568
rect 803 5516 809 5568
rect 510 5498 809 5516
rect 14249 5565 14371 5583
rect 14249 5513 14313 5565
rect 14365 5513 14371 5565
rect 14249 5495 14371 5513
rect 14974 5567 15068 5601
rect 15102 5567 15114 5601
rect 14974 5529 15114 5567
rect 14974 5495 15068 5529
rect 15102 5495 15114 5529
rect 435 5465 703 5471
rect 487 5413 507 5465
rect 559 5413 579 5465
rect 631 5413 651 5465
rect 742 5427 748 5479
rect 800 5427 811 5479
rect 14241 5465 14495 5471
rect 435 5400 703 5413
rect 487 5348 507 5400
rect 559 5348 579 5400
rect 631 5348 651 5400
rect 435 5335 703 5348
rect 487 5283 507 5335
rect 559 5283 579 5335
rect 631 5283 651 5335
rect 435 5270 703 5283
rect 487 5218 507 5270
rect 559 5218 579 5270
rect 631 5218 651 5270
rect 435 5205 703 5218
rect 487 5153 507 5205
rect 559 5153 579 5205
rect 631 5153 651 5205
rect 435 5140 703 5153
rect 487 5088 507 5140
rect 559 5088 579 5140
rect 631 5088 651 5140
rect 435 5075 703 5088
rect 487 5023 507 5075
rect 559 5023 579 5075
rect 631 5023 651 5075
rect 435 5010 703 5023
rect 487 4958 507 5010
rect 559 4958 579 5010
rect 631 4958 651 5010
rect 435 4945 703 4958
rect 487 4893 507 4945
rect 559 4893 579 4945
rect 631 4893 651 4945
rect 435 4880 703 4893
rect 487 4828 507 4880
rect 559 4828 579 4880
rect 631 4828 651 4880
rect 435 4815 703 4828
rect 487 4763 507 4815
rect 559 4763 579 4815
rect 631 4763 651 4815
rect 435 4750 703 4763
rect 487 4698 507 4750
rect 559 4698 579 4750
rect 631 4698 651 4750
rect 435 4685 703 4698
rect 487 4633 507 4685
rect 559 4633 579 4685
rect 631 4633 651 4685
rect 435 4620 703 4633
rect 487 4568 507 4620
rect 559 4568 579 4620
rect 631 4568 651 4620
rect 435 4555 703 4568
rect 487 4503 507 4555
rect 559 4503 579 4555
rect 631 4503 651 4555
rect 435 4490 703 4503
rect 487 4438 507 4490
rect 559 4438 579 4490
rect 631 4438 651 4490
rect 435 4425 703 4438
rect 487 4373 507 4425
rect 559 4373 579 4425
rect 631 4373 651 4425
rect 435 4360 703 4373
rect 487 4308 507 4360
rect 559 4308 579 4360
rect 631 4308 651 4360
rect 435 4295 703 4308
rect 487 4243 507 4295
rect 559 4243 579 4295
rect 631 4243 651 4295
rect 435 4230 703 4243
rect 487 4178 507 4230
rect 559 4178 579 4230
rect 631 4178 651 4230
rect 435 4165 703 4178
rect 487 4113 507 4165
rect 559 4113 579 4165
rect 631 4113 651 4165
rect 435 4099 703 4113
rect 487 4047 507 4099
rect 559 4047 579 4099
rect 631 4047 651 4099
rect 435 4033 703 4047
rect 487 3981 507 4033
rect 559 3981 579 4033
rect 631 3981 651 4033
rect 435 3967 703 3981
rect 487 3915 507 3967
rect 559 3915 579 3967
rect 631 3915 651 3967
rect 435 3901 703 3915
rect 487 3849 507 3901
rect 559 3849 579 3901
rect 631 3849 651 3901
rect 435 3835 703 3849
rect 487 3783 507 3835
rect 559 3783 579 3835
rect 631 3783 651 3835
rect 435 3769 703 3783
rect 487 3717 507 3769
rect 559 3717 579 3769
rect 631 3717 651 3769
rect 435 3703 703 3717
rect 487 3651 507 3703
rect 559 3651 579 3703
rect 631 3651 651 3703
rect 435 1923 703 3651
rect 14241 5413 14243 5465
rect 14295 5413 14309 5465
rect 14361 5413 14375 5465
rect 14427 5413 14441 5465
rect 14493 5413 14495 5465
rect 14241 5400 14495 5413
rect 14241 5348 14243 5400
rect 14295 5348 14309 5400
rect 14361 5348 14375 5400
rect 14427 5348 14441 5400
rect 14493 5348 14495 5400
rect 14241 5335 14495 5348
rect 14241 5283 14243 5335
rect 14295 5283 14309 5335
rect 14361 5283 14375 5335
rect 14427 5283 14441 5335
rect 14493 5283 14495 5335
rect 14241 5270 14495 5283
rect 14241 5218 14243 5270
rect 14295 5218 14309 5270
rect 14361 5218 14375 5270
rect 14427 5218 14441 5270
rect 14493 5218 14495 5270
rect 14241 5205 14495 5218
rect 14241 5153 14243 5205
rect 14295 5153 14309 5205
rect 14361 5153 14375 5205
rect 14427 5153 14441 5205
rect 14493 5153 14495 5205
rect 14241 5140 14495 5153
rect 14241 5088 14243 5140
rect 14295 5088 14309 5140
rect 14361 5088 14375 5140
rect 14427 5088 14441 5140
rect 14493 5088 14495 5140
rect 14241 5075 14495 5088
rect 14241 5023 14243 5075
rect 14295 5023 14309 5075
rect 14361 5023 14375 5075
rect 14427 5023 14441 5075
rect 14493 5023 14495 5075
rect 14241 5010 14495 5023
rect 14241 4958 14243 5010
rect 14295 4958 14309 5010
rect 14361 4958 14375 5010
rect 14427 4958 14441 5010
rect 14493 4958 14495 5010
rect 14241 4945 14495 4958
rect 14241 4893 14243 4945
rect 14295 4893 14309 4945
rect 14361 4893 14375 4945
rect 14427 4893 14441 4945
rect 14493 4893 14495 4945
rect 14241 4880 14495 4893
rect 14241 4828 14243 4880
rect 14295 4828 14309 4880
rect 14361 4828 14375 4880
rect 14427 4828 14441 4880
rect 14493 4828 14495 4880
rect 14241 4815 14495 4828
rect 14241 4763 14243 4815
rect 14295 4763 14309 4815
rect 14361 4763 14375 4815
rect 14427 4763 14441 4815
rect 14493 4763 14495 4815
rect 14241 4750 14495 4763
rect 14241 4698 14243 4750
rect 14295 4698 14309 4750
rect 14361 4698 14375 4750
rect 14427 4698 14441 4750
rect 14493 4698 14495 4750
rect 14241 4685 14495 4698
rect 14241 4633 14243 4685
rect 14295 4633 14309 4685
rect 14361 4633 14375 4685
rect 14427 4633 14441 4685
rect 14493 4633 14495 4685
rect 14241 4620 14495 4633
rect 14241 4568 14243 4620
rect 14295 4568 14309 4620
rect 14361 4568 14375 4620
rect 14427 4568 14441 4620
rect 14493 4568 14495 4620
rect 14241 4555 14495 4568
rect 14241 4503 14243 4555
rect 14295 4503 14309 4555
rect 14361 4503 14375 4555
rect 14427 4503 14441 4555
rect 14493 4503 14495 4555
rect 14241 4490 14495 4503
rect 14241 4438 14243 4490
rect 14295 4438 14309 4490
rect 14361 4438 14375 4490
rect 14427 4438 14441 4490
rect 14493 4438 14495 4490
rect 14241 4425 14495 4438
rect 14241 4373 14243 4425
rect 14295 4373 14309 4425
rect 14361 4373 14375 4425
rect 14427 4373 14441 4425
rect 14493 4373 14495 4425
rect 14241 4359 14495 4373
rect 14241 4307 14243 4359
rect 14295 4307 14309 4359
rect 14361 4307 14375 4359
rect 14427 4307 14441 4359
rect 14493 4307 14495 4359
rect 14241 4293 14495 4307
rect 14241 4241 14243 4293
rect 14295 4241 14309 4293
rect 14361 4241 14375 4293
rect 14427 4241 14441 4293
rect 14493 4241 14495 4293
rect 14241 4227 14495 4241
rect 14241 4175 14243 4227
rect 14295 4175 14309 4227
rect 14361 4175 14375 4227
rect 14427 4175 14441 4227
rect 14493 4175 14495 4227
rect 14241 4161 14495 4175
rect 14241 4109 14243 4161
rect 14295 4109 14309 4161
rect 14361 4109 14375 4161
rect 14427 4109 14441 4161
rect 14493 4109 14495 4161
rect 14241 4095 14495 4109
rect 14241 4043 14243 4095
rect 14295 4043 14309 4095
rect 14361 4043 14375 4095
rect 14427 4043 14441 4095
rect 14493 4043 14495 4095
rect 14241 4029 14495 4043
rect 14241 3977 14243 4029
rect 14295 3977 14309 4029
rect 14361 3977 14375 4029
rect 14427 3977 14441 4029
rect 14493 3977 14495 4029
rect 14241 3963 14495 3977
rect 14241 3911 14243 3963
rect 14295 3911 14309 3963
rect 14361 3911 14375 3963
rect 14427 3911 14441 3963
rect 14493 3911 14495 3963
rect 14241 3897 14495 3911
rect 14241 3845 14243 3897
rect 14295 3845 14309 3897
rect 14361 3845 14375 3897
rect 14427 3845 14441 3897
rect 14493 3845 14495 3897
rect 14241 3831 14495 3845
rect 14241 3779 14243 3831
rect 14295 3779 14309 3831
rect 14361 3779 14375 3831
rect 14427 3779 14441 3831
rect 14493 3779 14495 3831
rect 14241 3765 14495 3779
rect 14241 3713 14243 3765
rect 14295 3713 14309 3765
rect 14361 3713 14375 3765
rect 14427 3713 14441 3765
rect 14493 3713 14495 3765
rect 14241 3699 14495 3713
rect 14241 3647 14243 3699
rect 14295 3647 14309 3699
rect 14361 3647 14375 3699
rect 14427 3647 14441 3699
rect 14493 3647 14495 3699
rect 14241 3641 14495 3647
rect 14974 5457 15114 5495
rect 14974 5423 15068 5457
rect 15102 5423 15114 5457
rect 14974 5385 15114 5423
rect 14974 5351 15068 5385
rect 15102 5351 15114 5385
rect 14974 5313 15114 5351
rect 14974 5279 15068 5313
rect 15102 5279 15114 5313
rect 14974 5241 15114 5279
rect 14974 5207 15068 5241
rect 15102 5207 15114 5241
rect 14974 5169 15114 5207
rect 14974 5135 15068 5169
rect 15102 5135 15114 5169
rect 14974 5097 15114 5135
rect 14974 5063 15068 5097
rect 15102 5063 15114 5097
rect 14974 5025 15114 5063
rect 14974 4991 15068 5025
rect 15102 4991 15114 5025
rect 14974 4953 15114 4991
rect 14974 4919 15068 4953
rect 15102 4919 15114 4953
rect 14974 4881 15114 4919
rect 14974 4847 15068 4881
rect 15102 4847 15114 4881
rect 14974 4809 15114 4847
rect 14974 4775 15068 4809
rect 15102 4775 15114 4809
rect 14974 4737 15114 4775
rect 14974 4703 15068 4737
rect 15102 4703 15114 4737
rect 14974 4665 15114 4703
rect 14974 4631 15068 4665
rect 15102 4631 15114 4665
rect 14974 4593 15114 4631
rect 14974 4559 15068 4593
rect 15102 4559 15114 4593
rect 14974 4521 15114 4559
rect 14974 4487 15068 4521
rect 15102 4487 15114 4521
rect 14974 4449 15114 4487
rect 14974 4415 15068 4449
rect 15102 4415 15114 4449
rect 14974 4377 15114 4415
rect 14974 4343 15068 4377
rect 15102 4343 15114 4377
rect 14974 4305 15114 4343
rect 14974 4271 15068 4305
rect 15102 4271 15114 4305
rect 14974 4233 15114 4271
rect 14974 4199 15068 4233
rect 15102 4199 15114 4233
rect 14974 4161 15114 4199
rect 14974 4127 15068 4161
rect 15102 4127 15114 4161
rect 14974 4089 15114 4127
rect 14974 4055 15068 4089
rect 15102 4055 15114 4089
rect 14974 4017 15114 4055
rect 14974 3983 15068 4017
rect 15102 3983 15114 4017
rect 14974 3945 15114 3983
rect 14974 3911 15068 3945
rect 15102 3911 15114 3945
rect 14974 3873 15114 3911
rect 14974 3839 15068 3873
rect 15102 3839 15114 3873
rect 14974 3801 15114 3839
rect 14974 3767 15068 3801
rect 15102 3767 15114 3801
rect 14974 3729 15114 3767
rect 14974 3695 15068 3729
rect 15102 3695 15114 3729
rect 14974 3657 15114 3695
rect 14974 3623 15068 3657
rect 15102 3623 15114 3657
rect 14974 3585 15114 3623
rect 14974 3551 15068 3585
rect 15102 3551 15114 3585
rect 14974 3513 15114 3551
rect 14974 3479 15068 3513
rect 15102 3479 15114 3513
rect 14974 3441 15114 3479
rect 14974 3407 15068 3441
rect 15102 3407 15114 3441
rect 14974 3369 15114 3407
rect 14974 3335 15068 3369
rect 15102 3335 15114 3369
rect 14974 3297 15114 3335
rect 14974 3263 15068 3297
rect 15102 3263 15114 3297
rect 14974 3225 15114 3263
rect 14974 3191 15068 3225
rect 15102 3191 15114 3225
rect 14974 3153 15114 3191
rect 14974 3119 15068 3153
rect 15102 3119 15114 3153
rect 14974 3081 15114 3119
rect 14974 3047 15068 3081
rect 15102 3047 15114 3081
rect 14974 3009 15114 3047
rect 14974 2975 15068 3009
rect 15102 2975 15114 3009
rect 14974 2937 15114 2975
rect 14974 2903 15068 2937
rect 15102 2903 15114 2937
rect 14974 2865 15114 2903
rect 14974 2831 15068 2865
rect 15102 2831 15114 2865
rect 14974 2793 15114 2831
rect 14974 2759 15068 2793
rect 15102 2759 15114 2793
rect 14974 2721 15114 2759
rect 14974 2687 15068 2721
rect 15102 2687 15114 2721
rect 14974 2649 15114 2687
rect 14974 2615 15068 2649
rect 15102 2615 15114 2649
rect 14974 2577 15114 2615
rect 14974 2543 15068 2577
rect 15102 2543 15114 2577
rect 14974 2505 15114 2543
rect 14974 2471 15068 2505
rect 15102 2471 15114 2505
rect 14974 2433 15114 2471
rect 14974 2399 15068 2433
rect 15102 2399 15114 2433
rect 14974 2361 15114 2399
rect 14974 2327 15068 2361
rect 15102 2327 15114 2361
rect 14974 2289 15114 2327
rect 14974 2255 15068 2289
rect 15102 2255 15114 2289
rect 14974 2217 15114 2255
rect 14974 2183 15068 2217
rect 15102 2183 15114 2217
rect 14974 2145 15114 2183
rect 14974 2111 15068 2145
rect 15102 2111 15114 2145
rect 14974 2073 15114 2111
rect 14974 2039 15068 2073
rect 15102 2039 15114 2073
rect 14974 2001 15114 2039
rect 14974 1967 15068 2001
rect 15102 1967 15114 2001
rect 14974 1929 15114 1967
rect 14974 1895 15068 1929
rect 15102 1895 15114 1929
rect 14974 1857 15114 1895
rect 14974 1823 15068 1857
rect 15102 1823 15114 1857
rect 14974 1785 15114 1823
rect 14974 1751 15068 1785
rect 15102 1751 15114 1785
rect 14974 1713 15114 1751
rect 14974 1679 15068 1713
rect 15102 1679 15114 1713
rect 14974 1641 15114 1679
rect 14974 1607 15068 1641
rect 15102 1607 15114 1641
rect 14974 1569 15114 1607
rect 14974 1535 15068 1569
rect 15102 1535 15114 1569
rect 14974 1497 15114 1535
rect 14974 1463 15068 1497
rect 15102 1463 15114 1497
rect 14974 1425 15114 1463
rect 14974 1391 15068 1425
rect 15102 1391 15114 1425
rect 14974 1353 15114 1391
rect 14974 1319 15068 1353
rect 15102 1319 15114 1353
rect 14974 1300 15114 1319
rect 7031 1282 15114 1300
rect 3545 1281 15114 1282
rect 3545 1251 15068 1281
rect 3545 1217 3565 1251
rect 3599 1217 3637 1251
rect 3671 1217 3709 1251
rect 3743 1217 3781 1251
rect 3815 1217 3853 1251
rect 3887 1217 3925 1251
rect 3959 1217 3997 1251
rect 4031 1217 4069 1251
rect 4103 1217 4141 1251
rect 4175 1217 4213 1251
rect 4247 1217 4285 1251
rect 4319 1217 4357 1251
rect 4391 1217 4429 1251
rect 4463 1217 4501 1251
rect 4535 1217 4573 1251
rect 4607 1217 4645 1251
rect 4679 1217 4717 1251
rect 4751 1217 4789 1251
rect 4823 1217 4861 1251
rect 4895 1217 4933 1251
rect 4967 1217 5005 1251
rect 5039 1217 5077 1251
rect 5111 1217 5149 1251
rect 5183 1217 5221 1251
rect 5255 1217 5293 1251
rect 5327 1217 5365 1251
rect 5399 1217 5437 1251
rect 5471 1217 5509 1251
rect 5543 1217 5581 1251
rect 5615 1217 5653 1251
rect 5687 1217 5725 1251
rect 5759 1217 5797 1251
rect 5831 1217 5869 1251
rect 5903 1217 5941 1251
rect 5975 1217 6013 1251
rect 6047 1217 6085 1251
rect 6119 1217 6157 1251
rect 6191 1217 6229 1251
rect 6263 1217 6301 1251
rect 6335 1217 6373 1251
rect 6407 1217 6445 1251
rect 6479 1217 6517 1251
rect 6551 1217 6589 1251
rect 6623 1217 6661 1251
rect 6695 1217 6733 1251
rect 6767 1217 6805 1251
rect 6839 1217 6877 1251
rect 6911 1247 15068 1251
rect 15102 1247 15114 1281
rect 6911 1239 15114 1247
rect 6911 1217 6988 1239
rect 3545 1205 6988 1217
rect 7022 1217 15114 1239
rect 7022 1205 7069 1217
tri 6828 1183 6850 1205 ne
rect 6850 1183 7069 1205
rect 7103 1183 7142 1217
rect 7176 1183 7215 1217
rect 7249 1183 7288 1217
rect 7322 1183 7361 1217
rect 7395 1183 7434 1217
rect 7468 1183 7507 1217
rect 7541 1183 7580 1217
rect 7614 1183 7653 1217
rect 7687 1183 7726 1217
rect 7760 1183 7799 1217
rect 7833 1183 7872 1217
rect 7906 1183 7945 1217
rect 7979 1183 8018 1217
rect 8052 1183 8091 1217
rect 8125 1183 8164 1217
rect 8198 1183 8237 1217
rect 8271 1183 8310 1217
rect 8344 1183 8383 1217
rect 8417 1183 8456 1217
rect 8490 1183 8528 1217
rect 8562 1183 8600 1217
rect 8634 1183 8672 1217
rect 8706 1183 8744 1217
rect 8778 1183 8816 1217
rect 8850 1183 8888 1217
rect 8922 1183 8960 1217
rect 8994 1183 9032 1217
rect 9066 1183 9104 1217
rect 9138 1183 9176 1217
rect 9210 1183 9248 1217
rect 9282 1183 9320 1217
rect 9354 1183 9392 1217
rect 9426 1183 9464 1217
rect 9498 1183 9536 1217
rect 9570 1183 9608 1217
rect 9642 1183 9680 1217
rect 9714 1183 9752 1217
rect 9786 1183 9824 1217
rect 9858 1183 9896 1217
rect 9930 1183 9968 1217
rect 10002 1183 10040 1217
rect 10074 1183 10112 1217
rect 10146 1183 10184 1217
rect 10218 1183 10256 1217
rect 10290 1183 10328 1217
rect 10362 1183 10400 1217
rect 10434 1183 10472 1217
rect 10506 1183 10544 1217
rect 10578 1183 10616 1217
rect 10650 1183 10688 1217
rect 10722 1183 10760 1217
rect 10794 1183 10832 1217
rect 10866 1183 10904 1217
rect 10938 1183 10976 1217
rect 11010 1183 11048 1217
rect 11082 1183 11120 1217
rect 11154 1183 11192 1217
rect 11226 1183 11264 1217
rect 11298 1183 11336 1217
rect 11370 1183 11408 1217
rect 11442 1183 11480 1217
rect 11514 1183 11552 1217
rect 11586 1183 11624 1217
rect 11658 1183 11696 1217
rect 11730 1183 11768 1217
rect 11802 1183 11840 1217
rect 11874 1183 11912 1217
rect 11946 1183 11984 1217
rect 12018 1183 12056 1217
rect 12090 1183 12139 1217
rect 12173 1183 12212 1217
rect 12246 1183 12285 1217
rect 12319 1183 12358 1217
rect 12392 1183 12431 1217
rect 12465 1183 12504 1217
rect 12538 1183 12577 1217
rect 12611 1183 12650 1217
rect 12684 1183 12723 1217
rect 12757 1183 12796 1217
rect 12830 1183 12869 1217
rect 12903 1183 12942 1217
rect 12976 1183 13015 1217
rect 13049 1183 13088 1217
rect 13122 1183 13161 1217
rect 13195 1183 13234 1217
rect 13268 1183 13307 1217
rect 13341 1183 13380 1217
rect 13414 1183 13452 1217
rect 13486 1183 13524 1217
rect 13558 1183 13596 1217
rect 13630 1183 13668 1217
rect 13702 1183 13740 1217
rect 13774 1183 13812 1217
rect 13846 1183 13884 1217
rect 13918 1183 13956 1217
rect 13990 1183 14028 1217
rect 14062 1183 14100 1217
rect 14134 1183 14172 1217
rect 14206 1183 14244 1217
rect 14278 1183 14316 1217
rect 14350 1183 14388 1217
rect 14422 1183 14460 1217
rect 14494 1183 14532 1217
rect 14566 1183 14604 1217
rect 14638 1183 14676 1217
rect 14710 1183 14748 1217
rect 14782 1183 14820 1217
rect 14854 1183 14892 1217
rect 14926 1183 14964 1217
rect 14998 1209 15114 1217
rect 14998 1183 15068 1209
tri 6850 1175 6858 1183 ne
rect 6858 1175 15068 1183
rect 15102 1175 15114 1209
tri 6858 1167 6866 1175 ne
rect 6866 1167 15114 1175
tri 6866 1133 6900 1167 ne
rect 6900 1133 6988 1167
rect 7022 1139 15114 1167
rect 7022 1133 7069 1139
tri 6900 1105 6928 1133 ne
rect 6928 1105 7069 1133
rect 7103 1105 7142 1139
rect 7176 1105 7215 1139
rect 7249 1105 7288 1139
rect 7322 1105 7361 1139
rect 7395 1105 7434 1139
rect 7468 1105 7507 1139
rect 7541 1105 7580 1139
rect 7614 1105 7653 1139
rect 7687 1105 7726 1139
rect 7760 1105 7799 1139
rect 7833 1105 7872 1139
rect 7906 1105 7945 1139
rect 7979 1105 8018 1139
rect 8052 1105 8091 1139
rect 8125 1105 8164 1139
rect 8198 1105 8237 1139
rect 8271 1105 8310 1139
rect 8344 1105 8383 1139
rect 8417 1105 8456 1139
rect 8490 1105 8528 1139
rect 8562 1105 8600 1139
rect 8634 1105 8672 1139
rect 8706 1105 8744 1139
rect 8778 1105 8816 1139
rect 8850 1105 8888 1139
rect 8922 1105 8960 1139
rect 8994 1105 9032 1139
rect 9066 1105 9104 1139
rect 9138 1105 9176 1139
rect 9210 1105 9248 1139
rect 9282 1105 9320 1139
rect 9354 1105 9392 1139
rect 9426 1105 9464 1139
rect 9498 1105 9536 1139
rect 9570 1105 9608 1139
rect 9642 1105 9680 1139
rect 9714 1105 9752 1139
rect 9786 1105 9824 1139
rect 9858 1105 9896 1139
rect 9930 1105 9968 1139
rect 10002 1105 10040 1139
rect 10074 1105 10112 1139
rect 10146 1105 10184 1139
rect 10218 1105 10256 1139
rect 10290 1105 10328 1139
rect 10362 1105 10400 1139
rect 10434 1105 10472 1139
rect 10506 1105 10544 1139
rect 10578 1105 10616 1139
rect 10650 1105 10688 1139
rect 10722 1105 10760 1139
rect 10794 1105 10832 1139
rect 10866 1105 10904 1139
rect 10938 1105 10976 1139
rect 11010 1105 11048 1139
rect 11082 1105 11120 1139
rect 11154 1105 11192 1139
rect 11226 1105 11264 1139
rect 11298 1105 11336 1139
rect 11370 1105 11408 1139
rect 11442 1105 11480 1139
rect 11514 1105 11552 1139
rect 11586 1105 11624 1139
rect 11658 1105 11696 1139
rect 11730 1105 11768 1139
rect 11802 1105 11840 1139
rect 11874 1105 11912 1139
rect 11946 1105 11984 1139
rect 12018 1105 12056 1139
rect 12090 1105 12139 1139
rect 12173 1105 12212 1139
rect 12246 1105 12285 1139
rect 12319 1105 12358 1139
rect 12392 1105 12431 1139
rect 12465 1105 12504 1139
rect 12538 1105 12577 1139
rect 12611 1105 12650 1139
rect 12684 1105 12723 1139
rect 12757 1105 12796 1139
rect 12830 1105 12869 1139
rect 12903 1105 12942 1139
rect 12976 1105 13015 1139
rect 13049 1105 13088 1139
rect 13122 1105 13161 1139
rect 13195 1105 13234 1139
rect 13268 1105 13307 1139
rect 13341 1105 13380 1139
rect 13414 1105 13452 1139
rect 13486 1105 13524 1139
rect 13558 1105 13596 1139
rect 13630 1105 13668 1139
rect 13702 1105 13740 1139
rect 13774 1105 13812 1139
rect 13846 1105 13884 1139
rect 13918 1105 13956 1139
rect 13990 1105 14028 1139
rect 14062 1105 14100 1139
rect 14134 1105 14172 1139
rect 14206 1105 14244 1139
rect 14278 1105 14316 1139
rect 14350 1105 14388 1139
rect 14422 1105 14460 1139
rect 14494 1105 14532 1139
rect 14566 1105 14604 1139
rect 14638 1105 14676 1139
rect 14710 1105 14748 1139
rect 14782 1105 14820 1139
rect 14854 1105 14892 1139
rect 14926 1105 14964 1139
rect 14998 1137 15114 1139
rect 14998 1105 15068 1137
tri 6928 1103 6930 1105 ne
rect 6930 1103 15068 1105
rect 15102 1103 15114 1137
tri 6930 1095 6938 1103 ne
rect 6938 1095 15114 1103
tri 6938 1077 6956 1095 ne
rect 6956 1077 6988 1095
rect 451 932 1620 1077
tri 6956 1061 6972 1077 ne
rect 6972 1061 6988 1077
rect 7022 1065 15114 1095
rect 7022 1061 15068 1065
tri 6972 1057 6976 1061 ne
rect 6976 1027 7069 1061
rect 7103 1027 7142 1061
rect 7176 1027 7215 1061
rect 7249 1027 7288 1061
rect 7322 1027 7361 1061
rect 7395 1027 7434 1061
rect 7468 1027 7507 1061
rect 7541 1027 7580 1061
rect 7614 1027 7653 1061
rect 7687 1027 7726 1061
rect 7760 1027 7799 1061
rect 7833 1027 7872 1061
rect 7906 1027 7945 1061
rect 7979 1027 8018 1061
rect 8052 1027 8091 1061
rect 8125 1027 8164 1061
rect 8198 1027 8237 1061
rect 8271 1027 8310 1061
rect 8344 1027 8383 1061
rect 8417 1027 8456 1061
rect 8490 1027 8528 1061
rect 8562 1027 8600 1061
rect 8634 1027 8672 1061
rect 8706 1027 8744 1061
rect 8778 1027 8816 1061
rect 8850 1027 8888 1061
rect 8922 1027 8960 1061
rect 8994 1027 9032 1061
rect 9066 1027 9104 1061
rect 9138 1027 9176 1061
rect 9210 1027 9248 1061
rect 9282 1027 9320 1061
rect 9354 1027 9392 1061
rect 9426 1027 9464 1061
rect 9498 1027 9536 1061
rect 9570 1027 9608 1061
rect 9642 1027 9680 1061
rect 9714 1027 9752 1061
rect 9786 1027 9824 1061
rect 9858 1027 9896 1061
rect 9930 1027 9968 1061
rect 10002 1027 10040 1061
rect 10074 1027 10112 1061
rect 10146 1027 10184 1061
rect 10218 1027 10256 1061
rect 10290 1027 10328 1061
rect 10362 1027 10400 1061
rect 10434 1027 10472 1061
rect 10506 1027 10544 1061
rect 10578 1027 10616 1061
rect 10650 1027 10688 1061
rect 10722 1027 10760 1061
rect 10794 1027 10832 1061
rect 10866 1027 10904 1061
rect 10938 1027 10976 1061
rect 11010 1027 11048 1061
rect 11082 1027 11120 1061
rect 11154 1027 11192 1061
rect 11226 1027 11264 1061
rect 11298 1027 11336 1061
rect 11370 1027 11408 1061
rect 11442 1027 11480 1061
rect 11514 1027 11552 1061
rect 11586 1027 11624 1061
rect 11658 1027 11696 1061
rect 11730 1027 11768 1061
rect 11802 1027 11840 1061
rect 11874 1027 11912 1061
rect 11946 1027 11984 1061
rect 12018 1027 12056 1061
rect 12090 1027 12139 1061
rect 12173 1027 12212 1061
rect 12246 1027 12285 1061
rect 12319 1027 12358 1061
rect 12392 1027 12431 1061
rect 12465 1027 12504 1061
rect 12538 1027 12577 1061
rect 12611 1027 12650 1061
rect 12684 1027 12723 1061
rect 12757 1027 12796 1061
rect 12830 1027 12869 1061
rect 12903 1027 12942 1061
rect 12976 1027 13015 1061
rect 13049 1027 13088 1061
rect 13122 1027 13161 1061
rect 13195 1027 13234 1061
rect 13268 1027 13307 1061
rect 13341 1027 13380 1061
rect 13414 1027 13452 1061
rect 13486 1027 13524 1061
rect 13558 1027 13596 1061
rect 13630 1027 13668 1061
rect 13702 1027 13740 1061
rect 13774 1027 13812 1061
rect 13846 1027 13884 1061
rect 13918 1027 13956 1061
rect 13990 1027 14028 1061
rect 14062 1027 14100 1061
rect 14134 1027 14172 1061
rect 14206 1027 14244 1061
rect 14278 1027 14316 1061
rect 14350 1027 14388 1061
rect 14422 1027 14460 1061
rect 14494 1027 14532 1061
rect 14566 1027 14604 1061
rect 14638 1027 14676 1061
rect 14710 1027 14748 1061
rect 14782 1027 14820 1061
rect 14854 1027 14892 1061
rect 14926 1027 14964 1061
rect 14998 1031 15068 1061
rect 15102 1031 15114 1065
rect 14998 1027 15114 1031
rect 6976 1023 15114 1027
rect 6976 989 6988 1023
rect 7022 1020 15114 1023
rect 7022 993 7295 1020
tri 7295 993 7322 1020 nw
tri 14305 993 14332 1020 ne
rect 14332 993 15114 1020
rect 7022 989 7291 993
tri 7291 989 7295 993 nw
tri 14332 989 14336 993 ne
rect 14336 989 15068 993
rect 6976 966 7268 989
tri 7268 966 7291 989 nw
tri 14336 966 14359 989 ne
rect 14359 966 14576 989
rect 6976 955 7257 966
tri 7257 955 7268 966 nw
tri 14359 955 14370 966 ne
rect 14370 955 14576 966
rect 14610 955 14654 989
rect 14688 955 14732 989
rect 14766 955 14810 989
rect 14844 955 14888 989
rect 14922 955 14966 989
rect 15000 959 15068 989
rect 15102 959 15114 993
rect 15000 955 15114 959
rect 3522 944 3568 955
rect 3574 949 6836 955
rect 3574 944 3722 949
rect 3516 943 3722 944
rect 3516 909 3528 943
rect 3562 915 3722 943
rect 3756 915 3794 949
rect 3828 915 3866 949
rect 3900 915 3938 949
rect 3972 915 4010 949
rect 4044 915 4082 949
rect 4116 915 4154 949
rect 4188 915 4226 949
rect 4260 915 4298 949
rect 4332 915 4370 949
rect 4404 915 4442 949
rect 4476 915 4514 949
rect 4548 915 4586 949
rect 4620 915 4658 949
rect 4692 915 4730 949
rect 4764 915 4802 949
rect 4836 915 4874 949
rect 4908 915 4946 949
rect 4980 915 5018 949
rect 5052 915 5090 949
rect 5124 915 5252 949
rect 5286 915 5324 949
rect 5358 915 5396 949
rect 5430 915 5468 949
rect 5502 915 5540 949
rect 5574 915 5612 949
rect 5646 915 5684 949
rect 5718 915 5756 949
rect 5790 915 5828 949
rect 5862 915 5900 949
rect 5934 915 5972 949
rect 6006 915 6044 949
rect 6078 915 6116 949
rect 6150 915 6188 949
rect 6222 915 6260 949
rect 6294 915 6332 949
rect 6366 915 6404 949
rect 6438 915 6476 949
rect 6510 915 6548 949
rect 6582 915 6620 949
rect 6654 915 6836 949
rect 3562 909 6836 915
rect 3516 884 3608 909
tri 3608 884 3633 909 nw
tri 6752 884 6777 909 ne
rect 6777 884 6836 909
rect 3516 883 3607 884
tri 3607 883 3608 884 nw
tri 6777 883 6778 884 ne
rect 3516 882 3606 883
tri 3606 882 3607 883 nw
rect 3516 879 3603 882
tri 3603 879 3606 882 nw
rect 3516 872 3596 879
tri 3596 872 3603 879 nw
rect 574 820 580 872
rect 632 820 648 872
rect 700 820 706 872
rect 574 806 706 820
rect 574 754 580 806
rect 632 754 648 806
rect 700 754 706 806
rect 3516 871 3593 872
rect 3516 837 3528 871
rect 3562 869 3593 871
tri 3593 869 3596 872 nw
rect 3710 871 6666 872
rect 3562 837 3574 869
tri 3574 850 3593 869 nw
rect 3516 799 3574 837
rect 3516 765 3528 799
rect 3562 765 3574 799
rect 3516 727 3574 765
rect 3710 819 3716 871
rect 3768 819 3796 871
rect 3848 819 3876 871
rect 3928 819 6666 871
rect 3710 805 6666 819
rect 3710 753 3716 805
rect 3768 793 3796 805
rect 3848 793 3876 805
rect 3928 793 6666 805
rect 3768 759 3794 793
rect 3848 759 3866 793
rect 3928 759 3938 793
rect 3972 759 4010 793
rect 4044 759 4082 793
rect 4116 759 4154 793
rect 4188 759 4226 793
rect 4260 759 4298 793
rect 4332 759 4370 793
rect 4404 759 4442 793
rect 4476 759 4514 793
rect 4548 759 4586 793
rect 4620 759 4658 793
rect 4692 759 4730 793
rect 4764 759 4802 793
rect 4836 759 4874 793
rect 4908 759 4946 793
rect 4980 759 5018 793
rect 5052 759 5090 793
rect 5124 759 5252 793
rect 5286 759 5324 793
rect 5358 759 5396 793
rect 5430 759 5468 793
rect 5502 759 5540 793
rect 5574 759 5612 793
rect 5646 759 5684 793
rect 5718 759 5756 793
rect 5790 759 5828 793
rect 5862 759 5900 793
rect 5934 759 5972 793
rect 6006 759 6044 793
rect 6078 759 6116 793
rect 6150 759 6188 793
rect 6222 759 6260 793
rect 6294 759 6332 793
rect 6366 759 6404 793
rect 6438 759 6476 793
rect 6510 759 6548 793
rect 6582 759 6620 793
rect 6654 759 6666 793
rect 3768 753 3796 759
rect 3848 753 3876 759
rect 3928 753 6666 759
rect 6778 869 6836 884
rect 6778 835 6790 869
rect 6824 835 6836 869
rect 6778 797 6836 835
rect 6778 763 6790 797
rect 6824 763 6836 797
rect 761 683 794 715
rect 3516 693 3528 727
rect 3562 693 3574 727
rect 6778 725 6836 763
rect 3516 680 3574 693
rect 3633 714 6738 720
tri 3574 680 3584 690 sw
rect 3633 680 3645 714
rect 3679 680 3717 714
rect 3751 680 5115 714
rect 5149 680 5187 714
rect 5221 680 6620 714
rect 6654 680 6692 714
rect 6726 680 6738 714
rect 3516 674 3584 680
tri 3584 674 3590 680 sw
rect 3633 674 6738 680
rect 6778 691 6790 725
rect 6824 691 6836 725
rect 3516 672 3590 674
tri 3590 672 3592 674 sw
rect 3516 671 3592 672
tri 3592 671 3593 672 sw
tri 6777 671 6778 672 se
rect 6778 671 6836 691
rect 3516 663 3593 671
tri 3593 663 3601 671 sw
tri 6769 663 6777 671 se
rect 6777 663 6836 671
rect 3516 655 3601 663
rect 3516 621 3528 655
rect 3562 653 3601 655
tri 3601 653 3611 663 sw
tri 6759 653 6769 663 se
rect 6769 653 6836 663
rect 3562 643 3611 653
tri 3611 643 3621 653 sw
tri 6749 643 6759 653 se
rect 6759 643 6790 653
rect 3562 637 6790 643
rect 3562 621 3722 637
rect 3516 603 3722 621
rect 3756 603 3794 637
rect 3828 603 3866 637
rect 3900 603 3938 637
rect 3972 603 4010 637
rect 4044 603 4082 637
rect 4116 603 4154 637
rect 4188 603 4226 637
rect 4260 603 4298 637
rect 4332 603 4370 637
rect 4404 603 4442 637
rect 4476 603 4514 637
rect 4548 603 4586 637
rect 4620 603 4658 637
rect 4692 603 4730 637
rect 4764 603 4802 637
rect 4836 603 4874 637
rect 4908 603 4946 637
rect 4980 603 5018 637
rect 5052 603 5090 637
rect 5124 603 5252 637
rect 5286 603 5324 637
rect 5358 603 5396 637
rect 5430 603 5468 637
rect 5502 603 5540 637
rect 5574 603 5612 637
rect 5646 603 5684 637
rect 5718 603 5756 637
rect 5790 603 5828 637
rect 5862 603 5900 637
rect 5934 603 5972 637
rect 6006 603 6044 637
rect 6078 603 6116 637
rect 6150 603 6188 637
rect 6222 603 6260 637
rect 6294 603 6332 637
rect 6366 603 6404 637
rect 6438 603 6476 637
rect 6510 603 6548 637
rect 6582 603 6620 637
rect 6654 619 6790 637
rect 6824 619 6836 653
rect 6654 603 6836 619
rect 3516 583 6836 603
rect 3516 549 3528 583
rect 3562 581 6836 583
rect 3562 549 6790 581
rect 3516 547 6790 549
rect 6824 547 6836 581
rect 3516 524 6836 547
rect 3516 519 3619 524
tri 3619 519 3624 524 nw
tri 6747 519 6752 524 ne
rect 6752 519 6836 524
rect 3516 511 3609 519
rect 574 435 580 487
rect 632 435 648 487
rect 700 435 706 487
rect 574 421 706 435
rect 574 369 580 421
rect 632 369 648 421
rect 700 369 706 421
rect 3516 477 3528 511
rect 3562 509 3609 511
tri 3609 509 3619 519 nw
tri 6752 509 6762 519 ne
rect 6762 509 6836 519
rect 3562 493 3593 509
tri 3593 493 3609 509 nw
tri 6762 493 6778 509 ne
rect 3562 487 3587 493
tri 3587 487 3593 493 nw
rect 3562 481 3581 487
tri 3581 481 3587 487 nw
rect 3562 477 3574 481
rect 3516 439 3574 477
tri 3574 474 3581 481 nw
rect 3516 405 3528 439
rect 3562 405 3574 439
rect 3516 390 3574 405
rect 3710 435 3716 487
rect 3768 481 3796 487
rect 3848 481 3876 487
rect 3928 481 6666 487
rect 3768 447 3794 481
rect 3848 447 3866 481
rect 3928 447 3938 481
rect 3972 447 4010 481
rect 4044 447 4082 481
rect 4116 447 4154 481
rect 4188 447 4226 481
rect 4260 447 4298 481
rect 4332 447 4370 481
rect 4404 447 4442 481
rect 4476 447 4514 481
rect 4548 447 4586 481
rect 4620 447 4658 481
rect 4692 447 4730 481
rect 4764 447 4802 481
rect 4836 447 4874 481
rect 4908 447 4946 481
rect 4980 447 5018 481
rect 5052 447 5090 481
rect 5124 447 5252 481
rect 5286 447 5324 481
rect 5358 447 5396 481
rect 5430 447 5468 481
rect 5502 447 5540 481
rect 5574 447 5612 481
rect 5646 447 5684 481
rect 5718 447 5756 481
rect 5790 447 5828 481
rect 5862 447 5900 481
rect 5934 447 5972 481
rect 6006 447 6044 481
rect 6078 447 6116 481
rect 6150 447 6188 481
rect 6222 447 6260 481
rect 6294 447 6332 481
rect 6366 447 6404 481
rect 6438 447 6476 481
rect 6510 447 6548 481
rect 6582 447 6620 481
rect 6654 447 6666 481
rect 3768 435 3796 447
rect 3848 435 3876 447
rect 3928 435 6666 447
rect 3710 421 6666 435
tri 3574 390 3576 392 sw
rect 3516 375 3576 390
tri 3576 375 3591 390 sw
rect 3516 369 3591 375
tri 3591 369 3597 375 sw
rect 3710 369 3716 421
rect 3768 369 3796 421
rect 3848 369 3876 421
rect 3928 369 6666 421
rect 3516 368 3597 369
tri 3597 368 3598 369 sw
rect 3710 368 6666 369
rect 6778 475 6790 509
rect 6824 475 6836 509
rect 6778 437 6836 475
rect 6778 403 6790 437
rect 6824 403 6836 437
rect 3516 367 3598 368
rect 3516 333 3528 367
rect 3562 365 3598 367
tri 3598 365 3601 368 sw
tri 6775 365 6778 368 se
rect 6778 365 6836 403
rect 3562 333 3601 365
rect 3516 331 3601 333
tri 3601 331 3635 365 sw
tri 6741 331 6775 365 se
rect 6775 331 6790 365
rect 6824 331 6836 365
rect 3516 325 6836 331
rect 3516 294 3722 325
rect 3516 260 3528 294
rect 3562 291 3722 294
rect 3756 291 3794 325
rect 3828 291 3866 325
rect 3900 291 3938 325
rect 3972 291 4010 325
rect 4044 291 4082 325
rect 4116 291 4154 325
rect 4188 291 4226 325
rect 4260 291 4298 325
rect 4332 291 4370 325
rect 4404 291 4442 325
rect 4476 291 4514 325
rect 4548 291 4586 325
rect 4620 291 4658 325
rect 4692 291 4730 325
rect 4764 291 4802 325
rect 4836 291 4874 325
rect 4908 291 4946 325
rect 4980 291 5018 325
rect 5052 291 5090 325
rect 5124 291 5252 325
rect 5286 291 5324 325
rect 5358 291 5396 325
rect 5430 291 5468 325
rect 5502 291 5540 325
rect 5574 291 5612 325
rect 5646 291 5684 325
rect 5718 291 5756 325
rect 5790 291 5828 325
rect 5862 291 5900 325
rect 5934 291 5972 325
rect 6006 291 6044 325
rect 6078 291 6116 325
rect 6150 291 6188 325
rect 6222 291 6260 325
rect 6294 291 6332 325
rect 6366 291 6404 325
rect 6438 291 6476 325
rect 6510 291 6548 325
rect 6582 291 6620 325
rect 6654 293 6836 325
rect 6654 291 6790 293
rect 3562 260 6790 291
rect 3516 259 6790 260
rect 6824 259 6836 293
rect 3516 237 6836 259
rect 3493 221 6836 237
rect 3493 187 3528 221
rect 3562 209 6790 221
rect 3562 187 3632 209
rect 3493 175 3632 187
rect 3666 175 3704 209
rect 3738 175 3776 209
rect 3810 175 3848 209
rect 3882 175 3920 209
rect 3954 175 3992 209
rect 4026 175 4064 209
rect 4098 175 4136 209
rect 4170 175 4208 209
rect 4242 175 4280 209
rect 4314 175 4352 209
rect 4386 175 4424 209
rect 4458 175 4496 209
rect 4530 175 4568 209
rect 4602 175 4640 209
rect 4674 175 4712 209
rect 4746 175 4784 209
rect 4818 175 4856 209
rect 4890 175 4928 209
rect 4962 175 5000 209
rect 5034 175 5072 209
rect 5106 175 5144 209
rect 5178 175 5216 209
rect 5250 175 5288 209
rect 5322 175 5360 209
rect 5394 175 5432 209
rect 5466 175 5504 209
rect 5538 175 5576 209
rect 5610 175 5648 209
rect 5682 175 5720 209
rect 5754 175 5792 209
rect 5826 175 5864 209
rect 5898 175 5936 209
rect 5970 175 6008 209
rect 6042 175 6080 209
rect 6114 175 6152 209
rect 6186 175 6224 209
rect 6258 175 6296 209
rect 6330 175 6368 209
rect 6402 175 6440 209
rect 6474 175 6512 209
rect 6546 175 6584 209
rect 6618 175 6656 209
rect 6690 187 6790 209
rect 6824 187 6836 221
rect 6690 175 6836 187
rect 3493 163 6836 175
rect 6976 951 7232 955
rect 6976 917 6988 951
rect 7022 930 7232 951
tri 7232 930 7257 955 nw
tri 14370 930 14395 955 ne
rect 14395 930 15114 955
rect 7022 923 7225 930
tri 7225 923 7232 930 nw
rect 9784 923 11347 930
rect 7022 918 7191 923
rect 7022 917 7104 918
rect 6976 884 7104 917
rect 7138 889 7191 918
tri 7191 889 7225 923 nw
rect 9784 889 9796 923
rect 9830 889 9872 923
rect 9906 889 9948 923
rect 9982 889 10024 923
rect 10058 889 10100 923
rect 10134 889 10176 923
rect 10210 889 10251 923
rect 10285 889 10326 923
rect 10360 889 10401 923
rect 10435 889 10476 923
rect 10510 889 10551 923
rect 10585 889 10626 923
rect 10660 889 10701 923
rect 10735 889 10776 923
rect 10810 889 10851 923
rect 10885 889 10926 923
rect 10960 889 11001 923
rect 11035 889 11076 923
rect 11110 889 11151 923
rect 11185 889 11226 923
rect 11260 889 11301 923
rect 11335 889 11347 923
tri 14395 921 14404 930 ne
rect 14404 921 15114 930
tri 14404 916 14409 921 ne
rect 14409 916 15068 921
rect 7138 884 7184 889
rect 6976 882 7184 884
tri 7184 882 7191 889 nw
rect 6976 879 7174 882
rect 6976 845 6988 879
rect 7022 872 7174 879
tri 7174 872 7184 882 nw
rect 7022 871 7173 872
tri 7173 871 7174 872 nw
rect 7022 849 7151 871
tri 7151 849 7173 871 nw
rect 7022 845 7145 849
rect 6976 843 7145 845
tri 7145 843 7151 849 nw
rect 6976 839 7141 843
tri 7141 839 7145 843 nw
rect 9784 839 11347 889
tri 14409 882 14443 916 ne
rect 14443 882 14576 916
rect 14610 882 14654 916
rect 14688 882 14732 916
rect 14766 882 14810 916
rect 14844 882 14888 916
rect 14922 882 14966 916
rect 15000 887 15068 916
rect 15102 887 15114 921
rect 15000 882 15114 887
tri 14443 872 14453 882 ne
rect 14453 872 15114 882
tri 14453 871 14454 872 ne
rect 14454 871 15114 872
tri 14454 849 14476 871 ne
rect 14476 849 15114 871
tri 14476 843 14482 849 ne
rect 14482 843 15068 849
rect 6976 807 7107 839
rect 6976 773 6988 807
rect 7022 805 7107 807
tri 7107 805 7141 839 nw
rect 9784 805 9796 839
rect 9830 805 9872 839
rect 9906 805 9948 839
rect 9982 805 10024 839
rect 10058 805 10100 839
rect 10134 805 10176 839
rect 10210 805 10251 839
rect 10285 805 10326 839
rect 10360 805 10401 839
rect 10435 805 10476 839
rect 10510 805 10551 839
rect 10585 805 10626 839
rect 10660 805 10701 839
rect 10735 805 10776 839
rect 10810 805 10851 839
rect 10885 805 10926 839
rect 10960 805 11001 839
rect 11035 805 11076 839
rect 11110 805 11151 839
rect 11185 805 11226 839
rect 11260 805 11301 839
rect 11335 805 11347 839
tri 14482 809 14516 843 ne
rect 14516 809 14576 843
rect 14610 809 14654 843
rect 14688 809 14732 843
rect 14766 809 14810 843
rect 14844 809 14888 843
rect 14922 809 14966 843
rect 15000 815 15068 843
rect 15102 815 15114 849
rect 15000 809 15114 815
rect 7022 777 7079 805
tri 7079 777 7107 805 nw
rect 7022 773 7072 777
rect 6976 770 7072 773
tri 7072 770 7079 777 nw
rect 6976 755 7057 770
tri 7057 755 7072 770 nw
rect 9784 755 11347 805
tri 14516 794 14531 809 ne
rect 14531 794 15114 809
rect 6976 753 7055 755
tri 7055 753 7057 755 nw
rect 6976 735 7034 753
rect 6976 701 6988 735
rect 7022 701 7034 735
tri 7034 732 7055 753 nw
rect 6976 663 7034 701
rect 6976 629 6988 663
rect 7022 629 7034 663
rect 6976 591 7034 629
rect 6976 557 6988 591
rect 7022 557 7034 591
rect 6976 519 7034 557
rect 6976 485 6988 519
rect 7022 485 7034 519
rect 6976 447 7034 485
rect 9784 721 9796 755
rect 9830 721 9872 755
rect 9906 721 9948 755
rect 9982 721 10024 755
rect 10058 721 10100 755
rect 10134 721 10176 755
rect 10210 721 10251 755
rect 10285 721 10326 755
rect 10360 721 10401 755
rect 10435 721 10476 755
rect 10510 721 10551 755
rect 10585 721 10626 755
rect 10660 721 10701 755
rect 10735 721 10776 755
rect 10810 721 10851 755
rect 10885 721 10926 755
rect 10960 721 11001 755
rect 11035 721 11076 755
rect 11110 721 11151 755
rect 11185 721 11226 755
rect 11260 721 11301 755
rect 11335 721 11347 755
rect 11799 736 11831 794
tri 14531 777 14548 794 ne
rect 14548 777 15114 794
tri 14548 770 14555 777 ne
rect 14555 770 15068 777
tri 14555 759 14566 770 ne
rect 14566 736 14576 770
rect 14610 736 14654 770
rect 14688 736 14732 770
rect 14766 736 14810 770
rect 14844 736 14888 770
rect 14922 736 14966 770
rect 15000 743 15068 770
rect 15102 743 15114 777
rect 15000 736 15114 743
rect 9784 671 11347 721
rect 9784 637 9796 671
rect 9830 637 9872 671
rect 9906 637 9948 671
rect 9982 637 10024 671
rect 10058 637 10100 671
rect 10134 637 10176 671
rect 10210 637 10251 671
rect 10285 637 10326 671
rect 10360 637 10401 671
rect 10435 637 10476 671
rect 10510 637 10551 671
rect 10585 637 10626 671
rect 10660 637 10701 671
rect 10735 637 10776 671
rect 10810 637 10851 671
rect 10885 637 10926 671
rect 10960 637 11001 671
rect 11035 637 11076 671
rect 11110 637 11151 671
rect 11185 637 11226 671
rect 11260 637 11301 671
rect 11335 637 11347 671
rect 9784 587 11347 637
rect 9784 553 9796 587
rect 9830 553 9872 587
rect 9906 553 9948 587
rect 9982 553 10024 587
rect 10058 553 10100 587
rect 10134 553 10176 587
rect 10210 553 10251 587
rect 10285 553 10326 587
rect 10360 553 10401 587
rect 10435 553 10476 587
rect 10510 553 10551 587
rect 10585 553 10626 587
rect 10660 553 10701 587
rect 10735 553 10776 587
rect 10810 553 10851 587
rect 10885 553 10926 587
rect 10960 553 11001 587
rect 11035 553 11076 587
rect 11110 553 11151 587
rect 11185 553 11226 587
rect 11260 553 11301 587
rect 11335 553 11347 587
rect 9784 503 11347 553
rect 9784 469 9796 503
rect 9830 469 9872 503
rect 9906 469 9948 503
rect 9982 469 10024 503
rect 10058 469 10100 503
rect 10134 469 10176 503
rect 10210 469 10251 503
rect 10285 469 10326 503
rect 10360 469 10401 503
rect 10435 469 10476 503
rect 10510 469 10551 503
rect 10585 469 10626 503
rect 10660 469 10701 503
rect 10735 469 10776 503
rect 10810 469 10851 503
rect 10885 469 10926 503
rect 10960 469 11001 503
rect 11035 469 11076 503
rect 11110 469 11151 503
rect 11185 469 11226 503
rect 11260 469 11301 503
rect 11335 469 11347 503
rect 9784 462 11347 469
rect 14566 705 15114 736
rect 14566 697 15068 705
rect 14566 663 14576 697
rect 14610 663 14654 697
rect 14688 663 14732 697
rect 14766 663 14810 697
rect 14844 663 14888 697
rect 14922 663 14966 697
rect 15000 671 15068 697
rect 15102 671 15114 705
rect 15000 663 15114 671
rect 14566 633 15114 663
rect 14566 623 15068 633
rect 14566 589 14576 623
rect 14610 589 14654 623
rect 14688 589 14732 623
rect 14766 589 14810 623
rect 14844 589 14888 623
rect 14922 589 14966 623
rect 15000 599 15068 623
rect 15102 599 15114 633
rect 15000 589 15114 599
rect 14566 561 15114 589
rect 14566 549 15068 561
rect 14566 515 14576 549
rect 14610 515 14654 549
rect 14688 515 14732 549
rect 14766 515 14810 549
rect 14844 515 14888 549
rect 14922 515 14966 549
rect 15000 527 15068 549
rect 15102 527 15114 561
rect 15000 515 15114 527
rect 14566 489 15114 515
rect 14566 475 15068 489
rect 6976 413 6988 447
rect 7022 413 7034 447
rect 14566 441 14576 475
rect 14610 441 14654 475
rect 14688 441 14732 475
rect 14766 441 14810 475
rect 14844 441 14888 475
rect 14922 441 14966 475
rect 15000 455 15068 475
rect 15102 455 15114 489
rect 15000 441 15114 455
rect 14566 429 15114 441
tri 14566 417 14578 429 ne
rect 14578 417 15114 429
rect 6976 375 7034 413
tri 14578 402 14593 417 ne
rect 14593 402 15068 417
tri 14593 390 14605 402 ne
rect 14605 390 15068 402
rect 6976 341 6988 375
rect 7022 341 7034 375
tri 14605 369 14626 390 ne
rect 14626 369 14657 390
tri 14626 356 14639 369 ne
rect 14639 356 14657 369
rect 14691 356 14735 390
rect 14769 356 14813 390
rect 14847 356 14891 390
rect 14925 356 14969 390
rect 15003 383 15068 390
rect 15102 383 15114 417
rect 15003 356 15114 383
tri 14639 355 14640 356 ne
rect 6976 303 7034 341
rect 14640 345 15114 356
rect 6976 269 6988 303
rect 7022 269 7034 303
rect 14167 280 14252 332
rect 14640 312 15068 345
rect 6976 231 7034 269
rect 6976 197 6988 231
rect 7022 197 7034 231
rect 14640 278 14657 312
rect 14691 278 14735 312
rect 14769 278 14813 312
rect 14847 278 14891 312
rect 14925 278 14969 312
rect 15003 311 15068 312
rect 15102 311 15114 345
rect 15003 278 15114 311
rect 14640 272 15114 278
rect 14640 238 15068 272
rect 15102 238 15114 272
rect 14640 234 15114 238
rect 6976 159 7034 197
rect 13921 168 14073 220
rect 14640 200 14657 234
rect 14691 200 14735 234
rect 14769 200 14813 234
rect 14847 200 14891 234
rect 14925 200 14969 234
rect 15003 200 15114 234
rect 14640 199 15114 200
rect 278 83 284 135
rect 336 83 348 135
rect 400 83 3716 135
rect 3768 83 3796 135
rect 3848 83 3876 135
rect 3928 83 3934 135
rect 6976 125 6988 159
rect 7022 125 7034 159
rect 14640 165 15068 199
rect 15102 165 15114 199
rect 14640 156 15114 165
tri 6967 92 6976 101 se
rect 6976 92 7034 125
tri 6958 83 6967 92 se
rect 6967 83 7034 92
rect 14164 88 14240 140
rect 14640 122 14657 156
rect 14691 122 14735 156
rect 14769 122 14813 156
rect 14847 122 14891 156
rect 14925 122 14969 156
rect 15003 126 15114 156
rect 15003 122 15068 126
rect 14640 92 15068 122
rect 15102 92 15114 126
tri 6952 77 6958 83 se
rect 6958 77 7034 83
tri 6918 43 6952 77 se
rect 6952 43 7034 77
tri 6916 41 6918 43 se
rect 6918 41 7034 43
rect 3524 35 5844 41
tri 5844 35 5850 41 sw
tri 6910 35 6916 41 se
rect 6916 35 7034 41
rect 3524 1 3578 35
rect 3612 1 3652 35
rect 3686 1 3726 35
rect 3760 1 3800 35
rect 3834 1 3874 35
rect 3908 1 3948 35
rect 3982 1 4022 35
rect 4056 1 4096 35
rect 4130 1 4170 35
rect 4204 1 4244 35
rect 4278 1 4318 35
rect 4352 1 4392 35
rect 4426 1 4466 35
rect 4500 1 4540 35
rect 4574 1 4614 35
rect 4648 1 4688 35
rect 4722 1 4762 35
rect 4796 1 4836 35
rect 4870 1 4910 35
rect 4944 1 4984 35
rect 5018 1 5058 35
rect 5092 1 5132 35
rect 5166 1 5206 35
rect 5240 1 5280 35
rect 5314 1 5354 35
rect 5388 1 5428 35
rect 5462 1 5502 35
rect 5536 1 5576 35
rect 5610 1 5650 35
rect 5684 1 5724 35
rect 5758 1 5798 35
rect 5832 23 7034 35
rect 5832 1 5896 23
rect 3524 -5 5896 1
tri 5826 -11 5832 -5 ne
rect 5832 -11 5896 -5
rect 5930 -11 5968 23
rect 6002 -11 6040 23
rect 6074 -11 6112 23
rect 6146 -11 6184 23
rect 6218 -11 6256 23
rect 6290 -11 6328 23
rect 6362 -11 6400 23
rect 6434 -11 6472 23
rect 6506 -11 6544 23
rect 6578 -11 6616 23
rect 6650 -11 6688 23
rect 6722 -11 6760 23
rect 6794 -11 6832 23
rect 6866 -11 6904 23
rect 6938 -11 6976 23
rect 7010 -11 7034 23
tri 5832 -23 5844 -11 ne
rect 5844 -23 7034 -11
rect 14640 77 15114 92
rect 14640 43 14657 77
rect 14691 43 14735 77
rect 14769 43 14813 77
rect 14847 43 14891 77
rect 14925 43 14969 77
rect 15003 53 15114 77
rect 15003 43 15068 53
rect 14640 19 15068 43
rect 15102 19 15114 53
rect 14640 -23 15114 19
rect 49 -1067 83 -1013
rect 167 -1074 205 -1007
rect 258 -1075 313 -1023
rect 377 -1075 415 -1020
rect 5878 -9151 5930 -9145
rect 5878 -9223 5930 -9203
rect 5878 -9281 5930 -9275
rect 5247 -9994 5253 -9942
rect 5305 -9994 5328 -9942
rect 5380 -9994 5403 -9942
rect 5455 -9994 5478 -9942
rect 5530 -9994 5553 -9942
rect 5605 -9994 5627 -9942
rect 5679 -9994 5685 -9942
rect 5247 -10017 5685 -9994
rect 5247 -10069 5253 -10017
rect 5305 -10069 5328 -10017
rect 5380 -10069 5403 -10017
rect 5455 -10069 5478 -10017
rect 5530 -10069 5553 -10017
rect 5605 -10069 5627 -10017
rect 5679 -10069 5685 -10017
rect 5247 -10092 5685 -10069
rect 5247 -10144 5253 -10092
rect 5305 -10144 5328 -10092
rect 5380 -10144 5403 -10092
rect 5455 -10144 5478 -10092
rect 5530 -10144 5553 -10092
rect 5605 -10144 5627 -10092
rect 5679 -10144 5685 -10092
rect 5247 -10985 5253 -10933
rect 5305 -10985 5328 -10933
rect 5380 -10985 5403 -10933
rect 5455 -10985 5478 -10933
rect 5530 -10985 5553 -10933
rect 5605 -10985 5627 -10933
rect 5679 -10985 5685 -10933
rect 5247 -11011 5685 -10985
rect 5247 -11063 5253 -11011
rect 5305 -11063 5328 -11011
rect 5380 -11063 5403 -11011
rect 5455 -11063 5478 -11011
rect 5530 -11063 5553 -11011
rect 5605 -11063 5627 -11011
rect 5679 -11063 5685 -11011
<< rmetal1 >>
rect 9881 8258 9883 8259
rect 10183 8258 10185 8259
rect 9881 7996 9882 8258
rect 10184 7996 10185 8258
rect 9881 7995 9883 7996
rect 10183 7995 10185 7996
<< via1 >>
rect 2287 16493 2339 16505
rect 2287 16459 2303 16493
rect 2303 16459 2337 16493
rect 2337 16459 2339 16493
rect 2287 16453 2339 16459
rect 2369 16493 2421 16505
rect 14101 16493 14153 16505
rect 2369 16459 2375 16493
rect 2375 16459 2409 16493
rect 2409 16459 2421 16493
rect 14101 16459 14111 16493
rect 14111 16459 14145 16493
rect 14145 16459 14153 16493
rect 2369 16453 2421 16459
rect 14101 16453 14153 16459
rect 14175 16493 14227 16505
rect 14175 16459 14183 16493
rect 14183 16459 14217 16493
rect 14217 16459 14227 16493
rect 14175 16453 14227 16459
rect 14249 16493 14301 16505
rect 14249 16459 14255 16493
rect 14255 16459 14289 16493
rect 14289 16459 14301 16493
rect 14249 16453 14301 16459
rect 14323 16493 14375 16505
rect 14323 16459 14327 16493
rect 14327 16459 14361 16493
rect 14361 16459 14375 16493
rect 14323 16453 14375 16459
rect 14397 16493 14449 16505
rect 14397 16459 14399 16493
rect 14399 16459 14433 16493
rect 14433 16459 14449 16493
rect 14397 16453 14449 16459
rect 385 16366 437 16418
rect 506 16372 558 16424
rect 570 16372 622 16424
rect 1938 16372 1990 16424
rect 2002 16372 2054 16424
rect 3468 16372 3520 16424
rect 3532 16372 3584 16424
rect 7754 16372 7806 16424
rect 7818 16372 7870 16424
rect 9456 16372 9508 16424
rect 9520 16372 9572 16424
rect 10936 16372 10988 16424
rect 11000 16372 11052 16424
rect 12279 16372 12331 16424
rect 12343 16372 12395 16424
rect 13713 16372 13765 16424
rect 13777 16372 13829 16424
rect 14946 16372 14998 16424
rect 15010 16372 15062 16424
rect 385 16302 437 16354
rect 748 16292 800 16344
rect 812 16292 864 16344
rect 1655 16292 1707 16344
rect 1719 16292 1771 16344
rect 3185 16292 3237 16344
rect 3249 16292 3301 16344
rect 3960 16292 4012 16344
rect 4024 16292 4076 16344
rect 4088 16292 4140 16344
rect 4152 16292 4204 16344
rect 4216 16292 4268 16344
rect 7324 16292 7376 16344
rect 7388 16292 7440 16344
rect 9026 16292 9078 16344
rect 9090 16292 9142 16344
rect 10506 16292 10558 16344
rect 10570 16292 10622 16344
rect 11849 16292 11901 16344
rect 11913 16292 11965 16344
rect 13283 16292 13335 16344
rect 13347 16292 13399 16344
rect 14866 16292 14918 16344
rect 14930 16292 14982 16344
rect 989 16212 1041 16264
rect 1053 16212 1105 16264
rect 1351 16212 1403 16264
rect 1415 16212 1467 16264
rect 5738 16212 5790 16264
rect 5827 16212 5879 16264
rect 5916 16212 5968 16264
rect 6005 16212 6057 16264
rect 6894 16212 6946 16264
rect 6958 16212 7010 16264
rect 8596 16212 8648 16264
rect 8660 16212 8712 16264
rect 10076 16212 10128 16264
rect 10140 16212 10192 16264
rect 11419 16212 11471 16264
rect 11483 16212 11535 16264
rect 12853 16212 12905 16264
rect 12917 16212 12969 16264
rect 14786 16212 14838 16264
rect 14850 16212 14902 16264
rect 359 16093 411 16145
rect 2538 16103 2590 16155
rect 2602 16103 2654 16155
rect 14706 16103 14758 16155
rect 14770 16103 14822 16155
rect 359 16029 411 16081
rect 8191 16023 8243 16075
rect 8255 16023 8307 16075
rect 9861 16023 9913 16075
rect 9925 16023 9977 16075
rect 10258 16023 10310 16075
rect 10322 16023 10374 16075
rect 14626 16023 14678 16075
rect 14690 16023 14742 16075
rect 278 15937 330 15989
rect 278 15873 330 15925
rect 2162 15937 2214 15989
rect 3616 15943 3668 15995
rect 3680 15943 3732 15995
rect 4439 15980 4491 15985
rect 4506 15980 4558 15985
rect 4573 15980 4625 15985
rect 4640 15980 4692 15985
rect 4707 15980 4759 15985
rect 4774 15980 4826 15985
rect 4841 15980 4893 15985
rect 4908 15980 4960 15985
rect 4439 15946 4466 15980
rect 4466 15946 4491 15980
rect 4506 15946 4539 15980
rect 4539 15946 4558 15980
rect 4573 15946 4612 15980
rect 4612 15946 4625 15980
rect 4640 15946 4646 15980
rect 4646 15946 4685 15980
rect 4685 15946 4692 15980
rect 4707 15946 4719 15980
rect 4719 15946 4758 15980
rect 4758 15946 4759 15980
rect 4774 15946 4792 15980
rect 4792 15946 4826 15980
rect 4841 15946 4865 15980
rect 4865 15946 4893 15980
rect 4908 15946 4938 15980
rect 4938 15946 4960 15980
rect 2162 15873 2214 15925
rect 4439 15933 4491 15946
rect 4506 15933 4558 15946
rect 4573 15933 4625 15946
rect 4640 15933 4692 15946
rect 4707 15933 4759 15946
rect 4774 15933 4826 15946
rect 4841 15933 4893 15946
rect 4908 15933 4960 15946
rect 4975 15980 5027 15985
rect 4975 15946 4977 15980
rect 4977 15946 5011 15980
rect 5011 15946 5027 15980
rect 4975 15933 5027 15946
rect 5042 15980 5094 15985
rect 5042 15946 5050 15980
rect 5050 15946 5084 15980
rect 5084 15946 5094 15980
rect 5042 15933 5094 15946
rect 5108 15980 5160 15985
rect 5108 15946 5123 15980
rect 5123 15946 5157 15980
rect 5157 15946 5160 15980
rect 5108 15933 5160 15946
rect 5174 15980 5226 15985
rect 5240 15980 5292 15985
rect 5306 15980 5358 15985
rect 5372 15980 5424 15985
rect 5438 15980 5490 15985
rect 6198 15980 6250 15985
rect 6269 15980 6321 15985
rect 6339 15980 6391 15985
rect 6409 15980 6461 15985
rect 6479 15980 6531 15985
rect 6549 15980 6601 15985
rect 6619 15980 6671 15985
rect 6689 15980 6741 15985
rect 6759 15980 6811 15985
rect 14103 15980 14155 15985
rect 14201 15980 14253 15985
rect 14298 15980 14350 15985
rect 14395 15980 14447 15985
rect 5174 15946 5196 15980
rect 5196 15946 5226 15980
rect 5240 15946 5269 15980
rect 5269 15946 5292 15980
rect 5306 15946 5342 15980
rect 5342 15946 5358 15980
rect 5372 15946 5376 15980
rect 5376 15946 5415 15980
rect 5415 15946 5424 15980
rect 5438 15946 5449 15980
rect 5449 15946 5488 15980
rect 5488 15946 5490 15980
rect 6198 15946 6218 15980
rect 6218 15946 6250 15980
rect 6269 15946 6291 15980
rect 6291 15946 6321 15980
rect 6339 15946 6364 15980
rect 6364 15946 6391 15980
rect 6409 15946 6437 15980
rect 6437 15946 6461 15980
rect 6479 15946 6510 15980
rect 6510 15946 6531 15980
rect 6549 15946 6583 15980
rect 6583 15946 6601 15980
rect 6619 15946 6656 15980
rect 6656 15946 6671 15980
rect 6689 15946 6690 15980
rect 6690 15946 6729 15980
rect 6729 15946 6741 15980
rect 6759 15946 6763 15980
rect 6763 15946 6802 15980
rect 6802 15946 6811 15980
rect 12534 15946 12549 15980
rect 12549 15946 12586 15980
rect 14103 15946 14133 15980
rect 14133 15946 14155 15980
rect 14201 15946 14205 15980
rect 14205 15946 14243 15980
rect 14243 15946 14253 15980
rect 14298 15946 14315 15980
rect 14315 15946 14349 15980
rect 14349 15946 14350 15980
rect 14395 15946 14421 15980
rect 14421 15946 14447 15980
rect 5174 15933 5226 15946
rect 5240 15933 5292 15946
rect 5306 15933 5358 15946
rect 5372 15933 5424 15946
rect 5438 15933 5490 15946
rect 6198 15933 6250 15946
rect 6269 15933 6321 15946
rect 6339 15933 6391 15946
rect 6409 15933 6461 15946
rect 6479 15933 6531 15946
rect 6549 15933 6601 15946
rect 6619 15933 6671 15946
rect 6689 15933 6741 15946
rect 6759 15933 6811 15946
rect 12534 15928 12586 15946
rect 14103 15933 14155 15946
rect 14201 15933 14253 15946
rect 14298 15933 14350 15946
rect 14395 15933 14447 15946
rect 4439 15906 4491 15915
rect 4506 15906 4558 15915
rect 4573 15906 4625 15915
rect 4640 15906 4692 15915
rect 4707 15906 4759 15915
rect 4774 15906 4826 15915
rect 4841 15906 4893 15915
rect 4908 15906 4960 15915
rect 4439 15872 4466 15906
rect 4466 15872 4491 15906
rect 4506 15872 4539 15906
rect 4539 15872 4558 15906
rect 4573 15872 4612 15906
rect 4612 15872 4625 15906
rect 4640 15872 4646 15906
rect 4646 15872 4685 15906
rect 4685 15872 4692 15906
rect 4707 15872 4719 15906
rect 4719 15872 4758 15906
rect 4758 15872 4759 15906
rect 4774 15872 4792 15906
rect 4792 15872 4826 15906
rect 4841 15872 4865 15906
rect 4865 15872 4893 15906
rect 4908 15872 4938 15906
rect 4938 15872 4960 15906
rect 4439 15863 4491 15872
rect 4506 15863 4558 15872
rect 4573 15863 4625 15872
rect 4640 15863 4692 15872
rect 4707 15863 4759 15872
rect 4774 15863 4826 15872
rect 4841 15863 4893 15872
rect 4908 15863 4960 15872
rect 4975 15906 5027 15915
rect 4975 15872 4977 15906
rect 4977 15872 5011 15906
rect 5011 15872 5027 15906
rect 4975 15863 5027 15872
rect 5042 15906 5094 15915
rect 5042 15872 5050 15906
rect 5050 15872 5084 15906
rect 5084 15872 5094 15906
rect 5042 15863 5094 15872
rect 5108 15906 5160 15915
rect 5108 15872 5123 15906
rect 5123 15872 5157 15906
rect 5157 15872 5160 15906
rect 5108 15863 5160 15872
rect 5174 15906 5226 15915
rect 5240 15906 5292 15915
rect 5306 15906 5358 15915
rect 5372 15906 5424 15915
rect 5438 15906 5490 15915
rect 6198 15906 6250 15915
rect 6269 15906 6321 15915
rect 6339 15906 6391 15915
rect 6409 15906 6461 15915
rect 6479 15906 6531 15915
rect 6549 15906 6601 15915
rect 6619 15906 6671 15915
rect 6689 15906 6741 15915
rect 6759 15906 6811 15915
rect 12534 15906 12586 15915
rect 14103 15906 14155 15917
rect 14201 15906 14253 15917
rect 14298 15906 14350 15917
rect 14395 15906 14447 15917
rect 5174 15872 5196 15906
rect 5196 15872 5226 15906
rect 5240 15872 5269 15906
rect 5269 15872 5292 15906
rect 5306 15872 5342 15906
rect 5342 15872 5358 15906
rect 5372 15872 5376 15906
rect 5376 15872 5415 15906
rect 5415 15872 5424 15906
rect 5438 15872 5449 15906
rect 5449 15872 5488 15906
rect 5488 15872 5490 15906
rect 6198 15872 6218 15906
rect 6218 15872 6250 15906
rect 6269 15872 6291 15906
rect 6291 15872 6321 15906
rect 6339 15872 6364 15906
rect 6364 15872 6391 15906
rect 6409 15872 6437 15906
rect 6437 15872 6461 15906
rect 6479 15872 6510 15906
rect 6510 15872 6531 15906
rect 6549 15872 6583 15906
rect 6583 15872 6601 15906
rect 6619 15872 6656 15906
rect 6656 15872 6671 15906
rect 6689 15872 6690 15906
rect 6690 15872 6729 15906
rect 6729 15872 6741 15906
rect 6759 15872 6763 15906
rect 6763 15872 6802 15906
rect 6802 15872 6811 15906
rect 12534 15872 12549 15906
rect 12549 15872 12586 15906
rect 14103 15872 14133 15906
rect 14133 15872 14155 15906
rect 14201 15872 14205 15906
rect 14205 15872 14243 15906
rect 14243 15872 14253 15906
rect 14298 15872 14315 15906
rect 14315 15872 14349 15906
rect 14349 15872 14350 15906
rect 14395 15872 14421 15906
rect 14421 15872 14447 15906
rect 5174 15863 5226 15872
rect 5240 15863 5292 15872
rect 5306 15863 5358 15872
rect 5372 15863 5424 15872
rect 5438 15863 5490 15872
rect 6198 15863 6250 15872
rect 6269 15863 6321 15872
rect 6339 15863 6391 15872
rect 6409 15863 6461 15872
rect 6479 15863 6531 15872
rect 6549 15863 6601 15872
rect 6619 15863 6671 15872
rect 6689 15863 6741 15872
rect 6759 15863 6811 15872
rect 12534 15863 12586 15872
rect 14103 15865 14155 15872
rect 14201 15865 14253 15872
rect 14298 15865 14350 15872
rect 14395 15865 14447 15872
rect 4439 15832 4491 15845
rect 4506 15832 4558 15845
rect 4573 15832 4625 15845
rect 4640 15832 4692 15845
rect 4707 15832 4759 15845
rect 4774 15832 4826 15845
rect 4841 15832 4893 15845
rect 4908 15832 4960 15845
rect 4439 15798 4466 15832
rect 4466 15798 4491 15832
rect 4506 15798 4539 15832
rect 4539 15798 4558 15832
rect 4573 15798 4612 15832
rect 4612 15798 4625 15832
rect 4640 15798 4646 15832
rect 4646 15798 4685 15832
rect 4685 15798 4692 15832
rect 4707 15798 4719 15832
rect 4719 15798 4758 15832
rect 4758 15798 4759 15832
rect 4774 15798 4792 15832
rect 4792 15798 4826 15832
rect 4841 15798 4865 15832
rect 4865 15798 4893 15832
rect 4908 15798 4938 15832
rect 4938 15798 4960 15832
rect 4439 15793 4491 15798
rect 4506 15793 4558 15798
rect 4573 15793 4625 15798
rect 4640 15793 4692 15798
rect 4707 15793 4759 15798
rect 4774 15793 4826 15798
rect 4841 15793 4893 15798
rect 4908 15793 4960 15798
rect 4975 15832 5027 15845
rect 4975 15798 4977 15832
rect 4977 15798 5011 15832
rect 5011 15798 5027 15832
rect 4975 15793 5027 15798
rect 5042 15832 5094 15845
rect 5042 15798 5050 15832
rect 5050 15798 5084 15832
rect 5084 15798 5094 15832
rect 5042 15793 5094 15798
rect 5108 15832 5160 15845
rect 5108 15798 5123 15832
rect 5123 15798 5157 15832
rect 5157 15798 5160 15832
rect 5108 15793 5160 15798
rect 5174 15832 5226 15845
rect 5240 15832 5292 15845
rect 5306 15832 5358 15845
rect 5372 15832 5424 15845
rect 5438 15832 5490 15845
rect 6198 15832 6250 15845
rect 6269 15832 6321 15845
rect 6339 15832 6391 15845
rect 6409 15832 6461 15845
rect 6479 15832 6531 15845
rect 6549 15832 6601 15845
rect 6619 15832 6671 15845
rect 6689 15832 6741 15845
rect 6759 15832 6811 15845
rect 12534 15832 12586 15850
rect 14103 15832 14155 15849
rect 14201 15832 14253 15849
rect 14298 15832 14350 15849
rect 14395 15832 14447 15849
rect 5174 15798 5196 15832
rect 5196 15798 5226 15832
rect 5240 15798 5269 15832
rect 5269 15798 5292 15832
rect 5306 15798 5342 15832
rect 5342 15798 5358 15832
rect 5372 15798 5376 15832
rect 5376 15798 5415 15832
rect 5415 15798 5424 15832
rect 5438 15798 5449 15832
rect 5449 15798 5488 15832
rect 5488 15798 5490 15832
rect 6198 15798 6218 15832
rect 6218 15798 6250 15832
rect 6269 15798 6291 15832
rect 6291 15798 6321 15832
rect 6339 15798 6364 15832
rect 6364 15798 6391 15832
rect 6409 15798 6437 15832
rect 6437 15798 6461 15832
rect 6479 15798 6510 15832
rect 6510 15798 6531 15832
rect 6549 15798 6583 15832
rect 6583 15798 6601 15832
rect 6619 15798 6656 15832
rect 6656 15798 6671 15832
rect 6689 15798 6690 15832
rect 6690 15798 6729 15832
rect 6729 15798 6741 15832
rect 6759 15798 6763 15832
rect 6763 15798 6802 15832
rect 6802 15798 6811 15832
rect 12534 15798 12549 15832
rect 12549 15798 12586 15832
rect 14103 15798 14133 15832
rect 14133 15798 14155 15832
rect 14201 15798 14205 15832
rect 14205 15798 14243 15832
rect 14243 15798 14253 15832
rect 14298 15798 14315 15832
rect 14315 15798 14349 15832
rect 14349 15798 14350 15832
rect 14395 15798 14421 15832
rect 14421 15798 14447 15832
rect 5174 15793 5226 15798
rect 5240 15793 5292 15798
rect 5306 15793 5358 15798
rect 5372 15793 5424 15798
rect 5438 15793 5490 15798
rect 6198 15793 6250 15798
rect 6269 15793 6321 15798
rect 6339 15793 6391 15798
rect 6409 15793 6461 15798
rect 6479 15793 6531 15798
rect 6549 15793 6601 15798
rect 6619 15793 6671 15798
rect 6689 15793 6741 15798
rect 6759 15793 6811 15798
rect 14103 15797 14155 15798
rect 14201 15797 14253 15798
rect 14298 15797 14350 15798
rect 14395 15797 14447 15798
rect 4439 15737 4491 15743
rect 4506 15737 4558 15743
rect 4573 15737 4625 15743
rect 4640 15737 4692 15743
rect 4707 15737 4759 15743
rect 4439 15703 4446 15737
rect 4446 15703 4484 15737
rect 4484 15703 4491 15737
rect 4506 15703 4518 15737
rect 4518 15703 4557 15737
rect 4557 15703 4558 15737
rect 4573 15703 4591 15737
rect 4591 15703 4625 15737
rect 4640 15703 4664 15737
rect 4664 15703 4692 15737
rect 4707 15703 4737 15737
rect 4737 15703 4759 15737
rect 4439 15691 4491 15703
rect 4506 15691 4558 15703
rect 4573 15691 4625 15703
rect 4640 15691 4692 15703
rect 4707 15691 4759 15703
rect 4774 15737 4826 15743
rect 4774 15703 4776 15737
rect 4776 15703 4810 15737
rect 4810 15703 4826 15737
rect 4774 15691 4826 15703
rect 4841 15737 4893 15743
rect 4841 15703 4849 15737
rect 4849 15703 4883 15737
rect 4883 15703 4893 15737
rect 4841 15691 4893 15703
rect 4908 15737 4960 15743
rect 4908 15703 4922 15737
rect 4922 15703 4956 15737
rect 4956 15703 4960 15737
rect 4908 15691 4960 15703
rect 4975 15737 5027 15743
rect 5042 15737 5094 15743
rect 5108 15737 5160 15743
rect 5174 15737 5226 15743
rect 5240 15737 5292 15743
rect 5306 15737 5358 15743
rect 5372 15737 5424 15743
rect 4975 15703 4995 15737
rect 4995 15703 5027 15737
rect 5042 15703 5068 15737
rect 5068 15703 5094 15737
rect 5108 15703 5141 15737
rect 5141 15703 5160 15737
rect 5174 15703 5175 15737
rect 5175 15703 5214 15737
rect 5214 15703 5226 15737
rect 5240 15703 5248 15737
rect 5248 15703 5287 15737
rect 5287 15703 5292 15737
rect 5306 15703 5321 15737
rect 5321 15703 5358 15737
rect 5372 15703 5394 15737
rect 5394 15703 5424 15737
rect 4975 15691 5027 15703
rect 5042 15691 5094 15703
rect 5108 15691 5160 15703
rect 5174 15691 5226 15703
rect 5240 15691 5292 15703
rect 5306 15691 5358 15703
rect 5372 15691 5424 15703
rect 5438 15691 5490 15743
rect 6198 15691 6250 15743
rect 6269 15691 6321 15743
rect 6339 15691 6391 15743
rect 6409 15691 6461 15743
rect 6479 15691 6531 15743
rect 6549 15691 6601 15743
rect 6619 15691 6671 15743
rect 6689 15691 6741 15743
rect 6759 15691 6811 15743
rect 4591 15504 4643 15513
rect 4658 15504 4710 15513
rect 4725 15504 4777 15513
rect 4792 15504 4844 15513
rect 4591 15470 4632 15504
rect 4632 15470 4643 15504
rect 4658 15470 4666 15504
rect 4666 15470 4708 15504
rect 4708 15470 4710 15504
rect 4725 15470 4742 15504
rect 4742 15470 4777 15504
rect 4792 15470 4818 15504
rect 4818 15470 4844 15504
rect 4591 15461 4643 15470
rect 4658 15461 4710 15470
rect 4725 15461 4777 15470
rect 4792 15461 4844 15470
rect 4859 15504 4911 15513
rect 4859 15470 4860 15504
rect 4860 15470 4894 15504
rect 4894 15470 4911 15504
rect 4859 15461 4911 15470
rect 4926 15504 4978 15513
rect 4926 15470 4936 15504
rect 4936 15470 4970 15504
rect 4970 15470 4978 15504
rect 4926 15461 4978 15470
rect 4993 15504 5045 15513
rect 5059 15504 5111 15513
rect 4993 15470 5012 15504
rect 5012 15470 5045 15504
rect 5059 15470 5088 15504
rect 5088 15470 5111 15504
rect 4993 15461 5045 15470
rect 5059 15461 5111 15470
rect 4602 15357 4625 15381
rect 4625 15357 4654 15381
rect 4687 15357 4701 15381
rect 4701 15357 4739 15381
rect 4772 15357 4777 15381
rect 4777 15357 4819 15381
rect 4819 15357 4824 15381
rect 4856 15357 4894 15381
rect 4894 15357 4908 15381
rect 4940 15357 4969 15381
rect 4969 15357 4992 15381
rect 5024 15357 5044 15381
rect 5044 15357 5076 15381
rect 4602 15329 4654 15357
rect 4687 15329 4739 15357
rect 4772 15329 4824 15357
rect 4856 15329 4908 15357
rect 4940 15329 4992 15357
rect 5024 15329 5076 15357
rect 1942 15305 1994 15311
rect 2006 15305 2058 15311
rect 3616 15305 3668 15311
rect 3680 15305 3732 15311
rect 1942 15271 1967 15305
rect 1967 15271 1994 15305
rect 2006 15271 2039 15305
rect 2039 15271 2058 15305
rect 3616 15271 3642 15305
rect 3642 15271 3668 15305
rect 3680 15271 3715 15305
rect 3715 15271 3732 15305
rect 1942 15259 1994 15271
rect 2006 15259 2058 15271
rect 3616 15259 3668 15271
rect 3680 15259 3732 15271
rect 2487 15203 2539 15215
rect 2487 15169 2498 15203
rect 2498 15169 2532 15203
rect 2532 15169 2539 15203
rect 2487 15163 2539 15169
rect 2551 15203 2603 15215
rect 4602 15213 4654 15265
rect 4687 15213 4739 15265
rect 4772 15213 4824 15265
rect 4856 15213 4908 15265
rect 4940 15213 4992 15265
rect 5024 15213 5076 15265
rect 2551 15169 2572 15203
rect 2572 15169 2603 15203
rect 2551 15163 2603 15169
rect 4602 15136 4654 15149
rect 4687 15136 4739 15149
rect 4772 15136 4824 15149
rect 4856 15136 4908 15149
rect 4940 15136 4992 15149
rect 5024 15136 5076 15149
rect 4602 15102 4625 15136
rect 4625 15102 4654 15136
rect 4687 15102 4701 15136
rect 4701 15102 4739 15136
rect 4772 15102 4777 15136
rect 4777 15102 4819 15136
rect 4819 15102 4824 15136
rect 4856 15102 4894 15136
rect 4894 15102 4908 15136
rect 4940 15102 4969 15136
rect 4969 15102 4992 15136
rect 5024 15102 5044 15136
rect 5044 15102 5076 15136
rect 4602 15097 4654 15102
rect 4687 15097 4739 15102
rect 4772 15097 4824 15102
rect 4856 15097 4908 15102
rect 4940 15097 4992 15102
rect 5024 15097 5076 15102
rect 12534 15685 12586 15737
rect 12534 15615 12586 15667
rect 12534 15545 12586 15597
rect 12534 15475 12586 15527
rect 12534 15405 12586 15457
rect 12534 15334 12586 15386
rect 14101 15430 14118 15459
rect 14118 15430 14152 15459
rect 14152 15430 14153 15459
rect 14101 15407 14153 15430
rect 14175 15430 14191 15459
rect 14191 15430 14225 15459
rect 14225 15430 14227 15459
rect 14175 15407 14227 15430
rect 14249 15430 14264 15459
rect 14264 15430 14298 15459
rect 14298 15430 14301 15459
rect 14249 15407 14301 15430
rect 14323 15430 14337 15459
rect 14337 15430 14371 15459
rect 14371 15430 14375 15459
rect 14323 15407 14375 15430
rect 14397 15430 14410 15459
rect 14410 15430 14444 15459
rect 14444 15430 14449 15459
rect 14397 15407 14449 15430
rect 14101 15382 14153 15394
rect 14101 15348 14118 15382
rect 14118 15348 14152 15382
rect 14152 15348 14153 15382
rect 14101 15342 14153 15348
rect 14175 15382 14227 15394
rect 14175 15348 14191 15382
rect 14191 15348 14225 15382
rect 14225 15348 14227 15382
rect 14175 15342 14227 15348
rect 14249 15382 14301 15394
rect 14249 15348 14264 15382
rect 14264 15348 14298 15382
rect 14298 15348 14301 15382
rect 14249 15342 14301 15348
rect 14323 15382 14375 15394
rect 14323 15348 14337 15382
rect 14337 15348 14371 15382
rect 14371 15348 14375 15382
rect 14323 15342 14375 15348
rect 14397 15382 14449 15394
rect 14397 15348 14410 15382
rect 14410 15348 14444 15382
rect 14444 15348 14449 15382
rect 14397 15342 14449 15348
rect 8189 15259 8241 15311
rect 8255 15259 8307 15311
rect 9861 15259 9913 15311
rect 9927 15259 9979 15311
rect 14101 15300 14153 15328
rect 14101 15276 14118 15300
rect 14118 15276 14152 15300
rect 14152 15276 14153 15300
rect 14175 15300 14227 15328
rect 14175 15276 14191 15300
rect 14191 15276 14225 15300
rect 14225 15276 14227 15300
rect 14249 15300 14301 15328
rect 14249 15276 14264 15300
rect 14264 15276 14298 15300
rect 14298 15276 14301 15300
rect 14323 15300 14375 15328
rect 14323 15276 14337 15300
rect 14337 15276 14371 15300
rect 14371 15276 14375 15300
rect 14397 15300 14449 15328
rect 14397 15276 14410 15300
rect 14410 15276 14444 15300
rect 14444 15276 14449 15300
rect 14101 15218 14153 15262
rect 9666 15163 9718 15215
rect 9730 15163 9782 15215
rect 14101 15210 14118 15218
rect 14118 15210 14152 15218
rect 14152 15210 14153 15218
rect 14175 15218 14227 15262
rect 14175 15210 14191 15218
rect 14191 15210 14225 15218
rect 14225 15210 14227 15218
rect 14249 15218 14301 15262
rect 14249 15210 14264 15218
rect 14264 15210 14298 15218
rect 14298 15210 14301 15218
rect 14323 15218 14375 15262
rect 14323 15210 14337 15218
rect 14337 15210 14371 15218
rect 14371 15210 14375 15218
rect 14397 15218 14449 15262
rect 14397 15210 14410 15218
rect 14410 15210 14444 15218
rect 14444 15210 14449 15218
rect 14101 15184 14118 15196
rect 14118 15184 14152 15196
rect 14152 15184 14153 15196
rect 14101 15144 14153 15184
rect 14175 15184 14191 15196
rect 14191 15184 14225 15196
rect 14225 15184 14227 15196
rect 14175 15144 14227 15184
rect 14249 15184 14264 15196
rect 14264 15184 14298 15196
rect 14298 15184 14301 15196
rect 14249 15144 14301 15184
rect 14323 15184 14337 15196
rect 14337 15184 14371 15196
rect 14371 15184 14375 15196
rect 14323 15144 14375 15184
rect 14397 15184 14410 15196
rect 14410 15184 14444 15196
rect 14444 15184 14449 15196
rect 14397 15144 14449 15184
rect 14101 15102 14118 15130
rect 14118 15102 14152 15130
rect 14152 15102 14153 15130
rect 14101 15078 14153 15102
rect 14175 15102 14191 15130
rect 14191 15102 14225 15130
rect 14225 15102 14227 15130
rect 14175 15078 14227 15102
rect 14249 15102 14264 15130
rect 14264 15102 14298 15130
rect 14298 15102 14301 15130
rect 14249 15078 14301 15102
rect 14323 15102 14337 15130
rect 14337 15102 14371 15130
rect 14371 15102 14375 15130
rect 14323 15078 14375 15102
rect 14397 15102 14410 15130
rect 14410 15102 14444 15130
rect 14444 15102 14449 15130
rect 14397 15078 14449 15102
rect 14101 15054 14153 15064
rect 14101 15020 14118 15054
rect 14118 15020 14152 15054
rect 14152 15020 14153 15054
rect 14101 15012 14153 15020
rect 14175 15054 14227 15064
rect 14175 15020 14191 15054
rect 14191 15020 14225 15054
rect 14225 15020 14227 15054
rect 14175 15012 14227 15020
rect 14249 15054 14301 15064
rect 14249 15020 14264 15054
rect 14264 15020 14298 15054
rect 14298 15020 14301 15054
rect 14249 15012 14301 15020
rect 14323 15054 14375 15064
rect 14323 15020 14337 15054
rect 14337 15020 14371 15054
rect 14371 15020 14375 15054
rect 14323 15012 14375 15020
rect 14397 15054 14449 15064
rect 14397 15020 14410 15054
rect 14410 15020 14444 15054
rect 14444 15020 14449 15054
rect 14397 15012 14449 15020
rect 14101 14972 14153 14998
rect 14101 14946 14118 14972
rect 14118 14946 14152 14972
rect 14152 14946 14153 14972
rect 14175 14972 14227 14998
rect 14175 14946 14191 14972
rect 14191 14946 14225 14972
rect 14225 14946 14227 14972
rect 14249 14972 14301 14998
rect 14249 14946 14264 14972
rect 14264 14946 14298 14972
rect 14298 14946 14301 14972
rect 14323 14972 14375 14998
rect 14323 14946 14337 14972
rect 14337 14946 14371 14972
rect 14371 14946 14375 14972
rect 14397 14972 14449 14998
rect 14397 14946 14410 14972
rect 14410 14946 14444 14972
rect 14444 14946 14449 14972
rect 1861 14731 1913 14783
rect 1955 14731 2007 14783
rect 1861 14662 1913 14714
rect 1955 14662 2007 14714
rect 1861 14593 1913 14645
rect 1955 14593 2007 14645
rect 14101 14736 14153 14788
rect 14175 14736 14227 14788
rect 14249 14736 14301 14788
rect 14323 14736 14375 14788
rect 14397 14736 14449 14788
rect 14101 14662 14153 14714
rect 14175 14662 14227 14714
rect 14249 14662 14301 14714
rect 14323 14662 14375 14714
rect 14397 14662 14449 14714
rect 14101 14588 14153 14640
rect 14175 14588 14227 14640
rect 14249 14588 14301 14640
rect 14323 14588 14375 14640
rect 14397 14588 14449 14640
rect 876 13798 928 13850
rect 942 13798 994 13850
rect 876 13734 928 13786
rect 942 13734 994 13786
rect 2226 13805 2278 13857
rect 2292 13805 2344 13857
rect 2226 13727 2278 13779
rect 2292 13727 2344 13779
rect 2788 13798 2840 13850
rect 2854 13798 2906 13850
rect 2788 13734 2840 13786
rect 2854 13734 2906 13786
rect 3901 13798 3953 13850
rect 3980 13798 4032 13850
rect 4059 13798 4111 13850
rect 4138 13798 4190 13850
rect 4216 13798 4268 13850
rect 3901 13734 3953 13786
rect 3980 13734 4032 13786
rect 4059 13734 4111 13786
rect 4138 13734 4190 13786
rect 4216 13734 4268 13786
rect 6194 13799 6246 13851
rect 6259 13799 6311 13851
rect 6324 13799 6376 13851
rect 6389 13799 6441 13851
rect 6453 13799 6505 13851
rect 6517 13799 6569 13851
rect 6581 13799 6633 13851
rect 6645 13799 6697 13851
rect 6709 13799 6761 13851
rect 6773 13799 6825 13851
rect 6837 13799 6889 13851
rect 6194 13727 6246 13779
rect 6259 13727 6311 13779
rect 6324 13727 6376 13779
rect 6389 13727 6441 13779
rect 6453 13727 6505 13779
rect 6517 13727 6569 13779
rect 6581 13727 6633 13779
rect 6645 13727 6697 13779
rect 6709 13727 6761 13779
rect 6773 13727 6825 13779
rect 6837 13727 6889 13779
rect 7748 13805 7800 13857
rect 7814 13805 7866 13857
rect 7748 13727 7800 13779
rect 7814 13727 7866 13779
rect 8680 13801 8732 13853
rect 8745 13801 8797 13853
rect 8809 13801 8861 13853
rect 8873 13801 8925 13853
rect 8680 13727 8732 13779
rect 8745 13727 8797 13779
rect 8809 13727 8861 13779
rect 8873 13727 8925 13779
rect 10305 13769 10357 13821
rect 10371 13769 10423 13821
rect 10437 13769 10489 13821
rect 10503 13769 10555 13821
rect 10568 13769 10620 13821
rect 10633 13769 10685 13821
rect 10698 13769 10750 13821
rect 10763 13769 10815 13821
rect 11716 13768 11768 13820
rect 11781 13768 11833 13820
rect 11846 13768 11898 13820
rect 11911 13768 11963 13820
rect 11976 13768 12028 13820
rect 12041 13768 12093 13820
rect 12106 13768 12158 13820
rect 13138 13805 13190 13857
rect 13205 13805 13257 13857
rect 13272 13805 13324 13857
rect 13339 13805 13391 13857
rect 13406 13805 13458 13857
rect 13473 13805 13525 13857
rect 13540 13805 13592 13857
rect 13138 13727 13190 13779
rect 13205 13727 13257 13779
rect 13272 13727 13324 13779
rect 13339 13727 13391 13779
rect 13406 13727 13458 13779
rect 13473 13727 13525 13779
rect 13540 13727 13592 13779
rect 541 9978 593 10030
rect 616 9978 668 10030
rect 690 9978 742 10030
rect 764 9978 816 10030
rect 838 9978 890 10030
rect 912 9978 964 10030
rect 541 9904 593 9956
rect 616 9904 668 9956
rect 690 9904 742 9956
rect 764 9904 816 9956
rect 838 9904 890 9956
rect 912 9904 964 9956
rect 541 9830 593 9882
rect 616 9830 668 9882
rect 690 9830 742 9882
rect 764 9830 816 9882
rect 838 9830 890 9882
rect 912 9830 964 9882
rect 12258 9342 12310 9359
rect 12335 9342 12387 9359
rect 12412 9342 12464 9359
rect 12488 9342 12540 9359
rect 12258 9308 12287 9342
rect 12287 9308 12310 9342
rect 12335 9308 12359 9342
rect 12359 9308 12387 9342
rect 12412 9308 12431 9342
rect 12431 9308 12464 9342
rect 12488 9308 12503 9342
rect 12503 9308 12537 9342
rect 12537 9308 12540 9342
rect 12258 9307 12310 9308
rect 12335 9307 12387 9308
rect 12412 9307 12464 9308
rect 12488 9307 12540 9308
rect 12564 9342 12616 9359
rect 12564 9308 12575 9342
rect 12575 9308 12609 9342
rect 12609 9308 12616 9342
rect 12564 9307 12616 9308
rect 12258 9256 12310 9271
rect 12335 9256 12387 9271
rect 12412 9256 12464 9271
rect 12488 9256 12540 9271
rect 12258 9222 12287 9256
rect 12287 9222 12310 9256
rect 12335 9222 12359 9256
rect 12359 9222 12387 9256
rect 12412 9222 12431 9256
rect 12431 9222 12464 9256
rect 12488 9222 12503 9256
rect 12503 9222 12537 9256
rect 12537 9222 12540 9256
rect 12258 9219 12310 9222
rect 12335 9219 12387 9222
rect 12412 9219 12464 9222
rect 12488 9219 12540 9222
rect 12564 9256 12616 9271
rect 12564 9222 12575 9256
rect 12575 9222 12609 9256
rect 12609 9222 12616 9256
rect 12564 9219 12616 9222
rect 12258 9170 12310 9183
rect 12335 9170 12387 9183
rect 12412 9170 12464 9183
rect 12488 9170 12540 9183
rect 12258 9136 12287 9170
rect 12287 9136 12310 9170
rect 12335 9136 12359 9170
rect 12359 9136 12387 9170
rect 12412 9136 12431 9170
rect 12431 9136 12464 9170
rect 12488 9136 12503 9170
rect 12503 9136 12537 9170
rect 12537 9136 12540 9170
rect 12258 9131 12310 9136
rect 12335 9131 12387 9136
rect 12412 9131 12464 9136
rect 12488 9131 12540 9136
rect 12564 9170 12616 9183
rect 12564 9136 12575 9170
rect 12575 9136 12609 9170
rect 12609 9136 12616 9170
rect 12564 9131 12616 9136
rect 14240 9408 14292 9460
rect 14312 9408 14364 9460
rect 14384 9408 14436 9460
rect 14456 9408 14508 9460
rect 14528 9408 14580 9460
rect 14600 9408 14652 9460
rect 14240 9343 14292 9395
rect 14312 9343 14364 9395
rect 14384 9343 14436 9395
rect 14456 9343 14508 9395
rect 14528 9343 14580 9395
rect 14600 9343 14652 9395
rect 14240 9278 14292 9330
rect 14312 9278 14364 9330
rect 14384 9278 14436 9330
rect 14456 9278 14508 9330
rect 14528 9278 14580 9330
rect 14600 9278 14652 9330
rect 14240 9213 14292 9265
rect 14312 9213 14364 9265
rect 14384 9213 14436 9265
rect 14456 9213 14508 9265
rect 14528 9213 14580 9265
rect 14600 9213 14652 9265
rect 14240 9148 14292 9200
rect 14312 9148 14364 9200
rect 14384 9148 14436 9200
rect 14456 9148 14508 9200
rect 14528 9148 14580 9200
rect 14600 9148 14652 9200
rect 14240 9083 14292 9135
rect 14312 9083 14364 9135
rect 14384 9083 14436 9135
rect 14456 9083 14508 9135
rect 14528 9083 14580 9135
rect 14600 9083 14652 9135
rect 14240 9018 14292 9070
rect 14312 9018 14364 9070
rect 14384 9018 14436 9070
rect 14456 9018 14508 9070
rect 14528 9018 14580 9070
rect 14600 9018 14652 9070
rect 14240 8953 14292 9005
rect 14312 8953 14364 9005
rect 14384 8953 14436 9005
rect 14456 8953 14508 9005
rect 14528 8953 14580 9005
rect 14600 8953 14652 9005
rect 14240 8888 14292 8940
rect 14312 8888 14364 8940
rect 14384 8888 14436 8940
rect 14456 8888 14508 8940
rect 14528 8888 14580 8940
rect 14600 8888 14652 8940
rect 541 8775 593 8827
rect 616 8775 668 8827
rect 690 8775 742 8827
rect 764 8775 816 8827
rect 838 8775 890 8827
rect 912 8775 964 8827
rect 14240 8823 14292 8875
rect 14312 8823 14364 8875
rect 14384 8823 14436 8875
rect 14456 8823 14508 8875
rect 14528 8823 14580 8875
rect 14600 8823 14652 8875
rect 14240 8760 14292 8810
rect 14312 8760 14364 8810
rect 14384 8760 14436 8810
rect 14456 8760 14508 8810
rect 14528 8760 14580 8810
rect 14600 8760 14652 8810
rect 541 8719 544 8751
rect 544 8719 578 8751
rect 578 8719 593 8751
rect 541 8699 593 8719
rect 616 8719 618 8751
rect 618 8719 652 8751
rect 652 8719 668 8751
rect 616 8699 668 8719
rect 690 8719 691 8751
rect 691 8719 725 8751
rect 725 8719 742 8751
rect 690 8699 742 8719
rect 764 8719 798 8751
rect 798 8719 816 8751
rect 838 8719 871 8751
rect 871 8719 890 8751
rect 764 8699 816 8719
rect 838 8699 890 8719
rect 912 8726 946 8751
rect 946 8726 964 8751
rect 912 8699 964 8726
rect 14240 8758 14267 8760
rect 14267 8758 14292 8760
rect 14312 8758 14339 8760
rect 14339 8758 14364 8760
rect 14384 8758 14411 8760
rect 14411 8758 14436 8760
rect 14456 8758 14483 8760
rect 14483 8758 14508 8760
rect 14528 8758 14555 8760
rect 14555 8758 14580 8760
rect 14600 8758 14627 8760
rect 14627 8758 14652 8760
rect 14240 8726 14267 8745
rect 14267 8726 14292 8745
rect 14312 8726 14339 8745
rect 14339 8726 14364 8745
rect 14384 8726 14411 8745
rect 14411 8726 14436 8745
rect 14456 8726 14483 8745
rect 14483 8726 14508 8745
rect 14528 8726 14555 8745
rect 14555 8726 14580 8745
rect 14600 8726 14627 8745
rect 14627 8726 14652 8745
rect 842 8618 894 8670
rect 912 8636 964 8670
rect 14240 8693 14292 8726
rect 14312 8693 14364 8726
rect 14384 8693 14436 8726
rect 14456 8693 14508 8726
rect 14528 8693 14580 8726
rect 14600 8693 14652 8726
rect 14240 8636 14292 8680
rect 14312 8636 14364 8680
rect 14384 8636 14436 8680
rect 14456 8636 14508 8680
rect 14528 8636 14580 8680
rect 14600 8636 14652 8680
rect 912 8618 946 8636
rect 946 8618 964 8636
rect 14240 8628 14267 8636
rect 14267 8628 14292 8636
rect 14312 8628 14339 8636
rect 14339 8628 14364 8636
rect 14384 8628 14411 8636
rect 14411 8628 14436 8636
rect 14456 8628 14483 8636
rect 14483 8628 14508 8636
rect 14528 8628 14555 8636
rect 14555 8628 14580 8636
rect 14600 8628 14627 8636
rect 14627 8628 14652 8636
rect 14240 8602 14267 8615
rect 14267 8602 14292 8615
rect 14312 8602 14339 8615
rect 14339 8602 14364 8615
rect 14384 8602 14411 8615
rect 14411 8602 14436 8615
rect 14456 8602 14483 8615
rect 14483 8602 14508 8615
rect 14528 8602 14555 8615
rect 14555 8602 14580 8615
rect 14600 8602 14627 8615
rect 14627 8602 14652 8615
rect 14240 8563 14292 8602
rect 14312 8563 14364 8602
rect 14384 8563 14436 8602
rect 14456 8563 14508 8602
rect 14528 8563 14580 8602
rect 14600 8563 14652 8602
rect 14240 8512 14292 8550
rect 14240 8498 14257 8512
rect 14257 8498 14291 8512
rect 14291 8498 14292 8512
rect 14312 8512 14364 8550
rect 14312 8498 14329 8512
rect 14329 8498 14363 8512
rect 14363 8498 14364 8512
rect 14384 8512 14436 8550
rect 14384 8498 14401 8512
rect 14401 8498 14435 8512
rect 14435 8498 14436 8512
rect 14456 8512 14508 8550
rect 14456 8498 14473 8512
rect 14473 8498 14507 8512
rect 14507 8498 14508 8512
rect 14528 8498 14580 8550
rect 14600 8498 14652 8550
rect 14240 8478 14257 8485
rect 14257 8478 14291 8485
rect 14291 8478 14292 8485
rect 14240 8435 14292 8478
rect 14240 8433 14257 8435
rect 14257 8433 14291 8435
rect 14291 8433 14292 8435
rect 14312 8478 14329 8485
rect 14329 8478 14363 8485
rect 14363 8478 14364 8485
rect 14312 8435 14364 8478
rect 14312 8433 14329 8435
rect 14329 8433 14363 8435
rect 14363 8433 14364 8435
rect 14384 8478 14401 8485
rect 14401 8478 14435 8485
rect 14435 8478 14436 8485
rect 14384 8435 14436 8478
rect 14384 8433 14401 8435
rect 14401 8433 14435 8435
rect 14435 8433 14436 8435
rect 14456 8478 14473 8485
rect 14473 8478 14507 8485
rect 14507 8478 14508 8485
rect 14456 8435 14508 8478
rect 14456 8433 14473 8435
rect 14473 8433 14507 8435
rect 14507 8433 14508 8435
rect 14528 8433 14580 8485
rect 14600 8462 14652 8485
rect 14600 8433 14614 8462
rect 14614 8433 14648 8462
rect 14648 8433 14652 8462
rect 14240 8401 14257 8420
rect 14257 8401 14291 8420
rect 14291 8401 14292 8420
rect 406 8355 458 8359
rect 406 8321 426 8355
rect 426 8321 458 8355
rect 406 8307 458 8321
rect 406 8243 458 8295
rect 14240 8368 14292 8401
rect 14312 8401 14329 8420
rect 14329 8401 14363 8420
rect 14363 8401 14364 8420
rect 14312 8368 14364 8401
rect 14384 8401 14401 8420
rect 14401 8401 14435 8420
rect 14435 8401 14436 8420
rect 14384 8368 14436 8401
rect 14456 8401 14473 8420
rect 14473 8401 14507 8420
rect 14507 8401 14508 8420
rect 14456 8368 14508 8401
rect 14528 8368 14580 8420
rect 14600 8388 14652 8420
rect 14600 8368 14614 8388
rect 14614 8368 14648 8388
rect 14648 8368 14652 8388
rect 14240 8324 14257 8354
rect 14257 8324 14291 8354
rect 14291 8324 14292 8354
rect 14240 8302 14292 8324
rect 14312 8324 14329 8354
rect 14329 8324 14363 8354
rect 14363 8324 14364 8354
rect 14312 8302 14364 8324
rect 14384 8324 14401 8354
rect 14401 8324 14435 8354
rect 14435 8324 14436 8354
rect 14384 8302 14436 8324
rect 14456 8324 14473 8354
rect 14473 8324 14507 8354
rect 14507 8324 14508 8354
rect 14456 8302 14508 8324
rect 14528 8302 14580 8354
rect 14600 8314 14652 8354
rect 14600 8302 14614 8314
rect 14614 8302 14648 8314
rect 14648 8302 14652 8314
rect 10800 8254 10852 8281
rect 10800 8229 10804 8254
rect 10804 8229 10838 8254
rect 10838 8229 10852 8254
rect 10876 8254 10928 8281
rect 10876 8229 10898 8254
rect 10898 8229 10928 8254
rect 10952 8229 11004 8281
rect 11028 8229 11080 8281
rect 11104 8229 11156 8281
rect 10800 8179 10852 8214
rect 10800 8162 10804 8179
rect 10804 8162 10838 8179
rect 10838 8162 10852 8179
rect 10876 8179 10928 8214
rect 10876 8162 10898 8179
rect 10898 8162 10928 8179
rect 10952 8162 11004 8214
rect 11028 8162 11080 8214
rect 11104 8162 11156 8214
rect 10800 8145 10804 8147
rect 10804 8145 10838 8147
rect 10838 8145 10852 8147
rect 10800 8104 10852 8145
rect 10800 8095 10804 8104
rect 10804 8095 10838 8104
rect 10838 8095 10852 8104
rect 10876 8145 10898 8147
rect 10898 8145 10928 8147
rect 10876 8104 10928 8145
rect 10876 8095 10898 8104
rect 10898 8095 10928 8104
rect 10952 8095 11004 8147
rect 11028 8095 11080 8147
rect 11104 8095 11156 8147
rect 10800 8070 10804 8079
rect 10804 8070 10838 8079
rect 10838 8070 10852 8079
rect 10800 8028 10852 8070
rect 10800 8027 10804 8028
rect 10804 8027 10838 8028
rect 10838 8027 10852 8028
rect 10876 8070 10898 8079
rect 10898 8070 10928 8079
rect 10876 8028 10928 8070
rect 10876 8027 10898 8028
rect 10898 8027 10928 8028
rect 10952 8027 11004 8079
rect 11028 8027 11080 8079
rect 11104 8027 11156 8079
rect 10800 7994 10804 8011
rect 10804 7994 10838 8011
rect 10838 7994 10852 8011
rect 10800 7959 10852 7994
rect 10876 7994 10898 8011
rect 10898 7994 10928 8011
rect 10876 7959 10928 7994
rect 10952 7959 11004 8011
rect 11028 7959 11080 8011
rect 11104 7959 11156 8011
rect 10800 7918 10804 7943
rect 10804 7918 10838 7943
rect 10838 7918 10852 7943
rect 10800 7891 10852 7918
rect 10876 7918 10898 7943
rect 10898 7918 10928 7943
rect 10876 7891 10928 7918
rect 10952 7891 11004 7943
rect 11028 7891 11080 7943
rect 11104 7891 11156 7943
rect 12255 8229 12307 8281
rect 12333 8229 12385 8281
rect 12411 8229 12463 8281
rect 12489 8229 12541 8281
rect 12567 8229 12619 8281
rect 14240 8280 14292 8288
rect 12255 8158 12307 8210
rect 12333 8158 12385 8210
rect 12411 8158 12463 8210
rect 12489 8158 12541 8210
rect 12567 8158 12619 8210
rect 12255 8087 12307 8139
rect 12333 8087 12385 8139
rect 12411 8087 12463 8139
rect 12489 8087 12541 8139
rect 12567 8087 12619 8139
rect 12255 8016 12307 8068
rect 12333 8016 12385 8068
rect 12411 8016 12463 8068
rect 12489 8016 12541 8068
rect 12567 8016 12619 8068
rect 12255 7945 12307 7997
rect 12333 7945 12385 7997
rect 12411 7945 12463 7997
rect 12489 7945 12541 7997
rect 12567 7945 12619 7997
rect 12255 7873 12307 7925
rect 12333 7873 12385 7925
rect 12411 7873 12463 7925
rect 12489 7873 12541 7925
rect 12567 7873 12619 7925
rect 14240 8246 14257 8280
rect 14257 8246 14291 8280
rect 14291 8246 14292 8280
rect 14240 8236 14292 8246
rect 14312 8280 14364 8288
rect 14312 8246 14329 8280
rect 14329 8246 14363 8280
rect 14363 8246 14364 8280
rect 14312 8236 14364 8246
rect 14384 8280 14436 8288
rect 14384 8246 14401 8280
rect 14401 8246 14435 8280
rect 14435 8246 14436 8280
rect 14384 8236 14436 8246
rect 14456 8280 14508 8288
rect 14456 8246 14473 8280
rect 14473 8246 14507 8280
rect 14507 8246 14508 8280
rect 14456 8236 14508 8246
rect 14528 8236 14580 8288
rect 14600 8280 14614 8288
rect 14614 8280 14648 8288
rect 14648 8280 14652 8288
rect 14600 8240 14652 8280
rect 14600 8236 14614 8240
rect 14614 8236 14648 8240
rect 14648 8236 14652 8240
rect 14240 8202 14292 8222
rect 14240 8170 14257 8202
rect 14257 8170 14291 8202
rect 14291 8170 14292 8202
rect 14312 8202 14364 8222
rect 14312 8170 14329 8202
rect 14329 8170 14363 8202
rect 14363 8170 14364 8202
rect 14384 8202 14436 8222
rect 14384 8170 14401 8202
rect 14401 8170 14435 8202
rect 14435 8170 14436 8202
rect 14456 8202 14508 8222
rect 14456 8170 14473 8202
rect 14473 8170 14507 8202
rect 14507 8170 14508 8202
rect 14528 8170 14580 8222
rect 14600 8206 14614 8222
rect 14614 8206 14648 8222
rect 14648 8206 14652 8222
rect 14600 8170 14652 8206
rect 14240 8104 14292 8156
rect 14312 8104 14364 8156
rect 14384 8115 14436 8156
rect 14456 8115 14508 8156
rect 14528 8115 14580 8156
rect 14384 8104 14431 8115
rect 14431 8104 14436 8115
rect 14456 8104 14465 8115
rect 14465 8104 14508 8115
rect 14528 8104 14545 8115
rect 14545 8104 14580 8115
rect 14600 8132 14614 8156
rect 14614 8132 14648 8156
rect 14648 8132 14652 8156
rect 14600 8104 14652 8132
rect 278 7799 330 7851
rect 278 7733 330 7785
rect 278 7666 330 7718
rect 278 7599 330 7651
rect 278 7532 330 7584
rect 11135 7509 11187 7561
rect 11208 7509 11260 7561
rect 11280 7509 11332 7561
rect 11135 7429 11187 7481
rect 11208 7429 11260 7481
rect 11280 7429 11332 7481
rect 338 6822 390 6874
rect 338 6756 390 6808
rect 516 5516 568 5568
rect 634 5516 686 5568
rect 751 5516 803 5568
rect 14313 5513 14365 5565
rect 435 5413 487 5465
rect 507 5413 559 5465
rect 579 5413 631 5465
rect 651 5413 703 5465
rect 748 5427 800 5479
rect 435 5348 487 5400
rect 507 5348 559 5400
rect 579 5348 631 5400
rect 651 5348 703 5400
rect 435 5283 487 5335
rect 507 5283 559 5335
rect 579 5283 631 5335
rect 651 5283 703 5335
rect 435 5218 487 5270
rect 507 5218 559 5270
rect 579 5218 631 5270
rect 651 5218 703 5270
rect 435 5153 487 5205
rect 507 5153 559 5205
rect 579 5153 631 5205
rect 651 5153 703 5205
rect 435 5088 487 5140
rect 507 5088 559 5140
rect 579 5088 631 5140
rect 651 5088 703 5140
rect 435 5023 487 5075
rect 507 5023 559 5075
rect 579 5023 631 5075
rect 651 5023 703 5075
rect 435 4958 487 5010
rect 507 4958 559 5010
rect 579 4958 631 5010
rect 651 4958 703 5010
rect 435 4893 487 4945
rect 507 4893 559 4945
rect 579 4893 631 4945
rect 651 4893 703 4945
rect 435 4828 487 4880
rect 507 4828 559 4880
rect 579 4828 631 4880
rect 651 4828 703 4880
rect 435 4763 487 4815
rect 507 4763 559 4815
rect 579 4763 631 4815
rect 651 4763 703 4815
rect 435 4698 487 4750
rect 507 4698 559 4750
rect 579 4698 631 4750
rect 651 4698 703 4750
rect 435 4633 487 4685
rect 507 4633 559 4685
rect 579 4633 631 4685
rect 651 4633 703 4685
rect 435 4568 487 4620
rect 507 4568 559 4620
rect 579 4568 631 4620
rect 651 4568 703 4620
rect 435 4503 487 4555
rect 507 4503 559 4555
rect 579 4503 631 4555
rect 651 4503 703 4555
rect 435 4438 487 4490
rect 507 4438 559 4490
rect 579 4438 631 4490
rect 651 4438 703 4490
rect 435 4373 487 4425
rect 507 4373 559 4425
rect 579 4373 631 4425
rect 651 4373 703 4425
rect 435 4308 487 4360
rect 507 4308 559 4360
rect 579 4308 631 4360
rect 651 4308 703 4360
rect 435 4243 487 4295
rect 507 4243 559 4295
rect 579 4243 631 4295
rect 651 4243 703 4295
rect 435 4178 487 4230
rect 507 4178 559 4230
rect 579 4178 631 4230
rect 651 4178 703 4230
rect 435 4113 487 4165
rect 507 4113 559 4165
rect 579 4113 631 4165
rect 651 4113 703 4165
rect 435 4047 487 4099
rect 507 4047 559 4099
rect 579 4047 631 4099
rect 651 4047 703 4099
rect 435 3981 487 4033
rect 507 3981 559 4033
rect 579 3981 631 4033
rect 651 3981 703 4033
rect 435 3915 487 3967
rect 507 3915 559 3967
rect 579 3915 631 3967
rect 651 3915 703 3967
rect 435 3849 487 3901
rect 507 3849 559 3901
rect 579 3849 631 3901
rect 651 3849 703 3901
rect 435 3783 487 3835
rect 507 3783 559 3835
rect 579 3783 631 3835
rect 651 3783 703 3835
rect 435 3717 487 3769
rect 507 3717 559 3769
rect 579 3717 631 3769
rect 651 3717 703 3769
rect 435 3651 487 3703
rect 507 3651 559 3703
rect 579 3651 631 3703
rect 651 3651 703 3703
rect 14243 5413 14295 5465
rect 14309 5413 14361 5465
rect 14375 5413 14427 5465
rect 14441 5413 14493 5465
rect 14243 5348 14295 5400
rect 14309 5348 14361 5400
rect 14375 5348 14427 5400
rect 14441 5348 14493 5400
rect 14243 5283 14295 5335
rect 14309 5283 14361 5335
rect 14375 5283 14427 5335
rect 14441 5283 14493 5335
rect 14243 5218 14295 5270
rect 14309 5218 14361 5270
rect 14375 5218 14427 5270
rect 14441 5218 14493 5270
rect 14243 5153 14295 5205
rect 14309 5153 14361 5205
rect 14375 5153 14427 5205
rect 14441 5153 14493 5205
rect 14243 5088 14295 5140
rect 14309 5088 14361 5140
rect 14375 5088 14427 5140
rect 14441 5088 14493 5140
rect 14243 5023 14295 5075
rect 14309 5023 14361 5075
rect 14375 5023 14427 5075
rect 14441 5023 14493 5075
rect 14243 4958 14295 5010
rect 14309 4958 14361 5010
rect 14375 4958 14427 5010
rect 14441 4958 14493 5010
rect 14243 4893 14295 4945
rect 14309 4893 14361 4945
rect 14375 4893 14427 4945
rect 14441 4893 14493 4945
rect 14243 4828 14295 4880
rect 14309 4828 14361 4880
rect 14375 4828 14427 4880
rect 14441 4828 14493 4880
rect 14243 4763 14295 4815
rect 14309 4763 14361 4815
rect 14375 4763 14427 4815
rect 14441 4763 14493 4815
rect 14243 4698 14295 4750
rect 14309 4698 14361 4750
rect 14375 4698 14427 4750
rect 14441 4698 14493 4750
rect 14243 4633 14295 4685
rect 14309 4633 14361 4685
rect 14375 4633 14427 4685
rect 14441 4633 14493 4685
rect 14243 4568 14295 4620
rect 14309 4568 14361 4620
rect 14375 4568 14427 4620
rect 14441 4568 14493 4620
rect 14243 4503 14295 4555
rect 14309 4503 14361 4555
rect 14375 4503 14427 4555
rect 14441 4503 14493 4555
rect 14243 4438 14295 4490
rect 14309 4438 14361 4490
rect 14375 4438 14427 4490
rect 14441 4438 14493 4490
rect 14243 4373 14295 4425
rect 14309 4373 14361 4425
rect 14375 4373 14427 4425
rect 14441 4373 14493 4425
rect 14243 4307 14295 4359
rect 14309 4307 14361 4359
rect 14375 4307 14427 4359
rect 14441 4307 14493 4359
rect 14243 4241 14295 4293
rect 14309 4241 14361 4293
rect 14375 4241 14427 4293
rect 14441 4241 14493 4293
rect 14243 4175 14295 4227
rect 14309 4175 14361 4227
rect 14375 4175 14427 4227
rect 14441 4175 14493 4227
rect 14243 4109 14295 4161
rect 14309 4109 14361 4161
rect 14375 4109 14427 4161
rect 14441 4109 14493 4161
rect 14243 4043 14295 4095
rect 14309 4043 14361 4095
rect 14375 4043 14427 4095
rect 14441 4043 14493 4095
rect 14243 3977 14295 4029
rect 14309 3977 14361 4029
rect 14375 3977 14427 4029
rect 14441 3977 14493 4029
rect 14243 3911 14295 3963
rect 14309 3911 14361 3963
rect 14375 3911 14427 3963
rect 14441 3911 14493 3963
rect 14243 3845 14295 3897
rect 14309 3845 14361 3897
rect 14375 3845 14427 3897
rect 14441 3845 14493 3897
rect 14243 3779 14295 3831
rect 14309 3779 14361 3831
rect 14375 3779 14427 3831
rect 14441 3779 14493 3831
rect 14243 3713 14295 3765
rect 14309 3713 14361 3765
rect 14375 3713 14427 3765
rect 14441 3713 14493 3765
rect 14243 3647 14295 3699
rect 14309 3647 14361 3699
rect 14375 3647 14427 3699
rect 14441 3647 14493 3699
rect 580 820 632 872
rect 648 820 700 872
rect 580 754 632 806
rect 648 754 700 806
rect 3716 819 3768 871
rect 3796 819 3848 871
rect 3876 819 3928 871
rect 3716 793 3768 805
rect 3796 793 3848 805
rect 3876 793 3928 805
rect 3716 759 3722 793
rect 3722 759 3756 793
rect 3756 759 3768 793
rect 3796 759 3828 793
rect 3828 759 3848 793
rect 3876 759 3900 793
rect 3900 759 3928 793
rect 3716 753 3768 759
rect 3796 753 3848 759
rect 3876 753 3928 759
rect 580 435 632 487
rect 648 435 700 487
rect 580 369 632 421
rect 648 369 700 421
rect 3716 481 3768 487
rect 3796 481 3848 487
rect 3876 481 3928 487
rect 3716 447 3722 481
rect 3722 447 3756 481
rect 3756 447 3768 481
rect 3796 447 3828 481
rect 3828 447 3848 481
rect 3876 447 3900 481
rect 3900 447 3928 481
rect 3716 435 3768 447
rect 3796 435 3848 447
rect 3876 435 3928 447
rect 3716 369 3768 421
rect 3796 369 3848 421
rect 3876 369 3928 421
rect 284 83 336 135
rect 348 83 400 135
rect 3716 83 3768 135
rect 3796 83 3848 135
rect 3876 83 3928 135
rect 5878 -9157 5930 -9151
rect 5878 -9191 5884 -9157
rect 5884 -9191 5918 -9157
rect 5918 -9191 5930 -9157
rect 5878 -9203 5930 -9191
rect 5878 -9229 5930 -9223
rect 5878 -9263 5884 -9229
rect 5884 -9263 5918 -9229
rect 5918 -9263 5930 -9229
rect 5878 -9275 5930 -9263
rect 5253 -9994 5305 -9942
rect 5328 -9994 5380 -9942
rect 5403 -9994 5455 -9942
rect 5478 -9994 5530 -9942
rect 5553 -9994 5605 -9942
rect 5627 -9994 5679 -9942
rect 5253 -10069 5305 -10017
rect 5328 -10069 5380 -10017
rect 5403 -10069 5455 -10017
rect 5478 -10069 5530 -10017
rect 5553 -10069 5605 -10017
rect 5627 -10069 5679 -10017
rect 5253 -10144 5305 -10092
rect 5328 -10144 5380 -10092
rect 5403 -10144 5455 -10092
rect 5478 -10144 5530 -10092
rect 5553 -10144 5605 -10092
rect 5627 -10144 5679 -10092
rect 5253 -10985 5305 -10933
rect 5328 -10985 5380 -10933
rect 5403 -10985 5455 -10933
rect 5478 -10985 5530 -10933
rect 5553 -10985 5605 -10933
rect 5627 -10985 5679 -10933
rect 5253 -11063 5305 -11011
rect 5328 -11063 5380 -11011
rect 5403 -11063 5455 -11011
rect 5478 -11063 5530 -11011
rect 5553 -11063 5605 -11011
rect 5627 -11063 5679 -11011
<< metal2 >>
tri 14573 16601 14591 16619 se
rect 14591 16610 14647 16619
tri 3147 16549 3199 16601 se
rect 3199 16554 14591 16601
rect 3199 16549 14647 16554
tri 3103 16505 3147 16549 se
rect 3147 16513 3185 16549
tri 3185 16513 3221 16549 nw
tri 14555 16513 14591 16549 ne
rect 14591 16530 14647 16549
rect 3147 16505 3177 16513
tri 3177 16505 3185 16513 nw
rect 2281 16453 2287 16505
rect 2339 16453 2369 16505
rect 2421 16453 2427 16505
tri 3073 16475 3103 16505 se
rect 3103 16475 3147 16505
tri 3147 16475 3177 16505 nw
tri 3051 16453 3073 16475 se
rect 3073 16465 3137 16475
tri 3137 16465 3147 16475 nw
rect 3073 16453 3125 16465
tri 3125 16453 3137 16465 nw
rect 14095 16453 14101 16505
rect 14153 16453 14175 16505
rect 14227 16453 14249 16505
rect 14301 16453 14323 16505
rect 14375 16453 14397 16505
rect 14449 16453 14455 16505
rect 14591 16465 14647 16474
rect 385 16418 437 16424
rect 385 16354 437 16366
rect 385 16296 437 16302
tri 386 16292 390 16296 ne
rect 390 16292 437 16296
tri 390 16276 406 16292 ne
rect 406 16212 437 16292
rect 498 16372 506 16424
rect 558 16372 570 16424
rect 622 16372 628 16424
tri 437 16212 440 16215 sw
rect 406 16204 440 16212
tri 440 16204 448 16212 sw
tri 406 16183 427 16204 ne
rect 427 16183 448 16204
tri 448 16183 469 16204 sw
tri 427 16173 437 16183 ne
rect 437 16173 469 16183
tri 437 16171 439 16173 ne
rect 359 16145 411 16151
rect 359 16081 411 16093
rect 359 16023 411 16029
rect 278 15989 330 15995
rect 278 15925 330 15937
rect 278 15867 330 15873
rect 278 15863 326 15867
tri 326 15863 330 15867 nw
rect 278 15850 313 15863
tri 313 15850 326 15863 nw
rect 278 7873 310 15850
tri 310 15847 313 15850 nw
tri 356 15847 359 15850 se
rect 359 15847 399 16023
tri 399 16011 411 16023 nw
tri 354 15845 356 15847 se
rect 356 15845 399 15847
tri 341 15832 354 15845 se
rect 354 15832 399 15845
tri 338 15829 341 15832 se
rect 341 15829 378 15832
rect 338 7959 378 15829
tri 378 15811 399 15832 nw
tri 437 15800 439 15802 se
rect 439 15800 469 16173
rect 498 16119 628 16372
rect 1932 16372 1938 16424
rect 1990 16372 2002 16424
rect 2054 16372 2062 16424
rect 499 16117 627 16118
rect 740 16292 748 16344
rect 800 16292 812 16344
rect 864 16292 870 16344
rect 740 16119 870 16292
rect 1649 16292 1655 16344
rect 1707 16292 1719 16344
rect 1771 16292 1779 16344
rect 741 16117 869 16118
rect 981 16212 989 16264
rect 1041 16212 1053 16264
rect 1105 16212 1111 16264
rect 981 16119 1111 16212
rect 982 16117 1110 16118
rect 1345 16212 1351 16264
rect 1403 16212 1415 16264
rect 1467 16212 1475 16264
rect 1345 16119 1475 16212
rect 1346 16117 1474 16118
rect 1649 16119 1779 16292
rect 1650 16117 1778 16118
rect 1932 16119 2062 16372
rect 1933 16117 2061 16118
rect 740 15817 870 16117
rect 1345 15817 1475 16117
rect 2162 15989 2214 15995
rect 2162 15925 2214 15937
tri 436 15799 437 15800 se
rect 437 15799 469 15800
tri 434 15797 436 15799 se
rect 436 15797 469 15799
tri 430 15793 434 15797 se
rect 434 15793 469 15797
tri 427 15790 430 15793 se
rect 430 15790 469 15793
tri 406 15769 427 15790 se
rect 427 15769 448 15790
tri 448 15769 469 15790 nw
rect 499 15816 627 15817
rect 498 15793 628 15815
rect 741 15816 869 15817
tri 628 15793 632 15797 sw
tri 736 15793 740 15797 se
rect 740 15793 870 15815
rect 982 15816 1110 15817
tri 870 15793 874 15797 sw
tri 977 15793 981 15797 se
rect 981 15793 1111 15815
rect 406 15763 442 15769
tri 442 15763 448 15769 nw
rect 498 15763 632 15793
tri 632 15763 662 15793 sw
tri 706 15763 736 15793 se
rect 736 15763 874 15793
tri 874 15763 904 15793 sw
tri 947 15763 977 15793 se
rect 977 15763 1111 15793
rect 406 8380 437 15763
tri 437 15758 442 15763 nw
rect 498 15649 1111 15763
rect 1346 15816 1474 15817
rect 1345 15797 1475 15815
rect 1650 15816 1778 15817
tri 1475 15797 1477 15799 sw
tri 1647 15797 1649 15799 se
rect 1649 15797 1779 15815
rect 1933 15816 2061 15817
tri 1779 15797 1781 15799 sw
tri 1930 15797 1932 15799 se
rect 1932 15797 2062 15815
rect 1345 15793 1477 15797
tri 1477 15793 1481 15797 sw
tri 1643 15793 1647 15797 se
rect 1647 15793 1781 15797
tri 1781 15793 1785 15797 sw
tri 1926 15793 1930 15797 se
rect 1930 15793 2062 15797
rect 1345 15763 1481 15793
tri 1481 15763 1511 15793 sw
tri 1613 15763 1643 15793 se
rect 1643 15763 1785 15793
tri 1785 15763 1815 15793 sw
tri 1896 15763 1926 15793 se
rect 1926 15763 2062 15793
rect 1345 15649 2062 15763
tri 609 15615 643 15649 ne
rect 643 15615 819 15649
tri 819 15615 853 15649 nw
tri 1495 15615 1529 15649 ne
rect 1529 15615 1765 15649
tri 1765 15615 1799 15649 nw
tri 643 15597 661 15615 ne
rect 661 15597 801 15615
tri 801 15597 819 15615 nw
tri 1529 15597 1547 15615 ne
rect 1547 15597 1747 15615
tri 1747 15597 1765 15615 nw
tri 661 15589 669 15597 ne
rect 669 14498 799 15597
tri 799 15595 801 15597 nw
tri 1547 15595 1549 15597 ne
rect 1549 15595 1712 15597
tri 1549 15562 1582 15595 ne
tri 799 14498 869 14568 sw
rect 669 14368 1000 14498
tri 800 14298 870 14368 ne
rect 870 13850 1000 14368
rect 1582 14032 1712 15595
tri 1712 15562 1747 15597 nw
tri 2144 15562 2162 15580 se
rect 2162 15562 2214 15873
tri 2140 15558 2144 15562 se
rect 2144 15558 2214 15562
tri 2127 15545 2140 15558 se
rect 2140 15545 2201 15558
tri 2201 15545 2214 15558 nw
tri 2109 15527 2127 15545 se
rect 2127 15527 2183 15545
tri 2183 15527 2201 15545 nw
tri 2095 15513 2109 15527 se
rect 2109 15513 2169 15527
tri 2169 15513 2183 15527 nw
tri 2066 15484 2095 15513 se
rect 2095 15484 2140 15513
tri 2140 15484 2169 15513 nw
tri 2064 15482 2066 15484 se
rect 2066 15482 2117 15484
tri 2043 15461 2064 15482 se
rect 2064 15461 2117 15482
tri 2117 15461 2140 15484 nw
tri 2041 15459 2043 15461 se
rect 2043 15459 2115 15461
tri 2115 15459 2117 15461 nw
tri 2039 15457 2041 15459 se
rect 2041 15457 2113 15459
tri 2113 15457 2115 15459 nw
tri 1992 15410 2039 15457 se
rect 2039 15410 2066 15457
tri 2066 15410 2113 15457 nw
tri 1990 15408 1992 15410 se
rect 1992 15408 2064 15410
tri 2064 15408 2066 15410 nw
tri 1987 15405 1990 15408 se
rect 1990 15405 2064 15408
tri 1976 15394 1987 15405 se
rect 1987 15394 2064 15405
tri 1968 15386 1976 15394 se
rect 1976 15386 2064 15394
tri 1963 15381 1968 15386 se
rect 1968 15381 2064 15386
tri 1936 15354 1963 15381 se
rect 1963 15354 2064 15381
rect 1936 15311 2064 15354
tri 2262 15329 2281 15348 se
rect 2281 15329 2427 16453
tri 3022 16424 3051 16453 se
rect 3051 16440 3112 16453
tri 3112 16440 3125 16453 nw
rect 3051 16424 3096 16440
tri 3096 16424 3112 16440 nw
tri 9829 16424 9845 16440 se
rect 9845 16424 10262 16440
tri 10262 16424 10278 16440 sw
tri 3005 16407 3022 16424 se
rect 3022 16407 3078 16424
tri 3004 16406 3005 16407 se
rect 3005 16406 3078 16407
tri 3078 16406 3096 16424 nw
tri 2999 16401 3004 16406 se
rect 3004 16401 3073 16406
tri 3073 16401 3078 16406 nw
tri 2970 16372 2999 16401 se
rect 2999 16372 3044 16401
tri 3044 16372 3073 16401 nw
rect 3462 16372 3468 16424
rect 3520 16372 3532 16424
rect 3584 16372 3592 16424
tri 2942 16344 2970 16372 se
rect 2970 16344 3016 16372
tri 3016 16344 3044 16372 nw
tri 2931 16333 2942 16344 se
rect 2942 16333 3005 16344
tri 3005 16333 3016 16344 nw
tri 2924 16326 2931 16333 se
rect 2931 16326 3005 16333
tri 2890 16292 2924 16326 se
rect 2924 16292 3005 16326
tri 2875 16277 2890 16292 se
rect 2890 16277 3005 16292
tri 2261 15328 2262 15329 se
rect 2262 15328 2427 15329
tri 2244 15311 2261 15328 se
rect 2261 15311 2427 15328
rect 1936 15259 1942 15311
rect 1994 15259 2006 15311
rect 2058 15259 2064 15311
tri 2213 15280 2244 15311 se
rect 2244 15288 2427 15311
rect 2244 15280 2419 15288
tri 2419 15280 2427 15288 nw
rect 2532 16103 2538 16155
rect 2590 16103 2602 16155
rect 2654 16103 2660 16155
rect 2532 16075 2632 16103
tri 2632 16075 2660 16103 nw
rect 2532 16057 2614 16075
tri 2614 16057 2632 16075 nw
tri 2192 15259 2213 15280 se
rect 2213 15266 2405 15280
tri 2405 15266 2419 15280 nw
rect 2213 15259 2398 15266
tri 2398 15259 2405 15266 nw
tri 2525 15259 2532 15266 se
rect 2532 15259 2584 16057
tri 2584 16027 2614 16057 nw
rect 2875 15797 3005 16277
rect 3179 16292 3185 16344
rect 3237 16292 3249 16344
rect 3301 16292 3309 16344
rect 3179 16171 3309 16292
rect 3462 16171 3592 16372
rect 7748 16372 7754 16424
rect 7806 16372 7818 16424
rect 7870 16372 7878 16424
rect 3895 16292 3960 16344
rect 4012 16292 4024 16344
rect 4076 16292 4088 16344
rect 4140 16292 4152 16344
rect 4204 16292 4216 16344
rect 4268 16292 4274 16344
rect 3610 15943 3616 15995
rect 3668 15943 3680 15995
rect 3732 15943 3738 15995
tri 3005 15797 3007 15799 sw
rect 2875 15793 3007 15797
tri 3007 15793 3011 15797 sw
rect 2875 15763 3011 15793
tri 3011 15763 3041 15793 sw
rect 2875 15649 3305 15763
tri 3088 15615 3122 15649 ne
rect 3122 15615 3305 15649
tri 3122 15597 3140 15615 ne
rect 3140 15597 3305 15615
tri 3140 15562 3175 15597 ne
tri 2148 15215 2192 15259 se
rect 2192 15240 2379 15259
tri 2379 15240 2398 15259 nw
tri 2506 15240 2525 15259 se
rect 2525 15240 2584 15259
rect 2192 15215 2354 15240
tri 2354 15215 2379 15240 nw
tri 2481 15215 2506 15240 se
rect 2506 15215 2584 15240
tri 2584 15215 2609 15240 sw
tri 2096 15163 2148 15215 se
rect 2148 15163 2302 15215
tri 2302 15163 2354 15215 nw
rect 2481 15163 2487 15215
rect 2539 15163 2551 15215
rect 2603 15163 2609 15215
tri 2082 15149 2096 15163 se
rect 2096 15149 2288 15163
tri 2288 15149 2302 15163 nw
tri 2030 15097 2082 15149 se
rect 2082 15097 2236 15149
tri 2236 15097 2288 15149 nw
tri 2011 15078 2030 15097 se
rect 2030 15078 2217 15097
tri 2217 15078 2236 15097 nw
tri 2007 15074 2011 15078 se
rect 2011 15074 2213 15078
tri 2213 15074 2217 15078 nw
tri 1997 15064 2007 15074 se
rect 2007 15064 2203 15074
tri 2203 15064 2213 15074 nw
tri 1945 15012 1997 15064 se
rect 1997 15012 2151 15064
tri 2151 15012 2203 15064 nw
tri 1931 14998 1945 15012 se
rect 1945 14998 2137 15012
tri 2137 14998 2151 15012 nw
tri 1879 14946 1931 14998 se
rect 1931 14946 2085 14998
tri 2085 14946 2137 14998 nw
tri 1861 14928 1879 14946 se
rect 1879 14928 2007 14946
rect 1861 14783 2007 14928
tri 2007 14868 2085 14946 nw
tri 3121 14804 3175 14858 se
rect 3175 14804 3305 15597
rect 3610 15311 3738 15943
rect 3610 15259 3616 15311
rect 3668 15259 3680 15311
rect 3732 15259 3738 15311
tri 3105 14788 3121 14804 se
rect 3121 14788 3289 14804
tri 3289 14788 3305 14804 nw
rect 1913 14731 1955 14783
tri 3053 14736 3105 14788 se
rect 3105 14736 3237 14788
tri 3237 14736 3289 14788 nw
rect 1861 14714 2007 14731
tri 3031 14714 3053 14736 se
rect 3053 14714 3215 14736
tri 3215 14714 3237 14736 nw
rect 1913 14662 1955 14714
tri 2979 14662 3031 14714 se
rect 3031 14662 3163 14714
tri 3163 14662 3215 14714 nw
rect 1861 14645 2007 14662
rect 1913 14593 1955 14645
tri 2957 14640 2979 14662 se
rect 2979 14640 3141 14662
tri 3141 14640 3163 14662 nw
tri 2937 14620 2957 14640 se
rect 2957 14620 3121 14640
tri 3121 14620 3141 14640 nw
rect 1861 14587 2007 14593
tri 2905 14588 2937 14620 se
rect 2937 14588 3089 14620
tri 3089 14588 3121 14620 nw
tri 2904 14587 2905 14588 se
rect 2905 14587 2937 14588
tri 2782 14465 2904 14587 se
rect 2904 14465 2937 14587
rect 2782 14436 2937 14465
tri 2937 14436 3089 14588 nw
tri 1712 14032 1766 14086 sw
tri 1582 13911 1703 14032 ne
rect 1703 13911 1766 14032
tri 1766 13911 1887 14032 sw
tri 1703 13857 1757 13911 ne
rect 1757 13857 1887 13911
tri 1887 13857 1941 13911 sw
tri 1757 13853 1761 13857 ne
rect 1761 13853 2226 13857
rect 870 13798 876 13850
rect 928 13798 942 13850
rect 994 13798 1000 13850
tri 1761 13805 1809 13853 ne
rect 1809 13805 2226 13853
rect 2278 13805 2292 13857
rect 2344 13805 2350 13857
tri 1809 13798 1816 13805 ne
rect 1816 13798 2350 13805
rect 870 13786 1000 13798
tri 1816 13786 1828 13798 ne
rect 1828 13786 2350 13798
rect 870 13734 876 13786
rect 928 13734 942 13786
rect 994 13734 1000 13786
tri 1828 13779 1835 13786 ne
rect 1835 13779 2350 13786
rect 870 13727 1000 13734
tri 1835 13727 1887 13779 ne
rect 1887 13727 2226 13779
rect 2278 13727 2292 13779
rect 2344 13727 2350 13779
rect 2782 13850 2912 14436
tri 2912 14411 2937 14436 nw
rect 2782 13798 2788 13850
rect 2840 13798 2854 13850
rect 2906 13798 2912 13850
rect 2782 13786 2912 13798
rect 2782 13734 2788 13786
rect 2840 13734 2854 13786
rect 2906 13734 2912 13786
rect 2782 13727 2912 13734
rect 3895 13850 4274 16292
rect 7318 16292 7324 16344
rect 7376 16292 7388 16344
rect 7440 16292 7448 16344
rect 5732 16212 5738 16264
rect 5790 16212 5827 16264
rect 5879 16212 5916 16264
rect 5968 16212 6005 16264
rect 6057 16212 6063 16264
rect 4433 15985 5496 15986
rect 4433 15933 4439 15985
rect 4491 15933 4506 15985
rect 4558 15933 4573 15985
rect 4625 15933 4640 15985
rect 4692 15933 4707 15985
rect 4759 15933 4774 15985
rect 4826 15933 4841 15985
rect 4893 15933 4908 15985
rect 4960 15933 4975 15985
rect 5027 15933 5042 15985
rect 5094 15933 5108 15985
rect 5160 15933 5174 15985
rect 5226 15933 5240 15985
rect 5292 15933 5306 15985
rect 5358 15933 5372 15985
rect 5424 15933 5438 15985
rect 5490 15933 5496 15985
rect 4433 15915 5496 15933
rect 4433 15863 4439 15915
rect 4491 15863 4506 15915
rect 4558 15863 4573 15915
rect 4625 15863 4640 15915
rect 4692 15863 4707 15915
rect 4759 15863 4774 15915
rect 4826 15863 4841 15915
rect 4893 15863 4908 15915
rect 4960 15863 4975 15915
rect 5027 15863 5042 15915
rect 5094 15863 5108 15915
rect 5160 15863 5174 15915
rect 5226 15863 5240 15915
rect 5292 15863 5306 15915
rect 5358 15863 5372 15915
rect 5424 15863 5438 15915
rect 5490 15863 5496 15915
rect 4433 15845 5496 15863
rect 4433 15793 4439 15845
rect 4491 15793 4506 15845
rect 4558 15793 4573 15845
rect 4625 15793 4640 15845
rect 4692 15793 4707 15845
rect 4759 15793 4774 15845
rect 4826 15793 4841 15845
rect 4893 15793 4908 15845
rect 4960 15793 4975 15845
rect 5027 15793 5042 15845
rect 5094 15793 5108 15845
rect 5160 15793 5174 15845
rect 5226 15793 5240 15845
rect 5292 15793 5306 15845
rect 5358 15793 5372 15845
rect 5424 15793 5438 15845
rect 5490 15793 5496 15845
rect 4433 15743 5496 15793
rect 4433 15691 4439 15743
rect 4491 15691 4506 15743
rect 4558 15691 4573 15743
rect 4625 15691 4640 15743
rect 4692 15691 4707 15743
rect 4759 15691 4774 15743
rect 4826 15691 4841 15743
rect 4893 15691 4908 15743
rect 4960 15691 4975 15743
rect 5027 15691 5042 15743
rect 5094 15691 5108 15743
rect 5160 15691 5174 15743
rect 5226 15691 5240 15743
rect 5292 15691 5306 15743
rect 5358 15691 5372 15743
rect 5424 15691 5438 15743
rect 5490 15691 5496 15743
rect 4582 15513 5119 15527
rect 4582 15461 4591 15513
rect 4643 15461 4658 15513
rect 4710 15461 4725 15513
rect 4777 15461 4792 15513
rect 4844 15461 4859 15513
rect 4911 15461 4926 15513
rect 4978 15461 4993 15513
rect 5045 15461 5059 15513
rect 5111 15461 5119 15513
rect 4582 15388 5119 15461
rect 4582 15381 4605 15388
rect 4661 15381 4710 15388
rect 4766 15381 4815 15388
rect 4871 15381 4919 15388
rect 4975 15381 5023 15388
rect 4582 15329 4602 15381
rect 4661 15332 4687 15381
rect 4766 15332 4772 15381
rect 4908 15332 4919 15381
rect 4992 15332 5023 15381
rect 5079 15332 5119 15388
rect 4654 15329 4687 15332
rect 4739 15329 4772 15332
rect 4824 15329 4856 15332
rect 4908 15329 4940 15332
rect 4992 15329 5024 15332
rect 5076 15329 5119 15332
rect 4582 15268 5119 15329
rect 4582 15265 4605 15268
rect 4661 15265 4710 15268
rect 4766 15265 4815 15268
rect 4871 15265 4919 15268
rect 4975 15265 5023 15268
rect 4582 15213 4602 15265
rect 4661 15213 4687 15265
rect 4766 15213 4772 15265
rect 4908 15213 4919 15265
rect 4992 15213 5023 15265
rect 4582 15212 4605 15213
rect 4661 15212 4710 15213
rect 4766 15212 4815 15213
rect 4871 15212 4919 15213
rect 4975 15212 5023 15213
rect 5079 15212 5119 15268
rect 4582 15149 5119 15212
rect 4582 15097 4602 15149
rect 4654 15148 4687 15149
rect 4739 15148 4772 15149
rect 4824 15148 4856 15149
rect 4908 15148 4940 15149
rect 4992 15148 5024 15149
rect 5076 15148 5119 15149
rect 4661 15097 4687 15148
rect 4766 15097 4772 15148
rect 4908 15097 4919 15148
rect 4992 15097 5023 15148
rect 4582 15092 4605 15097
rect 4661 15092 4710 15097
rect 4766 15092 4815 15097
rect 4871 15092 4919 15097
rect 4975 15092 5023 15097
rect 5079 15092 5119 15148
rect 4582 15090 5119 15092
rect 3895 13798 3901 13850
rect 3953 13798 3980 13850
rect 4032 13798 4059 13850
rect 4111 13798 4138 13850
rect 4190 13798 4216 13850
rect 4268 13798 4274 13850
rect 3895 13786 4274 13798
rect 3895 13734 3901 13786
rect 3953 13734 3980 13786
rect 4032 13734 4059 13786
rect 4111 13734 4138 13786
rect 4190 13734 4216 13786
rect 4268 13734 4274 13786
rect 3895 13727 4274 13734
rect 5732 13857 6063 16212
rect 6888 16212 6894 16264
rect 6946 16212 6958 16264
rect 7010 16212 7018 16264
rect 6888 16119 7018 16212
rect 6889 16117 7017 16118
rect 7318 16119 7448 16292
rect 7319 16117 7447 16118
rect 7748 16119 7878 16372
rect 9450 16372 9456 16424
rect 9508 16372 9520 16424
rect 9572 16372 9580 16424
tri 9811 16406 9829 16424 se
rect 9829 16406 10278 16424
tri 10278 16406 10296 16424 sw
tri 9793 16388 9811 16406 se
rect 9811 16388 10296 16406
tri 10296 16388 10314 16406 sw
tri 9777 16372 9793 16388 se
rect 9793 16372 9851 16388
tri 9851 16372 9867 16388 nw
tri 10240 16372 10256 16388 ne
rect 10256 16372 10314 16388
tri 10314 16372 10330 16388 sw
rect 10930 16372 10936 16424
rect 10988 16372 11000 16424
rect 11052 16372 11060 16424
rect 9020 16292 9026 16344
rect 9078 16292 9090 16344
rect 9142 16292 9150 16344
rect 7749 16117 7877 16118
rect 8590 16212 8596 16264
rect 8648 16212 8660 16264
rect 8712 16212 8720 16264
rect 8590 16119 8720 16212
rect 8591 16117 8719 16118
rect 9020 16119 9150 16292
rect 9021 16117 9149 16118
rect 9450 16119 9580 16372
tri 9759 16354 9777 16372 se
rect 9777 16354 9823 16372
tri 9749 16344 9759 16354 se
rect 9759 16344 9823 16354
tri 9823 16344 9851 16372 nw
tri 10256 16344 10284 16372 ne
rect 10284 16351 10330 16372
tri 10330 16351 10351 16372 sw
rect 10284 16344 10351 16351
tri 9731 16326 9749 16344 se
rect 9749 16329 9808 16344
tri 9808 16329 9823 16344 nw
tri 10284 16329 10299 16344 ne
rect 9749 16326 9805 16329
tri 9805 16326 9808 16329 nw
tri 9719 16314 9731 16326 se
rect 9731 16314 9793 16326
tri 9793 16314 9805 16326 nw
rect 9451 16117 9579 16118
tri 9707 16302 9719 16314 se
rect 9719 16302 9771 16314
rect 9707 16292 9771 16302
tri 9771 16292 9793 16314 nw
rect 6192 15985 6817 15986
rect 6192 15933 6198 15985
rect 6250 15933 6269 15985
rect 6321 15933 6339 15985
rect 6391 15933 6409 15985
rect 6461 15933 6479 15985
rect 6531 15933 6549 15985
rect 6601 15933 6619 15985
rect 6671 15933 6689 15985
rect 6741 15933 6759 15985
rect 6811 15933 6817 15985
rect 6192 15915 6817 15933
rect 6192 15863 6198 15915
rect 6250 15863 6269 15915
rect 6321 15863 6339 15915
rect 6391 15863 6409 15915
rect 6461 15863 6479 15915
rect 6531 15863 6549 15915
rect 6601 15863 6619 15915
rect 6671 15863 6689 15915
rect 6741 15863 6759 15915
rect 6811 15863 6817 15915
rect 6192 15845 6817 15863
rect 6192 15793 6198 15845
rect 6250 15793 6269 15845
rect 6321 15793 6339 15845
rect 6391 15793 6409 15845
rect 6461 15793 6479 15845
rect 6531 15793 6549 15845
rect 6601 15793 6619 15845
rect 6671 15793 6689 15845
rect 6741 15793 6759 15845
rect 6811 15793 6817 15845
rect 7318 15817 7448 16117
rect 8183 16023 8191 16075
rect 8243 16023 8255 16075
rect 8307 16023 8313 16075
rect 6192 15743 6817 15793
rect 6192 15691 6198 15743
rect 6250 15691 6269 15743
rect 6321 15691 6339 15743
rect 6391 15691 6409 15743
rect 6461 15691 6479 15743
rect 6531 15691 6549 15743
rect 6601 15691 6619 15743
rect 6671 15691 6689 15743
rect 6741 15691 6759 15743
rect 6811 15691 6817 15743
rect 6889 15816 7017 15817
rect 6888 15798 7018 15815
rect 7319 15816 7447 15817
tri 7018 15798 7019 15799 sw
tri 7317 15798 7318 15799 se
rect 7318 15798 7448 15815
rect 7749 15816 7877 15817
tri 7448 15798 7449 15799 sw
tri 7747 15798 7748 15799 se
rect 7748 15798 7878 15815
rect 6888 15797 7019 15798
tri 7019 15797 7020 15798 sw
tri 7316 15797 7317 15798 se
rect 7317 15797 7449 15798
tri 7449 15797 7450 15798 sw
tri 7746 15797 7747 15798 se
rect 7747 15797 7878 15798
rect 6888 15763 7020 15797
tri 7020 15763 7054 15797 sw
tri 7282 15763 7316 15797 se
rect 7316 15763 7450 15797
tri 7450 15763 7484 15797 sw
tri 7712 15763 7746 15797 se
rect 7746 15763 7878 15797
rect 6888 15649 7878 15763
tri 7430 15615 7464 15649 ne
rect 7464 15615 7878 15649
tri 7464 15605 7474 15615 ne
rect 7474 15605 7878 15615
tri 7474 15597 7482 15605 ne
rect 7482 15597 7878 15605
tri 7482 15545 7534 15597 ne
rect 7534 15545 7878 15597
tri 7534 15537 7542 15545 ne
rect 7542 15537 7878 15545
tri 7542 15531 7548 15537 ne
rect 7548 15531 7872 15537
tri 7872 15531 7878 15537 nw
tri 7548 15527 7552 15531 ne
rect 7552 15527 7872 15531
tri 7552 15475 7604 15527 ne
rect 7604 15475 7872 15527
tri 7604 15459 7620 15475 ne
rect 7620 15459 7872 15475
tri 7620 15457 7622 15459 ne
rect 7622 15457 7872 15459
tri 7622 15405 7674 15457 ne
rect 7674 15405 7872 15457
tri 7674 15394 7685 15405 ne
rect 7685 15394 7872 15405
tri 7685 15386 7693 15394 ne
rect 7693 15386 7872 15394
tri 7693 15337 7742 15386 ne
tri 6063 13857 6192 13986 sw
rect 7742 13857 7872 15386
rect 8183 15311 8313 16023
rect 9020 15817 9150 16117
rect 8591 15816 8719 15817
rect 8590 15798 8720 15815
rect 9021 15816 9149 15817
tri 8720 15798 8721 15799 sw
tri 9019 15798 9020 15799 se
rect 9020 15798 9150 15815
rect 9451 15816 9579 15817
tri 9150 15798 9151 15799 sw
tri 9449 15798 9450 15799 se
rect 9450 15798 9580 15815
rect 8590 15797 8721 15798
tri 8721 15797 8722 15798 sw
tri 9018 15797 9019 15798 se
rect 9019 15797 9151 15798
tri 9151 15797 9152 15798 sw
tri 9448 15797 9449 15798 se
rect 9449 15797 9580 15798
rect 8590 15763 8722 15797
tri 8722 15763 8756 15797 sw
tri 8984 15763 9018 15797 se
rect 9018 15763 9152 15797
tri 9152 15763 9186 15797 sw
tri 9414 15763 9448 15797 se
rect 9448 15763 9580 15797
rect 8590 15689 9580 15763
tri 8590 15685 8594 15689 ne
rect 8594 15685 9017 15689
tri 9017 15685 9021 15689 nw
tri 8594 15667 8612 15685 ne
rect 8612 15667 8999 15685
tri 8999 15667 9017 15685 nw
tri 8612 15649 8630 15667 ne
rect 8630 15649 8981 15667
tri 8981 15649 8999 15667 nw
tri 8630 15615 8664 15649 ne
rect 8664 15615 8947 15649
tri 8947 15615 8981 15649 nw
tri 8664 15605 8674 15615 ne
rect 8183 15259 8189 15311
rect 8241 15259 8255 15311
rect 8307 15259 8313 15311
rect 5732 13851 6192 13857
tri 6192 13851 6198 13857 sw
rect 5732 13799 6194 13851
rect 6246 13799 6259 13851
rect 6311 13799 6324 13851
rect 6376 13799 6389 13851
rect 6441 13799 6453 13851
rect 6505 13799 6517 13851
rect 6569 13799 6581 13851
rect 6633 13799 6645 13851
rect 6697 13799 6709 13851
rect 6761 13799 6773 13851
rect 6825 13799 6837 13851
rect 6889 13799 6895 13851
rect 5732 13779 6895 13799
rect 5732 13727 6194 13779
rect 6246 13727 6259 13779
rect 6311 13727 6324 13779
rect 6376 13727 6389 13779
rect 6441 13727 6453 13779
rect 6505 13727 6517 13779
rect 6569 13727 6581 13779
rect 6633 13727 6645 13779
rect 6697 13727 6709 13779
rect 6761 13727 6773 13779
rect 6825 13727 6837 13779
rect 6889 13727 6895 13779
rect 7742 13805 7748 13857
rect 7800 13805 7814 13857
rect 7866 13805 7872 13857
rect 7742 13779 7872 13805
rect 7742 13727 7748 13779
rect 7800 13727 7814 13779
rect 7866 13727 7872 13779
rect 8674 13853 8931 15615
tri 8931 15599 8947 15615 nw
rect 9043 15332 9052 15388
rect 9108 15332 9169 15388
rect 9225 15332 9286 15388
rect 9342 15332 9351 15388
rect 9043 15268 9351 15332
rect 9043 15212 9052 15268
rect 9108 15212 9169 15268
rect 9225 15212 9286 15268
rect 9342 15212 9351 15268
tri 9704 15259 9707 15262 se
rect 9707 15259 9759 16292
tri 9759 16280 9771 16292 nw
rect 10070 16212 10076 16264
rect 10128 16212 10140 16264
rect 10192 16212 10200 16264
rect 10070 16119 10200 16212
rect 10071 16117 10199 16118
tri 10293 16103 10299 16109 se
rect 10299 16103 10351 16344
rect 10500 16292 10506 16344
rect 10558 16292 10570 16344
rect 10622 16292 10630 16344
rect 10500 16119 10630 16292
rect 10501 16117 10629 16118
rect 10930 16119 11060 16372
rect 12273 16372 12279 16424
rect 12331 16372 12343 16424
rect 12395 16372 12403 16424
rect 11843 16292 11849 16344
rect 11901 16292 11913 16344
rect 11965 16292 11973 16344
rect 10931 16117 11059 16118
rect 11413 16212 11419 16264
rect 11471 16212 11483 16264
rect 11535 16212 11543 16264
rect 11413 16119 11543 16212
rect 11414 16117 11542 16118
rect 11843 16119 11973 16292
rect 11844 16117 11972 16118
rect 12273 16119 12403 16372
rect 13707 16372 13713 16424
rect 13765 16372 13777 16424
rect 13829 16372 13837 16424
rect 13277 16292 13283 16344
rect 13335 16292 13347 16344
rect 13399 16292 13407 16344
rect 12274 16117 12402 16118
rect 12847 16212 12853 16264
rect 12905 16212 12917 16264
rect 12969 16212 12977 16264
rect 12847 16119 12977 16212
rect 12848 16117 12976 16118
rect 13277 16119 13407 16292
rect 13278 16117 13406 16118
rect 13707 16119 13837 16372
rect 13708 16117 13836 16118
tri 10351 16103 10352 16104 sw
tri 10265 16075 10293 16103 se
rect 10293 16075 10352 16103
tri 10352 16075 10380 16103 sw
rect 9855 16023 9861 16075
rect 9913 16023 9925 16075
rect 9977 16023 9985 16075
rect 10252 16023 10258 16075
rect 10310 16023 10322 16075
rect 10374 16023 10380 16075
rect 9855 15311 9985 16023
rect 10500 15817 10630 16117
rect 11843 15817 11973 16117
rect 12534 15980 12586 15986
rect 12534 15915 12586 15928
rect 12534 15850 12586 15863
rect 10071 15816 10199 15817
rect 10070 15798 10200 15815
rect 10501 15816 10629 15817
tri 10200 15798 10201 15799 sw
tri 10499 15798 10500 15799 se
rect 10500 15798 10630 15815
rect 10931 15816 11059 15817
tri 10630 15798 10631 15799 sw
tri 10929 15798 10930 15799 se
rect 10930 15798 11060 15815
rect 10070 15797 10201 15798
tri 10201 15797 10202 15798 sw
tri 10498 15797 10499 15798 se
rect 10499 15797 10631 15798
tri 10631 15797 10632 15798 sw
tri 10928 15797 10929 15798 se
rect 10929 15797 11060 15798
rect 10070 15763 10202 15797
tri 10202 15763 10236 15797 sw
tri 10464 15763 10498 15797 se
rect 10498 15763 10632 15797
tri 10632 15763 10666 15797 sw
tri 10894 15763 10928 15797 se
rect 10928 15763 11060 15797
rect 10070 15649 11060 15763
rect 11414 15816 11542 15817
rect 11413 15798 11543 15815
rect 11844 15816 11972 15817
tri 11543 15798 11544 15799 sw
tri 11842 15798 11843 15799 se
rect 11843 15798 11973 15815
rect 12274 15816 12402 15817
tri 11973 15798 11974 15799 sw
tri 12272 15798 12273 15799 se
rect 12273 15798 12403 15815
rect 11413 15797 11544 15798
tri 11544 15797 11545 15798 sw
tri 11841 15797 11842 15798 se
rect 11842 15797 11974 15798
tri 11974 15797 11975 15798 sw
tri 12271 15797 12272 15798 se
rect 12272 15797 12403 15798
rect 11413 15763 11545 15797
tri 11545 15763 11579 15797 sw
tri 11807 15763 11841 15797 se
rect 11841 15763 11975 15797
tri 11975 15763 12009 15797 sw
tri 12237 15763 12271 15797 se
rect 12271 15763 12403 15797
rect 11413 15649 12403 15763
rect 13707 15817 13837 16117
rect 12534 15737 12586 15798
rect 12534 15667 12586 15685
tri 10167 15615 10201 15649 ne
rect 10201 15615 10919 15649
tri 10919 15615 10953 15649 nw
tri 11510 15615 11544 15649 ne
rect 11544 15615 12262 15649
tri 12262 15615 12296 15649 nw
rect 12848 15816 12976 15817
rect 12847 15797 12977 15815
rect 13278 15816 13406 15817
tri 12977 15797 12979 15799 sw
tri 13275 15797 13277 15799 se
rect 13277 15797 13407 15815
rect 13708 15816 13836 15817
tri 13407 15797 13409 15799 sw
tri 13705 15797 13707 15799 se
rect 13707 15797 13837 15815
rect 12847 15763 12979 15797
tri 12979 15763 13013 15797 sw
tri 13241 15763 13275 15797 se
rect 13275 15763 13409 15797
tri 13409 15763 13443 15797 sw
tri 13671 15763 13705 15797 se
rect 13705 15763 13837 15797
rect 12847 15649 13837 15763
rect 14095 15985 14455 16453
rect 14940 16372 14946 16424
rect 14998 16372 15010 16424
rect 15062 16372 15068 16424
tri 15000 16344 15028 16372 ne
rect 14860 16292 14866 16344
rect 14918 16292 14930 16344
rect 14982 16292 14988 16344
tri 14920 16264 14948 16292 ne
rect 14780 16212 14786 16264
rect 14838 16212 14850 16264
rect 14902 16212 14908 16264
tri 14840 16184 14868 16212 ne
rect 14700 16103 14706 16155
rect 14758 16103 14770 16155
rect 14822 16103 14828 16155
tri 14760 16075 14788 16103 ne
rect 14620 16023 14626 16075
rect 14678 16023 14690 16075
rect 14742 16023 14748 16075
tri 14674 15989 14708 16023 ne
rect 14095 15933 14103 15985
rect 14155 15933 14201 15985
rect 14253 15933 14298 15985
rect 14350 15933 14395 15985
rect 14447 15933 14455 15985
rect 14095 15917 14455 15933
rect 14095 15865 14103 15917
rect 14155 15865 14201 15917
rect 14253 15865 14298 15917
rect 14350 15865 14395 15917
rect 14447 15865 14455 15917
rect 14095 15849 14455 15865
rect 14095 15797 14103 15849
rect 14155 15797 14201 15849
rect 14253 15797 14298 15849
rect 14350 15797 14395 15849
rect 14447 15797 14455 15849
tri 10201 15597 10219 15615 ne
rect 10219 15597 10901 15615
tri 10901 15597 10919 15615 nw
tri 11544 15597 11562 15615 ne
rect 11562 15597 12244 15615
tri 12244 15597 12262 15615 nw
rect 12534 15597 12586 15615
tri 10219 15545 10271 15597 ne
rect 10271 15545 10849 15597
tri 10849 15545 10901 15597 nw
tri 11562 15545 11614 15597 ne
rect 11614 15545 12192 15597
tri 12192 15545 12244 15597 nw
tri 10271 15527 10289 15545 ne
rect 10289 15527 10831 15545
tri 10831 15527 10849 15545 nw
tri 11614 15527 11632 15545 ne
rect 11632 15527 12174 15545
tri 12174 15527 12192 15545 nw
rect 12534 15527 12586 15545
tri 12970 15543 13076 15649 ne
rect 13076 15543 13598 15649
tri 13598 15543 13704 15649 nw
tri 10289 15517 10299 15527 ne
rect 9855 15259 9861 15311
rect 9913 15259 9927 15311
rect 9979 15259 9985 15311
tri 9689 15244 9704 15259 se
rect 9704 15244 9759 15259
rect 9043 15148 9351 15212
tri 9660 15215 9689 15244 se
rect 9689 15215 9759 15244
tri 9759 15215 9788 15244 sw
rect 9660 15163 9666 15215
rect 9718 15163 9730 15215
rect 9782 15163 9788 15215
rect 9043 15092 9052 15148
rect 9108 15092 9169 15148
rect 9225 15092 9286 15148
rect 9342 15092 9351 15148
rect 8674 13801 8680 13853
rect 8732 13801 8745 13853
rect 8797 13801 8809 13853
rect 8861 13801 8873 13853
rect 8925 13801 8931 13853
rect 8674 13779 8931 13801
rect 8674 13727 8680 13779
rect 8732 13727 8745 13779
rect 8797 13727 8809 13779
rect 8861 13727 8873 13779
rect 8925 13727 8931 13779
rect 10299 13821 10821 15527
tri 10821 15517 10831 15527 nw
tri 11632 15517 11642 15527 ne
rect 11642 15517 12164 15527
tri 12164 15517 12174 15527 nw
tri 11642 15475 11684 15517 ne
rect 11684 15475 12164 15517
tri 11684 15459 11700 15475 ne
rect 11700 15459 12164 15475
tri 11700 15457 11702 15459 ne
rect 11702 15457 12164 15459
tri 11702 15449 11710 15457 ne
rect 10299 13769 10305 13821
rect 10357 13769 10371 13821
rect 10423 13769 10437 13821
rect 10489 13769 10503 13821
rect 10555 13769 10568 13821
rect 10620 13769 10633 13821
rect 10685 13769 10698 13821
rect 10750 13769 10763 13821
rect 10815 13769 10821 13821
rect 10299 13738 10821 13769
rect 11710 13820 12164 15457
tri 13076 15517 13102 15543 ne
rect 13102 15517 13598 15543
tri 13102 15487 13132 15517 ne
rect 12534 15457 12586 15475
rect 12534 15386 12586 15405
rect 12534 15328 12586 15334
rect 11710 13768 11716 13820
rect 11768 13768 11781 13820
rect 11833 13768 11846 13820
rect 11898 13768 11911 13820
rect 11963 13768 11976 13820
rect 12028 13768 12041 13820
rect 12093 13768 12106 13820
rect 12158 13768 12164 13820
rect 11710 13737 12164 13768
rect 13132 13857 13598 15517
rect 14095 15459 14455 15797
rect 14095 15407 14101 15459
rect 14153 15407 14175 15459
rect 14227 15407 14249 15459
rect 14301 15407 14323 15459
rect 14375 15407 14397 15459
rect 14449 15407 14455 15459
rect 14095 15394 14455 15407
rect 14095 15342 14101 15394
rect 14153 15342 14175 15394
rect 14227 15342 14249 15394
rect 14301 15342 14323 15394
rect 14375 15342 14397 15394
rect 14449 15342 14455 15394
rect 14095 15328 14455 15342
rect 14095 15276 14101 15328
rect 14153 15276 14175 15328
rect 14227 15276 14249 15328
rect 14301 15276 14323 15328
rect 14375 15276 14397 15328
rect 14449 15276 14455 15328
rect 14095 15262 14455 15276
rect 14095 15210 14101 15262
rect 14153 15210 14175 15262
rect 14227 15210 14249 15262
rect 14301 15210 14323 15262
rect 14375 15210 14397 15262
rect 14449 15210 14455 15262
rect 14095 15196 14455 15210
rect 14095 15144 14101 15196
rect 14153 15144 14175 15196
rect 14227 15144 14249 15196
rect 14301 15144 14323 15196
rect 14375 15144 14397 15196
rect 14449 15144 14455 15196
rect 14095 15130 14455 15144
rect 14095 15078 14101 15130
rect 14153 15078 14175 15130
rect 14227 15078 14249 15130
rect 14301 15078 14323 15130
rect 14375 15078 14397 15130
rect 14449 15078 14455 15130
rect 14095 15064 14455 15078
rect 14095 15012 14101 15064
rect 14153 15012 14175 15064
rect 14227 15012 14249 15064
rect 14301 15012 14323 15064
rect 14375 15012 14397 15064
rect 14449 15012 14455 15064
rect 14095 14998 14455 15012
rect 14095 14946 14101 14998
rect 14153 14946 14175 14998
rect 14227 14946 14249 14998
rect 14301 14946 14323 14998
rect 14375 14946 14397 14998
rect 14449 14946 14455 14998
rect 14095 14788 14455 14946
rect 14095 14736 14101 14788
rect 14153 14736 14175 14788
rect 14227 14736 14249 14788
rect 14301 14736 14323 14788
rect 14375 14736 14397 14788
rect 14449 14736 14455 14788
rect 14095 14714 14455 14736
rect 14095 14662 14101 14714
rect 14153 14662 14175 14714
rect 14227 14662 14249 14714
rect 14301 14662 14323 14714
rect 14375 14662 14397 14714
rect 14449 14662 14455 14714
rect 14095 14640 14455 14662
rect 14095 14588 14101 14640
rect 14153 14588 14175 14640
rect 14227 14588 14249 14640
rect 14301 14588 14323 14640
rect 14375 14588 14397 14640
rect 14449 14588 14455 14640
rect 14095 14587 14455 14588
rect 13132 13805 13138 13857
rect 13190 13805 13205 13857
rect 13257 13805 13272 13857
rect 13324 13805 13339 13857
rect 13391 13805 13406 13857
rect 13458 13805 13473 13857
rect 13525 13805 13540 13857
rect 13592 13805 13598 13857
rect 13132 13779 13598 13805
rect 13132 13727 13138 13779
rect 13190 13727 13205 13779
rect 13257 13727 13272 13779
rect 13324 13727 13339 13779
rect 13391 13727 13406 13779
rect 13458 13727 13473 13779
rect 13525 13727 13540 13779
rect 13592 13727 13598 13779
rect 4395 12316 7294 13416
rect 10594 10828 12901 11953
rect 535 10030 970 10031
rect 535 9978 541 10030
rect 593 9978 616 10030
rect 668 9978 690 10030
rect 742 9978 764 10030
rect 816 9978 838 10030
rect 890 9978 912 10030
rect 964 9978 970 10030
rect 535 9956 970 9978
rect 535 9904 541 9956
rect 593 9904 616 9956
rect 668 9904 690 9956
rect 742 9904 764 9956
rect 816 9904 838 9956
rect 890 9904 912 9956
rect 964 9904 970 9956
rect 535 9882 970 9904
rect 535 9830 541 9882
rect 593 9830 616 9882
rect 668 9830 690 9882
rect 742 9830 764 9882
rect 816 9830 838 9882
rect 890 9830 912 9882
rect 964 9830 970 9882
rect 535 8827 970 9830
rect 14240 9460 14652 9466
rect 14292 9408 14312 9460
rect 14364 9408 14384 9460
rect 14436 9408 14456 9460
rect 14508 9408 14528 9460
rect 14580 9408 14600 9460
rect 14240 9395 14652 9408
rect 535 8775 541 8827
rect 593 8775 616 8827
rect 668 8775 690 8827
rect 742 8775 764 8827
rect 816 8775 838 8827
rect 890 8775 912 8827
rect 964 8775 970 8827
rect 535 8751 970 8775
rect 535 8699 541 8751
rect 593 8699 616 8751
rect 668 8699 690 8751
rect 742 8699 764 8751
rect 816 8699 838 8751
rect 890 8699 912 8751
rect 964 8699 970 8751
rect 535 8670 970 8699
rect 535 8618 842 8670
rect 894 8618 912 8670
rect 964 8618 970 8670
tri 437 8380 458 8401 sw
rect 406 8359 458 8380
rect 406 8295 458 8307
rect 406 8235 458 8243
tri 378 7959 383 7964 sw
rect 338 7945 383 7959
tri 383 7945 397 7959 sw
rect 338 7943 397 7945
tri 397 7943 399 7945 sw
rect 338 7942 399 7943
tri 399 7942 400 7943 sw
rect 338 7913 400 7942
tri 338 7891 360 7913 ne
tri 310 7873 314 7877 sw
rect 278 7857 314 7873
tri 314 7857 330 7873 sw
rect 278 7851 330 7857
rect 278 7785 330 7799
rect 278 7718 330 7733
rect 278 7651 330 7666
rect 278 7584 330 7599
rect 278 7526 330 7532
rect 278 135 310 7526
tri 310 7509 327 7526 nw
tri 338 7347 360 7369 se
rect 360 7347 400 7913
rect 338 7338 400 7347
rect 338 6880 378 7338
tri 378 7316 400 7338 nw
tri 435 7071 535 7171 se
rect 535 7071 970 8618
rect 12252 9359 12622 9360
rect 12252 9307 12258 9359
rect 12310 9307 12335 9359
rect 12387 9307 12412 9359
rect 12464 9307 12488 9359
rect 12540 9307 12564 9359
rect 12616 9307 12622 9359
rect 12252 9271 12622 9307
rect 12252 9219 12258 9271
rect 12310 9219 12335 9271
rect 12387 9219 12412 9271
rect 12464 9219 12488 9271
rect 12540 9219 12564 9271
rect 12616 9219 12622 9271
rect 12252 9183 12622 9219
rect 12252 9131 12258 9183
rect 12310 9131 12335 9183
rect 12387 9131 12412 9183
rect 12464 9131 12488 9183
rect 12540 9131 12564 9183
rect 12616 9131 12622 9183
rect 10800 8281 11156 8287
rect 10852 8229 10876 8281
rect 10928 8229 10952 8281
rect 11004 8229 11028 8281
rect 11080 8229 11104 8281
rect 10800 8214 11156 8229
rect 10852 8162 10876 8214
rect 10928 8162 10952 8214
rect 11004 8162 11028 8214
rect 11080 8162 11104 8214
rect 10800 8147 11156 8162
rect 10852 8095 10876 8147
rect 10928 8095 10952 8147
rect 11004 8095 11028 8147
rect 11080 8095 11104 8147
rect 10800 8079 11156 8095
rect 10852 8027 10876 8079
rect 10928 8027 10952 8079
rect 11004 8027 11028 8079
rect 11080 8027 11104 8079
rect 10800 8011 11156 8027
rect 10852 7959 10876 8011
rect 10928 7959 10952 8011
rect 11004 7959 11028 8011
rect 11080 7959 11104 8011
rect 10800 7943 11156 7959
rect 10852 7891 10876 7943
rect 10928 7891 10952 7943
rect 11004 7891 11028 7943
rect 11080 7891 11104 7943
rect 10800 7561 11156 7891
rect 12252 8281 12622 9131
rect 12252 8229 12255 8281
rect 12307 8229 12333 8281
rect 12385 8229 12411 8281
rect 12463 8229 12489 8281
rect 12541 8229 12567 8281
rect 12619 8229 12622 8281
rect 12252 8210 12622 8229
rect 12252 8158 12255 8210
rect 12307 8158 12333 8210
rect 12385 8158 12411 8210
rect 12463 8158 12489 8210
rect 12541 8158 12567 8210
rect 12619 8158 12622 8210
rect 12252 8139 12622 8158
rect 12252 8087 12255 8139
rect 12307 8087 12333 8139
rect 12385 8087 12411 8139
rect 12463 8087 12489 8139
rect 12541 8087 12567 8139
rect 12619 8087 12622 8139
rect 12252 8068 12622 8087
rect 12252 8016 12255 8068
rect 12307 8016 12333 8068
rect 12385 8016 12411 8068
rect 12463 8016 12489 8068
rect 12541 8016 12567 8068
rect 12619 8016 12622 8068
rect 12252 7997 12622 8016
rect 12252 7945 12255 7997
rect 12307 7945 12333 7997
rect 12385 7945 12411 7997
rect 12463 7945 12489 7997
rect 12541 7945 12567 7997
rect 12619 7945 12622 7997
rect 12252 7925 12622 7945
rect 12252 7873 12255 7925
rect 12307 7873 12333 7925
rect 12385 7873 12411 7925
rect 12463 7873 12489 7925
rect 12541 7873 12567 7925
rect 12619 7873 12622 7925
rect 12252 7867 12622 7873
rect 14292 9343 14312 9395
rect 14364 9343 14384 9395
rect 14436 9343 14456 9395
rect 14508 9343 14528 9395
rect 14580 9343 14600 9395
rect 14240 9330 14652 9343
rect 14292 9278 14312 9330
rect 14364 9278 14384 9330
rect 14436 9278 14456 9330
rect 14508 9278 14528 9330
rect 14580 9278 14600 9330
rect 14240 9265 14652 9278
rect 14292 9213 14312 9265
rect 14364 9213 14384 9265
rect 14436 9213 14456 9265
rect 14508 9213 14528 9265
rect 14580 9213 14600 9265
rect 14240 9200 14652 9213
rect 14292 9148 14312 9200
rect 14364 9148 14384 9200
rect 14436 9148 14456 9200
rect 14508 9148 14528 9200
rect 14580 9148 14600 9200
rect 14240 9135 14652 9148
rect 14292 9083 14312 9135
rect 14364 9083 14384 9135
rect 14436 9083 14456 9135
rect 14508 9083 14528 9135
rect 14580 9083 14600 9135
rect 14240 9070 14652 9083
rect 14292 9018 14312 9070
rect 14364 9018 14384 9070
rect 14436 9018 14456 9070
rect 14508 9018 14528 9070
rect 14580 9018 14600 9070
rect 14240 9005 14652 9018
rect 14292 8953 14312 9005
rect 14364 8953 14384 9005
rect 14436 8953 14456 9005
rect 14508 8953 14528 9005
rect 14580 8953 14600 9005
rect 14240 8940 14652 8953
rect 14292 8888 14312 8940
rect 14364 8888 14384 8940
rect 14436 8888 14456 8940
rect 14508 8888 14528 8940
rect 14580 8888 14600 8940
rect 14240 8875 14652 8888
rect 14292 8823 14312 8875
rect 14364 8823 14384 8875
rect 14436 8823 14456 8875
rect 14508 8823 14528 8875
rect 14580 8823 14600 8875
rect 14240 8810 14652 8823
rect 14292 8758 14312 8810
rect 14364 8758 14384 8810
rect 14436 8758 14456 8810
rect 14508 8758 14528 8810
rect 14580 8758 14600 8810
rect 14240 8745 14652 8758
rect 14292 8693 14312 8745
rect 14364 8693 14384 8745
rect 14436 8693 14456 8745
rect 14508 8693 14528 8745
rect 14580 8693 14600 8745
rect 14240 8680 14652 8693
rect 14292 8628 14312 8680
rect 14364 8628 14384 8680
rect 14436 8628 14456 8680
rect 14508 8628 14528 8680
rect 14580 8628 14600 8680
rect 14240 8615 14652 8628
rect 14292 8563 14312 8615
rect 14364 8563 14384 8615
rect 14436 8563 14456 8615
rect 14508 8563 14528 8615
rect 14580 8563 14600 8615
rect 14240 8550 14652 8563
rect 14292 8498 14312 8550
rect 14364 8498 14384 8550
rect 14436 8498 14456 8550
rect 14508 8498 14528 8550
rect 14580 8498 14600 8550
rect 14240 8485 14652 8498
rect 14292 8433 14312 8485
rect 14364 8433 14384 8485
rect 14436 8433 14456 8485
rect 14508 8433 14528 8485
rect 14580 8433 14600 8485
rect 14240 8420 14652 8433
rect 14292 8368 14312 8420
rect 14364 8368 14384 8420
rect 14436 8368 14456 8420
rect 14508 8368 14528 8420
rect 14580 8368 14600 8420
rect 14240 8354 14652 8368
rect 14292 8302 14312 8354
rect 14364 8302 14384 8354
rect 14436 8302 14456 8354
rect 14508 8302 14528 8354
rect 14580 8302 14600 8354
rect 14240 8288 14652 8302
rect 14292 8236 14312 8288
rect 14364 8236 14384 8288
rect 14436 8236 14456 8288
rect 14508 8236 14528 8288
rect 14580 8236 14600 8288
rect 14240 8222 14652 8236
rect 14292 8170 14312 8222
rect 14364 8170 14384 8222
rect 14436 8170 14456 8222
rect 14508 8170 14528 8222
rect 14580 8170 14600 8222
rect 14240 8156 14652 8170
rect 14292 8104 14312 8156
rect 14364 8104 14384 8156
rect 14436 8104 14456 8156
rect 14508 8104 14528 8156
rect 14580 8104 14600 8156
tri 11156 7561 11338 7743 sw
rect 10800 7509 11135 7561
rect 11187 7509 11208 7561
rect 11260 7509 11280 7561
rect 11332 7509 11338 7561
rect 10800 7481 11338 7509
rect 10800 7429 11135 7481
rect 11187 7429 11208 7481
rect 11260 7429 11280 7481
rect 11332 7429 11338 7481
rect 435 6992 970 7071
rect 435 6892 870 6992
tri 870 6892 970 6992 nw
tri 378 6880 390 6892 sw
rect 338 6874 390 6880
rect 338 6808 390 6822
rect 338 6750 390 6756
rect 338 872 378 6750
tri 378 6738 390 6750 nw
rect 435 5568 823 6892
tri 823 6845 870 6892 nw
rect 435 5516 516 5568
rect 568 5516 634 5568
rect 686 5516 751 5568
rect 803 5516 823 5568
rect 435 5479 823 5516
rect 435 5465 748 5479
rect 487 5413 507 5465
rect 559 5413 579 5465
rect 631 5413 651 5465
rect 703 5427 748 5465
rect 800 5427 823 5479
rect 703 5413 823 5427
rect 435 5400 823 5413
rect 487 5348 507 5400
rect 559 5348 579 5400
rect 631 5348 651 5400
rect 703 5348 823 5400
rect 435 5335 823 5348
rect 487 5283 507 5335
rect 559 5283 579 5335
rect 631 5283 651 5335
rect 703 5283 823 5335
rect 435 5270 823 5283
rect 487 5218 507 5270
rect 559 5218 579 5270
rect 631 5218 651 5270
rect 703 5218 823 5270
rect 435 5205 823 5218
rect 487 5153 507 5205
rect 559 5153 579 5205
rect 631 5153 651 5205
rect 703 5153 823 5205
rect 435 5140 823 5153
rect 487 5088 507 5140
rect 559 5088 579 5140
rect 631 5088 651 5140
rect 703 5088 823 5140
rect 14240 5565 14652 8104
rect 14240 5513 14313 5565
rect 14365 5513 14652 5565
rect 14240 5465 14652 5513
rect 14240 5413 14243 5465
rect 14295 5413 14309 5465
rect 14361 5413 14375 5465
rect 14427 5413 14441 5465
rect 14493 5413 14652 5465
rect 14240 5400 14652 5413
rect 14240 5348 14243 5400
rect 14295 5348 14309 5400
rect 14361 5348 14375 5400
rect 14427 5348 14441 5400
rect 14493 5348 14652 5400
rect 14240 5335 14652 5348
rect 14240 5283 14243 5335
rect 14295 5283 14309 5335
rect 14361 5283 14375 5335
rect 14427 5283 14441 5335
rect 14493 5283 14652 5335
rect 14240 5270 14652 5283
rect 14240 5218 14243 5270
rect 14295 5218 14309 5270
rect 14361 5218 14375 5270
rect 14427 5218 14441 5270
rect 14493 5218 14652 5270
rect 14240 5205 14652 5218
rect 14240 5153 14243 5205
rect 14295 5153 14309 5205
rect 14361 5153 14375 5205
rect 14427 5153 14441 5205
rect 14493 5153 14652 5205
rect 14240 5140 14652 5153
rect 14240 5088 14243 5140
rect 14295 5088 14309 5140
rect 14361 5088 14375 5140
rect 14427 5088 14441 5140
rect 14493 5088 14652 5140
rect 435 5075 823 5088
rect 487 5023 507 5075
rect 559 5023 579 5075
rect 631 5023 651 5075
rect 703 5023 823 5075
rect 435 5010 823 5023
rect 487 4958 507 5010
rect 559 4958 579 5010
rect 631 4958 651 5010
rect 703 4958 823 5010
rect 435 4945 823 4958
rect 487 4893 507 4945
rect 559 4893 579 4945
rect 631 4893 651 4945
rect 703 4893 823 4945
rect 435 4880 823 4893
rect 487 4828 507 4880
rect 559 4828 579 4880
rect 631 4828 651 4880
rect 703 4828 823 4880
rect 435 4815 823 4828
rect 487 4763 507 4815
rect 559 4763 579 4815
rect 631 4763 651 4815
rect 703 4763 823 4815
rect 435 4750 823 4763
rect 487 4698 507 4750
rect 559 4698 579 4750
rect 631 4698 651 4750
rect 703 4698 823 4750
rect 435 4685 823 4698
rect 487 4633 507 4685
rect 559 4633 579 4685
rect 631 4633 651 4685
rect 703 4633 823 4685
rect 435 4620 823 4633
rect 487 4568 507 4620
rect 559 4568 579 4620
rect 631 4568 651 4620
rect 703 4568 823 4620
rect 435 4555 823 4568
rect 487 4503 507 4555
rect 559 4503 579 4555
rect 631 4503 651 4555
rect 703 4503 823 4555
rect 435 4490 823 4503
rect 487 4438 507 4490
rect 559 4438 579 4490
rect 631 4438 651 4490
rect 703 4438 823 4490
rect 435 4425 823 4438
rect 487 4373 507 4425
rect 559 4373 579 4425
rect 631 4373 651 4425
rect 703 4373 823 4425
rect 435 4360 823 4373
rect 487 4308 507 4360
rect 559 4308 579 4360
rect 631 4308 651 4360
rect 703 4308 823 4360
rect 435 4295 823 4308
rect 487 4243 507 4295
rect 559 4243 579 4295
rect 631 4243 651 4295
rect 703 4243 823 4295
rect 435 4230 823 4243
rect 487 4178 507 4230
rect 559 4178 579 4230
rect 631 4178 651 4230
rect 703 4178 823 4230
rect 435 4165 823 4178
rect 487 4113 507 4165
rect 559 4113 579 4165
rect 631 4113 651 4165
rect 703 4113 823 4165
rect 435 4099 823 4113
rect 487 4047 507 4099
rect 559 4047 579 4099
rect 631 4047 651 4099
rect 703 4047 823 4099
rect 435 4033 823 4047
rect 487 3981 507 4033
rect 559 3981 579 4033
rect 631 3981 651 4033
rect 703 3981 823 4033
rect 11116 3995 12657 5088
rect 14240 5075 14652 5088
rect 14240 5023 14243 5075
rect 14295 5023 14309 5075
rect 14361 5023 14375 5075
rect 14427 5023 14441 5075
rect 14493 5023 14652 5075
rect 14240 5010 14652 5023
rect 14240 4958 14243 5010
rect 14295 4958 14309 5010
rect 14361 4958 14375 5010
rect 14427 4958 14441 5010
rect 14493 4958 14652 5010
rect 14240 4945 14652 4958
rect 14240 4893 14243 4945
rect 14295 4893 14309 4945
rect 14361 4893 14375 4945
rect 14427 4893 14441 4945
rect 14493 4893 14652 4945
rect 14240 4880 14652 4893
rect 14240 4828 14243 4880
rect 14295 4828 14309 4880
rect 14361 4828 14375 4880
rect 14427 4828 14441 4880
rect 14493 4828 14652 4880
rect 14240 4815 14652 4828
rect 14240 4763 14243 4815
rect 14295 4763 14309 4815
rect 14361 4763 14375 4815
rect 14427 4763 14441 4815
rect 14493 4763 14652 4815
rect 14240 4750 14652 4763
rect 14240 4698 14243 4750
rect 14295 4698 14309 4750
rect 14361 4698 14375 4750
rect 14427 4698 14441 4750
rect 14493 4698 14652 4750
rect 14240 4685 14652 4698
rect 14240 4633 14243 4685
rect 14295 4633 14309 4685
rect 14361 4633 14375 4685
rect 14427 4633 14441 4685
rect 14493 4633 14652 4685
rect 14240 4620 14652 4633
rect 14240 4568 14243 4620
rect 14295 4568 14309 4620
rect 14361 4568 14375 4620
rect 14427 4568 14441 4620
rect 14493 4568 14652 4620
rect 14240 4555 14652 4568
rect 14240 4503 14243 4555
rect 14295 4503 14309 4555
rect 14361 4503 14375 4555
rect 14427 4503 14441 4555
rect 14493 4503 14652 4555
rect 14240 4490 14652 4503
rect 14240 4438 14243 4490
rect 14295 4438 14309 4490
rect 14361 4438 14375 4490
rect 14427 4438 14441 4490
rect 14493 4438 14652 4490
rect 14240 4425 14652 4438
rect 14240 4373 14243 4425
rect 14295 4373 14309 4425
rect 14361 4373 14375 4425
rect 14427 4373 14441 4425
rect 14493 4373 14652 4425
rect 14240 4359 14652 4373
rect 14240 4307 14243 4359
rect 14295 4307 14309 4359
rect 14361 4307 14375 4359
rect 14427 4307 14441 4359
rect 14493 4307 14652 4359
rect 14240 4293 14652 4307
rect 14240 4241 14243 4293
rect 14295 4241 14309 4293
rect 14361 4241 14375 4293
rect 14427 4241 14441 4293
rect 14493 4241 14652 4293
rect 14240 4227 14652 4241
rect 14240 4175 14243 4227
rect 14295 4175 14309 4227
rect 14361 4175 14375 4227
rect 14427 4175 14441 4227
rect 14493 4175 14652 4227
rect 14240 4161 14652 4175
rect 14240 4109 14243 4161
rect 14295 4109 14309 4161
rect 14361 4109 14375 4161
rect 14427 4109 14441 4161
rect 14493 4109 14652 4161
rect 14240 4095 14652 4109
rect 14240 4043 14243 4095
rect 14295 4043 14309 4095
rect 14361 4043 14375 4095
rect 14427 4043 14441 4095
rect 14493 4043 14652 4095
rect 14240 4029 14652 4043
rect 435 3967 823 3981
rect 487 3915 507 3967
rect 559 3915 579 3967
rect 631 3915 651 3967
rect 703 3915 823 3967
rect 435 3901 823 3915
rect 487 3849 507 3901
rect 559 3849 579 3901
rect 631 3849 651 3901
rect 703 3849 823 3901
rect 14240 3977 14243 4029
rect 14295 3977 14309 4029
rect 14361 3977 14375 4029
rect 14427 3977 14441 4029
rect 14493 3977 14652 4029
rect 14240 3963 14652 3977
rect 14240 3911 14243 3963
rect 14295 3911 14309 3963
rect 14361 3911 14375 3963
rect 14427 3911 14441 3963
rect 14493 3911 14652 3963
rect 14240 3897 14652 3911
tri 14234 3883 14240 3889 se
rect 14240 3883 14243 3897
rect 435 3845 823 3849
tri 823 3845 861 3883 sw
tri 14196 3845 14234 3883 se
rect 14234 3845 14243 3883
rect 14295 3845 14309 3897
rect 14361 3845 14375 3897
rect 14427 3845 14441 3897
rect 14493 3845 14652 3897
rect 435 3835 861 3845
rect 487 3783 507 3835
rect 559 3783 579 3835
rect 631 3783 651 3835
rect 703 3831 861 3835
tri 861 3831 875 3845 sw
tri 14182 3831 14196 3845 se
rect 14196 3831 14652 3845
rect 703 3783 875 3831
rect 435 3779 875 3783
tri 875 3779 927 3831 sw
tri 14130 3779 14182 3831 se
rect 14182 3779 14243 3831
rect 14295 3779 14309 3831
rect 14361 3779 14375 3831
rect 14427 3779 14441 3831
rect 14493 3779 14652 3831
rect 435 3769 927 3779
rect 487 3717 507 3769
rect 559 3717 579 3769
rect 631 3717 651 3769
rect 703 3765 927 3769
tri 927 3765 941 3779 sw
tri 14116 3765 14130 3779 se
rect 14130 3765 14652 3779
rect 703 3717 941 3765
rect 435 3713 941 3717
tri 941 3713 993 3765 sw
tri 14064 3713 14116 3765 se
rect 14116 3713 14243 3765
rect 14295 3713 14309 3765
rect 14361 3713 14375 3765
rect 14427 3713 14441 3765
rect 14493 3713 14652 3765
rect 435 3703 993 3713
rect 487 3651 507 3703
rect 559 3651 579 3703
rect 631 3651 651 3703
rect 703 3699 993 3703
tri 993 3699 1007 3713 sw
tri 14050 3699 14064 3713 se
rect 14064 3699 14652 3713
rect 703 3651 1007 3699
rect 435 3647 1007 3651
tri 1007 3647 1059 3699 sw
tri 13998 3647 14050 3699 se
rect 14050 3647 14243 3699
rect 14295 3647 14309 3699
rect 14361 3647 14375 3699
rect 14427 3647 14441 3699
rect 14493 3647 14652 3699
rect 435 3645 1059 3647
tri 1059 3645 1061 3647 sw
tri 13996 3645 13998 3647 se
rect 13998 3645 14652 3647
rect 435 3631 1061 3645
tri 1061 3631 1075 3645 sw
tri 13992 3641 13996 3645 se
rect 13996 3641 14652 3645
tri 13982 3631 13992 3641 se
rect 13992 3631 14652 3641
rect 435 2530 1090 3631
rect 14439 3628 14652 3631
rect 13300 2554 14652 3628
rect 14439 2530 14652 2554
tri 378 872 412 906 sw
rect 338 820 580 872
rect 632 820 648 872
rect 700 820 707 872
rect 338 806 707 820
rect 338 754 580 806
rect 632 754 648 806
rect 700 754 707 806
rect 338 753 707 754
rect 3710 871 3934 872
rect 3710 819 3716 871
rect 3768 819 3796 871
rect 3848 819 3876 871
rect 3928 819 3934 871
rect 3710 805 3934 819
rect 3710 753 3716 805
rect 3768 753 3796 805
rect 3848 753 3876 805
rect 3928 753 3934 805
rect 338 487 486 753
tri 486 661 578 753 nw
tri 486 487 551 552 sw
rect 3710 487 3934 753
rect 338 435 580 487
rect 632 435 648 487
rect 700 435 708 487
rect 338 421 708 435
rect 338 369 580 421
rect 632 369 648 421
rect 700 369 708 421
rect 338 368 708 369
rect 3710 435 3716 487
rect 3768 435 3796 487
rect 3848 435 3876 487
rect 3928 435 3934 487
rect 3710 421 3934 435
rect 3710 369 3716 421
rect 3768 369 3796 421
rect 3848 369 3876 421
rect 3928 369 3934 421
tri 310 135 352 177 sw
rect 3710 135 3934 369
rect 278 83 284 135
rect 336 83 348 135
rect 400 83 406 135
rect 3710 83 3716 135
rect 3768 83 3796 135
rect 3848 83 3876 135
rect 3928 83 3934 135
rect 14708 -6 14748 16023
rect 14788 -6 14828 16103
rect 14868 -6 14908 16212
rect 14948 -6 14988 16292
rect 15028 -6 15068 16372
rect 5247 -9151 5930 -9145
rect 5247 -9203 5878 -9151
rect 5247 -9223 5930 -9203
rect 5247 -9275 5878 -9223
rect 5247 -9281 5930 -9275
rect 5247 -9942 5685 -9281
tri 5685 -9474 5878 -9281 nw
tri 13421 -9579 13477 -9523 se
rect 13477 -9579 14216 -9523
tri 14216 -9579 14272 -9523 sw
tri 13343 -9657 13421 -9579 se
rect 13421 -9644 13434 -9579
tri 13434 -9644 13499 -9579 nw
tri 14194 -9644 14259 -9579 ne
rect 14259 -9644 14272 -9579
tri 14272 -9644 14337 -9579 sw
tri 13421 -9657 13434 -9644 nw
tri 14259 -9657 14272 -9644 ne
rect 14272 -9657 14337 -9644
tri 13299 -9701 13343 -9657 se
rect 13343 -9701 13356 -9657
rect 5247 -9994 5253 -9942
rect 5305 -9994 5328 -9942
rect 5380 -9994 5403 -9942
rect 5455 -9994 5478 -9942
rect 5530 -9994 5553 -9942
rect 5605 -9994 5627 -9942
rect 5679 -9994 5685 -9942
rect 5247 -10017 5685 -9994
rect 5247 -10069 5253 -10017
rect 5305 -10069 5328 -10017
rect 5380 -10069 5403 -10017
rect 5455 -10069 5478 -10017
rect 5530 -10069 5553 -10017
rect 5605 -10069 5627 -10017
rect 5679 -10069 5685 -10017
rect 5247 -10092 5685 -10069
rect 5247 -10144 5253 -10092
rect 5305 -10144 5328 -10092
rect 5380 -10144 5403 -10092
rect 5455 -10144 5478 -10092
rect 5530 -10144 5553 -10092
rect 5605 -10144 5627 -10092
rect 5679 -10144 5685 -10092
rect 5247 -10933 5685 -10144
rect 8191 -10933 8667 -9701
tri 13273 -9727 13299 -9701 se
rect 13299 -9722 13356 -9701
tri 13356 -9722 13421 -9657 nw
tri 14272 -9722 14337 -9657 ne
tri 14337 -9722 14415 -9644 sw
rect 13299 -9727 13343 -9722
tri 13265 -9735 13273 -9727 se
rect 13273 -9735 13343 -9727
tri 13343 -9735 13356 -9722 nw
tri 14337 -9735 14350 -9722 ne
rect 14350 -9735 14415 -9722
tri 13217 -9783 13265 -9735 se
rect 13265 -9744 13334 -9735
tri 13334 -9744 13343 -9735 nw
tri 14350 -9744 14359 -9735 ne
rect 14359 -9744 14415 -9735
tri 14415 -9744 14437 -9722 sw
rect 13265 -9783 13278 -9744
rect 13217 -9800 13278 -9783
tri 13278 -9800 13334 -9744 nw
tri 14359 -9800 14415 -9744 ne
rect 14415 -9800 14485 -9744
rect 14541 -9800 14565 -9744
rect 14621 -9800 14630 -9744
tri 13195 -10328 13217 -10306 se
rect 13217 -10328 13273 -9800
tri 13273 -9805 13278 -9800 nw
tri 13117 -10406 13195 -10328 se
tri 13195 -10406 13273 -10328 nw
tri 13061 -10462 13117 -10406 se
tri 12501 -10484 12523 -10462 se
rect 12523 -10484 13117 -10462
tri 13117 -10484 13195 -10406 nw
tri 12467 -10518 12501 -10484 se
rect 12501 -10518 13083 -10484
tri 13083 -10518 13117 -10484 nw
tri 12389 -10596 12467 -10518 se
tri 12467 -10596 12545 -10518 nw
tri 12311 -10674 12389 -10596 se
tri 12389 -10674 12467 -10596 nw
tri 12235 -10750 12311 -10674 se
rect 12235 -10752 12311 -10750
tri 12311 -10752 12389 -10674 nw
tri 8667 -10933 8773 -10827 sw
rect 5247 -10985 5253 -10933
rect 5305 -10985 5328 -10933
rect 5380 -10985 5403 -10933
rect 5455 -10985 5478 -10933
rect 5530 -10985 5553 -10933
rect 5605 -10985 5627 -10933
rect 5679 -10985 5685 -10933
rect 5247 -11011 5685 -10985
rect 5247 -11063 5253 -11011
rect 5305 -11063 5328 -11011
rect 5380 -11063 5403 -11011
rect 5455 -11063 5478 -11011
rect 5530 -11063 5553 -11011
rect 5605 -11063 5627 -11011
rect 5679 -11063 5685 -11011
rect 12235 -13613 12291 -10752
tri 12291 -10772 12311 -10752 nw
<< rmetal2 >>
rect 498 16118 628 16119
rect 498 16117 499 16118
rect 627 16117 628 16118
rect 740 16118 870 16119
rect 740 16117 741 16118
rect 869 16117 870 16118
rect 981 16118 1111 16119
rect 981 16117 982 16118
rect 1110 16117 1111 16118
rect 1345 16118 1475 16119
rect 1345 16117 1346 16118
rect 1474 16117 1475 16118
rect 1649 16118 1779 16119
rect 1649 16117 1650 16118
rect 1778 16117 1779 16118
rect 1932 16118 2062 16119
rect 1932 16117 1933 16118
rect 2061 16117 2062 16118
rect 498 15816 499 15817
rect 627 15816 628 15817
rect 498 15815 628 15816
rect 740 15816 741 15817
rect 869 15816 870 15817
rect 740 15815 870 15816
rect 981 15816 982 15817
rect 1110 15816 1111 15817
rect 981 15815 1111 15816
rect 1345 15816 1346 15817
rect 1474 15816 1475 15817
rect 1345 15815 1475 15816
rect 1649 15816 1650 15817
rect 1778 15816 1779 15817
rect 1649 15815 1779 15816
rect 1932 15816 1933 15817
rect 2061 15816 2062 15817
rect 1932 15815 2062 15816
rect 6888 16118 7018 16119
rect 6888 16117 6889 16118
rect 7017 16117 7018 16118
rect 7318 16118 7448 16119
rect 7318 16117 7319 16118
rect 7447 16117 7448 16118
rect 7748 16118 7878 16119
rect 7748 16117 7749 16118
rect 7877 16117 7878 16118
rect 8590 16118 8720 16119
rect 8590 16117 8591 16118
rect 8719 16117 8720 16118
rect 9020 16118 9150 16119
rect 9020 16117 9021 16118
rect 9149 16117 9150 16118
rect 9450 16118 9580 16119
rect 9450 16117 9451 16118
rect 9579 16117 9580 16118
rect 6888 15816 6889 15817
rect 7017 15816 7018 15817
rect 6888 15815 7018 15816
rect 7318 15816 7319 15817
rect 7447 15816 7448 15817
rect 7318 15815 7448 15816
rect 7748 15816 7749 15817
rect 7877 15816 7878 15817
rect 7748 15815 7878 15816
rect 8590 15816 8591 15817
rect 8719 15816 8720 15817
rect 8590 15815 8720 15816
rect 9020 15816 9021 15817
rect 9149 15816 9150 15817
rect 9020 15815 9150 15816
rect 9450 15816 9451 15817
rect 9579 15816 9580 15817
rect 9450 15815 9580 15816
rect 10070 16118 10200 16119
rect 10070 16117 10071 16118
rect 10199 16117 10200 16118
rect 10500 16118 10630 16119
rect 10500 16117 10501 16118
rect 10629 16117 10630 16118
rect 10930 16118 11060 16119
rect 10930 16117 10931 16118
rect 11059 16117 11060 16118
rect 11413 16118 11543 16119
rect 11413 16117 11414 16118
rect 11542 16117 11543 16118
rect 11843 16118 11973 16119
rect 11843 16117 11844 16118
rect 11972 16117 11973 16118
rect 12273 16118 12403 16119
rect 12273 16117 12274 16118
rect 12402 16117 12403 16118
rect 12847 16118 12977 16119
rect 12847 16117 12848 16118
rect 12976 16117 12977 16118
rect 13277 16118 13407 16119
rect 13277 16117 13278 16118
rect 13406 16117 13407 16118
rect 13707 16118 13837 16119
rect 13707 16117 13708 16118
rect 13836 16117 13837 16118
rect 10070 15816 10071 15817
rect 10199 15816 10200 15817
rect 10070 15815 10200 15816
rect 10500 15816 10501 15817
rect 10629 15816 10630 15817
rect 10500 15815 10630 15816
rect 10930 15816 10931 15817
rect 11059 15816 11060 15817
rect 10930 15815 11060 15816
rect 11413 15816 11414 15817
rect 11542 15816 11543 15817
rect 11413 15815 11543 15816
rect 11843 15816 11844 15817
rect 11972 15816 11973 15817
rect 11843 15815 11973 15816
rect 12273 15816 12274 15817
rect 12402 15816 12403 15817
rect 12273 15815 12403 15816
rect 12847 15816 12848 15817
rect 12976 15816 12977 15817
rect 12847 15815 12977 15816
rect 13277 15816 13278 15817
rect 13406 15816 13407 15817
rect 13277 15815 13407 15816
rect 13707 15816 13708 15817
rect 13836 15816 13837 15817
rect 13707 15815 13837 15816
<< via2 >>
rect 14591 16554 14647 16610
rect 14591 16474 14647 16530
rect 4605 15381 4661 15388
rect 4710 15381 4766 15388
rect 4815 15381 4871 15388
rect 4919 15381 4975 15388
rect 5023 15381 5079 15388
rect 4605 15332 4654 15381
rect 4654 15332 4661 15381
rect 4710 15332 4739 15381
rect 4739 15332 4766 15381
rect 4815 15332 4824 15381
rect 4824 15332 4856 15381
rect 4856 15332 4871 15381
rect 4919 15332 4940 15381
rect 4940 15332 4975 15381
rect 5023 15332 5024 15381
rect 5024 15332 5076 15381
rect 5076 15332 5079 15381
rect 4605 15265 4661 15268
rect 4710 15265 4766 15268
rect 4815 15265 4871 15268
rect 4919 15265 4975 15268
rect 5023 15265 5079 15268
rect 4605 15213 4654 15265
rect 4654 15213 4661 15265
rect 4710 15213 4739 15265
rect 4739 15213 4766 15265
rect 4815 15213 4824 15265
rect 4824 15213 4856 15265
rect 4856 15213 4871 15265
rect 4919 15213 4940 15265
rect 4940 15213 4975 15265
rect 5023 15213 5024 15265
rect 5024 15213 5076 15265
rect 5076 15213 5079 15265
rect 4605 15212 4661 15213
rect 4710 15212 4766 15213
rect 4815 15212 4871 15213
rect 4919 15212 4975 15213
rect 5023 15212 5079 15213
rect 4605 15097 4654 15148
rect 4654 15097 4661 15148
rect 4710 15097 4739 15148
rect 4739 15097 4766 15148
rect 4815 15097 4824 15148
rect 4824 15097 4856 15148
rect 4856 15097 4871 15148
rect 4919 15097 4940 15148
rect 4940 15097 4975 15148
rect 5023 15097 5024 15148
rect 5024 15097 5076 15148
rect 5076 15097 5079 15148
rect 4605 15092 4661 15097
rect 4710 15092 4766 15097
rect 4815 15092 4871 15097
rect 4919 15092 4975 15097
rect 5023 15092 5079 15097
rect 9052 15332 9108 15388
rect 9169 15332 9225 15388
rect 9286 15332 9342 15388
rect 9052 15212 9108 15268
rect 9169 15212 9225 15268
rect 9286 15212 9342 15268
rect 9052 15092 9108 15148
rect 9169 15092 9225 15148
rect 9286 15092 9342 15148
rect 14485 -9800 14541 -9744
rect 14565 -9800 14621 -9744
<< metal3 >>
rect 14586 16610 14652 16615
rect 14586 16554 14591 16610
rect 14647 16554 14652 16610
rect 14586 16530 14652 16554
rect 14586 16474 14591 16530
rect 14647 16474 14652 16530
rect 4600 15388 5084 15393
rect 4600 15332 4605 15388
rect 4661 15332 4710 15388
rect 4766 15332 4815 15388
rect 4871 15332 4919 15388
rect 4975 15332 5023 15388
rect 5079 15332 5084 15388
rect 4600 15268 5084 15332
rect 4600 15212 4605 15268
rect 4661 15212 4710 15268
rect 4766 15212 4815 15268
rect 4871 15212 4919 15268
rect 4975 15212 5023 15268
rect 5079 15212 5084 15268
rect 4600 15148 5084 15212
rect 4600 15092 4605 15148
rect 4661 15092 4710 15148
rect 4766 15092 4815 15148
rect 4871 15092 4919 15148
rect 4975 15092 5023 15148
rect 5079 15092 5084 15148
rect 4600 13425 5084 15092
rect 9047 15388 9347 15393
rect 9047 15332 9052 15388
rect 9108 15332 9169 15388
rect 9225 15332 9286 15388
rect 9342 15332 9347 15388
rect 9047 15268 9347 15332
rect 9047 15212 9052 15268
rect 9108 15212 9169 15268
rect 9225 15212 9286 15268
rect 9342 15212 9347 15268
rect 9047 15148 9347 15212
rect 9047 15092 9052 15148
rect 9108 15092 9169 15148
rect 9225 15092 9286 15148
rect 9342 15092 9347 15148
rect 6107 13425 6811 15087
rect 9047 13425 9347 15092
tri 14480 -9739 14586 -9633 se
rect 14586 -9739 14652 16474
rect 14480 -9744 14652 -9739
rect 14480 -9800 14485 -9744
rect 14541 -9800 14565 -9744
rect 14621 -9800 14652 -9744
rect 14480 -9805 14652 -9800
use sky130_fd_io__com_pudrvr_strong_slowv2  sky130_fd_io__com_pudrvr_strong_slowv2_0
timestamp 1694700623
transform -1 0 7012 0 1 139
box 1755 196 3286 766
use sky130_fd_io__com_pudrvr_weakv2  sky130_fd_io__com_pudrvr_weakv2_0
timestamp 1694700623
transform 1 0 78 0 1 139
box -36 -176 3550 1143
use sky130_fd_io__com_res_weak  sky130_fd_io__com_res_weak_0
timestamp 1694700623
transform 0 1 1833 1 0 6897
box -160 1014 679 10611
use sky130_fd_io__gpio_pddrvr_strong_slowv2  sky130_fd_io__gpio_pddrvr_strong_slowv2_0
timestamp 1694700623
transform 0 1 420 -1 0 15675
box 414 362 536 4714
use sky130_fd_io__gpio_pddrvr_weakv2  sky130_fd_io__gpio_pddrvr_weakv2_0
timestamp 1694700623
transform 0 1 5329 -1 0 15675
box -202 0 1152 7520
use sky130_fd_io__gpio_pudrvr_strongv2  sky130_fd_io__gpio_pudrvr_strongv2_0
timestamp 1694700623
transform 1 0 -580 0 1 622
box 467 -902 15583 5464
use sky130_fd_io__gpiov2_pddrvr_strong  sky130_fd_io__gpiov2_pddrvr_strong_0
timestamp 1694700623
transform 1 0 85 0 -1 17755
box -85 1584 15088 9417
use sky130_fd_io__res250only_small  sky130_fd_io__res250only_small_0
timestamp 1694700623
transform -1 0 13372 0 -1 8288
box 0 0 2270 404
use sky130_fd_io__tk_em1s_cdns_5595914180852  sky130_fd_io__tk_em1s_cdns_5595914180852_0
timestamp 1694700623
transform -1 0 10237 0 -1 8259
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180853  sky130_fd_pr__res_generic_po__example_5595914180853_0
timestamp 1694700623
transform -1 0 10314 0 1 7886
box 15 31 585 32
use sky130_fd_pr__res_generic_po__example_5595914180855  sky130_fd_pr__res_generic_po__example_5595914180855_0
timestamp 1694700623
transform -1 0 9612 0 1 7886
box 15 31 985 32
use sky130_fd_pr__res_generic_po__example_5595914180856  sky130_fd_pr__res_generic_po__example_5595914180856_0
timestamp 1694700623
transform -1 0 10816 0 1 7886
box 15 31 385 32
use sky130_fd_pr__via_l1m1__example_5595914180832  sky130_fd_pr__via_l1m1__example_5595914180832_0
timestamp 1694700623
transform 1 0 8509 0 1 7932
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_0
timestamp 1694700623
transform 0 1 8561 1 0 8086
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_1
timestamp 1694700623
transform 0 -1 10867 1 0 8086
box 0 0 1 1
<< labels >>
flabel locali s 310 1322 402 1368 3 FreeSans 520 0 0 0 VGND
port 1 nsew
flabel comment s 1426 15454 1426 15454 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 6755 15452 6755 15452 0 FreeSans 440 0 0 0 CONDIODE
flabel metal2 s 14708 -6 14748 186 3 FreeSans 520 90 0 0 PD_H[0]
port 3 nsew
flabel metal2 s 14868 -6 14908 186 3 FreeSans 520 90 0 0 PD_H[2]
port 4 nsew
flabel metal2 s 14788 -6 14828 186 3 FreeSans 520 90 0 0 PD_H[1]
port 5 nsew
flabel metal2 s 14948 -6 14988 186 3 FreeSans 520 90 0 0 PD_H[3]
port 6 nsew
flabel metal2 s 13300 2554 14496 3628 3 FreeSans 520 0 0 0 VCC_IO
port 7 nsew
flabel metal2 s 11116 3995 12657 5088 3 FreeSans 520 0 0 0 PAD
port 8 nsew
flabel metal2 s 11116 10850 12657 11943 3 FreeSans 520 0 0 0 PAD
port 8 nsew
flabel metal2 s 15028 -6 15068 186 3 FreeSans 520 90 0 0 TIE_LO_ESD
port 9 nsew
flabel metal1 s 49 -1067 83 -1013 3 FreeSans 520 270 0 0 FORCE_HI_H_N
port 10 nsew
flabel metal1 s 377 -1075 415 -1020 3 FreeSans 520 270 0 0 FORCE_LO_H
port 11 nsew
flabel metal1 s 258 -1075 313 -1023 3 FreeSans 520 270 0 0 FORCE_LOVOL_H
port 12 nsew
flabel metal1 s 761 683 794 715 3 FreeSans 520 0 0 0 PU_H_N[0]
port 13 nsew
flabel metal1 s 6527 686 6583 719 3 FreeSans 520 0 0 0 PU_H_N[1]
port 14 nsew
flabel metal1 s 14167 280 14252 332 3 FreeSans 520 0 0 0 PU_H_N[2]
port 15 nsew
flabel metal1 s 13921 168 14073 220 3 FreeSans 520 0 0 0 PU_H_N[3]
port 16 nsew
flabel metal1 s 167 -1074 205 -1007 3 FreeSans 520 270 0 0 VSSIO_AMX
port 17 nsew
flabel metal1 s 2496 8314 2549 8360 3 FreeSans 520 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 14164 88 14240 140 3 FreeSans 520 0 0 0 TIE_HI_ESD
port 19 nsew
flabel metal1 s 13310 7924 13365 8257 3 FreeSans 520 0 0 0 PAD
port 8 nsew
flabel metal1 s 11799 736 11831 794 3 FreeSans 520 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 451 932 1620 1077 3 FreeSans 520 0 0 0 VCC_IO
port 7 nsew
flabel metal1 s 3948 909 5117 955 3 FreeSans 520 0 0 0 VCC_IO
port 7 nsew
<< properties >>
string GDS_END 6593872
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 5685286
<< end >>
