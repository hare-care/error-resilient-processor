magic
tech sky130A
timestamp 1694700623
<< properties >>
string GDS_END 7065550
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7064394
<< end >>
