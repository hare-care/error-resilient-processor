magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 355 47 385 177
rect 439 47 469 177
rect 627 47 657 177
<< scpmoshvt >>
rect 83 297 113 497
rect 174 297 204 497
rect 283 297 313 497
rect 433 297 463 497
rect 627 297 657 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 169 163 177
rect 109 135 119 169
rect 153 135 163 169
rect 109 47 163 135
rect 193 165 249 177
rect 193 131 207 165
rect 241 131 249 165
rect 193 47 249 131
rect 303 93 355 177
rect 303 59 311 93
rect 345 59 355 93
rect 303 47 355 59
rect 385 93 439 177
rect 385 59 395 93
rect 429 59 439 93
rect 385 47 439 59
rect 469 127 521 177
rect 469 93 479 127
rect 513 93 521 127
rect 469 47 521 93
rect 575 165 627 177
rect 575 131 583 165
rect 617 131 627 165
rect 575 97 627 131
rect 575 63 583 97
rect 617 63 627 97
rect 575 47 627 63
rect 657 93 709 177
rect 657 59 667 93
rect 701 59 709 93
rect 657 47 709 59
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 409 174 497
rect 113 375 123 409
rect 157 375 174 409
rect 113 341 174 375
rect 113 307 123 341
rect 157 307 174 341
rect 113 297 174 307
rect 204 297 283 497
rect 313 485 433 497
rect 313 451 349 485
rect 383 451 433 485
rect 313 417 433 451
rect 313 383 349 417
rect 383 383 433 417
rect 313 297 433 383
rect 463 481 515 497
rect 463 447 473 481
rect 507 447 515 481
rect 463 413 515 447
rect 463 379 473 413
rect 507 379 515 413
rect 463 345 515 379
rect 463 311 473 345
rect 507 311 515 345
rect 463 297 515 311
rect 569 477 627 497
rect 569 443 583 477
rect 617 443 627 477
rect 569 409 627 443
rect 569 375 583 409
rect 617 375 627 409
rect 569 341 627 375
rect 569 307 583 341
rect 617 307 627 341
rect 569 297 627 307
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 417 709 451
rect 657 383 667 417
rect 701 383 709 417
rect 657 297 709 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 135 153 169
rect 207 131 241 165
rect 311 59 345 93
rect 395 59 429 93
rect 479 93 513 127
rect 583 131 617 165
rect 583 63 617 97
rect 667 59 701 93
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 375 157 409
rect 123 307 157 341
rect 349 451 383 485
rect 349 383 383 417
rect 473 447 507 481
rect 473 379 507 413
rect 473 311 507 345
rect 583 443 617 477
rect 583 375 617 409
rect 583 307 617 341
rect 667 451 701 485
rect 667 383 701 417
<< poly >>
rect 83 497 113 523
rect 174 497 204 523
rect 283 497 313 523
rect 433 497 463 523
rect 627 497 657 523
rect 83 265 113 297
rect 174 265 204 297
rect 21 249 113 265
rect 21 215 34 249
rect 68 215 113 249
rect 21 200 113 215
rect 163 249 235 265
rect 163 215 191 249
rect 225 215 235 249
rect 21 199 109 200
rect 79 177 109 199
rect 163 199 235 215
rect 283 259 313 297
rect 433 270 463 297
rect 627 270 657 297
rect 433 265 657 270
rect 283 249 391 259
rect 283 215 299 249
rect 333 215 391 249
rect 433 249 715 265
rect 433 233 670 249
rect 283 205 391 215
rect 163 177 193 199
rect 355 177 385 205
rect 439 177 469 233
rect 627 215 670 233
rect 704 215 715 249
rect 627 198 715 215
rect 627 177 657 198
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 439 21 469 47
rect 627 21 657 47
<< polycont >>
rect 34 215 68 249
rect 191 215 225 249
rect 299 215 333 249
rect 670 215 704 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 24 477 315 493
rect 24 443 39 477
rect 73 459 315 477
rect 73 443 84 459
rect 24 409 84 443
rect 24 375 39 409
rect 73 375 84 409
rect 24 341 84 375
rect 24 307 39 341
rect 73 307 84 341
rect 24 291 84 307
rect 118 409 168 425
rect 118 375 123 409
rect 157 375 168 409
rect 118 341 168 375
rect 118 307 123 341
rect 157 307 168 341
rect 118 291 168 307
rect 17 249 84 257
rect 17 215 34 249
rect 68 215 84 249
rect 17 212 84 215
rect 17 161 69 177
rect 17 127 35 161
rect 17 93 69 127
rect 118 169 156 291
rect 207 289 247 422
rect 281 330 315 459
rect 349 485 395 527
rect 383 451 395 485
rect 349 417 395 451
rect 383 383 395 417
rect 349 367 395 383
rect 457 481 523 493
rect 457 447 473 481
rect 507 447 523 481
rect 457 413 523 447
rect 457 379 473 413
rect 507 379 523 413
rect 457 345 523 379
rect 457 330 473 345
rect 281 311 473 330
rect 507 311 523 345
rect 281 296 523 311
rect 572 477 617 493
rect 572 443 583 477
rect 572 409 617 443
rect 572 375 583 409
rect 572 341 617 375
rect 659 485 718 527
rect 659 451 667 485
rect 701 451 718 485
rect 659 417 718 451
rect 659 383 667 417
rect 701 383 718 417
rect 659 367 718 383
rect 572 307 583 341
rect 207 265 241 289
rect 191 249 241 265
rect 572 262 617 307
rect 225 231 241 249
rect 277 249 617 262
rect 277 215 299 249
rect 333 215 617 249
rect 191 199 225 215
rect 118 135 119 169
rect 153 135 156 169
rect 259 165 524 177
rect 118 119 156 135
rect 191 131 207 165
rect 241 143 524 165
rect 241 131 304 143
rect 477 127 524 143
rect 395 93 429 109
rect 17 59 35 93
rect 69 85 88 93
rect 193 85 311 93
rect 69 59 311 85
rect 345 59 361 93
rect 17 51 361 59
rect 395 17 429 59
rect 477 93 479 127
rect 513 93 524 127
rect 477 51 524 93
rect 560 165 617 215
rect 560 131 583 165
rect 652 249 719 324
rect 652 215 670 249
rect 704 215 719 249
rect 652 152 719 215
rect 560 97 617 131
rect 560 63 583 97
rect 617 63 633 97
rect 560 51 633 63
rect 667 93 711 109
rect 701 59 711 93
rect 667 17 711 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 213 357 247 391 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 672 153 706 187 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 672 289 706 323 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 121 357 155 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 mux2i_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1697552
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1690656
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
