magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< dnwell >>
rect 10767 4548 12349 4662
rect 7880 4441 12349 4548
rect 288 3528 12349 4441
rect 288 1264 12460 3528
rect 288 754 12410 1264
rect 288 362 8077 754
<< nwell >>
rect -568 4865 218 5007
rect -568 4633 324 4865
rect -568 4576 298 4633
rect 376 4576 1284 4770
rect 5946 4576 6819 4670
rect 10757 4646 12436 4666
rect 10757 4576 12453 4646
rect -568 4298 12603 4576
rect 204 4237 12603 4298
rect 204 3574 8268 4237
rect -310 3573 8268 3574
rect -567 3137 8268 3573
rect 9071 4117 12603 4237
rect 9071 3652 12781 4117
rect 9377 3187 10542 3652
rect 10943 3281 12781 3652
rect 10943 3239 11981 3281
rect -567 3037 6028 3137
rect -567 2967 4818 3037
rect -567 2835 494 2967
rect 1618 2959 4818 2967
rect -568 2134 494 2835
rect 9574 2872 10542 3187
rect 204 1647 494 2134
rect 204 1300 578 1647
rect 2236 1618 3400 1731
rect 12254 2714 12781 3281
rect 12254 1868 12603 2714
rect 2236 1586 10588 1618
rect 1185 1521 10588 1586
rect 1185 1415 11304 1521
rect 12254 1415 12626 1868
rect 1185 1300 12626 1415
rect 204 631 12626 1300
rect 204 282 12603 631
rect 7997 241 12603 282
rect 10044 239 10654 241
<< pwell >>
rect -487 4141 143 4193
rect -670 4001 143 4141
rect -670 3738 54 4001
rect -504 3735 54 3738
rect -224 3679 54 3735
rect 8725 4135 9011 4169
rect 8328 3227 9011 4135
rect 8328 3177 8608 3227
rect 7508 2744 9514 2996
rect 10826 3123 12160 3153
rect 7584 2676 9514 2744
rect 9722 2676 10394 2704
rect 7584 2398 10394 2676
rect 10718 2510 12160 3123
rect 7584 2333 7998 2398
rect -487 1837 143 2029
rect -459 1719 141 1837
rect 7544 1681 7998 2333
rect 8644 2334 10394 2398
rect 10750 2362 12160 2510
rect 8644 1739 10548 2334
rect 10750 1782 12193 2362
rect 10750 1746 12084 1782
rect 8644 1682 10436 1739
<< mvnmos >>
rect -408 4027 -288 4167
rect -232 4027 -112 4167
rect -56 4027 64 4167
rect -425 3761 -325 3845
rect -145 3705 -25 3845
rect 8354 3256 8438 4056
rect 8498 3256 8582 4056
rect 7587 2770 7707 2970
rect 7763 2770 7883 2970
rect 7939 2770 8059 2970
rect 8115 2770 8235 2970
rect 8291 2770 8411 2970
rect 8467 2770 8667 2970
rect 8723 2770 8923 2970
rect 8979 2770 9179 2970
rect 9235 2770 9435 2970
rect 7610 2477 8610 2597
rect -408 1863 -288 2003
rect -232 1863 -112 2003
rect -56 1863 64 2003
rect 7623 1707 7743 2307
rect 7799 1707 7919 2307
rect 8723 1708 8843 2708
rect 8956 2497 9556 2597
rect 9815 2478 9935 2678
rect 9991 2478 10111 2678
rect 10195 2478 10315 2678
rect 10905 2527 11025 3127
rect 11081 2527 11201 3127
rect 11257 2527 11377 3127
rect 11433 2527 11553 3127
rect 11609 2527 11729 3127
rect 11785 2527 11905 3127
rect 11961 2527 12081 3127
rect 9022 1708 9142 2308
rect 9198 1708 9318 2308
rect 9709 1708 9829 2308
rect 9885 1708 10005 2308
rect 10061 1708 10181 2308
rect 10237 1708 10357 2308
rect 10829 1772 10949 2372
rect 11005 1772 11125 2372
rect 11181 1772 11301 2372
rect 11357 1772 11477 2372
rect 11533 1772 11653 2372
rect 11709 1772 11829 2372
rect 11885 1772 12005 2372
<< mvpmos >>
rect -408 4633 -288 4833
rect -232 4633 -112 4833
rect -56 4633 64 4833
rect -408 4365 -288 4565
rect -232 4365 -112 4565
rect -56 4365 64 4565
rect -425 2907 -325 3507
rect -145 3307 -25 3507
rect -145 3039 -25 3239
rect 1159 3203 1259 4203
rect 1315 3203 1415 4203
rect 1581 3203 1681 4203
rect 1737 3203 1837 4203
rect 1893 3203 1993 4203
rect 2049 3203 2149 4203
rect 2205 3203 2305 4203
rect 2361 3203 2461 4203
rect 2517 3203 2617 4203
rect 2673 3203 2773 4203
rect 3025 3203 3125 4203
rect 3181 3203 3281 4203
rect 3337 3203 3437 4203
rect 3493 3203 3593 4203
rect 3649 3203 3749 4203
rect 3805 3203 3905 4203
rect 3961 3203 4061 4203
rect 4117 3203 4217 4203
rect 4469 3253 4569 4253
rect 4625 3253 4725 4253
rect 4781 3253 4881 4253
rect 4937 3253 5037 4253
rect 5093 3253 5193 4253
rect 5249 3253 5349 4253
rect 5405 3253 5505 4253
rect 5561 3253 5661 4253
rect 5913 3203 6013 4203
rect 6069 3203 6169 4203
rect 6225 3203 6325 4203
rect 6381 3203 6481 4203
rect 6537 3203 6637 4203
rect 6693 3203 6793 4203
rect 6849 3203 6949 4203
rect 7005 3203 7105 4203
rect 7161 3203 7261 4203
rect 7513 3603 7613 4203
rect 7655 3603 7755 4203
rect 7797 3603 7897 4203
rect 7513 3208 7613 3408
rect 7669 3208 7769 3408
rect 8026 3256 8110 4056
rect 9190 3718 9290 4318
rect 9346 3718 9446 4318
rect 9502 3718 9602 4318
rect 9782 3718 9882 4318
rect 9938 3718 10038 4318
rect 10094 3718 10194 4318
rect 10250 3718 10350 4318
rect 10530 3718 10630 4318
rect 10686 3718 10786 4318
rect 11062 4155 11862 4239
rect 12137 4036 12221 4236
rect 11062 3941 11862 4025
rect 11062 3747 11862 3831
rect 12137 3780 12221 3980
rect 1737 3025 3337 3109
rect 9815 2938 9935 3538
rect 9991 2938 10111 3538
rect 10195 2938 10315 3538
rect 11062 3521 11862 3605
rect 12137 3400 12221 3600
rect 11062 3305 11862 3389
rect -408 2469 -288 2669
rect -232 2469 -112 2669
rect -56 2469 64 2669
rect -408 2201 -288 2401
rect -232 2201 -112 2401
rect -56 2201 64 2401
rect 7467 544 7587 1544
rect 7643 544 7763 1544
rect 7819 544 7939 1544
rect 8929 944 9029 1544
rect 9085 944 9185 1544
rect 9241 944 9341 1544
rect 9397 944 9497 1544
rect 9801 944 9901 1544
rect 9957 944 10057 1544
rect 10113 944 10213 1544
rect 10269 944 10369 1544
rect 10617 1155 10717 1455
rect 10773 1155 10873 1455
rect 10929 1155 11029 1455
rect 11085 1155 11185 1455
rect 11414 1265 12214 1349
rect 10902 843 11302 927
rect 11358 843 11758 927
rect 11814 843 12214 927
rect 10451 443 10551 643
rect 10607 443 10707 643
rect 10953 559 11053 643
rect 11109 559 11209 643
rect 11389 559 11489 643
rect 11545 559 11645 643
<< pdiff >>
rect 6858 6772 12565 6784
rect 3004 5002 3020 5318
rect 4208 5002 4226 5318
rect 3004 4976 3008 5002
rect 2970 4738 3008 4976
rect 4228 4738 4260 4976
<< mvndiff >>
rect -461 4155 -408 4167
rect -461 4121 -453 4155
rect -419 4121 -408 4155
rect -461 4087 -408 4121
rect -461 4053 -453 4087
rect -419 4053 -408 4087
rect -461 4027 -408 4053
rect -288 4155 -232 4167
rect -288 4121 -277 4155
rect -243 4121 -232 4155
rect -288 4087 -232 4121
rect -288 4053 -277 4087
rect -243 4053 -232 4087
rect -288 4027 -232 4053
rect -112 4027 -56 4167
rect 64 4155 117 4167
rect 64 4121 75 4155
rect 109 4121 117 4155
rect 64 4087 117 4121
rect 64 4053 75 4087
rect 109 4053 117 4087
rect 64 4027 117 4053
rect -478 3807 -425 3845
rect -478 3773 -470 3807
rect -436 3773 -425 3807
rect -478 3761 -425 3773
rect -325 3807 -272 3845
rect -325 3773 -314 3807
rect -280 3773 -272 3807
rect -325 3761 -272 3773
rect -198 3819 -145 3845
rect -198 3785 -190 3819
rect -156 3785 -145 3819
rect -198 3751 -145 3785
rect -198 3717 -190 3751
rect -156 3717 -145 3751
rect -198 3705 -145 3717
rect -25 3819 28 3845
rect -25 3785 -14 3819
rect 20 3785 28 3819
rect -25 3751 28 3785
rect -25 3717 -14 3751
rect 20 3717 28 3751
rect -25 3705 28 3717
rect 8354 4101 8438 4109
rect 8354 4067 8366 4101
rect 8400 4067 8438 4101
rect 8354 4056 8438 4067
rect 8498 4101 8582 4109
rect 8498 4067 8510 4101
rect 8544 4067 8582 4101
rect 8498 4056 8582 4067
rect 8354 3245 8438 3256
rect 8354 3211 8366 3245
rect 8400 3211 8438 3245
rect 8354 3203 8438 3211
rect 8498 3245 8582 3256
rect 8498 3211 8510 3245
rect 8544 3211 8582 3245
rect 8498 3203 8582 3211
rect 7534 2958 7587 2970
rect 7534 2924 7542 2958
rect 7576 2924 7587 2958
rect 7534 2890 7587 2924
rect 7534 2856 7542 2890
rect 7576 2856 7587 2890
rect 7534 2822 7587 2856
rect 7534 2788 7542 2822
rect 7576 2788 7587 2822
rect 7534 2770 7587 2788
rect 7707 2958 7763 2970
rect 7707 2924 7718 2958
rect 7752 2924 7763 2958
rect 7707 2890 7763 2924
rect 7707 2856 7718 2890
rect 7752 2856 7763 2890
rect 7707 2822 7763 2856
rect 7707 2788 7718 2822
rect 7752 2788 7763 2822
rect 7707 2770 7763 2788
rect 7883 2958 7939 2970
rect 7883 2924 7894 2958
rect 7928 2924 7939 2958
rect 7883 2890 7939 2924
rect 7883 2856 7894 2890
rect 7928 2856 7939 2890
rect 7883 2822 7939 2856
rect 7883 2788 7894 2822
rect 7928 2788 7939 2822
rect 7883 2770 7939 2788
rect 8059 2958 8115 2970
rect 8059 2924 8070 2958
rect 8104 2924 8115 2958
rect 8059 2890 8115 2924
rect 8059 2856 8070 2890
rect 8104 2856 8115 2890
rect 8059 2822 8115 2856
rect 8059 2788 8070 2822
rect 8104 2788 8115 2822
rect 8059 2770 8115 2788
rect 8235 2958 8291 2970
rect 8235 2924 8246 2958
rect 8280 2924 8291 2958
rect 8235 2890 8291 2924
rect 8235 2856 8246 2890
rect 8280 2856 8291 2890
rect 8235 2822 8291 2856
rect 8235 2788 8246 2822
rect 8280 2788 8291 2822
rect 8235 2770 8291 2788
rect 8411 2958 8467 2970
rect 8411 2924 8422 2958
rect 8456 2924 8467 2958
rect 8411 2890 8467 2924
rect 8411 2856 8422 2890
rect 8456 2856 8467 2890
rect 8411 2822 8467 2856
rect 8411 2788 8422 2822
rect 8456 2788 8467 2822
rect 8411 2770 8467 2788
rect 8667 2958 8723 2970
rect 8667 2924 8678 2958
rect 8712 2924 8723 2958
rect 8667 2890 8723 2924
rect 8667 2856 8678 2890
rect 8712 2856 8723 2890
rect 8667 2822 8723 2856
rect 8667 2788 8678 2822
rect 8712 2788 8723 2822
rect 8667 2770 8723 2788
rect 8923 2958 8979 2970
rect 8923 2924 8934 2958
rect 8968 2924 8979 2958
rect 8923 2890 8979 2924
rect 8923 2856 8934 2890
rect 8968 2856 8979 2890
rect 8923 2822 8979 2856
rect 8923 2788 8934 2822
rect 8968 2788 8979 2822
rect 8923 2770 8979 2788
rect 9179 2958 9235 2970
rect 9179 2924 9190 2958
rect 9224 2924 9235 2958
rect 9179 2890 9235 2924
rect 9179 2856 9190 2890
rect 9224 2856 9235 2890
rect 9179 2822 9235 2856
rect 9179 2788 9190 2822
rect 9224 2788 9235 2822
rect 9179 2770 9235 2788
rect 9435 2958 9488 2970
rect 9435 2924 9446 2958
rect 9480 2924 9488 2958
rect 9435 2890 9488 2924
rect 9435 2856 9446 2890
rect 9480 2856 9488 2890
rect 9435 2822 9488 2856
rect 9435 2788 9446 2822
rect 9480 2788 9488 2822
rect 9435 2770 9488 2788
rect 8670 2696 8723 2708
rect 8670 2662 8678 2696
rect 8712 2662 8723 2696
rect 7610 2642 8610 2650
rect 7610 2608 7680 2642
rect 7714 2608 7748 2642
rect 7782 2608 7816 2642
rect 7850 2608 7884 2642
rect 7918 2608 7952 2642
rect 7986 2608 8020 2642
rect 8054 2608 8088 2642
rect 8122 2608 8156 2642
rect 8190 2608 8224 2642
rect 8258 2608 8292 2642
rect 8326 2608 8360 2642
rect 8394 2608 8428 2642
rect 8462 2608 8496 2642
rect 8530 2608 8564 2642
rect 8598 2608 8610 2642
rect 7610 2597 8610 2608
rect 8670 2628 8723 2662
rect 8670 2594 8678 2628
rect 8712 2594 8723 2628
rect 8670 2560 8723 2594
rect 8670 2526 8678 2560
rect 8712 2526 8723 2560
rect 8670 2492 8723 2526
rect 7610 2466 8610 2477
rect 7610 2432 7680 2466
rect 7714 2432 7748 2466
rect 7782 2432 7816 2466
rect 7850 2432 7884 2466
rect 7918 2432 7952 2466
rect 7986 2432 8020 2466
rect 8054 2432 8088 2466
rect 8122 2432 8156 2466
rect 8190 2432 8224 2466
rect 8258 2432 8292 2466
rect 8326 2432 8360 2466
rect 8394 2432 8428 2466
rect 8462 2432 8496 2466
rect 8530 2432 8564 2466
rect 8598 2432 8610 2466
rect 7610 2424 8610 2432
rect 8670 2458 8678 2492
rect 8712 2458 8723 2492
rect 8670 2424 8723 2458
rect 8670 2390 8678 2424
rect 8712 2390 8723 2424
rect 8670 2356 8723 2390
rect 8670 2322 8678 2356
rect 8712 2322 8723 2356
rect -461 1991 -408 2003
rect -461 1957 -453 1991
rect -419 1957 -408 1991
rect -461 1923 -408 1957
rect -461 1889 -453 1923
rect -419 1889 -408 1923
rect -461 1863 -408 1889
rect -288 1991 -232 2003
rect -288 1957 -277 1991
rect -243 1957 -232 1991
rect -288 1923 -232 1957
rect -288 1889 -277 1923
rect -243 1889 -232 1923
rect -288 1863 -232 1889
rect -112 1863 -56 2003
rect 64 1991 117 2003
rect 64 1957 75 1991
rect 109 1957 117 1991
rect 64 1923 117 1957
rect 64 1889 75 1923
rect 109 1889 117 1923
rect 64 1863 117 1889
rect 7570 2295 7623 2307
rect 7570 2261 7578 2295
rect 7612 2261 7623 2295
rect 7570 2227 7623 2261
rect 7570 2193 7578 2227
rect 7612 2193 7623 2227
rect 7570 2159 7623 2193
rect 7570 2125 7578 2159
rect 7612 2125 7623 2159
rect 7570 2091 7623 2125
rect 7570 2057 7578 2091
rect 7612 2057 7623 2091
rect 7570 2023 7623 2057
rect 7570 1989 7578 2023
rect 7612 1989 7623 2023
rect 7570 1955 7623 1989
rect 7570 1921 7578 1955
rect 7612 1921 7623 1955
rect 7570 1887 7623 1921
rect 7570 1853 7578 1887
rect 7612 1853 7623 1887
rect 7570 1819 7623 1853
rect 7570 1785 7578 1819
rect 7612 1785 7623 1819
rect 7570 1707 7623 1785
rect 7743 2295 7799 2307
rect 7743 2261 7754 2295
rect 7788 2261 7799 2295
rect 7743 2227 7799 2261
rect 7743 2193 7754 2227
rect 7788 2193 7799 2227
rect 7743 2159 7799 2193
rect 7743 2125 7754 2159
rect 7788 2125 7799 2159
rect 7743 2091 7799 2125
rect 7743 2057 7754 2091
rect 7788 2057 7799 2091
rect 7743 2023 7799 2057
rect 7743 1989 7754 2023
rect 7788 1989 7799 2023
rect 7743 1955 7799 1989
rect 7743 1921 7754 1955
rect 7788 1921 7799 1955
rect 7743 1887 7799 1921
rect 7743 1853 7754 1887
rect 7788 1853 7799 1887
rect 7743 1819 7799 1853
rect 7743 1785 7754 1819
rect 7788 1785 7799 1819
rect 7743 1707 7799 1785
rect 7919 2295 7972 2307
rect 7919 2261 7930 2295
rect 7964 2261 7972 2295
rect 7919 2227 7972 2261
rect 7919 2193 7930 2227
rect 7964 2193 7972 2227
rect 7919 2159 7972 2193
rect 7919 2125 7930 2159
rect 7964 2125 7972 2159
rect 7919 2091 7972 2125
rect 7919 2057 7930 2091
rect 7964 2057 7972 2091
rect 7919 2023 7972 2057
rect 7919 1989 7930 2023
rect 7964 1989 7972 2023
rect 7919 1955 7972 1989
rect 7919 1921 7930 1955
rect 7964 1921 7972 1955
rect 7919 1887 7972 1921
rect 7919 1853 7930 1887
rect 7964 1853 7972 1887
rect 7919 1819 7972 1853
rect 7919 1785 7930 1819
rect 7964 1785 7972 1819
rect 7919 1707 7972 1785
rect 8670 2288 8723 2322
rect 8670 2254 8678 2288
rect 8712 2254 8723 2288
rect 8670 2220 8723 2254
rect 8670 2186 8678 2220
rect 8712 2186 8723 2220
rect 8670 2152 8723 2186
rect 8670 2118 8678 2152
rect 8712 2118 8723 2152
rect 8670 2084 8723 2118
rect 8670 2050 8678 2084
rect 8712 2050 8723 2084
rect 8670 2016 8723 2050
rect 8670 1982 8678 2016
rect 8712 1982 8723 2016
rect 8670 1948 8723 1982
rect 8670 1914 8678 1948
rect 8712 1914 8723 1948
rect 8670 1880 8723 1914
rect 8670 1846 8678 1880
rect 8712 1846 8723 1880
rect 8670 1812 8723 1846
rect 8670 1778 8678 1812
rect 8712 1778 8723 1812
rect 8670 1708 8723 1778
rect 8843 2696 8896 2708
rect 8843 2662 8854 2696
rect 8888 2662 8896 2696
rect 8843 2628 8896 2662
rect 9748 2666 9815 2678
rect 8843 2594 8854 2628
rect 8888 2594 8896 2628
rect 8956 2642 9556 2650
rect 8956 2608 8968 2642
rect 9002 2608 9036 2642
rect 9070 2608 9104 2642
rect 9138 2608 9172 2642
rect 9206 2608 9240 2642
rect 9274 2608 9308 2642
rect 9342 2608 9376 2642
rect 9410 2608 9444 2642
rect 9478 2608 9556 2642
rect 9748 2632 9756 2666
rect 9790 2632 9815 2666
rect 8956 2597 9556 2608
rect 8843 2560 8896 2594
rect 8843 2526 8854 2560
rect 8888 2526 8896 2560
rect 8843 2492 8896 2526
rect 8843 2458 8854 2492
rect 8888 2458 8896 2492
rect 8843 2424 8896 2458
rect 8956 2486 9556 2497
rect 9748 2598 9815 2632
rect 9748 2564 9756 2598
rect 9790 2564 9815 2598
rect 9748 2530 9815 2564
rect 9748 2496 9756 2530
rect 9790 2496 9815 2530
rect 8956 2452 8968 2486
rect 9002 2452 9036 2486
rect 9070 2452 9104 2486
rect 9138 2452 9172 2486
rect 9206 2452 9240 2486
rect 9274 2452 9308 2486
rect 9342 2452 9376 2486
rect 9410 2452 9444 2486
rect 9478 2452 9556 2486
rect 9748 2478 9815 2496
rect 9935 2666 9991 2678
rect 9935 2632 9946 2666
rect 9980 2632 9991 2666
rect 9935 2598 9991 2632
rect 9935 2564 9946 2598
rect 9980 2564 9991 2598
rect 9935 2530 9991 2564
rect 9935 2496 9946 2530
rect 9980 2496 9991 2530
rect 9935 2478 9991 2496
rect 10111 2666 10195 2678
rect 10111 2632 10136 2666
rect 10170 2632 10195 2666
rect 10111 2598 10195 2632
rect 10111 2564 10136 2598
rect 10170 2564 10195 2598
rect 10111 2530 10195 2564
rect 10111 2496 10136 2530
rect 10170 2496 10195 2530
rect 10111 2478 10195 2496
rect 10315 2666 10368 2678
rect 10315 2632 10326 2666
rect 10360 2632 10368 2666
rect 10315 2598 10368 2632
rect 10315 2564 10326 2598
rect 10360 2564 10368 2598
rect 10315 2530 10368 2564
rect 10852 3049 10905 3127
rect 10852 3015 10860 3049
rect 10894 3015 10905 3049
rect 10852 2981 10905 3015
rect 10852 2947 10860 2981
rect 10894 2947 10905 2981
rect 10852 2913 10905 2947
rect 10852 2879 10860 2913
rect 10894 2879 10905 2913
rect 10852 2845 10905 2879
rect 10852 2811 10860 2845
rect 10894 2811 10905 2845
rect 10852 2777 10905 2811
rect 10852 2743 10860 2777
rect 10894 2743 10905 2777
rect 10852 2709 10905 2743
rect 10852 2675 10860 2709
rect 10894 2675 10905 2709
rect 10852 2641 10905 2675
rect 10852 2607 10860 2641
rect 10894 2607 10905 2641
rect 10852 2573 10905 2607
rect 10852 2539 10860 2573
rect 10894 2539 10905 2573
rect 10315 2496 10326 2530
rect 10360 2496 10368 2530
rect 10852 2527 10905 2539
rect 11025 3049 11081 3127
rect 11025 3015 11036 3049
rect 11070 3015 11081 3049
rect 11025 2981 11081 3015
rect 11025 2947 11036 2981
rect 11070 2947 11081 2981
rect 11025 2913 11081 2947
rect 11025 2879 11036 2913
rect 11070 2879 11081 2913
rect 11025 2845 11081 2879
rect 11025 2811 11036 2845
rect 11070 2811 11081 2845
rect 11025 2777 11081 2811
rect 11025 2743 11036 2777
rect 11070 2743 11081 2777
rect 11025 2709 11081 2743
rect 11025 2675 11036 2709
rect 11070 2675 11081 2709
rect 11025 2641 11081 2675
rect 11025 2607 11036 2641
rect 11070 2607 11081 2641
rect 11025 2573 11081 2607
rect 11025 2539 11036 2573
rect 11070 2539 11081 2573
rect 11025 2527 11081 2539
rect 11201 3049 11257 3127
rect 11201 3015 11212 3049
rect 11246 3015 11257 3049
rect 11201 2981 11257 3015
rect 11201 2947 11212 2981
rect 11246 2947 11257 2981
rect 11201 2913 11257 2947
rect 11201 2879 11212 2913
rect 11246 2879 11257 2913
rect 11201 2845 11257 2879
rect 11201 2811 11212 2845
rect 11246 2811 11257 2845
rect 11201 2777 11257 2811
rect 11201 2743 11212 2777
rect 11246 2743 11257 2777
rect 11201 2709 11257 2743
rect 11201 2675 11212 2709
rect 11246 2675 11257 2709
rect 11201 2641 11257 2675
rect 11201 2607 11212 2641
rect 11246 2607 11257 2641
rect 11201 2573 11257 2607
rect 11201 2539 11212 2573
rect 11246 2539 11257 2573
rect 11201 2527 11257 2539
rect 11377 3049 11433 3127
rect 11377 3015 11388 3049
rect 11422 3015 11433 3049
rect 11377 2981 11433 3015
rect 11377 2947 11388 2981
rect 11422 2947 11433 2981
rect 11377 2913 11433 2947
rect 11377 2879 11388 2913
rect 11422 2879 11433 2913
rect 11377 2845 11433 2879
rect 11377 2811 11388 2845
rect 11422 2811 11433 2845
rect 11377 2777 11433 2811
rect 11377 2743 11388 2777
rect 11422 2743 11433 2777
rect 11377 2709 11433 2743
rect 11377 2675 11388 2709
rect 11422 2675 11433 2709
rect 11377 2641 11433 2675
rect 11377 2607 11388 2641
rect 11422 2607 11433 2641
rect 11377 2573 11433 2607
rect 11377 2539 11388 2573
rect 11422 2539 11433 2573
rect 11377 2527 11433 2539
rect 11553 3049 11609 3127
rect 11553 3015 11564 3049
rect 11598 3015 11609 3049
rect 11553 2981 11609 3015
rect 11553 2947 11564 2981
rect 11598 2947 11609 2981
rect 11553 2913 11609 2947
rect 11553 2879 11564 2913
rect 11598 2879 11609 2913
rect 11553 2845 11609 2879
rect 11553 2811 11564 2845
rect 11598 2811 11609 2845
rect 11553 2777 11609 2811
rect 11553 2743 11564 2777
rect 11598 2743 11609 2777
rect 11553 2709 11609 2743
rect 11553 2675 11564 2709
rect 11598 2675 11609 2709
rect 11553 2641 11609 2675
rect 11553 2607 11564 2641
rect 11598 2607 11609 2641
rect 11553 2573 11609 2607
rect 11553 2539 11564 2573
rect 11598 2539 11609 2573
rect 11553 2527 11609 2539
rect 11729 3049 11785 3127
rect 11729 3015 11740 3049
rect 11774 3015 11785 3049
rect 11729 2981 11785 3015
rect 11729 2947 11740 2981
rect 11774 2947 11785 2981
rect 11729 2913 11785 2947
rect 11729 2879 11740 2913
rect 11774 2879 11785 2913
rect 11729 2845 11785 2879
rect 11729 2811 11740 2845
rect 11774 2811 11785 2845
rect 11729 2777 11785 2811
rect 11729 2743 11740 2777
rect 11774 2743 11785 2777
rect 11729 2709 11785 2743
rect 11729 2675 11740 2709
rect 11774 2675 11785 2709
rect 11729 2641 11785 2675
rect 11729 2607 11740 2641
rect 11774 2607 11785 2641
rect 11729 2573 11785 2607
rect 11729 2539 11740 2573
rect 11774 2539 11785 2573
rect 11729 2527 11785 2539
rect 11905 3049 11961 3127
rect 11905 3015 11916 3049
rect 11950 3015 11961 3049
rect 11905 2981 11961 3015
rect 11905 2947 11916 2981
rect 11950 2947 11961 2981
rect 11905 2913 11961 2947
rect 11905 2879 11916 2913
rect 11950 2879 11961 2913
rect 11905 2845 11961 2879
rect 11905 2811 11916 2845
rect 11950 2811 11961 2845
rect 11905 2777 11961 2811
rect 11905 2743 11916 2777
rect 11950 2743 11961 2777
rect 11905 2709 11961 2743
rect 11905 2675 11916 2709
rect 11950 2675 11961 2709
rect 11905 2641 11961 2675
rect 11905 2607 11916 2641
rect 11950 2607 11961 2641
rect 11905 2573 11961 2607
rect 11905 2539 11916 2573
rect 11950 2539 11961 2573
rect 11905 2527 11961 2539
rect 12081 3049 12134 3127
rect 12081 3015 12092 3049
rect 12126 3015 12134 3049
rect 12081 2981 12134 3015
rect 12081 2947 12092 2981
rect 12126 2947 12134 2981
rect 12081 2913 12134 2947
rect 12081 2879 12092 2913
rect 12126 2879 12134 2913
rect 12081 2845 12134 2879
rect 12081 2811 12092 2845
rect 12126 2811 12134 2845
rect 12081 2777 12134 2811
rect 12081 2743 12092 2777
rect 12126 2743 12134 2777
rect 12081 2709 12134 2743
rect 12081 2675 12092 2709
rect 12126 2675 12134 2709
rect 12081 2641 12134 2675
rect 12081 2607 12092 2641
rect 12126 2607 12134 2641
rect 12081 2573 12134 2607
rect 12081 2539 12092 2573
rect 12126 2539 12134 2573
rect 12081 2527 12134 2539
rect 10315 2478 10368 2496
rect 8956 2444 9556 2452
rect 8843 2390 8854 2424
rect 8888 2390 8896 2424
rect 8843 2356 8896 2390
rect 8843 2322 8854 2356
rect 8888 2322 8896 2356
rect 8843 2288 8896 2322
rect 10776 2360 10829 2372
rect 10776 2326 10784 2360
rect 10818 2326 10829 2360
rect 8843 2254 8854 2288
rect 8888 2254 8896 2288
rect 8843 2220 8896 2254
rect 8843 2186 8854 2220
rect 8888 2186 8896 2220
rect 8843 2152 8896 2186
rect 8843 2118 8854 2152
rect 8888 2118 8896 2152
rect 8843 2084 8896 2118
rect 8843 2050 8854 2084
rect 8888 2050 8896 2084
rect 8843 2016 8896 2050
rect 8843 1982 8854 2016
rect 8888 1982 8896 2016
rect 8843 1948 8896 1982
rect 8843 1914 8854 1948
rect 8888 1914 8896 1948
rect 8843 1880 8896 1914
rect 8843 1846 8854 1880
rect 8888 1846 8896 1880
rect 8843 1812 8896 1846
rect 8843 1778 8854 1812
rect 8888 1778 8896 1812
rect 8843 1708 8896 1778
rect 8969 2296 9022 2308
rect 8969 2262 8977 2296
rect 9011 2262 9022 2296
rect 8969 2228 9022 2262
rect 8969 2194 8977 2228
rect 9011 2194 9022 2228
rect 8969 2160 9022 2194
rect 8969 2126 8977 2160
rect 9011 2126 9022 2160
rect 8969 2092 9022 2126
rect 8969 2058 8977 2092
rect 9011 2058 9022 2092
rect 8969 2024 9022 2058
rect 8969 1990 8977 2024
rect 9011 1990 9022 2024
rect 8969 1956 9022 1990
rect 8969 1922 8977 1956
rect 9011 1922 9022 1956
rect 8969 1888 9022 1922
rect 8969 1854 8977 1888
rect 9011 1854 9022 1888
rect 8969 1820 9022 1854
rect 8969 1786 8977 1820
rect 9011 1786 9022 1820
rect 8969 1708 9022 1786
rect 9142 2296 9198 2308
rect 9142 2262 9153 2296
rect 9187 2262 9198 2296
rect 9142 2228 9198 2262
rect 9142 2194 9153 2228
rect 9187 2194 9198 2228
rect 9142 2160 9198 2194
rect 9142 2126 9153 2160
rect 9187 2126 9198 2160
rect 9142 2092 9198 2126
rect 9142 2058 9153 2092
rect 9187 2058 9198 2092
rect 9142 2024 9198 2058
rect 9142 1990 9153 2024
rect 9187 1990 9198 2024
rect 9142 1956 9198 1990
rect 9142 1922 9153 1956
rect 9187 1922 9198 1956
rect 9142 1888 9198 1922
rect 9142 1854 9153 1888
rect 9187 1854 9198 1888
rect 9142 1820 9198 1854
rect 9142 1786 9153 1820
rect 9187 1786 9198 1820
rect 9142 1708 9198 1786
rect 9318 2296 9371 2308
rect 9318 2262 9329 2296
rect 9363 2262 9371 2296
rect 9318 2228 9371 2262
rect 9318 2194 9329 2228
rect 9363 2194 9371 2228
rect 9318 2160 9371 2194
rect 9318 2126 9329 2160
rect 9363 2126 9371 2160
rect 9318 2092 9371 2126
rect 9318 2058 9329 2092
rect 9363 2058 9371 2092
rect 9318 2024 9371 2058
rect 9318 1990 9329 2024
rect 9363 1990 9371 2024
rect 9318 1956 9371 1990
rect 9318 1922 9329 1956
rect 9363 1922 9371 1956
rect 9318 1888 9371 1922
rect 9318 1854 9329 1888
rect 9363 1854 9371 1888
rect 9318 1820 9371 1854
rect 9318 1786 9329 1820
rect 9363 1786 9371 1820
rect 9318 1708 9371 1786
rect 9656 2296 9709 2308
rect 9656 2262 9664 2296
rect 9698 2262 9709 2296
rect 9656 2228 9709 2262
rect 9656 2194 9664 2228
rect 9698 2194 9709 2228
rect 9656 2160 9709 2194
rect 9656 2126 9664 2160
rect 9698 2126 9709 2160
rect 9656 2092 9709 2126
rect 9656 2058 9664 2092
rect 9698 2058 9709 2092
rect 9656 2024 9709 2058
rect 9656 1990 9664 2024
rect 9698 1990 9709 2024
rect 9656 1956 9709 1990
rect 9656 1922 9664 1956
rect 9698 1922 9709 1956
rect 9656 1888 9709 1922
rect 9656 1854 9664 1888
rect 9698 1854 9709 1888
rect 9656 1820 9709 1854
rect 9656 1786 9664 1820
rect 9698 1786 9709 1820
rect 9656 1708 9709 1786
rect 9829 2296 9885 2308
rect 9829 2262 9840 2296
rect 9874 2262 9885 2296
rect 9829 2228 9885 2262
rect 9829 2194 9840 2228
rect 9874 2194 9885 2228
rect 9829 2160 9885 2194
rect 9829 2126 9840 2160
rect 9874 2126 9885 2160
rect 9829 2092 9885 2126
rect 9829 2058 9840 2092
rect 9874 2058 9885 2092
rect 9829 2024 9885 2058
rect 9829 1990 9840 2024
rect 9874 1990 9885 2024
rect 9829 1956 9885 1990
rect 9829 1922 9840 1956
rect 9874 1922 9885 1956
rect 9829 1888 9885 1922
rect 9829 1854 9840 1888
rect 9874 1854 9885 1888
rect 9829 1820 9885 1854
rect 9829 1786 9840 1820
rect 9874 1786 9885 1820
rect 9829 1708 9885 1786
rect 10005 2296 10061 2308
rect 10005 2262 10016 2296
rect 10050 2262 10061 2296
rect 10005 2228 10061 2262
rect 10005 2194 10016 2228
rect 10050 2194 10061 2228
rect 10005 2160 10061 2194
rect 10005 2126 10016 2160
rect 10050 2126 10061 2160
rect 10005 2092 10061 2126
rect 10005 2058 10016 2092
rect 10050 2058 10061 2092
rect 10005 2024 10061 2058
rect 10005 1990 10016 2024
rect 10050 1990 10061 2024
rect 10005 1956 10061 1990
rect 10005 1922 10016 1956
rect 10050 1922 10061 1956
rect 10005 1888 10061 1922
rect 10005 1854 10016 1888
rect 10050 1854 10061 1888
rect 10005 1820 10061 1854
rect 10005 1786 10016 1820
rect 10050 1786 10061 1820
rect 10005 1708 10061 1786
rect 10181 2296 10237 2308
rect 10181 2262 10192 2296
rect 10226 2262 10237 2296
rect 10181 2228 10237 2262
rect 10181 2194 10192 2228
rect 10226 2194 10237 2228
rect 10181 2160 10237 2194
rect 10181 2126 10192 2160
rect 10226 2126 10237 2160
rect 10181 2092 10237 2126
rect 10181 2058 10192 2092
rect 10226 2058 10237 2092
rect 10181 2024 10237 2058
rect 10181 1990 10192 2024
rect 10226 1990 10237 2024
rect 10181 1956 10237 1990
rect 10181 1922 10192 1956
rect 10226 1922 10237 1956
rect 10181 1888 10237 1922
rect 10181 1854 10192 1888
rect 10226 1854 10237 1888
rect 10181 1820 10237 1854
rect 10181 1786 10192 1820
rect 10226 1786 10237 1820
rect 10181 1708 10237 1786
rect 10357 2296 10410 2308
rect 10357 2262 10368 2296
rect 10402 2262 10410 2296
rect 10357 2228 10410 2262
rect 10357 2194 10368 2228
rect 10402 2194 10410 2228
rect 10357 2160 10410 2194
rect 10357 2126 10368 2160
rect 10402 2126 10410 2160
rect 10357 2092 10410 2126
rect 10357 2058 10368 2092
rect 10402 2058 10410 2092
rect 10357 2024 10410 2058
rect 10357 1990 10368 2024
rect 10402 1990 10410 2024
rect 10357 1956 10410 1990
rect 10357 1922 10368 1956
rect 10402 1922 10410 1956
rect 10357 1888 10410 1922
rect 10357 1854 10368 1888
rect 10402 1854 10410 1888
rect 10357 1820 10410 1854
rect 10357 1786 10368 1820
rect 10402 1786 10410 1820
rect 10357 1708 10410 1786
rect 10776 2292 10829 2326
rect 10776 2258 10784 2292
rect 10818 2258 10829 2292
rect 10776 2224 10829 2258
rect 10776 2190 10784 2224
rect 10818 2190 10829 2224
rect 10776 2156 10829 2190
rect 10776 2122 10784 2156
rect 10818 2122 10829 2156
rect 10776 2088 10829 2122
rect 10776 2054 10784 2088
rect 10818 2054 10829 2088
rect 10776 2020 10829 2054
rect 10776 1986 10784 2020
rect 10818 1986 10829 2020
rect 10776 1952 10829 1986
rect 10776 1918 10784 1952
rect 10818 1918 10829 1952
rect 10776 1884 10829 1918
rect 10776 1850 10784 1884
rect 10818 1850 10829 1884
rect 10776 1772 10829 1850
rect 10949 2360 11005 2372
rect 10949 2326 10960 2360
rect 10994 2326 11005 2360
rect 10949 2292 11005 2326
rect 10949 2258 10960 2292
rect 10994 2258 11005 2292
rect 10949 2224 11005 2258
rect 10949 2190 10960 2224
rect 10994 2190 11005 2224
rect 10949 2156 11005 2190
rect 10949 2122 10960 2156
rect 10994 2122 11005 2156
rect 10949 2088 11005 2122
rect 10949 2054 10960 2088
rect 10994 2054 11005 2088
rect 10949 2020 11005 2054
rect 10949 1986 10960 2020
rect 10994 1986 11005 2020
rect 10949 1952 11005 1986
rect 10949 1918 10960 1952
rect 10994 1918 11005 1952
rect 10949 1884 11005 1918
rect 10949 1850 10960 1884
rect 10994 1850 11005 1884
rect 10949 1772 11005 1850
rect 11125 2360 11181 2372
rect 11125 2326 11136 2360
rect 11170 2326 11181 2360
rect 11125 2292 11181 2326
rect 11125 2258 11136 2292
rect 11170 2258 11181 2292
rect 11125 2224 11181 2258
rect 11125 2190 11136 2224
rect 11170 2190 11181 2224
rect 11125 2156 11181 2190
rect 11125 2122 11136 2156
rect 11170 2122 11181 2156
rect 11125 2088 11181 2122
rect 11125 2054 11136 2088
rect 11170 2054 11181 2088
rect 11125 2020 11181 2054
rect 11125 1986 11136 2020
rect 11170 1986 11181 2020
rect 11125 1952 11181 1986
rect 11125 1918 11136 1952
rect 11170 1918 11181 1952
rect 11125 1884 11181 1918
rect 11125 1850 11136 1884
rect 11170 1850 11181 1884
rect 11125 1772 11181 1850
rect 11301 2360 11357 2372
rect 11301 2326 11312 2360
rect 11346 2326 11357 2360
rect 11301 2292 11357 2326
rect 11301 2258 11312 2292
rect 11346 2258 11357 2292
rect 11301 2224 11357 2258
rect 11301 2190 11312 2224
rect 11346 2190 11357 2224
rect 11301 2156 11357 2190
rect 11301 2122 11312 2156
rect 11346 2122 11357 2156
rect 11301 2088 11357 2122
rect 11301 2054 11312 2088
rect 11346 2054 11357 2088
rect 11301 2020 11357 2054
rect 11301 1986 11312 2020
rect 11346 1986 11357 2020
rect 11301 1952 11357 1986
rect 11301 1918 11312 1952
rect 11346 1918 11357 1952
rect 11301 1884 11357 1918
rect 11301 1850 11312 1884
rect 11346 1850 11357 1884
rect 11301 1772 11357 1850
rect 11477 2360 11533 2372
rect 11477 2326 11488 2360
rect 11522 2326 11533 2360
rect 11477 2292 11533 2326
rect 11477 2258 11488 2292
rect 11522 2258 11533 2292
rect 11477 2224 11533 2258
rect 11477 2190 11488 2224
rect 11522 2190 11533 2224
rect 11477 2156 11533 2190
rect 11477 2122 11488 2156
rect 11522 2122 11533 2156
rect 11477 2088 11533 2122
rect 11477 2054 11488 2088
rect 11522 2054 11533 2088
rect 11477 2020 11533 2054
rect 11477 1986 11488 2020
rect 11522 1986 11533 2020
rect 11477 1952 11533 1986
rect 11477 1918 11488 1952
rect 11522 1918 11533 1952
rect 11477 1884 11533 1918
rect 11477 1850 11488 1884
rect 11522 1850 11533 1884
rect 11477 1772 11533 1850
rect 11653 2360 11709 2372
rect 11653 2326 11664 2360
rect 11698 2326 11709 2360
rect 11653 2292 11709 2326
rect 11653 2258 11664 2292
rect 11698 2258 11709 2292
rect 11653 2224 11709 2258
rect 11653 2190 11664 2224
rect 11698 2190 11709 2224
rect 11653 2156 11709 2190
rect 11653 2122 11664 2156
rect 11698 2122 11709 2156
rect 11653 2088 11709 2122
rect 11653 2054 11664 2088
rect 11698 2054 11709 2088
rect 11653 2020 11709 2054
rect 11653 1986 11664 2020
rect 11698 1986 11709 2020
rect 11653 1952 11709 1986
rect 11653 1918 11664 1952
rect 11698 1918 11709 1952
rect 11653 1884 11709 1918
rect 11653 1850 11664 1884
rect 11698 1850 11709 1884
rect 11653 1772 11709 1850
rect 11829 2360 11885 2372
rect 11829 2326 11840 2360
rect 11874 2326 11885 2360
rect 11829 2292 11885 2326
rect 11829 2258 11840 2292
rect 11874 2258 11885 2292
rect 11829 2224 11885 2258
rect 11829 2190 11840 2224
rect 11874 2190 11885 2224
rect 11829 2156 11885 2190
rect 11829 2122 11840 2156
rect 11874 2122 11885 2156
rect 11829 2088 11885 2122
rect 11829 2054 11840 2088
rect 11874 2054 11885 2088
rect 11829 2020 11885 2054
rect 11829 1986 11840 2020
rect 11874 1986 11885 2020
rect 11829 1952 11885 1986
rect 11829 1918 11840 1952
rect 11874 1918 11885 1952
rect 11829 1884 11885 1918
rect 11829 1850 11840 1884
rect 11874 1850 11885 1884
rect 11829 1772 11885 1850
rect 12005 2360 12058 2372
rect 12005 2326 12016 2360
rect 12050 2326 12058 2360
rect 12005 2292 12058 2326
rect 12005 2258 12016 2292
rect 12050 2258 12058 2292
rect 12005 2224 12058 2258
rect 12005 2190 12016 2224
rect 12050 2190 12058 2224
rect 12005 2156 12058 2190
rect 12005 2122 12016 2156
rect 12050 2122 12058 2156
rect 12005 2088 12058 2122
rect 12005 2054 12016 2088
rect 12050 2054 12058 2088
rect 12005 2020 12058 2054
rect 12005 1986 12016 2020
rect 12050 1986 12058 2020
rect 12005 1952 12058 1986
rect 12005 1918 12016 1952
rect 12050 1918 12058 1952
rect 12005 1884 12058 1918
rect 12005 1850 12016 1884
rect 12050 1850 12058 1884
rect 12005 1772 12058 1850
<< mvpdiff >>
rect -461 4815 -408 4833
rect -461 4781 -453 4815
rect -419 4781 -408 4815
rect -461 4747 -408 4781
rect -461 4713 -453 4747
rect -419 4713 -408 4747
rect -461 4679 -408 4713
rect -461 4645 -453 4679
rect -419 4645 -408 4679
rect -461 4633 -408 4645
rect -288 4815 -232 4833
rect -288 4781 -277 4815
rect -243 4781 -232 4815
rect -288 4747 -232 4781
rect -288 4713 -277 4747
rect -243 4713 -232 4747
rect -288 4679 -232 4713
rect -288 4645 -277 4679
rect -243 4645 -232 4679
rect -288 4633 -232 4645
rect -112 4815 -56 4833
rect -112 4781 -101 4815
rect -67 4781 -56 4815
rect -112 4747 -56 4781
rect -112 4713 -101 4747
rect -67 4713 -56 4747
rect -112 4679 -56 4713
rect -112 4645 -101 4679
rect -67 4645 -56 4679
rect -112 4633 -56 4645
rect 64 4815 117 4833
rect 64 4781 75 4815
rect 109 4781 117 4815
rect 64 4747 117 4781
rect 64 4713 75 4747
rect 109 4713 117 4747
rect 64 4679 117 4713
rect 64 4645 75 4679
rect 109 4645 117 4679
rect 64 4633 117 4645
rect -461 4553 -408 4565
rect -461 4519 -453 4553
rect -419 4519 -408 4553
rect -461 4485 -408 4519
rect -461 4451 -453 4485
rect -419 4451 -408 4485
rect -461 4417 -408 4451
rect -461 4383 -453 4417
rect -419 4383 -408 4417
rect -461 4365 -408 4383
rect -288 4553 -232 4565
rect -288 4519 -277 4553
rect -243 4519 -232 4553
rect -288 4485 -232 4519
rect -288 4451 -277 4485
rect -243 4451 -232 4485
rect -288 4417 -232 4451
rect -288 4383 -277 4417
rect -243 4383 -232 4417
rect -288 4365 -232 4383
rect -112 4553 -56 4565
rect -112 4519 -101 4553
rect -67 4519 -56 4553
rect -112 4485 -56 4519
rect -112 4451 -101 4485
rect -67 4451 -56 4485
rect -112 4417 -56 4451
rect -112 4383 -101 4417
rect -67 4383 -56 4417
rect -112 4365 -56 4383
rect 64 4553 117 4565
rect 64 4519 75 4553
rect 109 4519 117 4553
rect 64 4485 117 4519
rect 64 4451 75 4485
rect 109 4451 117 4485
rect 64 4417 117 4451
rect 64 4383 75 4417
rect 109 4383 117 4417
rect 64 4365 117 4383
rect 9137 4306 9190 4318
rect -478 3429 -425 3507
rect -478 3395 -470 3429
rect -436 3395 -425 3429
rect -478 3361 -425 3395
rect -478 3327 -470 3361
rect -436 3327 -425 3361
rect -478 3293 -425 3327
rect -478 3259 -470 3293
rect -436 3259 -425 3293
rect -478 3225 -425 3259
rect -478 3191 -470 3225
rect -436 3191 -425 3225
rect -478 3157 -425 3191
rect -478 3123 -470 3157
rect -436 3123 -425 3157
rect -478 3089 -425 3123
rect -478 3055 -470 3089
rect -436 3055 -425 3089
rect -478 3021 -425 3055
rect -478 2987 -470 3021
rect -436 2987 -425 3021
rect -478 2953 -425 2987
rect -478 2919 -470 2953
rect -436 2919 -425 2953
rect -478 2907 -425 2919
rect -325 3429 -272 3507
rect -325 3395 -314 3429
rect -280 3395 -272 3429
rect -325 3361 -272 3395
rect -325 3327 -314 3361
rect -280 3327 -272 3361
rect -325 3293 -272 3327
rect -198 3489 -145 3507
rect -198 3455 -190 3489
rect -156 3455 -145 3489
rect -198 3421 -145 3455
rect -198 3387 -190 3421
rect -156 3387 -145 3421
rect -198 3353 -145 3387
rect -198 3319 -190 3353
rect -156 3319 -145 3353
rect -198 3307 -145 3319
rect -25 3489 28 3507
rect -25 3455 -14 3489
rect 20 3455 28 3489
rect -25 3421 28 3455
rect -25 3387 -14 3421
rect 20 3387 28 3421
rect -25 3353 28 3387
rect -25 3319 -14 3353
rect 20 3319 28 3353
rect -25 3307 28 3319
rect -325 3259 -314 3293
rect -280 3259 -272 3293
rect -325 3225 -272 3259
rect -325 3191 -314 3225
rect -280 3191 -272 3225
rect -325 3157 -272 3191
rect -325 3123 -314 3157
rect -280 3123 -272 3157
rect -325 3089 -272 3123
rect -325 3055 -314 3089
rect -280 3055 -272 3089
rect -325 3021 -272 3055
rect -198 3227 -145 3239
rect -198 3193 -190 3227
rect -156 3193 -145 3227
rect -198 3159 -145 3193
rect -198 3125 -190 3159
rect -156 3125 -145 3159
rect -198 3091 -145 3125
rect -198 3057 -190 3091
rect -156 3057 -145 3091
rect -198 3039 -145 3057
rect -25 3227 28 3239
rect -25 3193 -14 3227
rect 20 3193 28 3227
rect -25 3159 28 3193
rect -25 3125 -14 3159
rect 20 3125 28 3159
rect -25 3091 28 3125
rect -25 3057 -14 3091
rect 20 3057 28 3091
rect -25 3039 28 3057
rect 1106 4133 1159 4203
rect 1106 4099 1114 4133
rect 1148 4099 1159 4133
rect 1106 4065 1159 4099
rect 1106 4031 1114 4065
rect 1148 4031 1159 4065
rect 1106 3997 1159 4031
rect 1106 3963 1114 3997
rect 1148 3963 1159 3997
rect 1106 3929 1159 3963
rect 1106 3895 1114 3929
rect 1148 3895 1159 3929
rect 1106 3861 1159 3895
rect 1106 3827 1114 3861
rect 1148 3827 1159 3861
rect 1106 3793 1159 3827
rect 1106 3759 1114 3793
rect 1148 3759 1159 3793
rect 1106 3725 1159 3759
rect 1106 3691 1114 3725
rect 1148 3691 1159 3725
rect 1106 3657 1159 3691
rect 1106 3623 1114 3657
rect 1148 3623 1159 3657
rect 1106 3589 1159 3623
rect 1106 3555 1114 3589
rect 1148 3555 1159 3589
rect 1106 3521 1159 3555
rect 1106 3487 1114 3521
rect 1148 3487 1159 3521
rect 1106 3453 1159 3487
rect 1106 3419 1114 3453
rect 1148 3419 1159 3453
rect 1106 3385 1159 3419
rect 1106 3351 1114 3385
rect 1148 3351 1159 3385
rect 1106 3317 1159 3351
rect 1106 3283 1114 3317
rect 1148 3283 1159 3317
rect 1106 3249 1159 3283
rect 1106 3215 1114 3249
rect 1148 3215 1159 3249
rect 1106 3203 1159 3215
rect 1259 4133 1315 4203
rect 1259 4099 1270 4133
rect 1304 4099 1315 4133
rect 1259 4065 1315 4099
rect 1259 4031 1270 4065
rect 1304 4031 1315 4065
rect 1259 3997 1315 4031
rect 1259 3963 1270 3997
rect 1304 3963 1315 3997
rect 1259 3929 1315 3963
rect 1259 3895 1270 3929
rect 1304 3895 1315 3929
rect 1259 3861 1315 3895
rect 1259 3827 1270 3861
rect 1304 3827 1315 3861
rect 1259 3793 1315 3827
rect 1259 3759 1270 3793
rect 1304 3759 1315 3793
rect 1259 3725 1315 3759
rect 1259 3691 1270 3725
rect 1304 3691 1315 3725
rect 1259 3657 1315 3691
rect 1259 3623 1270 3657
rect 1304 3623 1315 3657
rect 1259 3589 1315 3623
rect 1259 3555 1270 3589
rect 1304 3555 1315 3589
rect 1259 3521 1315 3555
rect 1259 3487 1270 3521
rect 1304 3487 1315 3521
rect 1259 3453 1315 3487
rect 1259 3419 1270 3453
rect 1304 3419 1315 3453
rect 1259 3385 1315 3419
rect 1259 3351 1270 3385
rect 1304 3351 1315 3385
rect 1259 3317 1315 3351
rect 1259 3283 1270 3317
rect 1304 3283 1315 3317
rect 1259 3249 1315 3283
rect 1259 3215 1270 3249
rect 1304 3215 1315 3249
rect 1259 3203 1315 3215
rect 1415 4133 1468 4203
rect 1415 4099 1426 4133
rect 1460 4099 1468 4133
rect 1415 4065 1468 4099
rect 1415 4031 1426 4065
rect 1460 4031 1468 4065
rect 1415 3997 1468 4031
rect 1415 3963 1426 3997
rect 1460 3963 1468 3997
rect 1415 3929 1468 3963
rect 1415 3895 1426 3929
rect 1460 3895 1468 3929
rect 1415 3861 1468 3895
rect 1415 3827 1426 3861
rect 1460 3827 1468 3861
rect 1415 3793 1468 3827
rect 1415 3759 1426 3793
rect 1460 3759 1468 3793
rect 1415 3725 1468 3759
rect 1415 3691 1426 3725
rect 1460 3691 1468 3725
rect 1415 3657 1468 3691
rect 1415 3623 1426 3657
rect 1460 3623 1468 3657
rect 1415 3589 1468 3623
rect 1415 3555 1426 3589
rect 1460 3555 1468 3589
rect 1415 3521 1468 3555
rect 1415 3487 1426 3521
rect 1460 3487 1468 3521
rect 1415 3453 1468 3487
rect 1415 3419 1426 3453
rect 1460 3419 1468 3453
rect 1415 3385 1468 3419
rect 1415 3351 1426 3385
rect 1460 3351 1468 3385
rect 1415 3317 1468 3351
rect 1415 3283 1426 3317
rect 1460 3283 1468 3317
rect 1415 3249 1468 3283
rect 1415 3215 1426 3249
rect 1460 3215 1468 3249
rect 1415 3203 1468 3215
rect 1528 4133 1581 4203
rect 1528 4099 1536 4133
rect 1570 4099 1581 4133
rect 1528 4065 1581 4099
rect 1528 4031 1536 4065
rect 1570 4031 1581 4065
rect 1528 3997 1581 4031
rect 1528 3963 1536 3997
rect 1570 3963 1581 3997
rect 1528 3929 1581 3963
rect 1528 3895 1536 3929
rect 1570 3895 1581 3929
rect 1528 3861 1581 3895
rect 1528 3827 1536 3861
rect 1570 3827 1581 3861
rect 1528 3793 1581 3827
rect 1528 3759 1536 3793
rect 1570 3759 1581 3793
rect 1528 3725 1581 3759
rect 1528 3691 1536 3725
rect 1570 3691 1581 3725
rect 1528 3657 1581 3691
rect 1528 3623 1536 3657
rect 1570 3623 1581 3657
rect 1528 3589 1581 3623
rect 1528 3555 1536 3589
rect 1570 3555 1581 3589
rect 1528 3521 1581 3555
rect 1528 3487 1536 3521
rect 1570 3487 1581 3521
rect 1528 3453 1581 3487
rect 1528 3419 1536 3453
rect 1570 3419 1581 3453
rect 1528 3385 1581 3419
rect 1528 3351 1536 3385
rect 1570 3351 1581 3385
rect 1528 3317 1581 3351
rect 1528 3283 1536 3317
rect 1570 3283 1581 3317
rect 1528 3249 1581 3283
rect 1528 3215 1536 3249
rect 1570 3215 1581 3249
rect 1528 3203 1581 3215
rect 1681 4133 1737 4203
rect 1681 4099 1692 4133
rect 1726 4099 1737 4133
rect 1681 4065 1737 4099
rect 1681 4031 1692 4065
rect 1726 4031 1737 4065
rect 1681 3997 1737 4031
rect 1681 3963 1692 3997
rect 1726 3963 1737 3997
rect 1681 3929 1737 3963
rect 1681 3895 1692 3929
rect 1726 3895 1737 3929
rect 1681 3861 1737 3895
rect 1681 3827 1692 3861
rect 1726 3827 1737 3861
rect 1681 3793 1737 3827
rect 1681 3759 1692 3793
rect 1726 3759 1737 3793
rect 1681 3725 1737 3759
rect 1681 3691 1692 3725
rect 1726 3691 1737 3725
rect 1681 3657 1737 3691
rect 1681 3623 1692 3657
rect 1726 3623 1737 3657
rect 1681 3589 1737 3623
rect 1681 3555 1692 3589
rect 1726 3555 1737 3589
rect 1681 3521 1737 3555
rect 1681 3487 1692 3521
rect 1726 3487 1737 3521
rect 1681 3453 1737 3487
rect 1681 3419 1692 3453
rect 1726 3419 1737 3453
rect 1681 3385 1737 3419
rect 1681 3351 1692 3385
rect 1726 3351 1737 3385
rect 1681 3317 1737 3351
rect 1681 3283 1692 3317
rect 1726 3283 1737 3317
rect 1681 3249 1737 3283
rect 1681 3215 1692 3249
rect 1726 3215 1737 3249
rect 1681 3203 1737 3215
rect 1837 4133 1893 4203
rect 1837 4099 1848 4133
rect 1882 4099 1893 4133
rect 1837 4065 1893 4099
rect 1837 4031 1848 4065
rect 1882 4031 1893 4065
rect 1837 3997 1893 4031
rect 1837 3963 1848 3997
rect 1882 3963 1893 3997
rect 1837 3929 1893 3963
rect 1837 3895 1848 3929
rect 1882 3895 1893 3929
rect 1837 3861 1893 3895
rect 1837 3827 1848 3861
rect 1882 3827 1893 3861
rect 1837 3793 1893 3827
rect 1837 3759 1848 3793
rect 1882 3759 1893 3793
rect 1837 3725 1893 3759
rect 1837 3691 1848 3725
rect 1882 3691 1893 3725
rect 1837 3657 1893 3691
rect 1837 3623 1848 3657
rect 1882 3623 1893 3657
rect 1837 3589 1893 3623
rect 1837 3555 1848 3589
rect 1882 3555 1893 3589
rect 1837 3521 1893 3555
rect 1837 3487 1848 3521
rect 1882 3487 1893 3521
rect 1837 3453 1893 3487
rect 1837 3419 1848 3453
rect 1882 3419 1893 3453
rect 1837 3385 1893 3419
rect 1837 3351 1848 3385
rect 1882 3351 1893 3385
rect 1837 3317 1893 3351
rect 1837 3283 1848 3317
rect 1882 3283 1893 3317
rect 1837 3249 1893 3283
rect 1837 3215 1848 3249
rect 1882 3215 1893 3249
rect 1837 3203 1893 3215
rect 1993 4133 2049 4203
rect 1993 4099 2004 4133
rect 2038 4099 2049 4133
rect 1993 4065 2049 4099
rect 1993 4031 2004 4065
rect 2038 4031 2049 4065
rect 1993 3997 2049 4031
rect 1993 3963 2004 3997
rect 2038 3963 2049 3997
rect 1993 3929 2049 3963
rect 1993 3895 2004 3929
rect 2038 3895 2049 3929
rect 1993 3861 2049 3895
rect 1993 3827 2004 3861
rect 2038 3827 2049 3861
rect 1993 3793 2049 3827
rect 1993 3759 2004 3793
rect 2038 3759 2049 3793
rect 1993 3725 2049 3759
rect 1993 3691 2004 3725
rect 2038 3691 2049 3725
rect 1993 3657 2049 3691
rect 1993 3623 2004 3657
rect 2038 3623 2049 3657
rect 1993 3589 2049 3623
rect 1993 3555 2004 3589
rect 2038 3555 2049 3589
rect 1993 3521 2049 3555
rect 1993 3487 2004 3521
rect 2038 3487 2049 3521
rect 1993 3453 2049 3487
rect 1993 3419 2004 3453
rect 2038 3419 2049 3453
rect 1993 3385 2049 3419
rect 1993 3351 2004 3385
rect 2038 3351 2049 3385
rect 1993 3317 2049 3351
rect 1993 3283 2004 3317
rect 2038 3283 2049 3317
rect 1993 3249 2049 3283
rect 1993 3215 2004 3249
rect 2038 3215 2049 3249
rect 1993 3203 2049 3215
rect 2149 4133 2205 4203
rect 2149 4099 2160 4133
rect 2194 4099 2205 4133
rect 2149 4065 2205 4099
rect 2149 4031 2160 4065
rect 2194 4031 2205 4065
rect 2149 3997 2205 4031
rect 2149 3963 2160 3997
rect 2194 3963 2205 3997
rect 2149 3929 2205 3963
rect 2149 3895 2160 3929
rect 2194 3895 2205 3929
rect 2149 3861 2205 3895
rect 2149 3827 2160 3861
rect 2194 3827 2205 3861
rect 2149 3793 2205 3827
rect 2149 3759 2160 3793
rect 2194 3759 2205 3793
rect 2149 3725 2205 3759
rect 2149 3691 2160 3725
rect 2194 3691 2205 3725
rect 2149 3657 2205 3691
rect 2149 3623 2160 3657
rect 2194 3623 2205 3657
rect 2149 3589 2205 3623
rect 2149 3555 2160 3589
rect 2194 3555 2205 3589
rect 2149 3521 2205 3555
rect 2149 3487 2160 3521
rect 2194 3487 2205 3521
rect 2149 3453 2205 3487
rect 2149 3419 2160 3453
rect 2194 3419 2205 3453
rect 2149 3385 2205 3419
rect 2149 3351 2160 3385
rect 2194 3351 2205 3385
rect 2149 3317 2205 3351
rect 2149 3283 2160 3317
rect 2194 3283 2205 3317
rect 2149 3249 2205 3283
rect 2149 3215 2160 3249
rect 2194 3215 2205 3249
rect 2149 3203 2205 3215
rect 2305 4133 2361 4203
rect 2305 4099 2316 4133
rect 2350 4099 2361 4133
rect 2305 4065 2361 4099
rect 2305 4031 2316 4065
rect 2350 4031 2361 4065
rect 2305 3997 2361 4031
rect 2305 3963 2316 3997
rect 2350 3963 2361 3997
rect 2305 3929 2361 3963
rect 2305 3895 2316 3929
rect 2350 3895 2361 3929
rect 2305 3861 2361 3895
rect 2305 3827 2316 3861
rect 2350 3827 2361 3861
rect 2305 3793 2361 3827
rect 2305 3759 2316 3793
rect 2350 3759 2361 3793
rect 2305 3725 2361 3759
rect 2305 3691 2316 3725
rect 2350 3691 2361 3725
rect 2305 3657 2361 3691
rect 2305 3623 2316 3657
rect 2350 3623 2361 3657
rect 2305 3589 2361 3623
rect 2305 3555 2316 3589
rect 2350 3555 2361 3589
rect 2305 3521 2361 3555
rect 2305 3487 2316 3521
rect 2350 3487 2361 3521
rect 2305 3453 2361 3487
rect 2305 3419 2316 3453
rect 2350 3419 2361 3453
rect 2305 3385 2361 3419
rect 2305 3351 2316 3385
rect 2350 3351 2361 3385
rect 2305 3317 2361 3351
rect 2305 3283 2316 3317
rect 2350 3283 2361 3317
rect 2305 3249 2361 3283
rect 2305 3215 2316 3249
rect 2350 3215 2361 3249
rect 2305 3203 2361 3215
rect 2461 4133 2517 4203
rect 2461 4099 2472 4133
rect 2506 4099 2517 4133
rect 2461 4065 2517 4099
rect 2461 4031 2472 4065
rect 2506 4031 2517 4065
rect 2461 3997 2517 4031
rect 2461 3963 2472 3997
rect 2506 3963 2517 3997
rect 2461 3929 2517 3963
rect 2461 3895 2472 3929
rect 2506 3895 2517 3929
rect 2461 3861 2517 3895
rect 2461 3827 2472 3861
rect 2506 3827 2517 3861
rect 2461 3793 2517 3827
rect 2461 3759 2472 3793
rect 2506 3759 2517 3793
rect 2461 3725 2517 3759
rect 2461 3691 2472 3725
rect 2506 3691 2517 3725
rect 2461 3657 2517 3691
rect 2461 3623 2472 3657
rect 2506 3623 2517 3657
rect 2461 3589 2517 3623
rect 2461 3555 2472 3589
rect 2506 3555 2517 3589
rect 2461 3521 2517 3555
rect 2461 3487 2472 3521
rect 2506 3487 2517 3521
rect 2461 3453 2517 3487
rect 2461 3419 2472 3453
rect 2506 3419 2517 3453
rect 2461 3385 2517 3419
rect 2461 3351 2472 3385
rect 2506 3351 2517 3385
rect 2461 3317 2517 3351
rect 2461 3283 2472 3317
rect 2506 3283 2517 3317
rect 2461 3249 2517 3283
rect 2461 3215 2472 3249
rect 2506 3215 2517 3249
rect 2461 3203 2517 3215
rect 2617 4133 2673 4203
rect 2617 4099 2628 4133
rect 2662 4099 2673 4133
rect 2617 4065 2673 4099
rect 2617 4031 2628 4065
rect 2662 4031 2673 4065
rect 2617 3997 2673 4031
rect 2617 3963 2628 3997
rect 2662 3963 2673 3997
rect 2617 3929 2673 3963
rect 2617 3895 2628 3929
rect 2662 3895 2673 3929
rect 2617 3861 2673 3895
rect 2617 3827 2628 3861
rect 2662 3827 2673 3861
rect 2617 3793 2673 3827
rect 2617 3759 2628 3793
rect 2662 3759 2673 3793
rect 2617 3725 2673 3759
rect 2617 3691 2628 3725
rect 2662 3691 2673 3725
rect 2617 3657 2673 3691
rect 2617 3623 2628 3657
rect 2662 3623 2673 3657
rect 2617 3589 2673 3623
rect 2617 3555 2628 3589
rect 2662 3555 2673 3589
rect 2617 3521 2673 3555
rect 2617 3487 2628 3521
rect 2662 3487 2673 3521
rect 2617 3453 2673 3487
rect 2617 3419 2628 3453
rect 2662 3419 2673 3453
rect 2617 3385 2673 3419
rect 2617 3351 2628 3385
rect 2662 3351 2673 3385
rect 2617 3317 2673 3351
rect 2617 3283 2628 3317
rect 2662 3283 2673 3317
rect 2617 3249 2673 3283
rect 2617 3215 2628 3249
rect 2662 3215 2673 3249
rect 2617 3203 2673 3215
rect 2773 4133 2826 4203
rect 2773 4099 2784 4133
rect 2818 4099 2826 4133
rect 2773 4065 2826 4099
rect 2773 4031 2784 4065
rect 2818 4031 2826 4065
rect 2773 3997 2826 4031
rect 2773 3963 2784 3997
rect 2818 3963 2826 3997
rect 2773 3929 2826 3963
rect 2773 3895 2784 3929
rect 2818 3895 2826 3929
rect 2773 3861 2826 3895
rect 2773 3827 2784 3861
rect 2818 3827 2826 3861
rect 2773 3793 2826 3827
rect 2773 3759 2784 3793
rect 2818 3759 2826 3793
rect 2773 3725 2826 3759
rect 2773 3691 2784 3725
rect 2818 3691 2826 3725
rect 2773 3657 2826 3691
rect 2773 3623 2784 3657
rect 2818 3623 2826 3657
rect 2773 3589 2826 3623
rect 2773 3555 2784 3589
rect 2818 3555 2826 3589
rect 2773 3521 2826 3555
rect 2773 3487 2784 3521
rect 2818 3487 2826 3521
rect 2773 3453 2826 3487
rect 2773 3419 2784 3453
rect 2818 3419 2826 3453
rect 2773 3385 2826 3419
rect 2773 3351 2784 3385
rect 2818 3351 2826 3385
rect 2773 3317 2826 3351
rect 2773 3283 2784 3317
rect 2818 3283 2826 3317
rect 2773 3249 2826 3283
rect 2773 3215 2784 3249
rect 2818 3215 2826 3249
rect 2773 3203 2826 3215
rect 2972 4133 3025 4203
rect 2972 4099 2980 4133
rect 3014 4099 3025 4133
rect 2972 4065 3025 4099
rect 2972 4031 2980 4065
rect 3014 4031 3025 4065
rect 2972 3997 3025 4031
rect 2972 3963 2980 3997
rect 3014 3963 3025 3997
rect 2972 3929 3025 3963
rect 2972 3895 2980 3929
rect 3014 3895 3025 3929
rect 2972 3861 3025 3895
rect 2972 3827 2980 3861
rect 3014 3827 3025 3861
rect 2972 3793 3025 3827
rect 2972 3759 2980 3793
rect 3014 3759 3025 3793
rect 2972 3725 3025 3759
rect 2972 3691 2980 3725
rect 3014 3691 3025 3725
rect 2972 3657 3025 3691
rect 2972 3623 2980 3657
rect 3014 3623 3025 3657
rect 2972 3589 3025 3623
rect 2972 3555 2980 3589
rect 3014 3555 3025 3589
rect 2972 3521 3025 3555
rect 2972 3487 2980 3521
rect 3014 3487 3025 3521
rect 2972 3453 3025 3487
rect 2972 3419 2980 3453
rect 3014 3419 3025 3453
rect 2972 3385 3025 3419
rect 2972 3351 2980 3385
rect 3014 3351 3025 3385
rect 2972 3317 3025 3351
rect 2972 3283 2980 3317
rect 3014 3283 3025 3317
rect 2972 3249 3025 3283
rect 2972 3215 2980 3249
rect 3014 3215 3025 3249
rect 2972 3203 3025 3215
rect 3125 4133 3181 4203
rect 3125 4099 3136 4133
rect 3170 4099 3181 4133
rect 3125 4065 3181 4099
rect 3125 4031 3136 4065
rect 3170 4031 3181 4065
rect 3125 3997 3181 4031
rect 3125 3963 3136 3997
rect 3170 3963 3181 3997
rect 3125 3929 3181 3963
rect 3125 3895 3136 3929
rect 3170 3895 3181 3929
rect 3125 3861 3181 3895
rect 3125 3827 3136 3861
rect 3170 3827 3181 3861
rect 3125 3793 3181 3827
rect 3125 3759 3136 3793
rect 3170 3759 3181 3793
rect 3125 3725 3181 3759
rect 3125 3691 3136 3725
rect 3170 3691 3181 3725
rect 3125 3657 3181 3691
rect 3125 3623 3136 3657
rect 3170 3623 3181 3657
rect 3125 3589 3181 3623
rect 3125 3555 3136 3589
rect 3170 3555 3181 3589
rect 3125 3521 3181 3555
rect 3125 3487 3136 3521
rect 3170 3487 3181 3521
rect 3125 3453 3181 3487
rect 3125 3419 3136 3453
rect 3170 3419 3181 3453
rect 3125 3385 3181 3419
rect 3125 3351 3136 3385
rect 3170 3351 3181 3385
rect 3125 3317 3181 3351
rect 3125 3283 3136 3317
rect 3170 3283 3181 3317
rect 3125 3249 3181 3283
rect 3125 3215 3136 3249
rect 3170 3215 3181 3249
rect 3125 3203 3181 3215
rect 3281 4133 3337 4203
rect 3281 4099 3292 4133
rect 3326 4099 3337 4133
rect 3281 4065 3337 4099
rect 3281 4031 3292 4065
rect 3326 4031 3337 4065
rect 3281 3997 3337 4031
rect 3281 3963 3292 3997
rect 3326 3963 3337 3997
rect 3281 3929 3337 3963
rect 3281 3895 3292 3929
rect 3326 3895 3337 3929
rect 3281 3861 3337 3895
rect 3281 3827 3292 3861
rect 3326 3827 3337 3861
rect 3281 3793 3337 3827
rect 3281 3759 3292 3793
rect 3326 3759 3337 3793
rect 3281 3725 3337 3759
rect 3281 3691 3292 3725
rect 3326 3691 3337 3725
rect 3281 3657 3337 3691
rect 3281 3623 3292 3657
rect 3326 3623 3337 3657
rect 3281 3589 3337 3623
rect 3281 3555 3292 3589
rect 3326 3555 3337 3589
rect 3281 3521 3337 3555
rect 3281 3487 3292 3521
rect 3326 3487 3337 3521
rect 3281 3453 3337 3487
rect 3281 3419 3292 3453
rect 3326 3419 3337 3453
rect 3281 3385 3337 3419
rect 3281 3351 3292 3385
rect 3326 3351 3337 3385
rect 3281 3317 3337 3351
rect 3281 3283 3292 3317
rect 3326 3283 3337 3317
rect 3281 3249 3337 3283
rect 3281 3215 3292 3249
rect 3326 3215 3337 3249
rect 3281 3203 3337 3215
rect 3437 4133 3493 4203
rect 3437 4099 3448 4133
rect 3482 4099 3493 4133
rect 3437 4065 3493 4099
rect 3437 4031 3448 4065
rect 3482 4031 3493 4065
rect 3437 3997 3493 4031
rect 3437 3963 3448 3997
rect 3482 3963 3493 3997
rect 3437 3929 3493 3963
rect 3437 3895 3448 3929
rect 3482 3895 3493 3929
rect 3437 3861 3493 3895
rect 3437 3827 3448 3861
rect 3482 3827 3493 3861
rect 3437 3793 3493 3827
rect 3437 3759 3448 3793
rect 3482 3759 3493 3793
rect 3437 3725 3493 3759
rect 3437 3691 3448 3725
rect 3482 3691 3493 3725
rect 3437 3657 3493 3691
rect 3437 3623 3448 3657
rect 3482 3623 3493 3657
rect 3437 3589 3493 3623
rect 3437 3555 3448 3589
rect 3482 3555 3493 3589
rect 3437 3521 3493 3555
rect 3437 3487 3448 3521
rect 3482 3487 3493 3521
rect 3437 3453 3493 3487
rect 3437 3419 3448 3453
rect 3482 3419 3493 3453
rect 3437 3385 3493 3419
rect 3437 3351 3448 3385
rect 3482 3351 3493 3385
rect 3437 3317 3493 3351
rect 3437 3283 3448 3317
rect 3482 3283 3493 3317
rect 3437 3249 3493 3283
rect 3437 3215 3448 3249
rect 3482 3215 3493 3249
rect 3437 3203 3493 3215
rect 3593 4133 3649 4203
rect 3593 4099 3604 4133
rect 3638 4099 3649 4133
rect 3593 4065 3649 4099
rect 3593 4031 3604 4065
rect 3638 4031 3649 4065
rect 3593 3997 3649 4031
rect 3593 3963 3604 3997
rect 3638 3963 3649 3997
rect 3593 3929 3649 3963
rect 3593 3895 3604 3929
rect 3638 3895 3649 3929
rect 3593 3861 3649 3895
rect 3593 3827 3604 3861
rect 3638 3827 3649 3861
rect 3593 3793 3649 3827
rect 3593 3759 3604 3793
rect 3638 3759 3649 3793
rect 3593 3725 3649 3759
rect 3593 3691 3604 3725
rect 3638 3691 3649 3725
rect 3593 3657 3649 3691
rect 3593 3623 3604 3657
rect 3638 3623 3649 3657
rect 3593 3589 3649 3623
rect 3593 3555 3604 3589
rect 3638 3555 3649 3589
rect 3593 3521 3649 3555
rect 3593 3487 3604 3521
rect 3638 3487 3649 3521
rect 3593 3453 3649 3487
rect 3593 3419 3604 3453
rect 3638 3419 3649 3453
rect 3593 3385 3649 3419
rect 3593 3351 3604 3385
rect 3638 3351 3649 3385
rect 3593 3317 3649 3351
rect 3593 3283 3604 3317
rect 3638 3283 3649 3317
rect 3593 3249 3649 3283
rect 3593 3215 3604 3249
rect 3638 3215 3649 3249
rect 3593 3203 3649 3215
rect 3749 4133 3805 4203
rect 3749 4099 3760 4133
rect 3794 4099 3805 4133
rect 3749 4065 3805 4099
rect 3749 4031 3760 4065
rect 3794 4031 3805 4065
rect 3749 3997 3805 4031
rect 3749 3963 3760 3997
rect 3794 3963 3805 3997
rect 3749 3929 3805 3963
rect 3749 3895 3760 3929
rect 3794 3895 3805 3929
rect 3749 3861 3805 3895
rect 3749 3827 3760 3861
rect 3794 3827 3805 3861
rect 3749 3793 3805 3827
rect 3749 3759 3760 3793
rect 3794 3759 3805 3793
rect 3749 3725 3805 3759
rect 3749 3691 3760 3725
rect 3794 3691 3805 3725
rect 3749 3657 3805 3691
rect 3749 3623 3760 3657
rect 3794 3623 3805 3657
rect 3749 3589 3805 3623
rect 3749 3555 3760 3589
rect 3794 3555 3805 3589
rect 3749 3521 3805 3555
rect 3749 3487 3760 3521
rect 3794 3487 3805 3521
rect 3749 3453 3805 3487
rect 3749 3419 3760 3453
rect 3794 3419 3805 3453
rect 3749 3385 3805 3419
rect 3749 3351 3760 3385
rect 3794 3351 3805 3385
rect 3749 3317 3805 3351
rect 3749 3283 3760 3317
rect 3794 3283 3805 3317
rect 3749 3249 3805 3283
rect 3749 3215 3760 3249
rect 3794 3215 3805 3249
rect 3749 3203 3805 3215
rect 3905 4133 3961 4203
rect 3905 4099 3916 4133
rect 3950 4099 3961 4133
rect 3905 4065 3961 4099
rect 3905 4031 3916 4065
rect 3950 4031 3961 4065
rect 3905 3997 3961 4031
rect 3905 3963 3916 3997
rect 3950 3963 3961 3997
rect 3905 3929 3961 3963
rect 3905 3895 3916 3929
rect 3950 3895 3961 3929
rect 3905 3861 3961 3895
rect 3905 3827 3916 3861
rect 3950 3827 3961 3861
rect 3905 3793 3961 3827
rect 3905 3759 3916 3793
rect 3950 3759 3961 3793
rect 3905 3725 3961 3759
rect 3905 3691 3916 3725
rect 3950 3691 3961 3725
rect 3905 3657 3961 3691
rect 3905 3623 3916 3657
rect 3950 3623 3961 3657
rect 3905 3589 3961 3623
rect 3905 3555 3916 3589
rect 3950 3555 3961 3589
rect 3905 3521 3961 3555
rect 3905 3487 3916 3521
rect 3950 3487 3961 3521
rect 3905 3453 3961 3487
rect 3905 3419 3916 3453
rect 3950 3419 3961 3453
rect 3905 3385 3961 3419
rect 3905 3351 3916 3385
rect 3950 3351 3961 3385
rect 3905 3317 3961 3351
rect 3905 3283 3916 3317
rect 3950 3283 3961 3317
rect 3905 3249 3961 3283
rect 3905 3215 3916 3249
rect 3950 3215 3961 3249
rect 3905 3203 3961 3215
rect 4061 4133 4117 4203
rect 4061 4099 4072 4133
rect 4106 4099 4117 4133
rect 4061 4065 4117 4099
rect 4061 4031 4072 4065
rect 4106 4031 4117 4065
rect 4061 3997 4117 4031
rect 4061 3963 4072 3997
rect 4106 3963 4117 3997
rect 4061 3929 4117 3963
rect 4061 3895 4072 3929
rect 4106 3895 4117 3929
rect 4061 3861 4117 3895
rect 4061 3827 4072 3861
rect 4106 3827 4117 3861
rect 4061 3793 4117 3827
rect 4061 3759 4072 3793
rect 4106 3759 4117 3793
rect 4061 3725 4117 3759
rect 4061 3691 4072 3725
rect 4106 3691 4117 3725
rect 4061 3657 4117 3691
rect 4061 3623 4072 3657
rect 4106 3623 4117 3657
rect 4061 3589 4117 3623
rect 4061 3555 4072 3589
rect 4106 3555 4117 3589
rect 4061 3521 4117 3555
rect 4061 3487 4072 3521
rect 4106 3487 4117 3521
rect 4061 3453 4117 3487
rect 4061 3419 4072 3453
rect 4106 3419 4117 3453
rect 4061 3385 4117 3419
rect 4061 3351 4072 3385
rect 4106 3351 4117 3385
rect 4061 3317 4117 3351
rect 4061 3283 4072 3317
rect 4106 3283 4117 3317
rect 4061 3249 4117 3283
rect 4061 3215 4072 3249
rect 4106 3215 4117 3249
rect 4061 3203 4117 3215
rect 4217 4133 4270 4203
rect 4217 4099 4228 4133
rect 4262 4099 4270 4133
rect 4217 4065 4270 4099
rect 4217 4031 4228 4065
rect 4262 4031 4270 4065
rect 4217 3997 4270 4031
rect 4217 3963 4228 3997
rect 4262 3963 4270 3997
rect 4217 3929 4270 3963
rect 4217 3895 4228 3929
rect 4262 3895 4270 3929
rect 4217 3861 4270 3895
rect 4217 3827 4228 3861
rect 4262 3827 4270 3861
rect 4217 3793 4270 3827
rect 4217 3759 4228 3793
rect 4262 3759 4270 3793
rect 4217 3725 4270 3759
rect 4217 3691 4228 3725
rect 4262 3691 4270 3725
rect 4217 3657 4270 3691
rect 4217 3623 4228 3657
rect 4262 3623 4270 3657
rect 4217 3589 4270 3623
rect 4217 3555 4228 3589
rect 4262 3555 4270 3589
rect 4217 3521 4270 3555
rect 4217 3487 4228 3521
rect 4262 3487 4270 3521
rect 4217 3453 4270 3487
rect 4217 3419 4228 3453
rect 4262 3419 4270 3453
rect 4217 3385 4270 3419
rect 4217 3351 4228 3385
rect 4262 3351 4270 3385
rect 4217 3317 4270 3351
rect 4217 3283 4228 3317
rect 4262 3283 4270 3317
rect 4217 3249 4270 3283
rect 4217 3215 4228 3249
rect 4262 3215 4270 3249
rect 4217 3203 4270 3215
rect 4416 4183 4469 4253
rect 4416 4149 4424 4183
rect 4458 4149 4469 4183
rect 4416 4115 4469 4149
rect 4416 4081 4424 4115
rect 4458 4081 4469 4115
rect 4416 4047 4469 4081
rect 4416 4013 4424 4047
rect 4458 4013 4469 4047
rect 4416 3979 4469 4013
rect 4416 3945 4424 3979
rect 4458 3945 4469 3979
rect 4416 3911 4469 3945
rect 4416 3877 4424 3911
rect 4458 3877 4469 3911
rect 4416 3843 4469 3877
rect 4416 3809 4424 3843
rect 4458 3809 4469 3843
rect 4416 3775 4469 3809
rect 4416 3741 4424 3775
rect 4458 3741 4469 3775
rect 4416 3707 4469 3741
rect 4416 3673 4424 3707
rect 4458 3673 4469 3707
rect 4416 3639 4469 3673
rect 4416 3605 4424 3639
rect 4458 3605 4469 3639
rect 4416 3571 4469 3605
rect 4416 3537 4424 3571
rect 4458 3537 4469 3571
rect 4416 3503 4469 3537
rect 4416 3469 4424 3503
rect 4458 3469 4469 3503
rect 4416 3435 4469 3469
rect 4416 3401 4424 3435
rect 4458 3401 4469 3435
rect 4416 3367 4469 3401
rect 4416 3333 4424 3367
rect 4458 3333 4469 3367
rect 4416 3299 4469 3333
rect 4416 3265 4424 3299
rect 4458 3265 4469 3299
rect 4416 3253 4469 3265
rect 4569 4183 4625 4253
rect 4569 4149 4580 4183
rect 4614 4149 4625 4183
rect 4569 4115 4625 4149
rect 4569 4081 4580 4115
rect 4614 4081 4625 4115
rect 4569 4047 4625 4081
rect 4569 4013 4580 4047
rect 4614 4013 4625 4047
rect 4569 3979 4625 4013
rect 4569 3945 4580 3979
rect 4614 3945 4625 3979
rect 4569 3911 4625 3945
rect 4569 3877 4580 3911
rect 4614 3877 4625 3911
rect 4569 3843 4625 3877
rect 4569 3809 4580 3843
rect 4614 3809 4625 3843
rect 4569 3775 4625 3809
rect 4569 3741 4580 3775
rect 4614 3741 4625 3775
rect 4569 3707 4625 3741
rect 4569 3673 4580 3707
rect 4614 3673 4625 3707
rect 4569 3639 4625 3673
rect 4569 3605 4580 3639
rect 4614 3605 4625 3639
rect 4569 3571 4625 3605
rect 4569 3537 4580 3571
rect 4614 3537 4625 3571
rect 4569 3503 4625 3537
rect 4569 3469 4580 3503
rect 4614 3469 4625 3503
rect 4569 3435 4625 3469
rect 4569 3401 4580 3435
rect 4614 3401 4625 3435
rect 4569 3367 4625 3401
rect 4569 3333 4580 3367
rect 4614 3333 4625 3367
rect 4569 3299 4625 3333
rect 4569 3265 4580 3299
rect 4614 3265 4625 3299
rect 4569 3253 4625 3265
rect 4725 4183 4781 4253
rect 4725 4149 4736 4183
rect 4770 4149 4781 4183
rect 4725 4115 4781 4149
rect 4725 4081 4736 4115
rect 4770 4081 4781 4115
rect 4725 4047 4781 4081
rect 4725 4013 4736 4047
rect 4770 4013 4781 4047
rect 4725 3979 4781 4013
rect 4725 3945 4736 3979
rect 4770 3945 4781 3979
rect 4725 3911 4781 3945
rect 4725 3877 4736 3911
rect 4770 3877 4781 3911
rect 4725 3843 4781 3877
rect 4725 3809 4736 3843
rect 4770 3809 4781 3843
rect 4725 3775 4781 3809
rect 4725 3741 4736 3775
rect 4770 3741 4781 3775
rect 4725 3707 4781 3741
rect 4725 3673 4736 3707
rect 4770 3673 4781 3707
rect 4725 3639 4781 3673
rect 4725 3605 4736 3639
rect 4770 3605 4781 3639
rect 4725 3571 4781 3605
rect 4725 3537 4736 3571
rect 4770 3537 4781 3571
rect 4725 3503 4781 3537
rect 4725 3469 4736 3503
rect 4770 3469 4781 3503
rect 4725 3435 4781 3469
rect 4725 3401 4736 3435
rect 4770 3401 4781 3435
rect 4725 3367 4781 3401
rect 4725 3333 4736 3367
rect 4770 3333 4781 3367
rect 4725 3299 4781 3333
rect 4725 3265 4736 3299
rect 4770 3265 4781 3299
rect 4725 3253 4781 3265
rect 4881 4183 4937 4253
rect 4881 4149 4892 4183
rect 4926 4149 4937 4183
rect 4881 4115 4937 4149
rect 4881 4081 4892 4115
rect 4926 4081 4937 4115
rect 4881 4047 4937 4081
rect 4881 4013 4892 4047
rect 4926 4013 4937 4047
rect 4881 3979 4937 4013
rect 4881 3945 4892 3979
rect 4926 3945 4937 3979
rect 4881 3911 4937 3945
rect 4881 3877 4892 3911
rect 4926 3877 4937 3911
rect 4881 3843 4937 3877
rect 4881 3809 4892 3843
rect 4926 3809 4937 3843
rect 4881 3775 4937 3809
rect 4881 3741 4892 3775
rect 4926 3741 4937 3775
rect 4881 3707 4937 3741
rect 4881 3673 4892 3707
rect 4926 3673 4937 3707
rect 4881 3639 4937 3673
rect 4881 3605 4892 3639
rect 4926 3605 4937 3639
rect 4881 3571 4937 3605
rect 4881 3537 4892 3571
rect 4926 3537 4937 3571
rect 4881 3503 4937 3537
rect 4881 3469 4892 3503
rect 4926 3469 4937 3503
rect 4881 3435 4937 3469
rect 4881 3401 4892 3435
rect 4926 3401 4937 3435
rect 4881 3367 4937 3401
rect 4881 3333 4892 3367
rect 4926 3333 4937 3367
rect 4881 3299 4937 3333
rect 4881 3265 4892 3299
rect 4926 3265 4937 3299
rect 4881 3253 4937 3265
rect 5037 4183 5093 4253
rect 5037 4149 5048 4183
rect 5082 4149 5093 4183
rect 5037 4115 5093 4149
rect 5037 4081 5048 4115
rect 5082 4081 5093 4115
rect 5037 4047 5093 4081
rect 5037 4013 5048 4047
rect 5082 4013 5093 4047
rect 5037 3979 5093 4013
rect 5037 3945 5048 3979
rect 5082 3945 5093 3979
rect 5037 3911 5093 3945
rect 5037 3877 5048 3911
rect 5082 3877 5093 3911
rect 5037 3843 5093 3877
rect 5037 3809 5048 3843
rect 5082 3809 5093 3843
rect 5037 3775 5093 3809
rect 5037 3741 5048 3775
rect 5082 3741 5093 3775
rect 5037 3707 5093 3741
rect 5037 3673 5048 3707
rect 5082 3673 5093 3707
rect 5037 3639 5093 3673
rect 5037 3605 5048 3639
rect 5082 3605 5093 3639
rect 5037 3571 5093 3605
rect 5037 3537 5048 3571
rect 5082 3537 5093 3571
rect 5037 3503 5093 3537
rect 5037 3469 5048 3503
rect 5082 3469 5093 3503
rect 5037 3435 5093 3469
rect 5037 3401 5048 3435
rect 5082 3401 5093 3435
rect 5037 3367 5093 3401
rect 5037 3333 5048 3367
rect 5082 3333 5093 3367
rect 5037 3299 5093 3333
rect 5037 3265 5048 3299
rect 5082 3265 5093 3299
rect 5037 3253 5093 3265
rect 5193 4183 5249 4253
rect 5193 4149 5204 4183
rect 5238 4149 5249 4183
rect 5193 4115 5249 4149
rect 5193 4081 5204 4115
rect 5238 4081 5249 4115
rect 5193 4047 5249 4081
rect 5193 4013 5204 4047
rect 5238 4013 5249 4047
rect 5193 3979 5249 4013
rect 5193 3945 5204 3979
rect 5238 3945 5249 3979
rect 5193 3911 5249 3945
rect 5193 3877 5204 3911
rect 5238 3877 5249 3911
rect 5193 3843 5249 3877
rect 5193 3809 5204 3843
rect 5238 3809 5249 3843
rect 5193 3775 5249 3809
rect 5193 3741 5204 3775
rect 5238 3741 5249 3775
rect 5193 3707 5249 3741
rect 5193 3673 5204 3707
rect 5238 3673 5249 3707
rect 5193 3639 5249 3673
rect 5193 3605 5204 3639
rect 5238 3605 5249 3639
rect 5193 3571 5249 3605
rect 5193 3537 5204 3571
rect 5238 3537 5249 3571
rect 5193 3503 5249 3537
rect 5193 3469 5204 3503
rect 5238 3469 5249 3503
rect 5193 3435 5249 3469
rect 5193 3401 5204 3435
rect 5238 3401 5249 3435
rect 5193 3367 5249 3401
rect 5193 3333 5204 3367
rect 5238 3333 5249 3367
rect 5193 3299 5249 3333
rect 5193 3265 5204 3299
rect 5238 3265 5249 3299
rect 5193 3253 5249 3265
rect 5349 4183 5405 4253
rect 5349 4149 5360 4183
rect 5394 4149 5405 4183
rect 5349 4115 5405 4149
rect 5349 4081 5360 4115
rect 5394 4081 5405 4115
rect 5349 4047 5405 4081
rect 5349 4013 5360 4047
rect 5394 4013 5405 4047
rect 5349 3979 5405 4013
rect 5349 3945 5360 3979
rect 5394 3945 5405 3979
rect 5349 3911 5405 3945
rect 5349 3877 5360 3911
rect 5394 3877 5405 3911
rect 5349 3843 5405 3877
rect 5349 3809 5360 3843
rect 5394 3809 5405 3843
rect 5349 3775 5405 3809
rect 5349 3741 5360 3775
rect 5394 3741 5405 3775
rect 5349 3707 5405 3741
rect 5349 3673 5360 3707
rect 5394 3673 5405 3707
rect 5349 3639 5405 3673
rect 5349 3605 5360 3639
rect 5394 3605 5405 3639
rect 5349 3571 5405 3605
rect 5349 3537 5360 3571
rect 5394 3537 5405 3571
rect 5349 3503 5405 3537
rect 5349 3469 5360 3503
rect 5394 3469 5405 3503
rect 5349 3435 5405 3469
rect 5349 3401 5360 3435
rect 5394 3401 5405 3435
rect 5349 3367 5405 3401
rect 5349 3333 5360 3367
rect 5394 3333 5405 3367
rect 5349 3299 5405 3333
rect 5349 3265 5360 3299
rect 5394 3265 5405 3299
rect 5349 3253 5405 3265
rect 5505 4183 5561 4253
rect 5505 4149 5516 4183
rect 5550 4149 5561 4183
rect 5505 4115 5561 4149
rect 5505 4081 5516 4115
rect 5550 4081 5561 4115
rect 5505 4047 5561 4081
rect 5505 4013 5516 4047
rect 5550 4013 5561 4047
rect 5505 3979 5561 4013
rect 5505 3945 5516 3979
rect 5550 3945 5561 3979
rect 5505 3911 5561 3945
rect 5505 3877 5516 3911
rect 5550 3877 5561 3911
rect 5505 3843 5561 3877
rect 5505 3809 5516 3843
rect 5550 3809 5561 3843
rect 5505 3775 5561 3809
rect 5505 3741 5516 3775
rect 5550 3741 5561 3775
rect 5505 3707 5561 3741
rect 5505 3673 5516 3707
rect 5550 3673 5561 3707
rect 5505 3639 5561 3673
rect 5505 3605 5516 3639
rect 5550 3605 5561 3639
rect 5505 3571 5561 3605
rect 5505 3537 5516 3571
rect 5550 3537 5561 3571
rect 5505 3503 5561 3537
rect 5505 3469 5516 3503
rect 5550 3469 5561 3503
rect 5505 3435 5561 3469
rect 5505 3401 5516 3435
rect 5550 3401 5561 3435
rect 5505 3367 5561 3401
rect 5505 3333 5516 3367
rect 5550 3333 5561 3367
rect 5505 3299 5561 3333
rect 5505 3265 5516 3299
rect 5550 3265 5561 3299
rect 5505 3253 5561 3265
rect 5661 4183 5714 4253
rect 9137 4272 9145 4306
rect 9179 4272 9190 4306
rect 9137 4238 9190 4272
rect 9137 4204 9145 4238
rect 9179 4204 9190 4238
rect 5661 4149 5672 4183
rect 5706 4149 5714 4183
rect 5661 4115 5714 4149
rect 5661 4081 5672 4115
rect 5706 4081 5714 4115
rect 5661 4047 5714 4081
rect 5661 4013 5672 4047
rect 5706 4013 5714 4047
rect 5661 3979 5714 4013
rect 5661 3945 5672 3979
rect 5706 3945 5714 3979
rect 5661 3911 5714 3945
rect 5661 3877 5672 3911
rect 5706 3877 5714 3911
rect 5661 3843 5714 3877
rect 5661 3809 5672 3843
rect 5706 3809 5714 3843
rect 5661 3775 5714 3809
rect 5661 3741 5672 3775
rect 5706 3741 5714 3775
rect 5661 3707 5714 3741
rect 5661 3673 5672 3707
rect 5706 3673 5714 3707
rect 5661 3639 5714 3673
rect 5661 3605 5672 3639
rect 5706 3605 5714 3639
rect 5661 3571 5714 3605
rect 5661 3537 5672 3571
rect 5706 3537 5714 3571
rect 5661 3503 5714 3537
rect 5661 3469 5672 3503
rect 5706 3469 5714 3503
rect 5661 3435 5714 3469
rect 5661 3401 5672 3435
rect 5706 3401 5714 3435
rect 5661 3367 5714 3401
rect 5661 3333 5672 3367
rect 5706 3333 5714 3367
rect 5661 3299 5714 3333
rect 5661 3265 5672 3299
rect 5706 3265 5714 3299
rect 5661 3253 5714 3265
rect 5860 4133 5913 4203
rect 5860 4099 5868 4133
rect 5902 4099 5913 4133
rect 5860 4065 5913 4099
rect 5860 4031 5868 4065
rect 5902 4031 5913 4065
rect 5860 3997 5913 4031
rect 5860 3963 5868 3997
rect 5902 3963 5913 3997
rect 5860 3929 5913 3963
rect 5860 3895 5868 3929
rect 5902 3895 5913 3929
rect 5860 3861 5913 3895
rect 5860 3827 5868 3861
rect 5902 3827 5913 3861
rect 5860 3793 5913 3827
rect 5860 3759 5868 3793
rect 5902 3759 5913 3793
rect 5860 3725 5913 3759
rect 5860 3691 5868 3725
rect 5902 3691 5913 3725
rect 5860 3657 5913 3691
rect 5860 3623 5868 3657
rect 5902 3623 5913 3657
rect 5860 3589 5913 3623
rect 5860 3555 5868 3589
rect 5902 3555 5913 3589
rect 5860 3521 5913 3555
rect 5860 3487 5868 3521
rect 5902 3487 5913 3521
rect 5860 3453 5913 3487
rect 5860 3419 5868 3453
rect 5902 3419 5913 3453
rect 5860 3385 5913 3419
rect 5860 3351 5868 3385
rect 5902 3351 5913 3385
rect 5860 3317 5913 3351
rect 5860 3283 5868 3317
rect 5902 3283 5913 3317
rect 5860 3249 5913 3283
rect 5860 3215 5868 3249
rect 5902 3215 5913 3249
rect 5860 3203 5913 3215
rect 6013 4133 6069 4203
rect 6013 4099 6024 4133
rect 6058 4099 6069 4133
rect 6013 4065 6069 4099
rect 6013 4031 6024 4065
rect 6058 4031 6069 4065
rect 6013 3997 6069 4031
rect 6013 3963 6024 3997
rect 6058 3963 6069 3997
rect 6013 3929 6069 3963
rect 6013 3895 6024 3929
rect 6058 3895 6069 3929
rect 6013 3861 6069 3895
rect 6013 3827 6024 3861
rect 6058 3827 6069 3861
rect 6013 3793 6069 3827
rect 6013 3759 6024 3793
rect 6058 3759 6069 3793
rect 6013 3725 6069 3759
rect 6013 3691 6024 3725
rect 6058 3691 6069 3725
rect 6013 3657 6069 3691
rect 6013 3623 6024 3657
rect 6058 3623 6069 3657
rect 6013 3589 6069 3623
rect 6013 3555 6024 3589
rect 6058 3555 6069 3589
rect 6013 3521 6069 3555
rect 6013 3487 6024 3521
rect 6058 3487 6069 3521
rect 6013 3453 6069 3487
rect 6013 3419 6024 3453
rect 6058 3419 6069 3453
rect 6013 3385 6069 3419
rect 6013 3351 6024 3385
rect 6058 3351 6069 3385
rect 6013 3317 6069 3351
rect 6013 3283 6024 3317
rect 6058 3283 6069 3317
rect 6013 3249 6069 3283
rect 6013 3215 6024 3249
rect 6058 3215 6069 3249
rect 6013 3203 6069 3215
rect 6169 4133 6225 4203
rect 6169 4099 6180 4133
rect 6214 4099 6225 4133
rect 6169 4065 6225 4099
rect 6169 4031 6180 4065
rect 6214 4031 6225 4065
rect 6169 3997 6225 4031
rect 6169 3963 6180 3997
rect 6214 3963 6225 3997
rect 6169 3929 6225 3963
rect 6169 3895 6180 3929
rect 6214 3895 6225 3929
rect 6169 3861 6225 3895
rect 6169 3827 6180 3861
rect 6214 3827 6225 3861
rect 6169 3793 6225 3827
rect 6169 3759 6180 3793
rect 6214 3759 6225 3793
rect 6169 3725 6225 3759
rect 6169 3691 6180 3725
rect 6214 3691 6225 3725
rect 6169 3657 6225 3691
rect 6169 3623 6180 3657
rect 6214 3623 6225 3657
rect 6169 3589 6225 3623
rect 6169 3555 6180 3589
rect 6214 3555 6225 3589
rect 6169 3521 6225 3555
rect 6169 3487 6180 3521
rect 6214 3487 6225 3521
rect 6169 3453 6225 3487
rect 6169 3419 6180 3453
rect 6214 3419 6225 3453
rect 6169 3385 6225 3419
rect 6169 3351 6180 3385
rect 6214 3351 6225 3385
rect 6169 3317 6225 3351
rect 6169 3283 6180 3317
rect 6214 3283 6225 3317
rect 6169 3249 6225 3283
rect 6169 3215 6180 3249
rect 6214 3215 6225 3249
rect 6169 3203 6225 3215
rect 6325 4133 6381 4203
rect 6325 4099 6336 4133
rect 6370 4099 6381 4133
rect 6325 4065 6381 4099
rect 6325 4031 6336 4065
rect 6370 4031 6381 4065
rect 6325 3997 6381 4031
rect 6325 3963 6336 3997
rect 6370 3963 6381 3997
rect 6325 3929 6381 3963
rect 6325 3895 6336 3929
rect 6370 3895 6381 3929
rect 6325 3861 6381 3895
rect 6325 3827 6336 3861
rect 6370 3827 6381 3861
rect 6325 3793 6381 3827
rect 6325 3759 6336 3793
rect 6370 3759 6381 3793
rect 6325 3725 6381 3759
rect 6325 3691 6336 3725
rect 6370 3691 6381 3725
rect 6325 3657 6381 3691
rect 6325 3623 6336 3657
rect 6370 3623 6381 3657
rect 6325 3589 6381 3623
rect 6325 3555 6336 3589
rect 6370 3555 6381 3589
rect 6325 3521 6381 3555
rect 6325 3487 6336 3521
rect 6370 3487 6381 3521
rect 6325 3453 6381 3487
rect 6325 3419 6336 3453
rect 6370 3419 6381 3453
rect 6325 3385 6381 3419
rect 6325 3351 6336 3385
rect 6370 3351 6381 3385
rect 6325 3317 6381 3351
rect 6325 3283 6336 3317
rect 6370 3283 6381 3317
rect 6325 3249 6381 3283
rect 6325 3215 6336 3249
rect 6370 3215 6381 3249
rect 6325 3203 6381 3215
rect 6481 4133 6537 4203
rect 6481 4099 6492 4133
rect 6526 4099 6537 4133
rect 6481 4065 6537 4099
rect 6481 4031 6492 4065
rect 6526 4031 6537 4065
rect 6481 3997 6537 4031
rect 6481 3963 6492 3997
rect 6526 3963 6537 3997
rect 6481 3929 6537 3963
rect 6481 3895 6492 3929
rect 6526 3895 6537 3929
rect 6481 3861 6537 3895
rect 6481 3827 6492 3861
rect 6526 3827 6537 3861
rect 6481 3793 6537 3827
rect 6481 3759 6492 3793
rect 6526 3759 6537 3793
rect 6481 3725 6537 3759
rect 6481 3691 6492 3725
rect 6526 3691 6537 3725
rect 6481 3657 6537 3691
rect 6481 3623 6492 3657
rect 6526 3623 6537 3657
rect 6481 3589 6537 3623
rect 6481 3555 6492 3589
rect 6526 3555 6537 3589
rect 6481 3521 6537 3555
rect 6481 3487 6492 3521
rect 6526 3487 6537 3521
rect 6481 3453 6537 3487
rect 6481 3419 6492 3453
rect 6526 3419 6537 3453
rect 6481 3385 6537 3419
rect 6481 3351 6492 3385
rect 6526 3351 6537 3385
rect 6481 3317 6537 3351
rect 6481 3283 6492 3317
rect 6526 3283 6537 3317
rect 6481 3249 6537 3283
rect 6481 3215 6492 3249
rect 6526 3215 6537 3249
rect 6481 3203 6537 3215
rect 6637 4133 6693 4203
rect 6637 4099 6648 4133
rect 6682 4099 6693 4133
rect 6637 4065 6693 4099
rect 6637 4031 6648 4065
rect 6682 4031 6693 4065
rect 6637 3997 6693 4031
rect 6637 3963 6648 3997
rect 6682 3963 6693 3997
rect 6637 3929 6693 3963
rect 6637 3895 6648 3929
rect 6682 3895 6693 3929
rect 6637 3861 6693 3895
rect 6637 3827 6648 3861
rect 6682 3827 6693 3861
rect 6637 3793 6693 3827
rect 6637 3759 6648 3793
rect 6682 3759 6693 3793
rect 6637 3725 6693 3759
rect 6637 3691 6648 3725
rect 6682 3691 6693 3725
rect 6637 3657 6693 3691
rect 6637 3623 6648 3657
rect 6682 3623 6693 3657
rect 6637 3589 6693 3623
rect 6637 3555 6648 3589
rect 6682 3555 6693 3589
rect 6637 3521 6693 3555
rect 6637 3487 6648 3521
rect 6682 3487 6693 3521
rect 6637 3453 6693 3487
rect 6637 3419 6648 3453
rect 6682 3419 6693 3453
rect 6637 3385 6693 3419
rect 6637 3351 6648 3385
rect 6682 3351 6693 3385
rect 6637 3317 6693 3351
rect 6637 3283 6648 3317
rect 6682 3283 6693 3317
rect 6637 3249 6693 3283
rect 6637 3215 6648 3249
rect 6682 3215 6693 3249
rect 6637 3203 6693 3215
rect 6793 4133 6849 4203
rect 6793 4099 6804 4133
rect 6838 4099 6849 4133
rect 6793 4065 6849 4099
rect 6793 4031 6804 4065
rect 6838 4031 6849 4065
rect 6793 3997 6849 4031
rect 6793 3963 6804 3997
rect 6838 3963 6849 3997
rect 6793 3929 6849 3963
rect 6793 3895 6804 3929
rect 6838 3895 6849 3929
rect 6793 3861 6849 3895
rect 6793 3827 6804 3861
rect 6838 3827 6849 3861
rect 6793 3793 6849 3827
rect 6793 3759 6804 3793
rect 6838 3759 6849 3793
rect 6793 3725 6849 3759
rect 6793 3691 6804 3725
rect 6838 3691 6849 3725
rect 6793 3657 6849 3691
rect 6793 3623 6804 3657
rect 6838 3623 6849 3657
rect 6793 3589 6849 3623
rect 6793 3555 6804 3589
rect 6838 3555 6849 3589
rect 6793 3521 6849 3555
rect 6793 3487 6804 3521
rect 6838 3487 6849 3521
rect 6793 3453 6849 3487
rect 6793 3419 6804 3453
rect 6838 3419 6849 3453
rect 6793 3385 6849 3419
rect 6793 3351 6804 3385
rect 6838 3351 6849 3385
rect 6793 3317 6849 3351
rect 6793 3283 6804 3317
rect 6838 3283 6849 3317
rect 6793 3249 6849 3283
rect 6793 3215 6804 3249
rect 6838 3215 6849 3249
rect 6793 3203 6849 3215
rect 6949 4133 7005 4203
rect 6949 4099 6960 4133
rect 6994 4099 7005 4133
rect 6949 4065 7005 4099
rect 6949 4031 6960 4065
rect 6994 4031 7005 4065
rect 6949 3997 7005 4031
rect 6949 3963 6960 3997
rect 6994 3963 7005 3997
rect 6949 3929 7005 3963
rect 6949 3895 6960 3929
rect 6994 3895 7005 3929
rect 6949 3861 7005 3895
rect 6949 3827 6960 3861
rect 6994 3827 7005 3861
rect 6949 3793 7005 3827
rect 6949 3759 6960 3793
rect 6994 3759 7005 3793
rect 6949 3725 7005 3759
rect 6949 3691 6960 3725
rect 6994 3691 7005 3725
rect 6949 3657 7005 3691
rect 6949 3623 6960 3657
rect 6994 3623 7005 3657
rect 6949 3589 7005 3623
rect 6949 3555 6960 3589
rect 6994 3555 7005 3589
rect 6949 3521 7005 3555
rect 6949 3487 6960 3521
rect 6994 3487 7005 3521
rect 6949 3453 7005 3487
rect 6949 3419 6960 3453
rect 6994 3419 7005 3453
rect 6949 3385 7005 3419
rect 6949 3351 6960 3385
rect 6994 3351 7005 3385
rect 6949 3317 7005 3351
rect 6949 3283 6960 3317
rect 6994 3283 7005 3317
rect 6949 3249 7005 3283
rect 6949 3215 6960 3249
rect 6994 3215 7005 3249
rect 6949 3203 7005 3215
rect 7105 4133 7161 4203
rect 7105 4099 7116 4133
rect 7150 4099 7161 4133
rect 7105 4065 7161 4099
rect 7105 4031 7116 4065
rect 7150 4031 7161 4065
rect 7105 3997 7161 4031
rect 7105 3963 7116 3997
rect 7150 3963 7161 3997
rect 7105 3929 7161 3963
rect 7105 3895 7116 3929
rect 7150 3895 7161 3929
rect 7105 3861 7161 3895
rect 7105 3827 7116 3861
rect 7150 3827 7161 3861
rect 7105 3793 7161 3827
rect 7105 3759 7116 3793
rect 7150 3759 7161 3793
rect 7105 3725 7161 3759
rect 7105 3691 7116 3725
rect 7150 3691 7161 3725
rect 7105 3657 7161 3691
rect 7105 3623 7116 3657
rect 7150 3623 7161 3657
rect 7105 3589 7161 3623
rect 7105 3555 7116 3589
rect 7150 3555 7161 3589
rect 7105 3521 7161 3555
rect 7105 3487 7116 3521
rect 7150 3487 7161 3521
rect 7105 3453 7161 3487
rect 7105 3419 7116 3453
rect 7150 3419 7161 3453
rect 7105 3385 7161 3419
rect 7105 3351 7116 3385
rect 7150 3351 7161 3385
rect 7105 3317 7161 3351
rect 7105 3283 7116 3317
rect 7150 3283 7161 3317
rect 7105 3249 7161 3283
rect 7105 3215 7116 3249
rect 7150 3215 7161 3249
rect 7105 3203 7161 3215
rect 7261 4133 7314 4203
rect 7261 4099 7272 4133
rect 7306 4099 7314 4133
rect 7261 4065 7314 4099
rect 7261 4031 7272 4065
rect 7306 4031 7314 4065
rect 7261 3997 7314 4031
rect 7261 3963 7272 3997
rect 7306 3963 7314 3997
rect 7261 3929 7314 3963
rect 7261 3895 7272 3929
rect 7306 3895 7314 3929
rect 7261 3861 7314 3895
rect 7261 3827 7272 3861
rect 7306 3827 7314 3861
rect 7261 3793 7314 3827
rect 7261 3759 7272 3793
rect 7306 3759 7314 3793
rect 7261 3725 7314 3759
rect 7261 3691 7272 3725
rect 7306 3691 7314 3725
rect 7261 3657 7314 3691
rect 7261 3623 7272 3657
rect 7306 3623 7314 3657
rect 7261 3589 7314 3623
rect 7261 3555 7272 3589
rect 7306 3555 7314 3589
rect 7261 3521 7314 3555
rect 7261 3487 7272 3521
rect 7306 3487 7314 3521
rect 7261 3453 7314 3487
rect 7261 3419 7272 3453
rect 7306 3419 7314 3453
rect 7261 3385 7314 3419
rect 7261 3351 7272 3385
rect 7306 3351 7314 3385
rect 7261 3317 7314 3351
rect 7261 3283 7272 3317
rect 7306 3283 7314 3317
rect 7261 3249 7314 3283
rect 7261 3215 7272 3249
rect 7306 3215 7314 3249
rect 7261 3203 7314 3215
rect 7460 4125 7513 4203
rect 7460 4091 7468 4125
rect 7502 4091 7513 4125
rect 7460 4057 7513 4091
rect 7460 4023 7468 4057
rect 7502 4023 7513 4057
rect 7460 3989 7513 4023
rect 7460 3955 7468 3989
rect 7502 3955 7513 3989
rect 7460 3921 7513 3955
rect 7460 3887 7468 3921
rect 7502 3887 7513 3921
rect 7460 3853 7513 3887
rect 7460 3819 7468 3853
rect 7502 3819 7513 3853
rect 7460 3785 7513 3819
rect 7460 3751 7468 3785
rect 7502 3751 7513 3785
rect 7460 3717 7513 3751
rect 7460 3683 7468 3717
rect 7502 3683 7513 3717
rect 7460 3649 7513 3683
rect 7460 3615 7468 3649
rect 7502 3615 7513 3649
rect 7460 3603 7513 3615
rect 7613 3603 7655 4203
rect 7755 3603 7797 4203
rect 7897 4125 7950 4203
rect 7897 4091 7908 4125
rect 7942 4091 7950 4125
rect 9137 4170 9190 4204
rect 7897 4057 7950 4091
rect 7897 4023 7908 4057
rect 7942 4023 7950 4057
rect 8026 4101 8110 4109
rect 8026 4067 8038 4101
rect 8072 4067 8110 4101
rect 8026 4056 8110 4067
rect 7897 3989 7950 4023
rect 7897 3955 7908 3989
rect 7942 3955 7950 3989
rect 7897 3921 7950 3955
rect 7897 3887 7908 3921
rect 7942 3887 7950 3921
rect 7897 3853 7950 3887
rect 7897 3819 7908 3853
rect 7942 3819 7950 3853
rect 7897 3785 7950 3819
rect 7897 3751 7908 3785
rect 7942 3751 7950 3785
rect 7897 3717 7950 3751
rect 7897 3683 7908 3717
rect 7942 3683 7950 3717
rect 7897 3649 7950 3683
rect 7897 3615 7908 3649
rect 7942 3615 7950 3649
rect 7897 3603 7950 3615
rect 7460 3390 7513 3408
rect 7460 3356 7468 3390
rect 7502 3356 7513 3390
rect 7460 3322 7513 3356
rect 7460 3288 7468 3322
rect 7502 3288 7513 3322
rect 7460 3254 7513 3288
rect 7460 3220 7468 3254
rect 7502 3220 7513 3254
rect 7460 3208 7513 3220
rect 7613 3390 7669 3408
rect 7613 3356 7624 3390
rect 7658 3356 7669 3390
rect 7613 3322 7669 3356
rect 7613 3288 7624 3322
rect 7658 3288 7669 3322
rect 7613 3254 7669 3288
rect 7613 3220 7624 3254
rect 7658 3220 7669 3254
rect 7613 3208 7669 3220
rect 7769 3390 7822 3408
rect 7769 3356 7780 3390
rect 7814 3356 7822 3390
rect 7769 3322 7822 3356
rect 7769 3288 7780 3322
rect 7814 3288 7822 3322
rect 7769 3254 7822 3288
rect 7769 3220 7780 3254
rect 7814 3220 7822 3254
rect 7769 3208 7822 3220
rect 8026 3245 8110 3256
rect 8026 3211 8038 3245
rect 8072 3211 8110 3245
rect 8026 3203 8110 3211
rect 9137 4136 9145 4170
rect 9179 4136 9190 4170
rect 9137 4102 9190 4136
rect 9137 4068 9145 4102
rect 9179 4068 9190 4102
rect 9137 4034 9190 4068
rect 9137 4000 9145 4034
rect 9179 4000 9190 4034
rect 9137 3966 9190 4000
rect 9137 3932 9145 3966
rect 9179 3932 9190 3966
rect 9137 3898 9190 3932
rect 9137 3864 9145 3898
rect 9179 3864 9190 3898
rect 9137 3830 9190 3864
rect 9137 3796 9145 3830
rect 9179 3796 9190 3830
rect 9137 3718 9190 3796
rect 9290 4306 9346 4318
rect 9290 4272 9301 4306
rect 9335 4272 9346 4306
rect 9290 4238 9346 4272
rect 9290 4204 9301 4238
rect 9335 4204 9346 4238
rect 9290 4170 9346 4204
rect 9290 4136 9301 4170
rect 9335 4136 9346 4170
rect 9290 4102 9346 4136
rect 9290 4068 9301 4102
rect 9335 4068 9346 4102
rect 9290 4034 9346 4068
rect 9290 4000 9301 4034
rect 9335 4000 9346 4034
rect 9290 3966 9346 4000
rect 9290 3932 9301 3966
rect 9335 3932 9346 3966
rect 9290 3898 9346 3932
rect 9290 3864 9301 3898
rect 9335 3864 9346 3898
rect 9290 3830 9346 3864
rect 9290 3796 9301 3830
rect 9335 3796 9346 3830
rect 9290 3718 9346 3796
rect 9446 4306 9502 4318
rect 9446 4272 9457 4306
rect 9491 4272 9502 4306
rect 9446 4238 9502 4272
rect 9446 4204 9457 4238
rect 9491 4204 9502 4238
rect 9446 4170 9502 4204
rect 9446 4136 9457 4170
rect 9491 4136 9502 4170
rect 9446 4102 9502 4136
rect 9446 4068 9457 4102
rect 9491 4068 9502 4102
rect 9446 4034 9502 4068
rect 9446 4000 9457 4034
rect 9491 4000 9502 4034
rect 9446 3966 9502 4000
rect 9446 3932 9457 3966
rect 9491 3932 9502 3966
rect 9446 3898 9502 3932
rect 9446 3864 9457 3898
rect 9491 3864 9502 3898
rect 9446 3830 9502 3864
rect 9446 3796 9457 3830
rect 9491 3796 9502 3830
rect 9446 3718 9502 3796
rect 9602 4306 9655 4318
rect 9602 4272 9613 4306
rect 9647 4272 9655 4306
rect 9602 4238 9655 4272
rect 9602 4204 9613 4238
rect 9647 4204 9655 4238
rect 9602 4170 9655 4204
rect 9602 4136 9613 4170
rect 9647 4136 9655 4170
rect 9602 4102 9655 4136
rect 9602 4068 9613 4102
rect 9647 4068 9655 4102
rect 9602 4034 9655 4068
rect 9602 4000 9613 4034
rect 9647 4000 9655 4034
rect 9602 3966 9655 4000
rect 9602 3932 9613 3966
rect 9647 3932 9655 3966
rect 9602 3898 9655 3932
rect 9602 3864 9613 3898
rect 9647 3864 9655 3898
rect 9602 3830 9655 3864
rect 9602 3796 9613 3830
rect 9647 3796 9655 3830
rect 9602 3718 9655 3796
rect 9729 4306 9782 4318
rect 9729 4272 9737 4306
rect 9771 4272 9782 4306
rect 9729 4238 9782 4272
rect 9729 4204 9737 4238
rect 9771 4204 9782 4238
rect 9729 4170 9782 4204
rect 9729 4136 9737 4170
rect 9771 4136 9782 4170
rect 9729 4102 9782 4136
rect 9729 4068 9737 4102
rect 9771 4068 9782 4102
rect 9729 4034 9782 4068
rect 9729 4000 9737 4034
rect 9771 4000 9782 4034
rect 9729 3966 9782 4000
rect 9729 3932 9737 3966
rect 9771 3932 9782 3966
rect 9729 3898 9782 3932
rect 9729 3864 9737 3898
rect 9771 3864 9782 3898
rect 9729 3830 9782 3864
rect 9729 3796 9737 3830
rect 9771 3796 9782 3830
rect 9729 3718 9782 3796
rect 9882 4306 9938 4318
rect 9882 4272 9893 4306
rect 9927 4272 9938 4306
rect 9882 4238 9938 4272
rect 9882 4204 9893 4238
rect 9927 4204 9938 4238
rect 9882 4170 9938 4204
rect 9882 4136 9893 4170
rect 9927 4136 9938 4170
rect 9882 4102 9938 4136
rect 9882 4068 9893 4102
rect 9927 4068 9938 4102
rect 9882 4034 9938 4068
rect 9882 4000 9893 4034
rect 9927 4000 9938 4034
rect 9882 3966 9938 4000
rect 9882 3932 9893 3966
rect 9927 3932 9938 3966
rect 9882 3898 9938 3932
rect 9882 3864 9893 3898
rect 9927 3864 9938 3898
rect 9882 3830 9938 3864
rect 9882 3796 9893 3830
rect 9927 3796 9938 3830
rect 9882 3718 9938 3796
rect 10038 4306 10094 4318
rect 10038 4272 10049 4306
rect 10083 4272 10094 4306
rect 10038 4238 10094 4272
rect 10038 4204 10049 4238
rect 10083 4204 10094 4238
rect 10038 4170 10094 4204
rect 10038 4136 10049 4170
rect 10083 4136 10094 4170
rect 10038 4102 10094 4136
rect 10038 4068 10049 4102
rect 10083 4068 10094 4102
rect 10038 4034 10094 4068
rect 10038 4000 10049 4034
rect 10083 4000 10094 4034
rect 10038 3966 10094 4000
rect 10038 3932 10049 3966
rect 10083 3932 10094 3966
rect 10038 3898 10094 3932
rect 10038 3864 10049 3898
rect 10083 3864 10094 3898
rect 10038 3830 10094 3864
rect 10038 3796 10049 3830
rect 10083 3796 10094 3830
rect 10038 3718 10094 3796
rect 10194 4306 10250 4318
rect 10194 4272 10205 4306
rect 10239 4272 10250 4306
rect 10194 4238 10250 4272
rect 10194 4204 10205 4238
rect 10239 4204 10250 4238
rect 10194 4170 10250 4204
rect 10194 4136 10205 4170
rect 10239 4136 10250 4170
rect 10194 4102 10250 4136
rect 10194 4068 10205 4102
rect 10239 4068 10250 4102
rect 10194 4034 10250 4068
rect 10194 4000 10205 4034
rect 10239 4000 10250 4034
rect 10194 3966 10250 4000
rect 10194 3932 10205 3966
rect 10239 3932 10250 3966
rect 10194 3898 10250 3932
rect 10194 3864 10205 3898
rect 10239 3864 10250 3898
rect 10194 3830 10250 3864
rect 10194 3796 10205 3830
rect 10239 3796 10250 3830
rect 10194 3718 10250 3796
rect 10350 4306 10403 4318
rect 10350 4272 10361 4306
rect 10395 4272 10403 4306
rect 10350 4238 10403 4272
rect 10350 4204 10361 4238
rect 10395 4204 10403 4238
rect 10350 4170 10403 4204
rect 10350 4136 10361 4170
rect 10395 4136 10403 4170
rect 10350 4102 10403 4136
rect 10350 4068 10361 4102
rect 10395 4068 10403 4102
rect 10350 4034 10403 4068
rect 10350 4000 10361 4034
rect 10395 4000 10403 4034
rect 10350 3966 10403 4000
rect 10350 3932 10361 3966
rect 10395 3932 10403 3966
rect 10350 3898 10403 3932
rect 10350 3864 10361 3898
rect 10395 3864 10403 3898
rect 10350 3830 10403 3864
rect 10350 3796 10361 3830
rect 10395 3796 10403 3830
rect 10350 3718 10403 3796
rect 10477 4306 10530 4318
rect 10477 4272 10485 4306
rect 10519 4272 10530 4306
rect 10477 4238 10530 4272
rect 10477 4204 10485 4238
rect 10519 4204 10530 4238
rect 10477 4170 10530 4204
rect 10477 4136 10485 4170
rect 10519 4136 10530 4170
rect 10477 4102 10530 4136
rect 10477 4068 10485 4102
rect 10519 4068 10530 4102
rect 10477 4034 10530 4068
rect 10477 4000 10485 4034
rect 10519 4000 10530 4034
rect 10477 3966 10530 4000
rect 10477 3932 10485 3966
rect 10519 3932 10530 3966
rect 10477 3898 10530 3932
rect 10477 3864 10485 3898
rect 10519 3864 10530 3898
rect 10477 3830 10530 3864
rect 10477 3796 10485 3830
rect 10519 3796 10530 3830
rect 10477 3718 10530 3796
rect 10630 4306 10686 4318
rect 10630 4272 10641 4306
rect 10675 4272 10686 4306
rect 10630 4238 10686 4272
rect 10630 4204 10641 4238
rect 10675 4204 10686 4238
rect 10630 4170 10686 4204
rect 10630 4136 10641 4170
rect 10675 4136 10686 4170
rect 10630 4102 10686 4136
rect 10630 4068 10641 4102
rect 10675 4068 10686 4102
rect 10630 4034 10686 4068
rect 10630 4000 10641 4034
rect 10675 4000 10686 4034
rect 10630 3966 10686 4000
rect 10630 3932 10641 3966
rect 10675 3932 10686 3966
rect 10630 3898 10686 3932
rect 10630 3864 10641 3898
rect 10675 3864 10686 3898
rect 10630 3830 10686 3864
rect 10630 3796 10641 3830
rect 10675 3796 10686 3830
rect 10630 3718 10686 3796
rect 10786 4306 10839 4318
rect 10786 4272 10797 4306
rect 10831 4272 10839 4306
rect 10786 4238 10839 4272
rect 12137 4281 12221 4289
rect 12137 4247 12149 4281
rect 12183 4247 12221 4281
rect 10786 4204 10797 4238
rect 10831 4204 10839 4238
rect 10786 4170 10839 4204
rect 10786 4136 10797 4170
rect 10831 4136 10839 4170
rect 11009 4201 11062 4239
rect 11009 4167 11017 4201
rect 11051 4167 11062 4201
rect 11009 4155 11062 4167
rect 11862 4201 11915 4239
rect 12137 4236 12221 4247
rect 11862 4167 11873 4201
rect 11907 4167 11915 4201
rect 11862 4155 11915 4167
rect 10786 4102 10839 4136
rect 10786 4068 10797 4102
rect 10831 4068 10839 4102
rect 10786 4034 10839 4068
rect 10786 4000 10797 4034
rect 10831 4000 10839 4034
rect 10786 3966 10839 4000
rect 10786 3932 10797 3966
rect 10831 3932 10839 3966
rect 11009 3987 11062 4025
rect 11009 3953 11017 3987
rect 11051 3953 11062 3987
rect 11009 3941 11062 3953
rect 11862 3987 11915 4025
rect 11862 3953 11873 3987
rect 11907 3953 11915 3987
rect 11862 3941 11915 3953
rect 12137 4025 12221 4036
rect 12137 3991 12149 4025
rect 12183 3991 12221 4025
rect 12137 3980 12221 3991
rect 10786 3898 10839 3932
rect 10786 3864 10797 3898
rect 10831 3864 10839 3898
rect 10786 3830 10839 3864
rect 10786 3796 10797 3830
rect 10831 3796 10839 3830
rect 10786 3718 10839 3796
rect 11009 3819 11062 3831
rect 11009 3785 11017 3819
rect 11051 3785 11062 3819
rect 11009 3747 11062 3785
rect 11862 3819 11915 3831
rect 11862 3785 11873 3819
rect 11907 3785 11915 3819
rect 11862 3747 11915 3785
rect 12137 3769 12221 3780
rect 12137 3735 12149 3769
rect 12183 3735 12221 3769
rect 12137 3727 12221 3735
rect 12137 3645 12221 3653
rect 12137 3611 12149 3645
rect 12183 3611 12221 3645
rect 11009 3567 11062 3605
rect -325 2987 -314 3021
rect -280 2987 -272 3021
rect 1684 3071 1737 3109
rect 1684 3037 1692 3071
rect 1726 3037 1737 3071
rect 1684 3025 1737 3037
rect 3337 3071 3390 3109
rect 3337 3037 3348 3071
rect 3382 3037 3390 3071
rect 3337 3025 3390 3037
rect -325 2953 -272 2987
rect -325 2919 -314 2953
rect -280 2919 -272 2953
rect -325 2907 -272 2919
rect 9748 3460 9815 3538
rect 9748 3426 9756 3460
rect 9790 3426 9815 3460
rect 9748 3392 9815 3426
rect 9748 3358 9756 3392
rect 9790 3358 9815 3392
rect 9748 3324 9815 3358
rect 9748 3290 9756 3324
rect 9790 3290 9815 3324
rect 9748 3256 9815 3290
rect 9748 3222 9756 3256
rect 9790 3222 9815 3256
rect 9748 3188 9815 3222
rect 9748 3154 9756 3188
rect 9790 3154 9815 3188
rect 9748 3120 9815 3154
rect 9748 3086 9756 3120
rect 9790 3086 9815 3120
rect 9748 3052 9815 3086
rect 9748 3018 9756 3052
rect 9790 3018 9815 3052
rect 9748 2984 9815 3018
rect 9748 2950 9756 2984
rect 9790 2950 9815 2984
rect 9748 2938 9815 2950
rect 9935 2938 9991 3538
rect 10111 3460 10195 3538
rect 10111 3426 10136 3460
rect 10170 3426 10195 3460
rect 10111 3392 10195 3426
rect 10111 3358 10136 3392
rect 10170 3358 10195 3392
rect 10111 3324 10195 3358
rect 10111 3290 10136 3324
rect 10170 3290 10195 3324
rect 10111 3256 10195 3290
rect 10111 3222 10136 3256
rect 10170 3222 10195 3256
rect 10111 3188 10195 3222
rect 10111 3154 10136 3188
rect 10170 3154 10195 3188
rect 10111 3120 10195 3154
rect 10111 3086 10136 3120
rect 10170 3086 10195 3120
rect 10111 3052 10195 3086
rect 10111 3018 10136 3052
rect 10170 3018 10195 3052
rect 10111 2984 10195 3018
rect 10111 2950 10136 2984
rect 10170 2950 10195 2984
rect 10111 2938 10195 2950
rect 10315 3460 10368 3538
rect 11009 3533 11017 3567
rect 11051 3533 11062 3567
rect 11009 3521 11062 3533
rect 11862 3567 11915 3605
rect 12137 3600 12221 3611
rect 11862 3533 11873 3567
rect 11907 3533 11915 3567
rect 11862 3521 11915 3533
rect 10315 3426 10326 3460
rect 10360 3426 10368 3460
rect 10315 3392 10368 3426
rect 10315 3358 10326 3392
rect 10360 3358 10368 3392
rect 10315 3324 10368 3358
rect 10315 3290 10326 3324
rect 10360 3290 10368 3324
rect 10315 3256 10368 3290
rect 10315 3222 10326 3256
rect 10360 3222 10368 3256
rect 10315 3188 10368 3222
rect 10315 3154 10326 3188
rect 10360 3154 10368 3188
rect 10315 3120 10368 3154
rect 10315 3086 10326 3120
rect 10360 3086 10368 3120
rect 10315 3052 10368 3086
rect 10315 3018 10326 3052
rect 10360 3018 10368 3052
rect 10315 2984 10368 3018
rect 10315 2950 10326 2984
rect 10360 2950 10368 2984
rect 10315 2938 10368 2950
rect 12137 3389 12221 3400
rect 11009 3351 11062 3389
rect 11009 3317 11017 3351
rect 11051 3317 11062 3351
rect 11009 3305 11062 3317
rect 11862 3351 11915 3389
rect 11862 3317 11873 3351
rect 11907 3317 11915 3351
rect 12137 3355 12149 3389
rect 12183 3355 12221 3389
rect 12137 3347 12221 3355
rect 11862 3305 11915 3317
rect -461 2651 -408 2669
rect -461 2617 -453 2651
rect -419 2617 -408 2651
rect -461 2583 -408 2617
rect -461 2549 -453 2583
rect -419 2549 -408 2583
rect -461 2515 -408 2549
rect -461 2481 -453 2515
rect -419 2481 -408 2515
rect -461 2469 -408 2481
rect -288 2651 -232 2669
rect -288 2617 -277 2651
rect -243 2617 -232 2651
rect -288 2583 -232 2617
rect -288 2549 -277 2583
rect -243 2549 -232 2583
rect -288 2515 -232 2549
rect -288 2481 -277 2515
rect -243 2481 -232 2515
rect -288 2469 -232 2481
rect -112 2651 -56 2669
rect -112 2617 -101 2651
rect -67 2617 -56 2651
rect -112 2583 -56 2617
rect -112 2549 -101 2583
rect -67 2549 -56 2583
rect -112 2515 -56 2549
rect -112 2481 -101 2515
rect -67 2481 -56 2515
rect -112 2469 -56 2481
rect 64 2651 117 2669
rect 64 2617 75 2651
rect 109 2617 117 2651
rect 64 2583 117 2617
rect 64 2549 75 2583
rect 109 2549 117 2583
rect 64 2515 117 2549
rect 64 2481 75 2515
rect 109 2481 117 2515
rect 64 2469 117 2481
rect -461 2389 -408 2401
rect -461 2355 -453 2389
rect -419 2355 -408 2389
rect -461 2321 -408 2355
rect -461 2287 -453 2321
rect -419 2287 -408 2321
rect -461 2253 -408 2287
rect -461 2219 -453 2253
rect -419 2219 -408 2253
rect -461 2201 -408 2219
rect -288 2389 -232 2401
rect -288 2355 -277 2389
rect -243 2355 -232 2389
rect -288 2321 -232 2355
rect -288 2287 -277 2321
rect -243 2287 -232 2321
rect -288 2253 -232 2287
rect -288 2219 -277 2253
rect -243 2219 -232 2253
rect -288 2201 -232 2219
rect -112 2389 -56 2401
rect -112 2355 -101 2389
rect -67 2355 -56 2389
rect -112 2321 -56 2355
rect -112 2287 -101 2321
rect -67 2287 -56 2321
rect -112 2253 -56 2287
rect -112 2219 -101 2253
rect -67 2219 -56 2253
rect -112 2201 -56 2219
rect 64 2389 117 2401
rect 64 2355 75 2389
rect 109 2355 117 2389
rect 64 2321 117 2355
rect 64 2287 75 2321
rect 109 2287 117 2321
rect 64 2253 117 2287
rect 64 2219 75 2253
rect 109 2219 117 2253
rect 64 2201 117 2219
rect 7414 1474 7467 1544
rect 7414 1440 7422 1474
rect 7456 1440 7467 1474
rect 7414 1406 7467 1440
rect 7414 1372 7422 1406
rect 7456 1372 7467 1406
rect 7414 1338 7467 1372
rect 7414 1304 7422 1338
rect 7456 1304 7467 1338
rect 7414 1270 7467 1304
rect 7414 1236 7422 1270
rect 7456 1236 7467 1270
rect 7414 1202 7467 1236
rect 7414 1168 7422 1202
rect 7456 1168 7467 1202
rect 7414 1134 7467 1168
rect 7414 1100 7422 1134
rect 7456 1100 7467 1134
rect 7414 1066 7467 1100
rect 7414 1032 7422 1066
rect 7456 1032 7467 1066
rect 7414 998 7467 1032
rect 7414 964 7422 998
rect 7456 964 7467 998
rect 7414 930 7467 964
rect 7414 896 7422 930
rect 7456 896 7467 930
rect 7414 862 7467 896
rect 7414 828 7422 862
rect 7456 828 7467 862
rect 7414 794 7467 828
rect 7414 760 7422 794
rect 7456 760 7467 794
rect 7414 726 7467 760
rect 7414 692 7422 726
rect 7456 692 7467 726
rect 7414 658 7467 692
rect 7414 624 7422 658
rect 7456 624 7467 658
rect 7414 590 7467 624
rect 7414 556 7422 590
rect 7456 556 7467 590
rect 7414 544 7467 556
rect 7587 1474 7643 1544
rect 7587 1440 7598 1474
rect 7632 1440 7643 1474
rect 7587 1406 7643 1440
rect 7587 1372 7598 1406
rect 7632 1372 7643 1406
rect 7587 1338 7643 1372
rect 7587 1304 7598 1338
rect 7632 1304 7643 1338
rect 7587 1270 7643 1304
rect 7587 1236 7598 1270
rect 7632 1236 7643 1270
rect 7587 1202 7643 1236
rect 7587 1168 7598 1202
rect 7632 1168 7643 1202
rect 7587 1134 7643 1168
rect 7587 1100 7598 1134
rect 7632 1100 7643 1134
rect 7587 1066 7643 1100
rect 7587 1032 7598 1066
rect 7632 1032 7643 1066
rect 7587 998 7643 1032
rect 7587 964 7598 998
rect 7632 964 7643 998
rect 7587 930 7643 964
rect 7587 896 7598 930
rect 7632 896 7643 930
rect 7587 862 7643 896
rect 7587 828 7598 862
rect 7632 828 7643 862
rect 7587 794 7643 828
rect 7587 760 7598 794
rect 7632 760 7643 794
rect 7587 726 7643 760
rect 7587 692 7598 726
rect 7632 692 7643 726
rect 7587 658 7643 692
rect 7587 624 7598 658
rect 7632 624 7643 658
rect 7587 590 7643 624
rect 7587 556 7598 590
rect 7632 556 7643 590
rect 7587 544 7643 556
rect 7763 1474 7819 1544
rect 7763 1440 7774 1474
rect 7808 1440 7819 1474
rect 7763 1406 7819 1440
rect 7763 1372 7774 1406
rect 7808 1372 7819 1406
rect 7763 1338 7819 1372
rect 7763 1304 7774 1338
rect 7808 1304 7819 1338
rect 7763 1270 7819 1304
rect 7763 1236 7774 1270
rect 7808 1236 7819 1270
rect 7763 1202 7819 1236
rect 7763 1168 7774 1202
rect 7808 1168 7819 1202
rect 7763 1134 7819 1168
rect 7763 1100 7774 1134
rect 7808 1100 7819 1134
rect 7763 1066 7819 1100
rect 7763 1032 7774 1066
rect 7808 1032 7819 1066
rect 7763 998 7819 1032
rect 7763 964 7774 998
rect 7808 964 7819 998
rect 7763 930 7819 964
rect 7763 896 7774 930
rect 7808 896 7819 930
rect 7763 862 7819 896
rect 7763 828 7774 862
rect 7808 828 7819 862
rect 7763 794 7819 828
rect 7763 760 7774 794
rect 7808 760 7819 794
rect 7763 726 7819 760
rect 7763 692 7774 726
rect 7808 692 7819 726
rect 7763 658 7819 692
rect 7763 624 7774 658
rect 7808 624 7819 658
rect 7763 590 7819 624
rect 7763 556 7774 590
rect 7808 556 7819 590
rect 7763 544 7819 556
rect 7939 1474 7992 1544
rect 7939 1440 7950 1474
rect 7984 1440 7992 1474
rect 7939 1406 7992 1440
rect 7939 1372 7950 1406
rect 7984 1372 7992 1406
rect 7939 1338 7992 1372
rect 7939 1304 7950 1338
rect 7984 1304 7992 1338
rect 7939 1270 7992 1304
rect 7939 1236 7950 1270
rect 7984 1236 7992 1270
rect 7939 1202 7992 1236
rect 7939 1168 7950 1202
rect 7984 1168 7992 1202
rect 7939 1134 7992 1168
rect 7939 1100 7950 1134
rect 7984 1100 7992 1134
rect 7939 1066 7992 1100
rect 7939 1032 7950 1066
rect 7984 1032 7992 1066
rect 7939 998 7992 1032
rect 7939 964 7950 998
rect 7984 964 7992 998
rect 7939 930 7992 964
rect 8876 1466 8929 1544
rect 8876 1432 8884 1466
rect 8918 1432 8929 1466
rect 8876 1398 8929 1432
rect 8876 1364 8884 1398
rect 8918 1364 8929 1398
rect 8876 1330 8929 1364
rect 8876 1296 8884 1330
rect 8918 1296 8929 1330
rect 8876 1262 8929 1296
rect 8876 1228 8884 1262
rect 8918 1228 8929 1262
rect 8876 1194 8929 1228
rect 8876 1160 8884 1194
rect 8918 1160 8929 1194
rect 8876 1126 8929 1160
rect 8876 1092 8884 1126
rect 8918 1092 8929 1126
rect 8876 1058 8929 1092
rect 8876 1024 8884 1058
rect 8918 1024 8929 1058
rect 8876 990 8929 1024
rect 8876 956 8884 990
rect 8918 956 8929 990
rect 8876 944 8929 956
rect 9029 1466 9085 1544
rect 9029 1432 9040 1466
rect 9074 1432 9085 1466
rect 9029 1398 9085 1432
rect 9029 1364 9040 1398
rect 9074 1364 9085 1398
rect 9029 1330 9085 1364
rect 9029 1296 9040 1330
rect 9074 1296 9085 1330
rect 9029 1262 9085 1296
rect 9029 1228 9040 1262
rect 9074 1228 9085 1262
rect 9029 1194 9085 1228
rect 9029 1160 9040 1194
rect 9074 1160 9085 1194
rect 9029 1126 9085 1160
rect 9029 1092 9040 1126
rect 9074 1092 9085 1126
rect 9029 1058 9085 1092
rect 9029 1024 9040 1058
rect 9074 1024 9085 1058
rect 9029 990 9085 1024
rect 9029 956 9040 990
rect 9074 956 9085 990
rect 9029 944 9085 956
rect 9185 1466 9241 1544
rect 9185 1432 9196 1466
rect 9230 1432 9241 1466
rect 9185 1398 9241 1432
rect 9185 1364 9196 1398
rect 9230 1364 9241 1398
rect 9185 1330 9241 1364
rect 9185 1296 9196 1330
rect 9230 1296 9241 1330
rect 9185 1262 9241 1296
rect 9185 1228 9196 1262
rect 9230 1228 9241 1262
rect 9185 1194 9241 1228
rect 9185 1160 9196 1194
rect 9230 1160 9241 1194
rect 9185 1126 9241 1160
rect 9185 1092 9196 1126
rect 9230 1092 9241 1126
rect 9185 1058 9241 1092
rect 9185 1024 9196 1058
rect 9230 1024 9241 1058
rect 9185 990 9241 1024
rect 9185 956 9196 990
rect 9230 956 9241 990
rect 9185 944 9241 956
rect 9341 1466 9397 1544
rect 9341 1432 9352 1466
rect 9386 1432 9397 1466
rect 9341 1398 9397 1432
rect 9341 1364 9352 1398
rect 9386 1364 9397 1398
rect 9341 1330 9397 1364
rect 9341 1296 9352 1330
rect 9386 1296 9397 1330
rect 9341 1262 9397 1296
rect 9341 1228 9352 1262
rect 9386 1228 9397 1262
rect 9341 1194 9397 1228
rect 9341 1160 9352 1194
rect 9386 1160 9397 1194
rect 9341 1126 9397 1160
rect 9341 1092 9352 1126
rect 9386 1092 9397 1126
rect 9341 1058 9397 1092
rect 9341 1024 9352 1058
rect 9386 1024 9397 1058
rect 9341 990 9397 1024
rect 9341 956 9352 990
rect 9386 956 9397 990
rect 9341 944 9397 956
rect 9497 1466 9550 1544
rect 9497 1432 9508 1466
rect 9542 1432 9550 1466
rect 9497 1398 9550 1432
rect 9497 1364 9508 1398
rect 9542 1364 9550 1398
rect 9497 1330 9550 1364
rect 9497 1296 9508 1330
rect 9542 1296 9550 1330
rect 9497 1262 9550 1296
rect 9497 1228 9508 1262
rect 9542 1228 9550 1262
rect 9497 1194 9550 1228
rect 9497 1160 9508 1194
rect 9542 1160 9550 1194
rect 9497 1126 9550 1160
rect 9497 1092 9508 1126
rect 9542 1092 9550 1126
rect 9497 1058 9550 1092
rect 9497 1024 9508 1058
rect 9542 1024 9550 1058
rect 9497 990 9550 1024
rect 9497 956 9508 990
rect 9542 956 9550 990
rect 9497 944 9550 956
rect 9748 1466 9801 1544
rect 9748 1432 9756 1466
rect 9790 1432 9801 1466
rect 9748 1398 9801 1432
rect 9748 1364 9756 1398
rect 9790 1364 9801 1398
rect 9748 1330 9801 1364
rect 9748 1296 9756 1330
rect 9790 1296 9801 1330
rect 9748 1262 9801 1296
rect 9748 1228 9756 1262
rect 9790 1228 9801 1262
rect 9748 1194 9801 1228
rect 9748 1160 9756 1194
rect 9790 1160 9801 1194
rect 9748 1126 9801 1160
rect 9748 1092 9756 1126
rect 9790 1092 9801 1126
rect 9748 1058 9801 1092
rect 9748 1024 9756 1058
rect 9790 1024 9801 1058
rect 9748 990 9801 1024
rect 9748 956 9756 990
rect 9790 956 9801 990
rect 9748 944 9801 956
rect 9901 1466 9957 1544
rect 9901 1432 9912 1466
rect 9946 1432 9957 1466
rect 9901 1398 9957 1432
rect 9901 1364 9912 1398
rect 9946 1364 9957 1398
rect 9901 1330 9957 1364
rect 9901 1296 9912 1330
rect 9946 1296 9957 1330
rect 9901 1262 9957 1296
rect 9901 1228 9912 1262
rect 9946 1228 9957 1262
rect 9901 1194 9957 1228
rect 9901 1160 9912 1194
rect 9946 1160 9957 1194
rect 9901 1126 9957 1160
rect 9901 1092 9912 1126
rect 9946 1092 9957 1126
rect 9901 1058 9957 1092
rect 9901 1024 9912 1058
rect 9946 1024 9957 1058
rect 9901 990 9957 1024
rect 9901 956 9912 990
rect 9946 956 9957 990
rect 9901 944 9957 956
rect 10057 1466 10113 1544
rect 10057 1432 10068 1466
rect 10102 1432 10113 1466
rect 10057 1398 10113 1432
rect 10057 1364 10068 1398
rect 10102 1364 10113 1398
rect 10057 1330 10113 1364
rect 10057 1296 10068 1330
rect 10102 1296 10113 1330
rect 10057 1262 10113 1296
rect 10057 1228 10068 1262
rect 10102 1228 10113 1262
rect 10057 1194 10113 1228
rect 10057 1160 10068 1194
rect 10102 1160 10113 1194
rect 10057 1126 10113 1160
rect 10057 1092 10068 1126
rect 10102 1092 10113 1126
rect 10057 1058 10113 1092
rect 10057 1024 10068 1058
rect 10102 1024 10113 1058
rect 10057 990 10113 1024
rect 10057 956 10068 990
rect 10102 956 10113 990
rect 10057 944 10113 956
rect 10213 1466 10269 1544
rect 10213 1432 10224 1466
rect 10258 1432 10269 1466
rect 10213 1398 10269 1432
rect 10213 1364 10224 1398
rect 10258 1364 10269 1398
rect 10213 1330 10269 1364
rect 10213 1296 10224 1330
rect 10258 1296 10269 1330
rect 10213 1262 10269 1296
rect 10213 1228 10224 1262
rect 10258 1228 10269 1262
rect 10213 1194 10269 1228
rect 10213 1160 10224 1194
rect 10258 1160 10269 1194
rect 10213 1126 10269 1160
rect 10213 1092 10224 1126
rect 10258 1092 10269 1126
rect 10213 1058 10269 1092
rect 10213 1024 10224 1058
rect 10258 1024 10269 1058
rect 10213 990 10269 1024
rect 10213 956 10224 990
rect 10258 956 10269 990
rect 10213 944 10269 956
rect 10369 1466 10422 1544
rect 10369 1432 10380 1466
rect 10414 1432 10422 1466
rect 10369 1398 10422 1432
rect 10369 1364 10380 1398
rect 10414 1364 10422 1398
rect 10369 1330 10422 1364
rect 10369 1296 10380 1330
rect 10414 1296 10422 1330
rect 10369 1262 10422 1296
rect 10369 1228 10380 1262
rect 10414 1228 10422 1262
rect 10369 1194 10422 1228
rect 10369 1160 10380 1194
rect 10414 1160 10422 1194
rect 10369 1126 10422 1160
rect 10564 1443 10617 1455
rect 10564 1409 10572 1443
rect 10606 1409 10617 1443
rect 10564 1375 10617 1409
rect 10564 1341 10572 1375
rect 10606 1341 10617 1375
rect 10564 1307 10617 1341
rect 10564 1273 10572 1307
rect 10606 1273 10617 1307
rect 10564 1239 10617 1273
rect 10564 1205 10572 1239
rect 10606 1205 10617 1239
rect 10564 1155 10617 1205
rect 10717 1443 10773 1455
rect 10717 1409 10728 1443
rect 10762 1409 10773 1443
rect 10717 1375 10773 1409
rect 10717 1341 10728 1375
rect 10762 1341 10773 1375
rect 10717 1307 10773 1341
rect 10717 1273 10728 1307
rect 10762 1273 10773 1307
rect 10717 1239 10773 1273
rect 10717 1205 10728 1239
rect 10762 1205 10773 1239
rect 10717 1155 10773 1205
rect 10873 1443 10929 1455
rect 10873 1409 10884 1443
rect 10918 1409 10929 1443
rect 10873 1375 10929 1409
rect 10873 1341 10884 1375
rect 10918 1341 10929 1375
rect 10873 1307 10929 1341
rect 10873 1273 10884 1307
rect 10918 1273 10929 1307
rect 10873 1239 10929 1273
rect 10873 1205 10884 1239
rect 10918 1205 10929 1239
rect 10873 1155 10929 1205
rect 11029 1443 11085 1455
rect 11029 1409 11040 1443
rect 11074 1409 11085 1443
rect 11029 1375 11085 1409
rect 11029 1341 11040 1375
rect 11074 1341 11085 1375
rect 11029 1307 11085 1341
rect 11029 1273 11040 1307
rect 11074 1273 11085 1307
rect 11029 1239 11085 1273
rect 11029 1205 11040 1239
rect 11074 1205 11085 1239
rect 11029 1155 11085 1205
rect 11185 1443 11238 1455
rect 11185 1409 11196 1443
rect 11230 1409 11238 1443
rect 11185 1375 11238 1409
rect 11185 1341 11196 1375
rect 11230 1341 11238 1375
rect 11185 1307 11238 1341
rect 11185 1273 11196 1307
rect 11230 1273 11238 1307
rect 11185 1239 11238 1273
rect 11361 1337 11414 1349
rect 11361 1303 11369 1337
rect 11403 1303 11414 1337
rect 11361 1265 11414 1303
rect 12214 1337 12267 1349
rect 12214 1303 12225 1337
rect 12259 1303 12267 1337
rect 12214 1265 12267 1303
rect 11185 1205 11196 1239
rect 11230 1205 11238 1239
rect 11185 1155 11238 1205
rect 10369 1092 10380 1126
rect 10414 1092 10422 1126
rect 10369 1058 10422 1092
rect 10369 1024 10380 1058
rect 10414 1024 10422 1058
rect 10369 990 10422 1024
rect 10369 956 10380 990
rect 10414 956 10422 990
rect 10369 944 10422 956
rect 7939 896 7950 930
rect 7984 896 7992 930
rect 7939 862 7992 896
rect 7939 828 7950 862
rect 7984 828 7992 862
rect 10849 915 10902 927
rect 10849 881 10857 915
rect 10891 881 10902 915
rect 10849 843 10902 881
rect 11302 915 11358 927
rect 11302 881 11313 915
rect 11347 881 11358 915
rect 11302 843 11358 881
rect 11758 915 11814 927
rect 11758 881 11769 915
rect 11803 881 11814 915
rect 11758 843 11814 881
rect 12214 915 12267 927
rect 12214 881 12225 915
rect 12259 881 12267 915
rect 12214 843 12267 881
rect 7939 794 7992 828
rect 7939 760 7950 794
rect 7984 760 7992 794
rect 7939 726 7992 760
rect 7939 692 7950 726
rect 7984 692 7992 726
rect 7939 658 7992 692
rect 7939 624 7950 658
rect 7984 624 7992 658
rect 7939 590 7992 624
rect 7939 556 7950 590
rect 7984 556 7992 590
rect 7939 544 7992 556
rect 10398 631 10451 643
rect 10398 597 10406 631
rect 10440 597 10451 631
rect 10398 563 10451 597
rect 10398 529 10406 563
rect 10440 529 10451 563
rect 10398 495 10451 529
rect 10398 461 10406 495
rect 10440 461 10451 495
rect 10398 443 10451 461
rect 10551 631 10607 643
rect 10551 597 10562 631
rect 10596 597 10607 631
rect 10551 563 10607 597
rect 10551 529 10562 563
rect 10596 529 10607 563
rect 10551 495 10607 529
rect 10551 461 10562 495
rect 10596 461 10607 495
rect 10551 443 10607 461
rect 10707 631 10760 643
rect 10707 597 10718 631
rect 10752 597 10760 631
rect 10707 563 10760 597
rect 10707 529 10718 563
rect 10752 529 10760 563
rect 10900 631 10953 643
rect 10900 597 10908 631
rect 10942 597 10953 631
rect 10900 559 10953 597
rect 11053 631 11109 643
rect 11053 597 11064 631
rect 11098 597 11109 631
rect 11053 559 11109 597
rect 11209 631 11262 643
rect 11209 597 11220 631
rect 11254 597 11262 631
rect 11209 559 11262 597
rect 11336 631 11389 643
rect 11336 597 11344 631
rect 11378 597 11389 631
rect 11336 559 11389 597
rect 11489 631 11545 643
rect 11489 597 11500 631
rect 11534 597 11545 631
rect 11489 559 11545 597
rect 11645 631 11698 643
rect 11645 597 11656 631
rect 11690 597 11698 631
rect 11645 559 11698 597
rect 10707 495 10760 529
rect 10707 461 10718 495
rect 10752 461 10760 495
rect 10707 443 10760 461
<< mvndiffc >>
rect -453 4121 -419 4155
rect -453 4053 -419 4087
rect -277 4121 -243 4155
rect -277 4053 -243 4087
rect 75 4121 109 4155
rect 75 4053 109 4087
rect -470 3773 -436 3807
rect -314 3773 -280 3807
rect -190 3785 -156 3819
rect -190 3717 -156 3751
rect -14 3785 20 3819
rect -14 3717 20 3751
rect 8366 4067 8400 4101
rect 8510 4067 8544 4101
rect 8366 3211 8400 3245
rect 8510 3211 8544 3245
rect 7542 2924 7576 2958
rect 7542 2856 7576 2890
rect 7542 2788 7576 2822
rect 7718 2924 7752 2958
rect 7718 2856 7752 2890
rect 7718 2788 7752 2822
rect 7894 2924 7928 2958
rect 7894 2856 7928 2890
rect 7894 2788 7928 2822
rect 8070 2924 8104 2958
rect 8070 2856 8104 2890
rect 8070 2788 8104 2822
rect 8246 2924 8280 2958
rect 8246 2856 8280 2890
rect 8246 2788 8280 2822
rect 8422 2924 8456 2958
rect 8422 2856 8456 2890
rect 8422 2788 8456 2822
rect 8678 2924 8712 2958
rect 8678 2856 8712 2890
rect 8678 2788 8712 2822
rect 8934 2924 8968 2958
rect 8934 2856 8968 2890
rect 8934 2788 8968 2822
rect 9190 2924 9224 2958
rect 9190 2856 9224 2890
rect 9190 2788 9224 2822
rect 9446 2924 9480 2958
rect 9446 2856 9480 2890
rect 9446 2788 9480 2822
rect 8678 2662 8712 2696
rect 7680 2608 7714 2642
rect 7748 2608 7782 2642
rect 7816 2608 7850 2642
rect 7884 2608 7918 2642
rect 7952 2608 7986 2642
rect 8020 2608 8054 2642
rect 8088 2608 8122 2642
rect 8156 2608 8190 2642
rect 8224 2608 8258 2642
rect 8292 2608 8326 2642
rect 8360 2608 8394 2642
rect 8428 2608 8462 2642
rect 8496 2608 8530 2642
rect 8564 2608 8598 2642
rect 8678 2594 8712 2628
rect 8678 2526 8712 2560
rect 7680 2432 7714 2466
rect 7748 2432 7782 2466
rect 7816 2432 7850 2466
rect 7884 2432 7918 2466
rect 7952 2432 7986 2466
rect 8020 2432 8054 2466
rect 8088 2432 8122 2466
rect 8156 2432 8190 2466
rect 8224 2432 8258 2466
rect 8292 2432 8326 2466
rect 8360 2432 8394 2466
rect 8428 2432 8462 2466
rect 8496 2432 8530 2466
rect 8564 2432 8598 2466
rect 8678 2458 8712 2492
rect 8678 2390 8712 2424
rect 8678 2322 8712 2356
rect -453 1957 -419 1991
rect -453 1889 -419 1923
rect -277 1957 -243 1991
rect -277 1889 -243 1923
rect 75 1957 109 1991
rect 75 1889 109 1923
rect 7578 2261 7612 2295
rect 7578 2193 7612 2227
rect 7578 2125 7612 2159
rect 7578 2057 7612 2091
rect 7578 1989 7612 2023
rect 7578 1921 7612 1955
rect 7578 1853 7612 1887
rect 7578 1785 7612 1819
rect 7754 2261 7788 2295
rect 7754 2193 7788 2227
rect 7754 2125 7788 2159
rect 7754 2057 7788 2091
rect 7754 1989 7788 2023
rect 7754 1921 7788 1955
rect 7754 1853 7788 1887
rect 7754 1785 7788 1819
rect 7930 2261 7964 2295
rect 7930 2193 7964 2227
rect 7930 2125 7964 2159
rect 7930 2057 7964 2091
rect 7930 1989 7964 2023
rect 7930 1921 7964 1955
rect 7930 1853 7964 1887
rect 7930 1785 7964 1819
rect 8678 2254 8712 2288
rect 8678 2186 8712 2220
rect 8678 2118 8712 2152
rect 8678 2050 8712 2084
rect 8678 1982 8712 2016
rect 8678 1914 8712 1948
rect 8678 1846 8712 1880
rect 8678 1778 8712 1812
rect 8854 2662 8888 2696
rect 8854 2594 8888 2628
rect 8968 2608 9002 2642
rect 9036 2608 9070 2642
rect 9104 2608 9138 2642
rect 9172 2608 9206 2642
rect 9240 2608 9274 2642
rect 9308 2608 9342 2642
rect 9376 2608 9410 2642
rect 9444 2608 9478 2642
rect 9756 2632 9790 2666
rect 8854 2526 8888 2560
rect 8854 2458 8888 2492
rect 9756 2564 9790 2598
rect 9756 2496 9790 2530
rect 8968 2452 9002 2486
rect 9036 2452 9070 2486
rect 9104 2452 9138 2486
rect 9172 2452 9206 2486
rect 9240 2452 9274 2486
rect 9308 2452 9342 2486
rect 9376 2452 9410 2486
rect 9444 2452 9478 2486
rect 9946 2632 9980 2666
rect 9946 2564 9980 2598
rect 9946 2496 9980 2530
rect 10136 2632 10170 2666
rect 10136 2564 10170 2598
rect 10136 2496 10170 2530
rect 10326 2632 10360 2666
rect 10326 2564 10360 2598
rect 10860 3015 10894 3049
rect 10860 2947 10894 2981
rect 10860 2879 10894 2913
rect 10860 2811 10894 2845
rect 10860 2743 10894 2777
rect 10860 2675 10894 2709
rect 10860 2607 10894 2641
rect 10860 2539 10894 2573
rect 10326 2496 10360 2530
rect 11036 3015 11070 3049
rect 11036 2947 11070 2981
rect 11036 2879 11070 2913
rect 11036 2811 11070 2845
rect 11036 2743 11070 2777
rect 11036 2675 11070 2709
rect 11036 2607 11070 2641
rect 11036 2539 11070 2573
rect 11212 3015 11246 3049
rect 11212 2947 11246 2981
rect 11212 2879 11246 2913
rect 11212 2811 11246 2845
rect 11212 2743 11246 2777
rect 11212 2675 11246 2709
rect 11212 2607 11246 2641
rect 11212 2539 11246 2573
rect 11388 3015 11422 3049
rect 11388 2947 11422 2981
rect 11388 2879 11422 2913
rect 11388 2811 11422 2845
rect 11388 2743 11422 2777
rect 11388 2675 11422 2709
rect 11388 2607 11422 2641
rect 11388 2539 11422 2573
rect 11564 3015 11598 3049
rect 11564 2947 11598 2981
rect 11564 2879 11598 2913
rect 11564 2811 11598 2845
rect 11564 2743 11598 2777
rect 11564 2675 11598 2709
rect 11564 2607 11598 2641
rect 11564 2539 11598 2573
rect 11740 3015 11774 3049
rect 11740 2947 11774 2981
rect 11740 2879 11774 2913
rect 11740 2811 11774 2845
rect 11740 2743 11774 2777
rect 11740 2675 11774 2709
rect 11740 2607 11774 2641
rect 11740 2539 11774 2573
rect 11916 3015 11950 3049
rect 11916 2947 11950 2981
rect 11916 2879 11950 2913
rect 11916 2811 11950 2845
rect 11916 2743 11950 2777
rect 11916 2675 11950 2709
rect 11916 2607 11950 2641
rect 11916 2539 11950 2573
rect 12092 3015 12126 3049
rect 12092 2947 12126 2981
rect 12092 2879 12126 2913
rect 12092 2811 12126 2845
rect 12092 2743 12126 2777
rect 12092 2675 12126 2709
rect 12092 2607 12126 2641
rect 12092 2539 12126 2573
rect 8854 2390 8888 2424
rect 8854 2322 8888 2356
rect 10784 2326 10818 2360
rect 8854 2254 8888 2288
rect 8854 2186 8888 2220
rect 8854 2118 8888 2152
rect 8854 2050 8888 2084
rect 8854 1982 8888 2016
rect 8854 1914 8888 1948
rect 8854 1846 8888 1880
rect 8854 1778 8888 1812
rect 8977 2262 9011 2296
rect 8977 2194 9011 2228
rect 8977 2126 9011 2160
rect 8977 2058 9011 2092
rect 8977 1990 9011 2024
rect 8977 1922 9011 1956
rect 8977 1854 9011 1888
rect 8977 1786 9011 1820
rect 9153 2262 9187 2296
rect 9153 2194 9187 2228
rect 9153 2126 9187 2160
rect 9153 2058 9187 2092
rect 9153 1990 9187 2024
rect 9153 1922 9187 1956
rect 9153 1854 9187 1888
rect 9153 1786 9187 1820
rect 9329 2262 9363 2296
rect 9329 2194 9363 2228
rect 9329 2126 9363 2160
rect 9329 2058 9363 2092
rect 9329 1990 9363 2024
rect 9329 1922 9363 1956
rect 9329 1854 9363 1888
rect 9329 1786 9363 1820
rect 9664 2262 9698 2296
rect 9664 2194 9698 2228
rect 9664 2126 9698 2160
rect 9664 2058 9698 2092
rect 9664 1990 9698 2024
rect 9664 1922 9698 1956
rect 9664 1854 9698 1888
rect 9664 1786 9698 1820
rect 9840 2262 9874 2296
rect 9840 2194 9874 2228
rect 9840 2126 9874 2160
rect 9840 2058 9874 2092
rect 9840 1990 9874 2024
rect 9840 1922 9874 1956
rect 9840 1854 9874 1888
rect 9840 1786 9874 1820
rect 10016 2262 10050 2296
rect 10016 2194 10050 2228
rect 10016 2126 10050 2160
rect 10016 2058 10050 2092
rect 10016 1990 10050 2024
rect 10016 1922 10050 1956
rect 10016 1854 10050 1888
rect 10016 1786 10050 1820
rect 10192 2262 10226 2296
rect 10192 2194 10226 2228
rect 10192 2126 10226 2160
rect 10192 2058 10226 2092
rect 10192 1990 10226 2024
rect 10192 1922 10226 1956
rect 10192 1854 10226 1888
rect 10192 1786 10226 1820
rect 10368 2262 10402 2296
rect 10368 2194 10402 2228
rect 10368 2126 10402 2160
rect 10368 2058 10402 2092
rect 10368 1990 10402 2024
rect 10368 1922 10402 1956
rect 10368 1854 10402 1888
rect 10368 1786 10402 1820
rect 10784 2258 10818 2292
rect 10784 2190 10818 2224
rect 10784 2122 10818 2156
rect 10784 2054 10818 2088
rect 10784 1986 10818 2020
rect 10784 1918 10818 1952
rect 10784 1850 10818 1884
rect 10960 2326 10994 2360
rect 10960 2258 10994 2292
rect 10960 2190 10994 2224
rect 10960 2122 10994 2156
rect 10960 2054 10994 2088
rect 10960 1986 10994 2020
rect 10960 1918 10994 1952
rect 10960 1850 10994 1884
rect 11136 2326 11170 2360
rect 11136 2258 11170 2292
rect 11136 2190 11170 2224
rect 11136 2122 11170 2156
rect 11136 2054 11170 2088
rect 11136 1986 11170 2020
rect 11136 1918 11170 1952
rect 11136 1850 11170 1884
rect 11312 2326 11346 2360
rect 11312 2258 11346 2292
rect 11312 2190 11346 2224
rect 11312 2122 11346 2156
rect 11312 2054 11346 2088
rect 11312 1986 11346 2020
rect 11312 1918 11346 1952
rect 11312 1850 11346 1884
rect 11488 2326 11522 2360
rect 11488 2258 11522 2292
rect 11488 2190 11522 2224
rect 11488 2122 11522 2156
rect 11488 2054 11522 2088
rect 11488 1986 11522 2020
rect 11488 1918 11522 1952
rect 11488 1850 11522 1884
rect 11664 2326 11698 2360
rect 11664 2258 11698 2292
rect 11664 2190 11698 2224
rect 11664 2122 11698 2156
rect 11664 2054 11698 2088
rect 11664 1986 11698 2020
rect 11664 1918 11698 1952
rect 11664 1850 11698 1884
rect 11840 2326 11874 2360
rect 11840 2258 11874 2292
rect 11840 2190 11874 2224
rect 11840 2122 11874 2156
rect 11840 2054 11874 2088
rect 11840 1986 11874 2020
rect 11840 1918 11874 1952
rect 11840 1850 11874 1884
rect 12016 2326 12050 2360
rect 12016 2258 12050 2292
rect 12016 2190 12050 2224
rect 12016 2122 12050 2156
rect 12016 2054 12050 2088
rect 12016 1986 12050 2020
rect 12016 1918 12050 1952
rect 12016 1850 12050 1884
<< mvpdiffc >>
rect -453 4781 -419 4815
rect -453 4713 -419 4747
rect -453 4645 -419 4679
rect -277 4781 -243 4815
rect -277 4713 -243 4747
rect -277 4645 -243 4679
rect -101 4781 -67 4815
rect -101 4713 -67 4747
rect -101 4645 -67 4679
rect 75 4781 109 4815
rect 75 4713 109 4747
rect 75 4645 109 4679
rect -453 4519 -419 4553
rect -453 4451 -419 4485
rect -453 4383 -419 4417
rect -277 4519 -243 4553
rect -277 4451 -243 4485
rect -277 4383 -243 4417
rect -101 4519 -67 4553
rect -101 4451 -67 4485
rect -101 4383 -67 4417
rect 75 4519 109 4553
rect 75 4451 109 4485
rect 75 4383 109 4417
rect -470 3395 -436 3429
rect -470 3327 -436 3361
rect -470 3259 -436 3293
rect -470 3191 -436 3225
rect -470 3123 -436 3157
rect -470 3055 -436 3089
rect -470 2987 -436 3021
rect -470 2919 -436 2953
rect -314 3395 -280 3429
rect -314 3327 -280 3361
rect -190 3455 -156 3489
rect -190 3387 -156 3421
rect -190 3319 -156 3353
rect -14 3455 20 3489
rect -14 3387 20 3421
rect -14 3319 20 3353
rect -314 3259 -280 3293
rect -314 3191 -280 3225
rect -314 3123 -280 3157
rect -314 3055 -280 3089
rect -190 3193 -156 3227
rect -190 3125 -156 3159
rect -190 3057 -156 3091
rect -14 3193 20 3227
rect -14 3125 20 3159
rect -14 3057 20 3091
rect 1114 4099 1148 4133
rect 1114 4031 1148 4065
rect 1114 3963 1148 3997
rect 1114 3895 1148 3929
rect 1114 3827 1148 3861
rect 1114 3759 1148 3793
rect 1114 3691 1148 3725
rect 1114 3623 1148 3657
rect 1114 3555 1148 3589
rect 1114 3487 1148 3521
rect 1114 3419 1148 3453
rect 1114 3351 1148 3385
rect 1114 3283 1148 3317
rect 1114 3215 1148 3249
rect 1270 4099 1304 4133
rect 1270 4031 1304 4065
rect 1270 3963 1304 3997
rect 1270 3895 1304 3929
rect 1270 3827 1304 3861
rect 1270 3759 1304 3793
rect 1270 3691 1304 3725
rect 1270 3623 1304 3657
rect 1270 3555 1304 3589
rect 1270 3487 1304 3521
rect 1270 3419 1304 3453
rect 1270 3351 1304 3385
rect 1270 3283 1304 3317
rect 1270 3215 1304 3249
rect 1426 4099 1460 4133
rect 1426 4031 1460 4065
rect 1426 3963 1460 3997
rect 1426 3895 1460 3929
rect 1426 3827 1460 3861
rect 1426 3759 1460 3793
rect 1426 3691 1460 3725
rect 1426 3623 1460 3657
rect 1426 3555 1460 3589
rect 1426 3487 1460 3521
rect 1426 3419 1460 3453
rect 1426 3351 1460 3385
rect 1426 3283 1460 3317
rect 1426 3215 1460 3249
rect 1536 4099 1570 4133
rect 1536 4031 1570 4065
rect 1536 3963 1570 3997
rect 1536 3895 1570 3929
rect 1536 3827 1570 3861
rect 1536 3759 1570 3793
rect 1536 3691 1570 3725
rect 1536 3623 1570 3657
rect 1536 3555 1570 3589
rect 1536 3487 1570 3521
rect 1536 3419 1570 3453
rect 1536 3351 1570 3385
rect 1536 3283 1570 3317
rect 1536 3215 1570 3249
rect 1692 4099 1726 4133
rect 1692 4031 1726 4065
rect 1692 3963 1726 3997
rect 1692 3895 1726 3929
rect 1692 3827 1726 3861
rect 1692 3759 1726 3793
rect 1692 3691 1726 3725
rect 1692 3623 1726 3657
rect 1692 3555 1726 3589
rect 1692 3487 1726 3521
rect 1692 3419 1726 3453
rect 1692 3351 1726 3385
rect 1692 3283 1726 3317
rect 1692 3215 1726 3249
rect 1848 4099 1882 4133
rect 1848 4031 1882 4065
rect 1848 3963 1882 3997
rect 1848 3895 1882 3929
rect 1848 3827 1882 3861
rect 1848 3759 1882 3793
rect 1848 3691 1882 3725
rect 1848 3623 1882 3657
rect 1848 3555 1882 3589
rect 1848 3487 1882 3521
rect 1848 3419 1882 3453
rect 1848 3351 1882 3385
rect 1848 3283 1882 3317
rect 1848 3215 1882 3249
rect 2004 4099 2038 4133
rect 2004 4031 2038 4065
rect 2004 3963 2038 3997
rect 2004 3895 2038 3929
rect 2004 3827 2038 3861
rect 2004 3759 2038 3793
rect 2004 3691 2038 3725
rect 2004 3623 2038 3657
rect 2004 3555 2038 3589
rect 2004 3487 2038 3521
rect 2004 3419 2038 3453
rect 2004 3351 2038 3385
rect 2004 3283 2038 3317
rect 2004 3215 2038 3249
rect 2160 4099 2194 4133
rect 2160 4031 2194 4065
rect 2160 3963 2194 3997
rect 2160 3895 2194 3929
rect 2160 3827 2194 3861
rect 2160 3759 2194 3793
rect 2160 3691 2194 3725
rect 2160 3623 2194 3657
rect 2160 3555 2194 3589
rect 2160 3487 2194 3521
rect 2160 3419 2194 3453
rect 2160 3351 2194 3385
rect 2160 3283 2194 3317
rect 2160 3215 2194 3249
rect 2316 4099 2350 4133
rect 2316 4031 2350 4065
rect 2316 3963 2350 3997
rect 2316 3895 2350 3929
rect 2316 3827 2350 3861
rect 2316 3759 2350 3793
rect 2316 3691 2350 3725
rect 2316 3623 2350 3657
rect 2316 3555 2350 3589
rect 2316 3487 2350 3521
rect 2316 3419 2350 3453
rect 2316 3351 2350 3385
rect 2316 3283 2350 3317
rect 2316 3215 2350 3249
rect 2472 4099 2506 4133
rect 2472 4031 2506 4065
rect 2472 3963 2506 3997
rect 2472 3895 2506 3929
rect 2472 3827 2506 3861
rect 2472 3759 2506 3793
rect 2472 3691 2506 3725
rect 2472 3623 2506 3657
rect 2472 3555 2506 3589
rect 2472 3487 2506 3521
rect 2472 3419 2506 3453
rect 2472 3351 2506 3385
rect 2472 3283 2506 3317
rect 2472 3215 2506 3249
rect 2628 4099 2662 4133
rect 2628 4031 2662 4065
rect 2628 3963 2662 3997
rect 2628 3895 2662 3929
rect 2628 3827 2662 3861
rect 2628 3759 2662 3793
rect 2628 3691 2662 3725
rect 2628 3623 2662 3657
rect 2628 3555 2662 3589
rect 2628 3487 2662 3521
rect 2628 3419 2662 3453
rect 2628 3351 2662 3385
rect 2628 3283 2662 3317
rect 2628 3215 2662 3249
rect 2784 4099 2818 4133
rect 2784 4031 2818 4065
rect 2784 3963 2818 3997
rect 2784 3895 2818 3929
rect 2784 3827 2818 3861
rect 2784 3759 2818 3793
rect 2784 3691 2818 3725
rect 2784 3623 2818 3657
rect 2784 3555 2818 3589
rect 2784 3487 2818 3521
rect 2784 3419 2818 3453
rect 2784 3351 2818 3385
rect 2784 3283 2818 3317
rect 2784 3215 2818 3249
rect 2980 4099 3014 4133
rect 2980 4031 3014 4065
rect 2980 3963 3014 3997
rect 2980 3895 3014 3929
rect 2980 3827 3014 3861
rect 2980 3759 3014 3793
rect 2980 3691 3014 3725
rect 2980 3623 3014 3657
rect 2980 3555 3014 3589
rect 2980 3487 3014 3521
rect 2980 3419 3014 3453
rect 2980 3351 3014 3385
rect 2980 3283 3014 3317
rect 2980 3215 3014 3249
rect 3136 4099 3170 4133
rect 3136 4031 3170 4065
rect 3136 3963 3170 3997
rect 3136 3895 3170 3929
rect 3136 3827 3170 3861
rect 3136 3759 3170 3793
rect 3136 3691 3170 3725
rect 3136 3623 3170 3657
rect 3136 3555 3170 3589
rect 3136 3487 3170 3521
rect 3136 3419 3170 3453
rect 3136 3351 3170 3385
rect 3136 3283 3170 3317
rect 3136 3215 3170 3249
rect 3292 4099 3326 4133
rect 3292 4031 3326 4065
rect 3292 3963 3326 3997
rect 3292 3895 3326 3929
rect 3292 3827 3326 3861
rect 3292 3759 3326 3793
rect 3292 3691 3326 3725
rect 3292 3623 3326 3657
rect 3292 3555 3326 3589
rect 3292 3487 3326 3521
rect 3292 3419 3326 3453
rect 3292 3351 3326 3385
rect 3292 3283 3326 3317
rect 3292 3215 3326 3249
rect 3448 4099 3482 4133
rect 3448 4031 3482 4065
rect 3448 3963 3482 3997
rect 3448 3895 3482 3929
rect 3448 3827 3482 3861
rect 3448 3759 3482 3793
rect 3448 3691 3482 3725
rect 3448 3623 3482 3657
rect 3448 3555 3482 3589
rect 3448 3487 3482 3521
rect 3448 3419 3482 3453
rect 3448 3351 3482 3385
rect 3448 3283 3482 3317
rect 3448 3215 3482 3249
rect 3604 4099 3638 4133
rect 3604 4031 3638 4065
rect 3604 3963 3638 3997
rect 3604 3895 3638 3929
rect 3604 3827 3638 3861
rect 3604 3759 3638 3793
rect 3604 3691 3638 3725
rect 3604 3623 3638 3657
rect 3604 3555 3638 3589
rect 3604 3487 3638 3521
rect 3604 3419 3638 3453
rect 3604 3351 3638 3385
rect 3604 3283 3638 3317
rect 3604 3215 3638 3249
rect 3760 4099 3794 4133
rect 3760 4031 3794 4065
rect 3760 3963 3794 3997
rect 3760 3895 3794 3929
rect 3760 3827 3794 3861
rect 3760 3759 3794 3793
rect 3760 3691 3794 3725
rect 3760 3623 3794 3657
rect 3760 3555 3794 3589
rect 3760 3487 3794 3521
rect 3760 3419 3794 3453
rect 3760 3351 3794 3385
rect 3760 3283 3794 3317
rect 3760 3215 3794 3249
rect 3916 4099 3950 4133
rect 3916 4031 3950 4065
rect 3916 3963 3950 3997
rect 3916 3895 3950 3929
rect 3916 3827 3950 3861
rect 3916 3759 3950 3793
rect 3916 3691 3950 3725
rect 3916 3623 3950 3657
rect 3916 3555 3950 3589
rect 3916 3487 3950 3521
rect 3916 3419 3950 3453
rect 3916 3351 3950 3385
rect 3916 3283 3950 3317
rect 3916 3215 3950 3249
rect 4072 4099 4106 4133
rect 4072 4031 4106 4065
rect 4072 3963 4106 3997
rect 4072 3895 4106 3929
rect 4072 3827 4106 3861
rect 4072 3759 4106 3793
rect 4072 3691 4106 3725
rect 4072 3623 4106 3657
rect 4072 3555 4106 3589
rect 4072 3487 4106 3521
rect 4072 3419 4106 3453
rect 4072 3351 4106 3385
rect 4072 3283 4106 3317
rect 4072 3215 4106 3249
rect 4228 4099 4262 4133
rect 4228 4031 4262 4065
rect 4228 3963 4262 3997
rect 4228 3895 4262 3929
rect 4228 3827 4262 3861
rect 4228 3759 4262 3793
rect 4228 3691 4262 3725
rect 4228 3623 4262 3657
rect 4228 3555 4262 3589
rect 4228 3487 4262 3521
rect 4228 3419 4262 3453
rect 4228 3351 4262 3385
rect 4228 3283 4262 3317
rect 4228 3215 4262 3249
rect 4424 4149 4458 4183
rect 4424 4081 4458 4115
rect 4424 4013 4458 4047
rect 4424 3945 4458 3979
rect 4424 3877 4458 3911
rect 4424 3809 4458 3843
rect 4424 3741 4458 3775
rect 4424 3673 4458 3707
rect 4424 3605 4458 3639
rect 4424 3537 4458 3571
rect 4424 3469 4458 3503
rect 4424 3401 4458 3435
rect 4424 3333 4458 3367
rect 4424 3265 4458 3299
rect 4580 4149 4614 4183
rect 4580 4081 4614 4115
rect 4580 4013 4614 4047
rect 4580 3945 4614 3979
rect 4580 3877 4614 3911
rect 4580 3809 4614 3843
rect 4580 3741 4614 3775
rect 4580 3673 4614 3707
rect 4580 3605 4614 3639
rect 4580 3537 4614 3571
rect 4580 3469 4614 3503
rect 4580 3401 4614 3435
rect 4580 3333 4614 3367
rect 4580 3265 4614 3299
rect 4736 4149 4770 4183
rect 4736 4081 4770 4115
rect 4736 4013 4770 4047
rect 4736 3945 4770 3979
rect 4736 3877 4770 3911
rect 4736 3809 4770 3843
rect 4736 3741 4770 3775
rect 4736 3673 4770 3707
rect 4736 3605 4770 3639
rect 4736 3537 4770 3571
rect 4736 3469 4770 3503
rect 4736 3401 4770 3435
rect 4736 3333 4770 3367
rect 4736 3265 4770 3299
rect 4892 4149 4926 4183
rect 4892 4081 4926 4115
rect 4892 4013 4926 4047
rect 4892 3945 4926 3979
rect 4892 3877 4926 3911
rect 4892 3809 4926 3843
rect 4892 3741 4926 3775
rect 4892 3673 4926 3707
rect 4892 3605 4926 3639
rect 4892 3537 4926 3571
rect 4892 3469 4926 3503
rect 4892 3401 4926 3435
rect 4892 3333 4926 3367
rect 4892 3265 4926 3299
rect 5048 4149 5082 4183
rect 5048 4081 5082 4115
rect 5048 4013 5082 4047
rect 5048 3945 5082 3979
rect 5048 3877 5082 3911
rect 5048 3809 5082 3843
rect 5048 3741 5082 3775
rect 5048 3673 5082 3707
rect 5048 3605 5082 3639
rect 5048 3537 5082 3571
rect 5048 3469 5082 3503
rect 5048 3401 5082 3435
rect 5048 3333 5082 3367
rect 5048 3265 5082 3299
rect 5204 4149 5238 4183
rect 5204 4081 5238 4115
rect 5204 4013 5238 4047
rect 5204 3945 5238 3979
rect 5204 3877 5238 3911
rect 5204 3809 5238 3843
rect 5204 3741 5238 3775
rect 5204 3673 5238 3707
rect 5204 3605 5238 3639
rect 5204 3537 5238 3571
rect 5204 3469 5238 3503
rect 5204 3401 5238 3435
rect 5204 3333 5238 3367
rect 5204 3265 5238 3299
rect 5360 4149 5394 4183
rect 5360 4081 5394 4115
rect 5360 4013 5394 4047
rect 5360 3945 5394 3979
rect 5360 3877 5394 3911
rect 5360 3809 5394 3843
rect 5360 3741 5394 3775
rect 5360 3673 5394 3707
rect 5360 3605 5394 3639
rect 5360 3537 5394 3571
rect 5360 3469 5394 3503
rect 5360 3401 5394 3435
rect 5360 3333 5394 3367
rect 5360 3265 5394 3299
rect 5516 4149 5550 4183
rect 5516 4081 5550 4115
rect 5516 4013 5550 4047
rect 5516 3945 5550 3979
rect 5516 3877 5550 3911
rect 5516 3809 5550 3843
rect 5516 3741 5550 3775
rect 5516 3673 5550 3707
rect 5516 3605 5550 3639
rect 5516 3537 5550 3571
rect 5516 3469 5550 3503
rect 5516 3401 5550 3435
rect 5516 3333 5550 3367
rect 5516 3265 5550 3299
rect 9145 4272 9179 4306
rect 9145 4204 9179 4238
rect 5672 4149 5706 4183
rect 5672 4081 5706 4115
rect 5672 4013 5706 4047
rect 5672 3945 5706 3979
rect 5672 3877 5706 3911
rect 5672 3809 5706 3843
rect 5672 3741 5706 3775
rect 5672 3673 5706 3707
rect 5672 3605 5706 3639
rect 5672 3537 5706 3571
rect 5672 3469 5706 3503
rect 5672 3401 5706 3435
rect 5672 3333 5706 3367
rect 5672 3265 5706 3299
rect 5868 4099 5902 4133
rect 5868 4031 5902 4065
rect 5868 3963 5902 3997
rect 5868 3895 5902 3929
rect 5868 3827 5902 3861
rect 5868 3759 5902 3793
rect 5868 3691 5902 3725
rect 5868 3623 5902 3657
rect 5868 3555 5902 3589
rect 5868 3487 5902 3521
rect 5868 3419 5902 3453
rect 5868 3351 5902 3385
rect 5868 3283 5902 3317
rect 5868 3215 5902 3249
rect 6024 4099 6058 4133
rect 6024 4031 6058 4065
rect 6024 3963 6058 3997
rect 6024 3895 6058 3929
rect 6024 3827 6058 3861
rect 6024 3759 6058 3793
rect 6024 3691 6058 3725
rect 6024 3623 6058 3657
rect 6024 3555 6058 3589
rect 6024 3487 6058 3521
rect 6024 3419 6058 3453
rect 6024 3351 6058 3385
rect 6024 3283 6058 3317
rect 6024 3215 6058 3249
rect 6180 4099 6214 4133
rect 6180 4031 6214 4065
rect 6180 3963 6214 3997
rect 6180 3895 6214 3929
rect 6180 3827 6214 3861
rect 6180 3759 6214 3793
rect 6180 3691 6214 3725
rect 6180 3623 6214 3657
rect 6180 3555 6214 3589
rect 6180 3487 6214 3521
rect 6180 3419 6214 3453
rect 6180 3351 6214 3385
rect 6180 3283 6214 3317
rect 6180 3215 6214 3249
rect 6336 4099 6370 4133
rect 6336 4031 6370 4065
rect 6336 3963 6370 3997
rect 6336 3895 6370 3929
rect 6336 3827 6370 3861
rect 6336 3759 6370 3793
rect 6336 3691 6370 3725
rect 6336 3623 6370 3657
rect 6336 3555 6370 3589
rect 6336 3487 6370 3521
rect 6336 3419 6370 3453
rect 6336 3351 6370 3385
rect 6336 3283 6370 3317
rect 6336 3215 6370 3249
rect 6492 4099 6526 4133
rect 6492 4031 6526 4065
rect 6492 3963 6526 3997
rect 6492 3895 6526 3929
rect 6492 3827 6526 3861
rect 6492 3759 6526 3793
rect 6492 3691 6526 3725
rect 6492 3623 6526 3657
rect 6492 3555 6526 3589
rect 6492 3487 6526 3521
rect 6492 3419 6526 3453
rect 6492 3351 6526 3385
rect 6492 3283 6526 3317
rect 6492 3215 6526 3249
rect 6648 4099 6682 4133
rect 6648 4031 6682 4065
rect 6648 3963 6682 3997
rect 6648 3895 6682 3929
rect 6648 3827 6682 3861
rect 6648 3759 6682 3793
rect 6648 3691 6682 3725
rect 6648 3623 6682 3657
rect 6648 3555 6682 3589
rect 6648 3487 6682 3521
rect 6648 3419 6682 3453
rect 6648 3351 6682 3385
rect 6648 3283 6682 3317
rect 6648 3215 6682 3249
rect 6804 4099 6838 4133
rect 6804 4031 6838 4065
rect 6804 3963 6838 3997
rect 6804 3895 6838 3929
rect 6804 3827 6838 3861
rect 6804 3759 6838 3793
rect 6804 3691 6838 3725
rect 6804 3623 6838 3657
rect 6804 3555 6838 3589
rect 6804 3487 6838 3521
rect 6804 3419 6838 3453
rect 6804 3351 6838 3385
rect 6804 3283 6838 3317
rect 6804 3215 6838 3249
rect 6960 4099 6994 4133
rect 6960 4031 6994 4065
rect 6960 3963 6994 3997
rect 6960 3895 6994 3929
rect 6960 3827 6994 3861
rect 6960 3759 6994 3793
rect 6960 3691 6994 3725
rect 6960 3623 6994 3657
rect 6960 3555 6994 3589
rect 6960 3487 6994 3521
rect 6960 3419 6994 3453
rect 6960 3351 6994 3385
rect 6960 3283 6994 3317
rect 6960 3215 6994 3249
rect 7116 4099 7150 4133
rect 7116 4031 7150 4065
rect 7116 3963 7150 3997
rect 7116 3895 7150 3929
rect 7116 3827 7150 3861
rect 7116 3759 7150 3793
rect 7116 3691 7150 3725
rect 7116 3623 7150 3657
rect 7116 3555 7150 3589
rect 7116 3487 7150 3521
rect 7116 3419 7150 3453
rect 7116 3351 7150 3385
rect 7116 3283 7150 3317
rect 7116 3215 7150 3249
rect 7272 4099 7306 4133
rect 7272 4031 7306 4065
rect 7272 3963 7306 3997
rect 7272 3895 7306 3929
rect 7272 3827 7306 3861
rect 7272 3759 7306 3793
rect 7272 3691 7306 3725
rect 7272 3623 7306 3657
rect 7272 3555 7306 3589
rect 7272 3487 7306 3521
rect 7272 3419 7306 3453
rect 7272 3351 7306 3385
rect 7272 3283 7306 3317
rect 7272 3215 7306 3249
rect 7468 4091 7502 4125
rect 7468 4023 7502 4057
rect 7468 3955 7502 3989
rect 7468 3887 7502 3921
rect 7468 3819 7502 3853
rect 7468 3751 7502 3785
rect 7468 3683 7502 3717
rect 7468 3615 7502 3649
rect 7908 4091 7942 4125
rect 7908 4023 7942 4057
rect 8038 4067 8072 4101
rect 7908 3955 7942 3989
rect 7908 3887 7942 3921
rect 7908 3819 7942 3853
rect 7908 3751 7942 3785
rect 7908 3683 7942 3717
rect 7908 3615 7942 3649
rect 7468 3356 7502 3390
rect 7468 3288 7502 3322
rect 7468 3220 7502 3254
rect 7624 3356 7658 3390
rect 7624 3288 7658 3322
rect 7624 3220 7658 3254
rect 7780 3356 7814 3390
rect 7780 3288 7814 3322
rect 7780 3220 7814 3254
rect 8038 3211 8072 3245
rect 9145 4136 9179 4170
rect 9145 4068 9179 4102
rect 9145 4000 9179 4034
rect 9145 3932 9179 3966
rect 9145 3864 9179 3898
rect 9145 3796 9179 3830
rect 9301 4272 9335 4306
rect 9301 4204 9335 4238
rect 9301 4136 9335 4170
rect 9301 4068 9335 4102
rect 9301 4000 9335 4034
rect 9301 3932 9335 3966
rect 9301 3864 9335 3898
rect 9301 3796 9335 3830
rect 9457 4272 9491 4306
rect 9457 4204 9491 4238
rect 9457 4136 9491 4170
rect 9457 4068 9491 4102
rect 9457 4000 9491 4034
rect 9457 3932 9491 3966
rect 9457 3864 9491 3898
rect 9457 3796 9491 3830
rect 9613 4272 9647 4306
rect 9613 4204 9647 4238
rect 9613 4136 9647 4170
rect 9613 4068 9647 4102
rect 9613 4000 9647 4034
rect 9613 3932 9647 3966
rect 9613 3864 9647 3898
rect 9613 3796 9647 3830
rect 9737 4272 9771 4306
rect 9737 4204 9771 4238
rect 9737 4136 9771 4170
rect 9737 4068 9771 4102
rect 9737 4000 9771 4034
rect 9737 3932 9771 3966
rect 9737 3864 9771 3898
rect 9737 3796 9771 3830
rect 9893 4272 9927 4306
rect 9893 4204 9927 4238
rect 9893 4136 9927 4170
rect 9893 4068 9927 4102
rect 9893 4000 9927 4034
rect 9893 3932 9927 3966
rect 9893 3864 9927 3898
rect 9893 3796 9927 3830
rect 10049 4272 10083 4306
rect 10049 4204 10083 4238
rect 10049 4136 10083 4170
rect 10049 4068 10083 4102
rect 10049 4000 10083 4034
rect 10049 3932 10083 3966
rect 10049 3864 10083 3898
rect 10049 3796 10083 3830
rect 10205 4272 10239 4306
rect 10205 4204 10239 4238
rect 10205 4136 10239 4170
rect 10205 4068 10239 4102
rect 10205 4000 10239 4034
rect 10205 3932 10239 3966
rect 10205 3864 10239 3898
rect 10205 3796 10239 3830
rect 10361 4272 10395 4306
rect 10361 4204 10395 4238
rect 10361 4136 10395 4170
rect 10361 4068 10395 4102
rect 10361 4000 10395 4034
rect 10361 3932 10395 3966
rect 10361 3864 10395 3898
rect 10361 3796 10395 3830
rect 10485 4272 10519 4306
rect 10485 4204 10519 4238
rect 10485 4136 10519 4170
rect 10485 4068 10519 4102
rect 10485 4000 10519 4034
rect 10485 3932 10519 3966
rect 10485 3864 10519 3898
rect 10485 3796 10519 3830
rect 10641 4272 10675 4306
rect 10641 4204 10675 4238
rect 10641 4136 10675 4170
rect 10641 4068 10675 4102
rect 10641 4000 10675 4034
rect 10641 3932 10675 3966
rect 10641 3864 10675 3898
rect 10641 3796 10675 3830
rect 10797 4272 10831 4306
rect 12149 4247 12183 4281
rect 10797 4204 10831 4238
rect 10797 4136 10831 4170
rect 11017 4167 11051 4201
rect 11873 4167 11907 4201
rect 10797 4068 10831 4102
rect 10797 4000 10831 4034
rect 10797 3932 10831 3966
rect 11017 3953 11051 3987
rect 11873 3953 11907 3987
rect 12149 3991 12183 4025
rect 10797 3864 10831 3898
rect 10797 3796 10831 3830
rect 11017 3785 11051 3819
rect 11873 3785 11907 3819
rect 12149 3735 12183 3769
rect 12149 3611 12183 3645
rect -314 2987 -280 3021
rect 1692 3037 1726 3071
rect 3348 3037 3382 3071
rect -314 2919 -280 2953
rect 9756 3426 9790 3460
rect 9756 3358 9790 3392
rect 9756 3290 9790 3324
rect 9756 3222 9790 3256
rect 9756 3154 9790 3188
rect 9756 3086 9790 3120
rect 9756 3018 9790 3052
rect 9756 2950 9790 2984
rect 10136 3426 10170 3460
rect 10136 3358 10170 3392
rect 10136 3290 10170 3324
rect 10136 3222 10170 3256
rect 10136 3154 10170 3188
rect 10136 3086 10170 3120
rect 10136 3018 10170 3052
rect 10136 2950 10170 2984
rect 11017 3533 11051 3567
rect 11873 3533 11907 3567
rect 10326 3426 10360 3460
rect 10326 3358 10360 3392
rect 10326 3290 10360 3324
rect 10326 3222 10360 3256
rect 10326 3154 10360 3188
rect 10326 3086 10360 3120
rect 10326 3018 10360 3052
rect 10326 2950 10360 2984
rect 11017 3317 11051 3351
rect 11873 3317 11907 3351
rect 12149 3355 12183 3389
rect -453 2617 -419 2651
rect -453 2549 -419 2583
rect -453 2481 -419 2515
rect -277 2617 -243 2651
rect -277 2549 -243 2583
rect -277 2481 -243 2515
rect -101 2617 -67 2651
rect -101 2549 -67 2583
rect -101 2481 -67 2515
rect 75 2617 109 2651
rect 75 2549 109 2583
rect 75 2481 109 2515
rect -453 2355 -419 2389
rect -453 2287 -419 2321
rect -453 2219 -419 2253
rect -277 2355 -243 2389
rect -277 2287 -243 2321
rect -277 2219 -243 2253
rect -101 2355 -67 2389
rect -101 2287 -67 2321
rect -101 2219 -67 2253
rect 75 2355 109 2389
rect 75 2287 109 2321
rect 75 2219 109 2253
rect 7422 1440 7456 1474
rect 7422 1372 7456 1406
rect 7422 1304 7456 1338
rect 7422 1236 7456 1270
rect 7422 1168 7456 1202
rect 7422 1100 7456 1134
rect 7422 1032 7456 1066
rect 7422 964 7456 998
rect 7422 896 7456 930
rect 7422 828 7456 862
rect 7422 760 7456 794
rect 7422 692 7456 726
rect 7422 624 7456 658
rect 7422 556 7456 590
rect 7598 1440 7632 1474
rect 7598 1372 7632 1406
rect 7598 1304 7632 1338
rect 7598 1236 7632 1270
rect 7598 1168 7632 1202
rect 7598 1100 7632 1134
rect 7598 1032 7632 1066
rect 7598 964 7632 998
rect 7598 896 7632 930
rect 7598 828 7632 862
rect 7598 760 7632 794
rect 7598 692 7632 726
rect 7598 624 7632 658
rect 7598 556 7632 590
rect 7774 1440 7808 1474
rect 7774 1372 7808 1406
rect 7774 1304 7808 1338
rect 7774 1236 7808 1270
rect 7774 1168 7808 1202
rect 7774 1100 7808 1134
rect 7774 1032 7808 1066
rect 7774 964 7808 998
rect 7774 896 7808 930
rect 7774 828 7808 862
rect 7774 760 7808 794
rect 7774 692 7808 726
rect 7774 624 7808 658
rect 7774 556 7808 590
rect 7950 1440 7984 1474
rect 7950 1372 7984 1406
rect 7950 1304 7984 1338
rect 7950 1236 7984 1270
rect 7950 1168 7984 1202
rect 7950 1100 7984 1134
rect 7950 1032 7984 1066
rect 7950 964 7984 998
rect 8884 1432 8918 1466
rect 8884 1364 8918 1398
rect 8884 1296 8918 1330
rect 8884 1228 8918 1262
rect 8884 1160 8918 1194
rect 8884 1092 8918 1126
rect 8884 1024 8918 1058
rect 8884 956 8918 990
rect 9040 1432 9074 1466
rect 9040 1364 9074 1398
rect 9040 1296 9074 1330
rect 9040 1228 9074 1262
rect 9040 1160 9074 1194
rect 9040 1092 9074 1126
rect 9040 1024 9074 1058
rect 9040 956 9074 990
rect 9196 1432 9230 1466
rect 9196 1364 9230 1398
rect 9196 1296 9230 1330
rect 9196 1228 9230 1262
rect 9196 1160 9230 1194
rect 9196 1092 9230 1126
rect 9196 1024 9230 1058
rect 9196 956 9230 990
rect 9352 1432 9386 1466
rect 9352 1364 9386 1398
rect 9352 1296 9386 1330
rect 9352 1228 9386 1262
rect 9352 1160 9386 1194
rect 9352 1092 9386 1126
rect 9352 1024 9386 1058
rect 9352 956 9386 990
rect 9508 1432 9542 1466
rect 9508 1364 9542 1398
rect 9508 1296 9542 1330
rect 9508 1228 9542 1262
rect 9508 1160 9542 1194
rect 9508 1092 9542 1126
rect 9508 1024 9542 1058
rect 9508 956 9542 990
rect 9756 1432 9790 1466
rect 9756 1364 9790 1398
rect 9756 1296 9790 1330
rect 9756 1228 9790 1262
rect 9756 1160 9790 1194
rect 9756 1092 9790 1126
rect 9756 1024 9790 1058
rect 9756 956 9790 990
rect 9912 1432 9946 1466
rect 9912 1364 9946 1398
rect 9912 1296 9946 1330
rect 9912 1228 9946 1262
rect 9912 1160 9946 1194
rect 9912 1092 9946 1126
rect 9912 1024 9946 1058
rect 9912 956 9946 990
rect 10068 1432 10102 1466
rect 10068 1364 10102 1398
rect 10068 1296 10102 1330
rect 10068 1228 10102 1262
rect 10068 1160 10102 1194
rect 10068 1092 10102 1126
rect 10068 1024 10102 1058
rect 10068 956 10102 990
rect 10224 1432 10258 1466
rect 10224 1364 10258 1398
rect 10224 1296 10258 1330
rect 10224 1228 10258 1262
rect 10224 1160 10258 1194
rect 10224 1092 10258 1126
rect 10224 1024 10258 1058
rect 10224 956 10258 990
rect 10380 1432 10414 1466
rect 10380 1364 10414 1398
rect 10380 1296 10414 1330
rect 10380 1228 10414 1262
rect 10380 1160 10414 1194
rect 10572 1409 10606 1443
rect 10572 1341 10606 1375
rect 10572 1273 10606 1307
rect 10572 1205 10606 1239
rect 10728 1409 10762 1443
rect 10728 1341 10762 1375
rect 10728 1273 10762 1307
rect 10728 1205 10762 1239
rect 10884 1409 10918 1443
rect 10884 1341 10918 1375
rect 10884 1273 10918 1307
rect 10884 1205 10918 1239
rect 11040 1409 11074 1443
rect 11040 1341 11074 1375
rect 11040 1273 11074 1307
rect 11040 1205 11074 1239
rect 11196 1409 11230 1443
rect 11196 1341 11230 1375
rect 11196 1273 11230 1307
rect 11369 1303 11403 1337
rect 12225 1303 12259 1337
rect 11196 1205 11230 1239
rect 10380 1092 10414 1126
rect 10380 1024 10414 1058
rect 10380 956 10414 990
rect 7950 896 7984 930
rect 7950 828 7984 862
rect 10857 881 10891 915
rect 11313 881 11347 915
rect 11769 881 11803 915
rect 12225 881 12259 915
rect 7950 760 7984 794
rect 7950 692 7984 726
rect 7950 624 7984 658
rect 7950 556 7984 590
rect 10406 597 10440 631
rect 10406 529 10440 563
rect 10406 461 10440 495
rect 10562 597 10596 631
rect 10562 529 10596 563
rect 10562 461 10596 495
rect 10718 597 10752 631
rect 10718 529 10752 563
rect 10908 597 10942 631
rect 11064 597 11098 631
rect 11220 597 11254 631
rect 11344 597 11378 631
rect 11500 597 11534 631
rect 11656 597 11690 631
rect 10718 461 10752 495
<< psubdiff >>
rect -644 4091 -574 4115
rect -644 4057 -615 4091
rect -581 4057 -574 4091
rect -644 4002 -574 4057
rect -644 3968 -615 4002
rect -581 3968 -574 4002
rect -644 3912 -574 3968
rect -644 3878 -615 3912
rect -581 3878 -574 3912
rect -644 3822 -574 3878
rect -644 3788 -615 3822
rect -581 3788 -574 3822
rect -644 3764 -574 3788
<< mvpsubdiff >>
rect -574 3764 -552 4115
rect 8751 4119 8985 4143
rect 8785 4085 8851 4119
rect 8885 4085 8951 4119
rect 8751 4046 8985 4085
rect 8785 4012 8851 4046
rect 8885 4012 8951 4046
rect 8751 3973 8985 4012
rect 8785 3939 8851 3973
rect 8885 3939 8951 3973
rect 8751 3900 8985 3939
rect 8785 3866 8851 3900
rect 8885 3866 8951 3900
rect 8751 3827 8985 3866
rect 8785 3793 8851 3827
rect 8885 3793 8951 3827
rect 8751 3754 8985 3793
rect 8785 3720 8851 3754
rect 8885 3720 8951 3754
rect 8751 3681 8985 3720
rect 8785 3647 8851 3681
rect 8885 3647 8951 3681
rect 8751 3607 8985 3647
rect 8785 3573 8851 3607
rect 8885 3573 8951 3607
rect 8751 3533 8985 3573
rect 8785 3499 8851 3533
rect 8885 3499 8951 3533
rect 8751 3459 8985 3499
rect 8785 3425 8851 3459
rect 8885 3425 8951 3459
rect 8751 3385 8985 3425
rect 8785 3351 8851 3385
rect 8885 3351 8951 3385
rect 8751 3311 8985 3351
rect 8785 3277 8851 3311
rect 8885 3277 8951 3311
rect 8751 3253 8985 3277
rect 10744 3073 10778 3097
rect 10744 3005 10778 3039
rect -433 1745 -409 1779
rect -375 1745 -331 1779
rect -297 1745 -253 1779
rect -219 1745 -175 1779
rect -141 1745 -97 1779
rect -63 1745 -20 1779
rect 14 1745 57 1779
rect 91 1745 115 1779
rect 10744 2937 10778 2971
rect 10744 2869 10778 2903
rect 10744 2801 10778 2835
rect 10744 2732 10778 2767
rect 10744 2663 10778 2698
rect 10744 2594 10778 2629
rect 10744 2536 10778 2560
rect 9445 2284 9547 2308
rect 9479 2250 9513 2284
rect 9445 2210 9547 2250
rect 9479 2176 9513 2210
rect 9445 2136 9547 2176
rect 9479 2102 9513 2136
rect 9445 2062 9547 2102
rect 9479 2028 9513 2062
rect 9445 1988 9547 2028
rect 9479 1954 9513 1988
rect 9445 1914 9547 1954
rect 9479 1880 9513 1914
rect 9445 1840 9547 1880
rect 9479 1806 9513 1840
rect 9445 1766 9547 1806
rect 9479 1732 9513 1766
rect 9445 1708 9547 1732
rect 10484 2255 10522 2308
rect 10484 2221 10486 2255
rect 10520 2221 10522 2255
rect 10484 2187 10522 2221
rect 10484 2153 10486 2187
rect 10520 2153 10522 2187
rect 10484 2119 10522 2153
rect 10484 2085 10486 2119
rect 10520 2085 10522 2119
rect 10484 2051 10522 2085
rect 10484 2017 10486 2051
rect 10520 2017 10522 2051
rect 10484 1983 10522 2017
rect 10484 1949 10486 1983
rect 10520 1949 10522 1983
rect 10484 1915 10522 1949
rect 10484 1881 10486 1915
rect 10520 1881 10522 1915
rect 10484 1847 10522 1881
rect 10484 1813 10486 1847
rect 10520 1813 10522 1847
rect 10484 1765 10522 1813
rect 12133 2312 12167 2336
rect 12133 2237 12167 2278
rect 12133 2162 12167 2203
rect 12133 2088 12167 2128
rect 12133 2014 12167 2054
rect 12133 1940 12167 1980
rect 12133 1866 12167 1906
rect 12133 1808 12167 1832
<< mvnsubdiff >>
rect -502 4907 -478 4941
rect -444 4907 -406 4941
rect -372 4907 -334 4941
rect -300 4907 -262 4941
rect -228 4907 -190 4941
rect -156 4907 -119 4941
rect -85 4907 -48 4941
rect -14 4907 23 4941
rect 57 4907 94 4941
rect 128 4907 152 4941
rect 10793 4580 12400 4642
rect 10793 4546 10909 4580
rect 10943 4546 10980 4580
rect 11014 4546 11051 4580
rect 11085 4546 11122 4580
rect 11156 4546 11193 4580
rect 11227 4546 11264 4580
rect 11298 4546 11335 4580
rect 11369 4546 11406 4580
rect 11440 4546 11477 4580
rect 11511 4546 11548 4580
rect 11582 4546 11619 4580
rect 11653 4546 11690 4580
rect 11724 4546 11761 4580
rect 11795 4546 11832 4580
rect 11866 4546 11903 4580
rect 11937 4546 11974 4580
rect 12008 4546 12045 4580
rect 12079 4546 12116 4580
rect 12150 4546 12187 4580
rect 12221 4546 12258 4580
rect 12292 4546 12329 4580
rect 12363 4546 12400 4580
rect 10793 4530 12400 4546
rect 10793 4506 10893 4530
rect 10793 4493 10839 4506
rect 271 4472 10839 4493
rect 10873 4472 10893 4506
rect 271 4460 10893 4472
rect 271 4426 409 4460
rect 443 4426 477 4460
rect 511 4426 545 4460
rect 579 4426 613 4460
rect 647 4426 681 4460
rect 715 4426 749 4460
rect 783 4426 817 4460
rect 851 4426 885 4460
rect 919 4426 953 4460
rect 987 4426 1021 4460
rect 1055 4426 1089 4460
rect 1123 4426 1157 4460
rect 1191 4426 1225 4460
rect 1259 4426 1293 4460
rect 1327 4426 1361 4460
rect 1395 4426 1429 4460
rect 1463 4426 1497 4460
rect 1531 4426 1565 4460
rect 1599 4426 1633 4460
rect 1667 4426 1701 4460
rect 1735 4426 1769 4460
rect 1803 4426 1837 4460
rect 1871 4426 1905 4460
rect 1939 4426 1973 4460
rect 2007 4426 2041 4460
rect 2075 4426 2109 4460
rect 2143 4426 2177 4460
rect 2211 4426 2245 4460
rect 2279 4426 2313 4460
rect 2347 4426 2381 4460
rect 2415 4426 2449 4460
rect 2483 4426 2517 4460
rect 2551 4426 2585 4460
rect 2619 4426 2653 4460
rect 2687 4426 2721 4460
rect 2755 4426 2789 4460
rect 2823 4426 2857 4460
rect 2891 4426 2925 4460
rect 2959 4426 2993 4460
rect 3027 4426 3061 4460
rect 3095 4426 3129 4460
rect 3163 4426 3197 4460
rect 3231 4426 3265 4460
rect 3299 4426 3333 4460
rect 3367 4426 3401 4460
rect 3435 4426 3469 4460
rect 3503 4426 3537 4460
rect 3571 4426 3605 4460
rect 3639 4426 3673 4460
rect 3707 4426 3741 4460
rect 3775 4426 3809 4460
rect 3843 4426 3877 4460
rect 3911 4426 3945 4460
rect 3979 4426 4013 4460
rect 4047 4426 4081 4460
rect 4115 4426 4149 4460
rect 4183 4426 4217 4460
rect 4251 4426 4285 4460
rect 4319 4426 4353 4460
rect 4387 4426 4421 4460
rect 4455 4426 4489 4460
rect 4523 4426 4557 4460
rect 4591 4426 4625 4460
rect 4659 4426 4693 4460
rect 4727 4426 4761 4460
rect 4795 4426 4829 4460
rect 4863 4426 4897 4460
rect 4931 4426 4965 4460
rect 4999 4426 5033 4460
rect 5067 4426 5101 4460
rect 5135 4426 5169 4460
rect 5203 4426 5237 4460
rect 5271 4426 5305 4460
rect 5339 4426 5373 4460
rect 5407 4426 5441 4460
rect 5475 4426 5509 4460
rect 5543 4426 5577 4460
rect 5611 4426 5645 4460
rect 5679 4426 5713 4460
rect 5747 4426 5781 4460
rect 5815 4426 5849 4460
rect 5883 4426 5917 4460
rect 5951 4426 5985 4460
rect 6019 4426 6053 4460
rect 6087 4426 6121 4460
rect 6155 4426 6189 4460
rect 6223 4426 6257 4460
rect 6291 4426 6325 4460
rect 6359 4426 6393 4460
rect 6427 4426 6461 4460
rect 6495 4426 6529 4460
rect 6563 4426 6597 4460
rect 6631 4426 6665 4460
rect 6699 4426 6733 4460
rect 6767 4426 6801 4460
rect 6835 4426 6869 4460
rect 6903 4426 6937 4460
rect 6971 4426 7005 4460
rect 7039 4426 7073 4460
rect 7107 4426 7141 4460
rect 7175 4426 7209 4460
rect 7243 4426 7277 4460
rect 7311 4426 7345 4460
rect 7379 4426 7413 4460
rect 7447 4426 7481 4460
rect 7515 4426 7549 4460
rect 7583 4426 7617 4460
rect 7651 4426 7685 4460
rect 7719 4426 7753 4460
rect 7787 4426 7821 4460
rect 7855 4426 7889 4460
rect 7923 4426 7957 4460
rect 7991 4426 8025 4460
rect 8059 4426 8093 4460
rect 8127 4426 8161 4460
rect 8195 4426 8229 4460
rect 8263 4426 8297 4460
rect 8331 4426 8365 4460
rect 8399 4426 8433 4460
rect 8467 4426 8501 4460
rect 8535 4426 8569 4460
rect 8603 4426 8637 4460
rect 8671 4426 8705 4460
rect 8739 4426 8773 4460
rect 8807 4426 8841 4460
rect 8875 4426 8909 4460
rect 8943 4426 8977 4460
rect 9011 4426 9045 4460
rect 9079 4426 9113 4460
rect 9147 4426 9181 4460
rect 9215 4426 9249 4460
rect 9283 4426 9317 4460
rect 9351 4426 9385 4460
rect 9419 4426 9453 4460
rect 9487 4426 9521 4460
rect 9555 4426 9589 4460
rect 9623 4426 9657 4460
rect 9691 4426 9725 4460
rect 9759 4426 9793 4460
rect 9827 4426 9861 4460
rect 9895 4426 9929 4460
rect 9963 4426 9997 4460
rect 10031 4426 10065 4460
rect 10099 4426 10133 4460
rect 10167 4426 10201 4460
rect 10235 4426 10269 4460
rect 10303 4426 10337 4460
rect 10371 4426 10405 4460
rect 10439 4426 10473 4460
rect 10507 4426 10541 4460
rect 10575 4426 10609 4460
rect 10643 4431 10893 4460
rect 10643 4426 10760 4431
rect 271 4409 10760 4426
rect 305 4397 10760 4409
rect 10794 4397 10893 4431
rect 305 4393 10893 4397
rect 12366 4496 12400 4530
rect 12366 4428 12400 4462
rect 271 4341 305 4375
rect 12366 4360 12400 4394
rect 271 4273 305 4307
rect 271 4205 305 4239
rect 271 4137 305 4171
rect 271 4069 305 4103
rect 271 4001 305 4035
rect 271 3933 305 3967
rect 271 3865 305 3899
rect 271 3797 305 3831
rect 271 3729 305 3763
rect 271 3661 305 3695
rect 271 3593 305 3627
rect 271 3525 305 3559
rect 271 3457 305 3491
rect 271 3389 305 3423
rect 271 3321 305 3355
rect 271 3253 305 3287
rect 271 3185 305 3219
rect 1014 4164 1052 4203
rect 1014 4130 1016 4164
rect 1050 4130 1052 4164
rect 1014 4096 1052 4130
rect 1014 4062 1016 4096
rect 1050 4062 1052 4096
rect 1014 4028 1052 4062
rect 1014 3994 1016 4028
rect 1050 3994 1052 4028
rect 1014 3960 1052 3994
rect 1014 3926 1016 3960
rect 1050 3926 1052 3960
rect 1014 3892 1052 3926
rect 1014 3858 1016 3892
rect 1050 3858 1052 3892
rect 1014 3824 1052 3858
rect 1014 3790 1016 3824
rect 1050 3790 1052 3824
rect 1014 3756 1052 3790
rect 1014 3722 1016 3756
rect 1050 3722 1052 3756
rect 1014 3688 1052 3722
rect 1014 3654 1016 3688
rect 1050 3654 1052 3688
rect 1014 3620 1052 3654
rect 1014 3586 1016 3620
rect 1050 3586 1052 3620
rect 1014 3552 1052 3586
rect 1014 3518 1016 3552
rect 1050 3518 1052 3552
rect 1014 3484 1052 3518
rect 1014 3450 1016 3484
rect 1050 3450 1052 3484
rect 1014 3416 1052 3450
rect 1014 3382 1016 3416
rect 1050 3382 1052 3416
rect 1014 3348 1052 3382
rect 1014 3314 1016 3348
rect 1050 3314 1052 3348
rect 1014 3280 1052 3314
rect 1014 3246 1016 3280
rect 1050 3246 1052 3280
rect 1014 3203 1052 3246
rect 2880 4164 2918 4203
rect 2880 4130 2882 4164
rect 2916 4130 2918 4164
rect 2880 4096 2918 4130
rect 2880 4062 2882 4096
rect 2916 4062 2918 4096
rect 2880 4028 2918 4062
rect 2880 3994 2882 4028
rect 2916 3994 2918 4028
rect 2880 3960 2918 3994
rect 2880 3926 2882 3960
rect 2916 3926 2918 3960
rect 2880 3892 2918 3926
rect 2880 3858 2882 3892
rect 2916 3858 2918 3892
rect 2880 3824 2918 3858
rect 2880 3790 2882 3824
rect 2916 3790 2918 3824
rect 2880 3756 2918 3790
rect 2880 3722 2882 3756
rect 2916 3722 2918 3756
rect 2880 3688 2918 3722
rect 2880 3654 2882 3688
rect 2916 3654 2918 3688
rect 2880 3620 2918 3654
rect 2880 3586 2882 3620
rect 2916 3586 2918 3620
rect 2880 3552 2918 3586
rect 2880 3518 2882 3552
rect 2916 3518 2918 3552
rect 2880 3484 2918 3518
rect 2880 3450 2882 3484
rect 2916 3450 2918 3484
rect 2880 3416 2918 3450
rect 2880 3382 2882 3416
rect 2916 3382 2918 3416
rect 2880 3348 2918 3382
rect 2880 3314 2882 3348
rect 2916 3314 2918 3348
rect 2880 3280 2918 3314
rect 2880 3246 2882 3280
rect 2916 3246 2918 3280
rect 2880 3203 2918 3246
rect 4324 4164 4362 4203
rect 4324 4130 4326 4164
rect 4360 4130 4362 4164
rect 4324 4096 4362 4130
rect 4324 4062 4326 4096
rect 4360 4062 4362 4096
rect 4324 4028 4362 4062
rect 4324 3994 4326 4028
rect 4360 3994 4362 4028
rect 4324 3960 4362 3994
rect 4324 3926 4326 3960
rect 4360 3926 4362 3960
rect 4324 3892 4362 3926
rect 4324 3858 4326 3892
rect 4360 3858 4362 3892
rect 4324 3824 4362 3858
rect 4324 3790 4326 3824
rect 4360 3790 4362 3824
rect 4324 3756 4362 3790
rect 4324 3722 4326 3756
rect 4360 3722 4362 3756
rect 4324 3688 4362 3722
rect 4324 3654 4326 3688
rect 4360 3654 4362 3688
rect 4324 3620 4362 3654
rect 4324 3586 4326 3620
rect 4360 3586 4362 3620
rect 4324 3552 4362 3586
rect 4324 3518 4326 3552
rect 4360 3518 4362 3552
rect 4324 3484 4362 3518
rect 4324 3450 4326 3484
rect 4360 3450 4362 3484
rect 4324 3416 4362 3450
rect 4324 3382 4326 3416
rect 4360 3382 4362 3416
rect 4324 3348 4362 3382
rect 4324 3314 4326 3348
rect 4360 3314 4362 3348
rect 4324 3280 4362 3314
rect 4324 3246 4326 3280
rect 4360 3246 4362 3280
rect 5768 4164 5806 4203
rect 5768 4130 5770 4164
rect 5804 4130 5806 4164
rect 5768 4096 5806 4130
rect 5768 4062 5770 4096
rect 5804 4062 5806 4096
rect 5768 4028 5806 4062
rect 5768 3994 5770 4028
rect 5804 3994 5806 4028
rect 5768 3960 5806 3994
rect 5768 3926 5770 3960
rect 5804 3926 5806 3960
rect 5768 3892 5806 3926
rect 5768 3858 5770 3892
rect 5804 3858 5806 3892
rect 5768 3824 5806 3858
rect 5768 3790 5770 3824
rect 5804 3790 5806 3824
rect 5768 3756 5806 3790
rect 5768 3722 5770 3756
rect 5804 3722 5806 3756
rect 5768 3688 5806 3722
rect 5768 3654 5770 3688
rect 5804 3654 5806 3688
rect 5768 3620 5806 3654
rect 5768 3586 5770 3620
rect 5804 3586 5806 3620
rect 5768 3552 5806 3586
rect 5768 3518 5770 3552
rect 5804 3518 5806 3552
rect 5768 3484 5806 3518
rect 5768 3450 5770 3484
rect 5804 3450 5806 3484
rect 5768 3416 5806 3450
rect 5768 3382 5770 3416
rect 5804 3382 5806 3416
rect 5768 3348 5806 3382
rect 5768 3314 5770 3348
rect 5804 3314 5806 3348
rect 5768 3280 5806 3314
rect 4324 3203 4362 3246
rect 5768 3246 5770 3280
rect 5804 3246 5806 3280
rect 5768 3203 5806 3246
rect 7368 4164 7406 4203
rect 7368 4130 7370 4164
rect 7404 4130 7406 4164
rect 7368 4096 7406 4130
rect 7368 4062 7370 4096
rect 7404 4062 7406 4096
rect 7368 4028 7406 4062
rect 7368 3994 7370 4028
rect 7404 3994 7406 4028
rect 7368 3960 7406 3994
rect 7368 3926 7370 3960
rect 7404 3926 7406 3960
rect 7368 3892 7406 3926
rect 7368 3858 7370 3892
rect 7404 3858 7406 3892
rect 7368 3824 7406 3858
rect 7368 3790 7370 3824
rect 7404 3790 7406 3824
rect 7368 3756 7406 3790
rect 7368 3722 7370 3756
rect 7404 3722 7406 3756
rect 7368 3688 7406 3722
rect 7368 3654 7370 3688
rect 7404 3654 7406 3688
rect 7368 3620 7406 3654
rect 7368 3586 7370 3620
rect 7404 3586 7406 3620
rect 8164 4164 8202 4203
rect 8164 4130 8166 4164
rect 8200 4130 8202 4164
rect 8164 4096 8202 4130
rect 8164 4062 8166 4096
rect 8200 4062 8202 4096
rect 7368 3552 7406 3586
rect 7368 3518 7370 3552
rect 7404 3518 7406 3552
rect 7368 3484 7406 3518
rect 7368 3450 7370 3484
rect 7404 3450 7406 3484
rect 7368 3416 7406 3450
rect 7368 3382 7370 3416
rect 7404 3382 7406 3416
rect 7368 3348 7406 3382
rect 7368 3314 7370 3348
rect 7404 3314 7406 3348
rect 7368 3280 7406 3314
rect 7368 3246 7370 3280
rect 7404 3246 7406 3280
rect 7368 3203 7406 3246
rect 8164 4028 8202 4062
rect 8164 3994 8166 4028
rect 8200 3994 8202 4028
rect 8164 3960 8202 3994
rect 8164 3926 8166 3960
rect 8200 3926 8202 3960
rect 8164 3892 8202 3926
rect 8164 3858 8166 3892
rect 8200 3858 8202 3892
rect 8164 3824 8202 3858
rect 8164 3790 8166 3824
rect 8200 3790 8202 3824
rect 8164 3756 8202 3790
rect 8164 3722 8166 3756
rect 8200 3722 8202 3756
rect 8164 3688 8202 3722
rect 8164 3654 8166 3688
rect 8200 3654 8202 3688
rect 8164 3620 8202 3654
rect 8164 3586 8166 3620
rect 8200 3586 8202 3620
rect 8164 3552 8202 3586
rect 8164 3518 8166 3552
rect 8200 3518 8202 3552
rect 8164 3484 8202 3518
rect 8164 3450 8166 3484
rect 8200 3450 8202 3484
rect 8164 3416 8202 3450
rect 8164 3382 8166 3416
rect 8200 3382 8202 3416
rect 8164 3348 8202 3382
rect 8164 3314 8166 3348
rect 8200 3314 8202 3348
rect 8164 3280 8202 3314
rect 271 3117 305 3151
rect 8164 3246 8166 3280
rect 8200 3246 8202 3280
rect 12366 4292 12400 4326
rect 12366 4224 12400 4258
rect 12366 4156 12400 4190
rect 12366 4088 12400 4122
rect 12366 4020 12400 4054
rect 12366 3952 12400 3986
rect 12366 3884 12400 3918
rect 12366 3816 12400 3850
rect 12366 3748 12400 3782
rect 12366 3680 12400 3714
rect 8164 3203 8202 3246
rect 9443 3513 9509 3537
rect 9443 3479 9459 3513
rect 9493 3479 9509 3513
rect 9443 3412 9509 3479
rect 9443 3378 9459 3412
rect 9493 3378 9509 3412
rect 9443 3311 9509 3378
rect 9443 3277 9459 3311
rect 9493 3277 9509 3311
rect 9443 3253 9509 3277
rect 9640 3514 9674 3538
rect 9640 3440 9674 3480
rect 9640 3366 9674 3406
rect 9640 3292 9674 3332
rect 9640 3218 9674 3258
rect 9640 3144 9674 3184
rect 271 3049 305 3083
rect 3464 3067 4752 3075
rect 3464 3033 3488 3067
rect 3522 3033 3559 3067
rect 3593 3033 3630 3067
rect 3664 3033 3701 3067
rect 3735 3033 3772 3067
rect 3806 3033 3843 3067
rect 3877 3033 3914 3067
rect 3948 3033 3985 3067
rect 4019 3033 4056 3067
rect 4090 3033 4127 3067
rect 4161 3033 4198 3067
rect 4232 3033 4269 3067
rect 4303 3033 4340 3067
rect 4374 3033 4411 3067
rect 4445 3033 4482 3067
rect 4516 3033 4553 3067
rect 4587 3033 4624 3067
rect 4658 3033 4694 3067
rect 4728 3033 4752 3067
rect 3464 3025 4752 3033
rect 9640 3070 9674 3110
rect 271 2981 305 3015
rect 271 2913 305 2947
rect 9640 2996 9674 3036
rect -135 2837 -111 2871
rect -77 2837 6 2871
rect 40 2837 64 2871
rect 271 2845 305 2879
rect 271 2777 305 2811
rect 9640 2938 9674 2962
rect 12366 3612 12400 3646
rect 10442 3404 10476 3428
rect 12366 3544 12400 3578
rect 12366 3476 12400 3510
rect 12366 3408 12400 3442
rect 10442 3336 10476 3370
rect 12366 3340 12400 3374
rect 10442 3268 10476 3302
rect 10442 3200 10476 3234
rect 10442 3132 10476 3166
rect 12366 3272 12400 3306
rect 12366 3204 12400 3238
rect 12366 3136 12400 3170
rect 10442 3064 10476 3098
rect 10442 2996 10476 3030
rect 10442 2938 10476 2962
rect 271 2709 305 2743
rect 271 2641 305 2675
rect 271 2573 305 2607
rect 271 2505 305 2539
rect 271 2437 305 2471
rect 271 2369 305 2403
rect 271 2301 305 2335
rect 271 2233 305 2267
rect 271 2165 305 2199
rect 271 2097 305 2131
rect 271 2029 305 2063
rect 271 1961 305 1995
rect 271 1893 305 1927
rect 271 1825 305 1859
rect 271 1757 305 1791
rect 271 1689 305 1723
rect 12366 3068 12400 3102
rect 12366 3000 12400 3034
rect 12366 2932 12400 2966
rect 12366 2864 12400 2898
rect 12366 2796 12400 2830
rect 12366 2728 12400 2762
rect 12366 2660 12400 2694
rect 12366 2592 12400 2626
rect 12366 2524 12400 2558
rect 12366 2456 12400 2490
rect 12366 2388 12400 2422
rect 12366 2320 12400 2354
rect 12366 2252 12400 2286
rect 12366 2184 12400 2218
rect 12366 2116 12400 2150
rect 12366 2048 12400 2082
rect 12366 1980 12400 2014
rect 12366 1912 12400 1946
rect 12366 1844 12400 1878
rect 12366 1776 12400 1810
rect 271 1621 305 1655
rect 271 1553 305 1587
rect 12366 1708 12400 1742
rect 12366 1640 12400 1674
rect 271 1485 305 1519
rect 271 1417 305 1451
rect 271 1349 305 1383
rect 271 1281 305 1315
rect 271 1213 305 1247
rect 271 1145 305 1179
rect 271 1077 305 1111
rect 271 1009 305 1043
rect 271 941 305 975
rect 271 873 305 907
rect 271 805 305 839
rect 271 737 305 771
rect 271 669 305 703
rect 271 601 305 635
rect 609 626 633 796
rect 1075 626 1099 796
rect 271 533 305 567
rect 9656 1514 9694 1544
rect 9656 1480 9658 1514
rect 9692 1480 9694 1514
rect 9656 1446 9694 1480
rect 9656 1412 9658 1446
rect 9692 1412 9694 1446
rect 9656 1378 9694 1412
rect 9656 1344 9658 1378
rect 9692 1344 9694 1378
rect 9656 1310 9694 1344
rect 9656 1276 9658 1310
rect 9692 1276 9694 1310
rect 9656 1235 9694 1276
rect 9656 1201 9658 1235
rect 9692 1201 9694 1235
rect 9656 1167 9694 1201
rect 9656 1133 9658 1167
rect 9692 1133 9694 1167
rect 9656 1099 9694 1133
rect 9656 1065 9658 1099
rect 9692 1065 9694 1099
rect 9656 1031 9694 1065
rect 9656 997 9658 1031
rect 9692 997 9694 1031
rect 9656 948 9694 997
rect 12366 1572 12400 1606
rect 12366 1504 12400 1538
rect 12366 1436 12400 1470
rect 12366 1368 12400 1402
rect 12366 1300 12400 1334
rect 10496 1054 10530 1078
rect 10496 986 10530 1020
rect 10496 928 10530 952
rect 12366 1232 12400 1266
rect 12366 1164 12400 1198
rect 12366 1096 12400 1130
rect 12366 1028 12400 1062
rect 12366 960 12400 994
rect 12366 892 12400 926
rect 12366 824 12400 858
rect 12366 763 12400 790
rect 12366 729 12427 763
rect 12393 661 12427 695
rect 10286 618 10320 642
rect 10286 550 10320 584
rect 271 465 305 499
rect 10286 492 10320 516
rect 12393 593 12427 627
rect 12393 525 12427 559
rect 12393 457 12427 491
rect 271 349 305 431
rect 339 349 449 383
rect 483 349 517 383
rect 551 349 585 383
rect 619 349 653 383
rect 687 349 721 383
rect 755 349 789 383
rect 823 349 857 383
rect 891 349 925 383
rect 959 349 993 383
rect 1027 349 1061 383
rect 1095 349 1129 383
rect 1163 349 1197 383
rect 1231 349 1265 383
rect 1299 349 1333 383
rect 1367 349 1401 383
rect 1435 349 1469 383
rect 1503 349 1537 383
rect 1571 349 1605 383
rect 1639 349 1673 383
rect 1707 349 1741 383
rect 1775 349 1809 383
rect 1843 349 1877 383
rect 1911 349 1945 383
rect 1979 349 2013 383
rect 2047 349 2081 383
rect 2115 349 2149 383
rect 2183 349 2217 383
rect 2251 349 2285 383
rect 2319 349 2353 383
rect 2387 349 2421 383
rect 2455 349 2489 383
rect 2523 349 2557 383
rect 2591 349 2625 383
rect 2659 349 2693 383
rect 2727 349 2761 383
rect 2795 349 2829 383
rect 2863 349 2897 383
rect 2931 349 2965 383
rect 2999 349 3033 383
rect 3067 349 3101 383
rect 3135 349 3169 383
rect 3203 349 3237 383
rect 3271 349 3305 383
rect 3339 349 3373 383
rect 3407 349 3441 383
rect 3475 349 3509 383
rect 3543 349 3577 383
rect 3611 349 3645 383
rect 3679 349 3713 383
rect 3747 349 3781 383
rect 3815 349 3849 383
rect 3883 349 3917 383
rect 3951 349 3985 383
rect 4019 349 4053 383
rect 4087 349 4121 383
rect 4155 349 4189 383
rect 4223 349 4257 383
rect 4291 349 4325 383
rect 4359 349 4393 383
rect 4427 349 4461 383
rect 4495 349 4529 383
rect 4563 349 4597 383
rect 4631 349 4665 383
rect 4699 349 4733 383
rect 4767 349 4801 383
rect 4835 349 4869 383
rect 4903 349 4937 383
rect 4971 349 5005 383
rect 5039 349 5073 383
rect 5107 349 5141 383
rect 5175 349 5209 383
rect 5243 349 5277 383
rect 5311 349 5345 383
rect 5379 349 5413 383
rect 5447 349 5481 383
rect 5515 349 5549 383
rect 5583 349 5617 383
rect 5651 349 5685 383
rect 5719 349 5753 383
rect 5787 349 5821 383
rect 5855 349 5889 383
rect 5923 349 5957 383
rect 5991 349 6025 383
rect 6059 349 6093 383
rect 6127 349 6161 383
rect 6195 349 6229 383
rect 6263 349 6297 383
rect 6331 349 6365 383
rect 6399 349 6433 383
rect 6467 349 6501 383
rect 6535 349 6569 383
rect 6603 349 6637 383
rect 6671 349 6705 383
rect 6739 349 6773 383
rect 6807 349 6841 383
rect 6875 349 6909 383
rect 6943 349 6977 383
rect 7011 349 7045 383
rect 7079 349 7113 383
rect 7147 349 7181 383
rect 7215 349 7249 383
rect 7283 349 7317 383
rect 7351 349 7385 383
rect 7419 349 7453 383
rect 7487 349 7521 383
rect 7555 349 7589 383
rect 7623 349 7657 383
rect 7691 349 7725 383
rect 7759 349 7793 383
rect 7827 349 7861 383
rect 7895 349 7929 383
rect 7963 349 7997 383
rect 8031 349 8098 383
rect 8064 308 8098 349
rect 8132 308 8166 342
rect 8200 308 8234 342
rect 8268 308 8302 342
rect 8336 308 8370 342
rect 8404 308 8438 342
rect 8472 308 8506 342
rect 8540 308 8574 342
rect 8608 308 8642 342
rect 8676 308 8710 342
rect 8744 308 8778 342
rect 8812 308 8846 342
rect 8880 308 8914 342
rect 8948 308 8982 342
rect 9016 308 9050 342
rect 9084 308 9118 342
rect 9152 308 9186 342
rect 9220 308 9254 342
rect 9288 308 9322 342
rect 9356 308 9390 342
rect 9424 308 9458 342
rect 9492 308 9526 342
rect 9560 308 9594 342
rect 9628 308 9662 342
rect 9696 308 9730 342
rect 9764 308 9798 342
rect 9832 308 9866 342
rect 9900 308 9934 342
rect 9968 308 10002 342
rect 10036 308 10070 342
rect 10104 308 10138 342
rect 10172 308 10206 342
rect 10240 308 10274 342
rect 10308 308 10342 342
rect 10376 308 10410 342
rect 10444 308 10478 342
rect 10512 308 10546 342
rect 10580 308 10614 342
rect 10648 308 10682 342
rect 10716 308 10750 342
rect 10784 308 10818 342
rect 10852 308 10886 342
rect 10920 308 10954 342
rect 10988 308 11022 342
rect 11056 308 11090 342
rect 11124 308 11158 342
rect 11192 308 11226 342
rect 11260 308 11294 342
rect 11328 308 11362 342
rect 11396 308 11430 342
rect 11464 308 11498 342
rect 11532 308 11566 342
rect 11600 308 11634 342
rect 11668 308 11702 342
rect 11736 308 11770 342
rect 11804 308 11838 342
rect 11872 308 11906 342
rect 11940 308 11974 342
rect 12008 308 12042 342
rect 12076 308 12110 342
rect 12144 308 12178 342
rect 12212 308 12359 342
rect 12393 308 12427 423
<< psubdiffcont >>
rect -615 4057 -581 4091
rect -615 3968 -581 4002
rect -615 3878 -581 3912
rect -615 3788 -581 3822
<< mvpsubdiffcont >>
rect 8751 4085 8785 4119
rect 8851 4085 8885 4119
rect 8951 4085 8985 4119
rect 8751 4012 8785 4046
rect 8851 4012 8885 4046
rect 8951 4012 8985 4046
rect 8751 3939 8785 3973
rect 8851 3939 8885 3973
rect 8951 3939 8985 3973
rect 8751 3866 8785 3900
rect 8851 3866 8885 3900
rect 8951 3866 8985 3900
rect 8751 3793 8785 3827
rect 8851 3793 8885 3827
rect 8951 3793 8985 3827
rect 8751 3720 8785 3754
rect 8851 3720 8885 3754
rect 8951 3720 8985 3754
rect 8751 3647 8785 3681
rect 8851 3647 8885 3681
rect 8951 3647 8985 3681
rect 8751 3573 8785 3607
rect 8851 3573 8885 3607
rect 8951 3573 8985 3607
rect 8751 3499 8785 3533
rect 8851 3499 8885 3533
rect 8951 3499 8985 3533
rect 8751 3425 8785 3459
rect 8851 3425 8885 3459
rect 8951 3425 8985 3459
rect 8751 3351 8785 3385
rect 8851 3351 8885 3385
rect 8951 3351 8985 3385
rect 8751 3277 8785 3311
rect 8851 3277 8885 3311
rect 8951 3277 8985 3311
rect 10744 3039 10778 3073
rect 10744 2971 10778 3005
rect -409 1745 -375 1779
rect -331 1745 -297 1779
rect -253 1745 -219 1779
rect -175 1745 -141 1779
rect -97 1745 -63 1779
rect -20 1745 14 1779
rect 57 1745 91 1779
rect 10744 2903 10778 2937
rect 10744 2835 10778 2869
rect 10744 2767 10778 2801
rect 10744 2698 10778 2732
rect 10744 2629 10778 2663
rect 10744 2560 10778 2594
rect 9445 2250 9479 2284
rect 9513 2250 9547 2284
rect 9445 2176 9479 2210
rect 9513 2176 9547 2210
rect 9445 2102 9479 2136
rect 9513 2102 9547 2136
rect 9445 2028 9479 2062
rect 9513 2028 9547 2062
rect 9445 1954 9479 1988
rect 9513 1954 9547 1988
rect 9445 1880 9479 1914
rect 9513 1880 9547 1914
rect 9445 1806 9479 1840
rect 9513 1806 9547 1840
rect 9445 1732 9479 1766
rect 9513 1732 9547 1766
rect 10486 2221 10520 2255
rect 10486 2153 10520 2187
rect 10486 2085 10520 2119
rect 10486 2017 10520 2051
rect 10486 1949 10520 1983
rect 10486 1881 10520 1915
rect 10486 1813 10520 1847
rect 12133 2278 12167 2312
rect 12133 2203 12167 2237
rect 12133 2128 12167 2162
rect 12133 2054 12167 2088
rect 12133 1980 12167 2014
rect 12133 1906 12167 1940
rect 12133 1832 12167 1866
<< mvnsubdiffcont >>
rect -478 4907 -444 4941
rect -406 4907 -372 4941
rect -334 4907 -300 4941
rect -262 4907 -228 4941
rect -190 4907 -156 4941
rect -119 4907 -85 4941
rect -48 4907 -14 4941
rect 23 4907 57 4941
rect 94 4907 128 4941
rect 10909 4546 10943 4580
rect 10980 4546 11014 4580
rect 11051 4546 11085 4580
rect 11122 4546 11156 4580
rect 11193 4546 11227 4580
rect 11264 4546 11298 4580
rect 11335 4546 11369 4580
rect 11406 4546 11440 4580
rect 11477 4546 11511 4580
rect 11548 4546 11582 4580
rect 11619 4546 11653 4580
rect 11690 4546 11724 4580
rect 11761 4546 11795 4580
rect 11832 4546 11866 4580
rect 11903 4546 11937 4580
rect 11974 4546 12008 4580
rect 12045 4546 12079 4580
rect 12116 4546 12150 4580
rect 12187 4546 12221 4580
rect 12258 4546 12292 4580
rect 12329 4546 12363 4580
rect 10839 4472 10873 4506
rect 409 4426 443 4460
rect 477 4426 511 4460
rect 545 4426 579 4460
rect 613 4426 647 4460
rect 681 4426 715 4460
rect 749 4426 783 4460
rect 817 4426 851 4460
rect 885 4426 919 4460
rect 953 4426 987 4460
rect 1021 4426 1055 4460
rect 1089 4426 1123 4460
rect 1157 4426 1191 4460
rect 1225 4426 1259 4460
rect 1293 4426 1327 4460
rect 1361 4426 1395 4460
rect 1429 4426 1463 4460
rect 1497 4426 1531 4460
rect 1565 4426 1599 4460
rect 1633 4426 1667 4460
rect 1701 4426 1735 4460
rect 1769 4426 1803 4460
rect 1837 4426 1871 4460
rect 1905 4426 1939 4460
rect 1973 4426 2007 4460
rect 2041 4426 2075 4460
rect 2109 4426 2143 4460
rect 2177 4426 2211 4460
rect 2245 4426 2279 4460
rect 2313 4426 2347 4460
rect 2381 4426 2415 4460
rect 2449 4426 2483 4460
rect 2517 4426 2551 4460
rect 2585 4426 2619 4460
rect 2653 4426 2687 4460
rect 2721 4426 2755 4460
rect 2789 4426 2823 4460
rect 2857 4426 2891 4460
rect 2925 4426 2959 4460
rect 2993 4426 3027 4460
rect 3061 4426 3095 4460
rect 3129 4426 3163 4460
rect 3197 4426 3231 4460
rect 3265 4426 3299 4460
rect 3333 4426 3367 4460
rect 3401 4426 3435 4460
rect 3469 4426 3503 4460
rect 3537 4426 3571 4460
rect 3605 4426 3639 4460
rect 3673 4426 3707 4460
rect 3741 4426 3775 4460
rect 3809 4426 3843 4460
rect 3877 4426 3911 4460
rect 3945 4426 3979 4460
rect 4013 4426 4047 4460
rect 4081 4426 4115 4460
rect 4149 4426 4183 4460
rect 4217 4426 4251 4460
rect 4285 4426 4319 4460
rect 4353 4426 4387 4460
rect 4421 4426 4455 4460
rect 4489 4426 4523 4460
rect 4557 4426 4591 4460
rect 4625 4426 4659 4460
rect 4693 4426 4727 4460
rect 4761 4426 4795 4460
rect 4829 4426 4863 4460
rect 4897 4426 4931 4460
rect 4965 4426 4999 4460
rect 5033 4426 5067 4460
rect 5101 4426 5135 4460
rect 5169 4426 5203 4460
rect 5237 4426 5271 4460
rect 5305 4426 5339 4460
rect 5373 4426 5407 4460
rect 5441 4426 5475 4460
rect 5509 4426 5543 4460
rect 5577 4426 5611 4460
rect 5645 4426 5679 4460
rect 5713 4426 5747 4460
rect 5781 4426 5815 4460
rect 5849 4426 5883 4460
rect 5917 4426 5951 4460
rect 5985 4426 6019 4460
rect 6053 4426 6087 4460
rect 6121 4426 6155 4460
rect 6189 4426 6223 4460
rect 6257 4426 6291 4460
rect 6325 4426 6359 4460
rect 6393 4426 6427 4460
rect 6461 4426 6495 4460
rect 6529 4426 6563 4460
rect 6597 4426 6631 4460
rect 6665 4426 6699 4460
rect 6733 4426 6767 4460
rect 6801 4426 6835 4460
rect 6869 4426 6903 4460
rect 6937 4426 6971 4460
rect 7005 4426 7039 4460
rect 7073 4426 7107 4460
rect 7141 4426 7175 4460
rect 7209 4426 7243 4460
rect 7277 4426 7311 4460
rect 7345 4426 7379 4460
rect 7413 4426 7447 4460
rect 7481 4426 7515 4460
rect 7549 4426 7583 4460
rect 7617 4426 7651 4460
rect 7685 4426 7719 4460
rect 7753 4426 7787 4460
rect 7821 4426 7855 4460
rect 7889 4426 7923 4460
rect 7957 4426 7991 4460
rect 8025 4426 8059 4460
rect 8093 4426 8127 4460
rect 8161 4426 8195 4460
rect 8229 4426 8263 4460
rect 8297 4426 8331 4460
rect 8365 4426 8399 4460
rect 8433 4426 8467 4460
rect 8501 4426 8535 4460
rect 8569 4426 8603 4460
rect 8637 4426 8671 4460
rect 8705 4426 8739 4460
rect 8773 4426 8807 4460
rect 8841 4426 8875 4460
rect 8909 4426 8943 4460
rect 8977 4426 9011 4460
rect 9045 4426 9079 4460
rect 9113 4426 9147 4460
rect 9181 4426 9215 4460
rect 9249 4426 9283 4460
rect 9317 4426 9351 4460
rect 9385 4426 9419 4460
rect 9453 4426 9487 4460
rect 9521 4426 9555 4460
rect 9589 4426 9623 4460
rect 9657 4426 9691 4460
rect 9725 4426 9759 4460
rect 9793 4426 9827 4460
rect 9861 4426 9895 4460
rect 9929 4426 9963 4460
rect 9997 4426 10031 4460
rect 10065 4426 10099 4460
rect 10133 4426 10167 4460
rect 10201 4426 10235 4460
rect 10269 4426 10303 4460
rect 10337 4426 10371 4460
rect 10405 4426 10439 4460
rect 10473 4426 10507 4460
rect 10541 4426 10575 4460
rect 10609 4426 10643 4460
rect 271 4375 305 4409
rect 10760 4397 10794 4431
rect 12366 4462 12400 4496
rect 12366 4394 12400 4428
rect 271 4307 305 4341
rect 12366 4326 12400 4360
rect 271 4239 305 4273
rect 271 4171 305 4205
rect 271 4103 305 4137
rect 271 4035 305 4069
rect 271 3967 305 4001
rect 271 3899 305 3933
rect 271 3831 305 3865
rect 271 3763 305 3797
rect 271 3695 305 3729
rect 271 3627 305 3661
rect 271 3559 305 3593
rect 271 3491 305 3525
rect 271 3423 305 3457
rect 271 3355 305 3389
rect 271 3287 305 3321
rect 271 3219 305 3253
rect 1016 4130 1050 4164
rect 1016 4062 1050 4096
rect 1016 3994 1050 4028
rect 1016 3926 1050 3960
rect 1016 3858 1050 3892
rect 1016 3790 1050 3824
rect 1016 3722 1050 3756
rect 1016 3654 1050 3688
rect 1016 3586 1050 3620
rect 1016 3518 1050 3552
rect 1016 3450 1050 3484
rect 1016 3382 1050 3416
rect 1016 3314 1050 3348
rect 1016 3246 1050 3280
rect 2882 4130 2916 4164
rect 2882 4062 2916 4096
rect 2882 3994 2916 4028
rect 2882 3926 2916 3960
rect 2882 3858 2916 3892
rect 2882 3790 2916 3824
rect 2882 3722 2916 3756
rect 2882 3654 2916 3688
rect 2882 3586 2916 3620
rect 2882 3518 2916 3552
rect 2882 3450 2916 3484
rect 2882 3382 2916 3416
rect 2882 3314 2916 3348
rect 2882 3246 2916 3280
rect 4326 4130 4360 4164
rect 4326 4062 4360 4096
rect 4326 3994 4360 4028
rect 4326 3926 4360 3960
rect 4326 3858 4360 3892
rect 4326 3790 4360 3824
rect 4326 3722 4360 3756
rect 4326 3654 4360 3688
rect 4326 3586 4360 3620
rect 4326 3518 4360 3552
rect 4326 3450 4360 3484
rect 4326 3382 4360 3416
rect 4326 3314 4360 3348
rect 4326 3246 4360 3280
rect 5770 4130 5804 4164
rect 5770 4062 5804 4096
rect 5770 3994 5804 4028
rect 5770 3926 5804 3960
rect 5770 3858 5804 3892
rect 5770 3790 5804 3824
rect 5770 3722 5804 3756
rect 5770 3654 5804 3688
rect 5770 3586 5804 3620
rect 5770 3518 5804 3552
rect 5770 3450 5804 3484
rect 5770 3382 5804 3416
rect 5770 3314 5804 3348
rect 5770 3246 5804 3280
rect 7370 4130 7404 4164
rect 7370 4062 7404 4096
rect 7370 3994 7404 4028
rect 7370 3926 7404 3960
rect 7370 3858 7404 3892
rect 7370 3790 7404 3824
rect 7370 3722 7404 3756
rect 7370 3654 7404 3688
rect 7370 3586 7404 3620
rect 8166 4130 8200 4164
rect 8166 4062 8200 4096
rect 7370 3518 7404 3552
rect 7370 3450 7404 3484
rect 7370 3382 7404 3416
rect 7370 3314 7404 3348
rect 7370 3246 7404 3280
rect 8166 3994 8200 4028
rect 8166 3926 8200 3960
rect 8166 3858 8200 3892
rect 8166 3790 8200 3824
rect 8166 3722 8200 3756
rect 8166 3654 8200 3688
rect 8166 3586 8200 3620
rect 8166 3518 8200 3552
rect 8166 3450 8200 3484
rect 8166 3382 8200 3416
rect 8166 3314 8200 3348
rect 271 3151 305 3185
rect 271 3083 305 3117
rect 8166 3246 8200 3280
rect 12366 4258 12400 4292
rect 12366 4190 12400 4224
rect 12366 4122 12400 4156
rect 12366 4054 12400 4088
rect 12366 3986 12400 4020
rect 12366 3918 12400 3952
rect 12366 3850 12400 3884
rect 12366 3782 12400 3816
rect 12366 3714 12400 3748
rect 9459 3479 9493 3513
rect 9459 3378 9493 3412
rect 9459 3277 9493 3311
rect 9640 3480 9674 3514
rect 9640 3406 9674 3440
rect 9640 3332 9674 3366
rect 9640 3258 9674 3292
rect 9640 3184 9674 3218
rect 9640 3110 9674 3144
rect 271 3015 305 3049
rect 3488 3033 3522 3067
rect 3559 3033 3593 3067
rect 3630 3033 3664 3067
rect 3701 3033 3735 3067
rect 3772 3033 3806 3067
rect 3843 3033 3877 3067
rect 3914 3033 3948 3067
rect 3985 3033 4019 3067
rect 4056 3033 4090 3067
rect 4127 3033 4161 3067
rect 4198 3033 4232 3067
rect 4269 3033 4303 3067
rect 4340 3033 4374 3067
rect 4411 3033 4445 3067
rect 4482 3033 4516 3067
rect 4553 3033 4587 3067
rect 4624 3033 4658 3067
rect 4694 3033 4728 3067
rect 271 2947 305 2981
rect 9640 3036 9674 3070
rect 271 2879 305 2913
rect -111 2837 -77 2871
rect 6 2837 40 2871
rect 271 2811 305 2845
rect 271 2743 305 2777
rect 9640 2962 9674 2996
rect 12366 3646 12400 3680
rect 10442 3370 10476 3404
rect 12366 3578 12400 3612
rect 12366 3510 12400 3544
rect 12366 3442 12400 3476
rect 10442 3302 10476 3336
rect 12366 3374 12400 3408
rect 12366 3306 12400 3340
rect 10442 3234 10476 3268
rect 10442 3166 10476 3200
rect 10442 3098 10476 3132
rect 12366 3238 12400 3272
rect 12366 3170 12400 3204
rect 10442 3030 10476 3064
rect 10442 2962 10476 2996
rect 271 2675 305 2709
rect 271 2607 305 2641
rect 271 2539 305 2573
rect 271 2471 305 2505
rect 271 2403 305 2437
rect 271 2335 305 2369
rect 271 2267 305 2301
rect 271 2199 305 2233
rect 271 2131 305 2165
rect 271 2063 305 2097
rect 271 1995 305 2029
rect 271 1927 305 1961
rect 271 1859 305 1893
rect 271 1791 305 1825
rect 271 1723 305 1757
rect 12366 3102 12400 3136
rect 12366 3034 12400 3068
rect 12366 2966 12400 3000
rect 12366 2898 12400 2932
rect 12366 2830 12400 2864
rect 12366 2762 12400 2796
rect 12366 2694 12400 2728
rect 12366 2626 12400 2660
rect 12366 2558 12400 2592
rect 12366 2490 12400 2524
rect 12366 2422 12400 2456
rect 12366 2354 12400 2388
rect 12366 2286 12400 2320
rect 12366 2218 12400 2252
rect 12366 2150 12400 2184
rect 12366 2082 12400 2116
rect 12366 2014 12400 2048
rect 12366 1946 12400 1980
rect 12366 1878 12400 1912
rect 12366 1810 12400 1844
rect 271 1655 305 1689
rect 271 1587 305 1621
rect 12366 1742 12400 1776
rect 12366 1674 12400 1708
rect 271 1519 305 1553
rect 271 1451 305 1485
rect 271 1383 305 1417
rect 271 1315 305 1349
rect 271 1247 305 1281
rect 271 1179 305 1213
rect 271 1111 305 1145
rect 271 1043 305 1077
rect 271 975 305 1009
rect 271 907 305 941
rect 271 839 305 873
rect 271 771 305 805
rect 271 703 305 737
rect 271 635 305 669
rect 633 626 1075 796
rect 271 567 305 601
rect 9658 1480 9692 1514
rect 9658 1412 9692 1446
rect 9658 1344 9692 1378
rect 9658 1276 9692 1310
rect 9658 1201 9692 1235
rect 9658 1133 9692 1167
rect 9658 1065 9692 1099
rect 9658 997 9692 1031
rect 12366 1606 12400 1640
rect 12366 1538 12400 1572
rect 12366 1470 12400 1504
rect 12366 1402 12400 1436
rect 12366 1334 12400 1368
rect 12366 1266 12400 1300
rect 10496 1020 10530 1054
rect 10496 952 10530 986
rect 12366 1198 12400 1232
rect 12366 1130 12400 1164
rect 12366 1062 12400 1096
rect 12366 994 12400 1028
rect 12366 926 12400 960
rect 12366 858 12400 892
rect 12366 790 12400 824
rect 12393 695 12427 729
rect 10286 584 10320 618
rect 271 499 305 533
rect 271 431 305 465
rect 10286 516 10320 550
rect 12393 627 12427 661
rect 12393 559 12427 593
rect 12393 491 12427 525
rect 12393 423 12427 457
rect 305 349 339 383
rect 449 349 483 383
rect 517 349 551 383
rect 585 349 619 383
rect 653 349 687 383
rect 721 349 755 383
rect 789 349 823 383
rect 857 349 891 383
rect 925 349 959 383
rect 993 349 1027 383
rect 1061 349 1095 383
rect 1129 349 1163 383
rect 1197 349 1231 383
rect 1265 349 1299 383
rect 1333 349 1367 383
rect 1401 349 1435 383
rect 1469 349 1503 383
rect 1537 349 1571 383
rect 1605 349 1639 383
rect 1673 349 1707 383
rect 1741 349 1775 383
rect 1809 349 1843 383
rect 1877 349 1911 383
rect 1945 349 1979 383
rect 2013 349 2047 383
rect 2081 349 2115 383
rect 2149 349 2183 383
rect 2217 349 2251 383
rect 2285 349 2319 383
rect 2353 349 2387 383
rect 2421 349 2455 383
rect 2489 349 2523 383
rect 2557 349 2591 383
rect 2625 349 2659 383
rect 2693 349 2727 383
rect 2761 349 2795 383
rect 2829 349 2863 383
rect 2897 349 2931 383
rect 2965 349 2999 383
rect 3033 349 3067 383
rect 3101 349 3135 383
rect 3169 349 3203 383
rect 3237 349 3271 383
rect 3305 349 3339 383
rect 3373 349 3407 383
rect 3441 349 3475 383
rect 3509 349 3543 383
rect 3577 349 3611 383
rect 3645 349 3679 383
rect 3713 349 3747 383
rect 3781 349 3815 383
rect 3849 349 3883 383
rect 3917 349 3951 383
rect 3985 349 4019 383
rect 4053 349 4087 383
rect 4121 349 4155 383
rect 4189 349 4223 383
rect 4257 349 4291 383
rect 4325 349 4359 383
rect 4393 349 4427 383
rect 4461 349 4495 383
rect 4529 349 4563 383
rect 4597 349 4631 383
rect 4665 349 4699 383
rect 4733 349 4767 383
rect 4801 349 4835 383
rect 4869 349 4903 383
rect 4937 349 4971 383
rect 5005 349 5039 383
rect 5073 349 5107 383
rect 5141 349 5175 383
rect 5209 349 5243 383
rect 5277 349 5311 383
rect 5345 349 5379 383
rect 5413 349 5447 383
rect 5481 349 5515 383
rect 5549 349 5583 383
rect 5617 349 5651 383
rect 5685 349 5719 383
rect 5753 349 5787 383
rect 5821 349 5855 383
rect 5889 349 5923 383
rect 5957 349 5991 383
rect 6025 349 6059 383
rect 6093 349 6127 383
rect 6161 349 6195 383
rect 6229 349 6263 383
rect 6297 349 6331 383
rect 6365 349 6399 383
rect 6433 349 6467 383
rect 6501 349 6535 383
rect 6569 349 6603 383
rect 6637 349 6671 383
rect 6705 349 6739 383
rect 6773 349 6807 383
rect 6841 349 6875 383
rect 6909 349 6943 383
rect 6977 349 7011 383
rect 7045 349 7079 383
rect 7113 349 7147 383
rect 7181 349 7215 383
rect 7249 349 7283 383
rect 7317 349 7351 383
rect 7385 349 7419 383
rect 7453 349 7487 383
rect 7521 349 7555 383
rect 7589 349 7623 383
rect 7657 349 7691 383
rect 7725 349 7759 383
rect 7793 349 7827 383
rect 7861 349 7895 383
rect 7929 349 7963 383
rect 7997 349 8031 383
rect 8098 308 8132 342
rect 8166 308 8200 342
rect 8234 308 8268 342
rect 8302 308 8336 342
rect 8370 308 8404 342
rect 8438 308 8472 342
rect 8506 308 8540 342
rect 8574 308 8608 342
rect 8642 308 8676 342
rect 8710 308 8744 342
rect 8778 308 8812 342
rect 8846 308 8880 342
rect 8914 308 8948 342
rect 8982 308 9016 342
rect 9050 308 9084 342
rect 9118 308 9152 342
rect 9186 308 9220 342
rect 9254 308 9288 342
rect 9322 308 9356 342
rect 9390 308 9424 342
rect 9458 308 9492 342
rect 9526 308 9560 342
rect 9594 308 9628 342
rect 9662 308 9696 342
rect 9730 308 9764 342
rect 9798 308 9832 342
rect 9866 308 9900 342
rect 9934 308 9968 342
rect 10002 308 10036 342
rect 10070 308 10104 342
rect 10138 308 10172 342
rect 10206 308 10240 342
rect 10274 308 10308 342
rect 10342 308 10376 342
rect 10410 308 10444 342
rect 10478 308 10512 342
rect 10546 308 10580 342
rect 10614 308 10648 342
rect 10682 308 10716 342
rect 10750 308 10784 342
rect 10818 308 10852 342
rect 10886 308 10920 342
rect 10954 308 10988 342
rect 11022 308 11056 342
rect 11090 308 11124 342
rect 11158 308 11192 342
rect 11226 308 11260 342
rect 11294 308 11328 342
rect 11362 308 11396 342
rect 11430 308 11464 342
rect 11498 308 11532 342
rect 11566 308 11600 342
rect 11634 308 11668 342
rect 11702 308 11736 342
rect 11770 308 11804 342
rect 11838 308 11872 342
rect 11906 308 11940 342
rect 11974 308 12008 342
rect 12042 308 12076 342
rect 12110 308 12144 342
rect 12178 308 12212 342
rect 12359 308 12393 342
<< poly >>
rect -408 4833 -288 4859
rect -232 4833 -112 4859
rect -56 4833 64 4859
rect -408 4565 -288 4633
rect -232 4565 -112 4633
rect -56 4565 64 4633
rect 13335 4597 13469 4613
rect 13335 4563 13351 4597
rect 13385 4563 13419 4597
rect 13453 4563 13469 4597
rect 13335 4547 13469 4563
rect 13335 4479 13455 4547
rect -408 4317 -288 4365
rect -408 4283 -366 4317
rect -332 4283 -288 4317
rect -408 4249 -288 4283
rect -408 4215 -366 4249
rect -332 4215 -288 4249
rect -408 4167 -288 4215
rect -232 4317 -112 4365
rect -232 4283 -186 4317
rect -152 4283 -112 4317
rect -232 4249 -112 4283
rect -232 4215 -186 4249
rect -152 4215 -112 4249
rect -232 4167 -112 4215
rect -56 4317 64 4365
rect -56 4283 -15 4317
rect 19 4283 64 4317
rect -56 4249 64 4283
rect -56 4215 -15 4249
rect 19 4215 64 4249
rect -56 4167 64 4215
rect 4469 4335 5661 4351
rect 4469 4301 4505 4335
rect 4539 4301 4573 4335
rect 4607 4301 4641 4335
rect 4675 4301 4709 4335
rect 4743 4301 4777 4335
rect 4811 4301 4845 4335
rect 4879 4301 4913 4335
rect 4947 4301 4981 4335
rect 5015 4301 5049 4335
rect 5083 4301 5117 4335
rect 5151 4301 5185 4335
rect 5219 4301 5253 4335
rect 5287 4301 5321 4335
rect 5355 4301 5389 4335
rect 5423 4301 5457 4335
rect 5491 4301 5525 4335
rect 5559 4301 5593 4335
rect 5627 4301 5661 4335
rect 9190 4318 9290 4350
rect 9346 4318 9446 4350
rect 9502 4318 9602 4350
rect 9782 4318 9882 4350
rect 9938 4318 10038 4350
rect 10094 4318 10194 4350
rect 10250 4318 10350 4350
rect 10530 4318 10630 4350
rect 10686 4318 10786 4350
rect 1581 4285 2148 4301
rect 1581 4251 1609 4285
rect 1643 4251 1677 4285
rect 1711 4251 1745 4285
rect 1779 4251 1813 4285
rect 1847 4251 1881 4285
rect 1915 4251 1949 4285
rect 1983 4251 2017 4285
rect 2051 4251 2085 4285
rect 2119 4251 2148 4285
rect 1581 4229 2148 4251
rect 2205 4285 2772 4301
rect 2205 4251 2233 4285
rect 2267 4251 2301 4285
rect 2335 4251 2369 4285
rect 2403 4251 2437 4285
rect 2471 4251 2505 4285
rect 2539 4251 2573 4285
rect 2607 4251 2641 4285
rect 2675 4251 2709 4285
rect 2743 4251 2772 4285
rect 2205 4229 2772 4251
rect 3025 4285 4217 4301
rect 3025 4251 3061 4285
rect 3095 4251 3129 4285
rect 3163 4251 3197 4285
rect 3231 4251 3265 4285
rect 3299 4251 3333 4285
rect 3367 4251 3401 4285
rect 3435 4251 3469 4285
rect 3503 4251 3537 4285
rect 3571 4251 3605 4285
rect 3639 4251 3673 4285
rect 3707 4251 3741 4285
rect 3775 4251 3809 4285
rect 3843 4251 3877 4285
rect 3911 4251 3945 4285
rect 3979 4251 4013 4285
rect 4047 4251 4081 4285
rect 4115 4251 4149 4285
rect 4183 4251 4217 4285
rect 4469 4279 5661 4301
rect 4469 4253 4569 4279
rect 4625 4253 4725 4279
rect 4781 4253 4881 4279
rect 4937 4253 5037 4279
rect 5093 4253 5193 4279
rect 5249 4253 5349 4279
rect 5405 4253 5505 4279
rect 5561 4253 5661 4279
rect 5913 4285 7105 4301
rect 3025 4229 4217 4251
rect 1159 4203 1259 4229
rect 1315 4203 1415 4229
rect 1581 4203 1681 4229
rect 1737 4203 1837 4229
rect 1893 4203 1993 4229
rect 2049 4203 2149 4229
rect 2205 4203 2305 4229
rect 2361 4203 2461 4229
rect 2517 4203 2617 4229
rect 2673 4203 2773 4229
rect 3025 4203 3125 4229
rect 3181 4203 3281 4229
rect 3337 4203 3437 4229
rect 3493 4203 3593 4229
rect 3649 4203 3749 4229
rect 3805 4203 3905 4229
rect 3961 4203 4061 4229
rect 4117 4203 4217 4229
rect -408 4001 -288 4027
rect -232 4001 -112 4027
rect -56 4001 64 4027
rect -425 3845 -325 3871
rect -145 3845 -25 3871
rect -425 3700 -325 3761
rect -425 3666 -394 3700
rect -360 3666 -325 3700
rect -425 3632 -325 3666
rect -425 3598 -394 3632
rect -360 3598 -325 3632
rect -425 3507 -325 3598
rect -145 3657 -25 3705
rect -145 3623 -101 3657
rect -67 3623 -25 3657
rect -145 3589 -25 3623
rect -145 3555 -101 3589
rect -67 3555 -25 3589
rect -145 3507 -25 3555
rect -145 3239 -25 3307
rect 5913 4251 5950 4285
rect 5984 4251 6018 4285
rect 6052 4251 6086 4285
rect 6120 4251 6154 4285
rect 6188 4251 6222 4285
rect 6256 4251 6290 4285
rect 6324 4251 6358 4285
rect 6392 4251 6426 4285
rect 6460 4251 6494 4285
rect 6528 4251 6562 4285
rect 6596 4251 6630 4285
rect 6664 4251 6698 4285
rect 6732 4251 6766 4285
rect 6800 4251 6834 4285
rect 6868 4251 6902 4285
rect 6936 4251 6970 4285
rect 7004 4251 7038 4285
rect 7072 4251 7105 4285
rect 5913 4229 7105 4251
rect 5913 4203 6013 4229
rect 6069 4203 6169 4229
rect 6225 4203 6325 4229
rect 6381 4203 6481 4229
rect 6537 4203 6637 4229
rect 6693 4203 6793 4229
rect 6849 4203 6949 4229
rect 7005 4203 7105 4229
rect 7161 4285 7295 4301
rect 7161 4251 7177 4285
rect 7211 4251 7245 4285
rect 7279 4251 7295 4285
rect 7161 4229 7295 4251
rect 7462 4285 7596 4301
rect 7462 4251 7478 4285
rect 7512 4251 7546 4285
rect 7580 4251 7596 4285
rect 7462 4229 7596 4251
rect 7814 4285 7948 4301
rect 7814 4251 7830 4285
rect 7864 4251 7898 4285
rect 7932 4251 7948 4285
rect 7814 4229 7948 4251
rect 7161 4203 7261 4229
rect 7513 4203 7613 4229
rect 7655 4203 7755 4229
rect 7797 4203 7897 4229
rect 4469 3227 4569 3253
rect 4625 3227 4725 3253
rect 4781 3227 4881 3253
rect 4937 3227 5037 3253
rect 5093 3227 5193 3253
rect 5249 3227 5349 3253
rect 5405 3227 5505 3253
rect 5561 3227 5661 3253
rect 7513 3577 7613 3603
rect 7655 3542 7755 3603
rect 7797 3577 7897 3603
rect 7638 3526 7772 3542
rect 8000 3526 8026 4056
rect 7638 3492 7654 3526
rect 7688 3492 7722 3526
rect 7756 3492 7772 3526
rect 7638 3476 7772 3492
rect 7928 3510 8026 3526
rect 7928 3476 7944 3510
rect 7978 3476 8026 3510
rect 7928 3442 8026 3476
rect 7513 3408 7613 3434
rect 7669 3408 7769 3434
rect 7928 3408 7944 3442
rect 7978 3408 8026 3442
rect 7928 3374 8026 3408
rect 7928 3340 7944 3374
rect 7978 3340 8026 3374
rect 7928 3306 8026 3340
rect 7928 3272 7944 3306
rect 7978 3272 8026 3306
rect 7928 3256 8026 3272
rect 8110 3256 8136 4056
rect 1159 3177 1259 3203
rect 1315 3177 1415 3203
rect 1581 3177 1681 3203
rect 1737 3177 1837 3203
rect 1893 3177 1993 3203
rect 2049 3177 2149 3203
rect 2205 3177 2305 3203
rect 2361 3177 2461 3203
rect 2517 3177 2617 3203
rect 2673 3177 2773 3203
rect 3025 3177 3125 3203
rect 3181 3177 3281 3203
rect 3337 3177 3437 3203
rect 3493 3177 3593 3203
rect 3649 3177 3749 3203
rect 3805 3177 3905 3203
rect 3961 3177 4061 3203
rect 4117 3177 4217 3203
rect 5913 3177 6013 3203
rect 6069 3177 6169 3203
rect 6225 3177 6325 3203
rect 6381 3177 6481 3203
rect 6537 3177 6637 3203
rect 6693 3177 6793 3203
rect 6849 3177 6949 3203
rect 7005 3177 7105 3203
rect 7161 3177 7261 3203
rect 7513 3182 7613 3208
rect 7669 3182 7769 3208
rect 8262 4017 8354 4056
rect 8262 3983 8278 4017
rect 8312 3983 8354 4017
rect 8262 3948 8354 3983
rect 8262 3914 8278 3948
rect 8312 3914 8354 3948
rect 8262 3879 8354 3914
rect 8262 3845 8278 3879
rect 8312 3845 8354 3879
rect 8262 3809 8354 3845
rect 8262 3775 8278 3809
rect 8312 3775 8354 3809
rect 8262 3739 8354 3775
rect 8262 3705 8278 3739
rect 8312 3705 8354 3739
rect 8262 3669 8354 3705
rect 8262 3635 8278 3669
rect 8312 3635 8354 3669
rect 8262 3599 8354 3635
rect 8262 3565 8278 3599
rect 8312 3565 8354 3599
rect 8262 3529 8354 3565
rect 8262 3495 8278 3529
rect 8312 3495 8354 3529
rect 8262 3459 8354 3495
rect 8262 3425 8278 3459
rect 8312 3425 8354 3459
rect 8262 3389 8354 3425
rect 8262 3355 8278 3389
rect 8312 3355 8354 3389
rect 8262 3319 8354 3355
rect 8262 3285 8278 3319
rect 8312 3285 8354 3319
rect 8262 3256 8354 3285
rect 8438 3256 8498 4056
rect 8582 4013 8680 4056
rect 8582 3979 8630 4013
rect 8664 3979 8680 4013
rect 8582 3945 8680 3979
rect 8582 3911 8630 3945
rect 8664 3911 8680 3945
rect 8582 3877 8680 3911
rect 8582 3843 8630 3877
rect 8664 3843 8680 3877
rect 8582 3809 8680 3843
rect 8582 3775 8630 3809
rect 8664 3775 8680 3809
rect 8582 3741 8680 3775
rect 8582 3707 8630 3741
rect 8664 3707 8680 3741
rect 8582 3673 8680 3707
rect 8582 3639 8630 3673
rect 8664 3639 8680 3673
rect 8582 3605 8680 3639
rect 8582 3571 8630 3605
rect 8664 3571 8680 3605
rect 8582 3537 8680 3571
rect 8582 3503 8630 3537
rect 8664 3503 8680 3537
rect 8582 3469 8680 3503
rect 8582 3435 8630 3469
rect 8664 3435 8680 3469
rect 8582 3401 8680 3435
rect 8582 3367 8630 3401
rect 8664 3367 8680 3401
rect 8582 3333 8680 3367
rect 8582 3299 8630 3333
rect 8664 3299 8680 3333
rect 8582 3256 8680 3299
rect 11062 4239 11862 4271
rect 12039 4220 12137 4236
rect 12039 4186 12055 4220
rect 12089 4186 12137 4220
rect 11062 4107 11862 4155
rect 11062 4073 11078 4107
rect 11112 4073 11152 4107
rect 11186 4073 11226 4107
rect 11260 4073 11300 4107
rect 11334 4073 11374 4107
rect 11408 4073 11447 4107
rect 11481 4073 11520 4107
rect 11554 4073 11593 4107
rect 11627 4073 11666 4107
rect 11700 4073 11739 4107
rect 11773 4073 11812 4107
rect 11846 4073 11862 4107
rect 11062 4025 11862 4073
rect 12039 4148 12137 4186
rect 12039 4114 12055 4148
rect 12089 4114 12137 4148
rect 12039 4076 12137 4114
rect 12039 4042 12055 4076
rect 12089 4042 12137 4076
rect 12039 4036 12137 4042
rect 12221 4036 12253 4236
rect 12039 4003 12105 4036
rect 12039 3969 12055 4003
rect 12089 3980 12105 4003
rect 12089 3969 12137 3980
rect 11062 3909 11862 3941
rect 12039 3930 12137 3969
rect 12039 3896 12055 3930
rect 12089 3896 12137 3930
rect 11062 3831 11862 3863
rect 12039 3857 12137 3896
rect 12039 3823 12055 3857
rect 12089 3823 12137 3857
rect 12039 3780 12137 3823
rect 12221 3780 12253 3980
rect 9190 3686 9290 3718
rect 9346 3686 9446 3718
rect 9502 3686 9602 3718
rect 9190 3670 9602 3686
rect 9190 3636 9206 3670
rect 9240 3636 9276 3670
rect 9310 3636 9345 3670
rect 9379 3636 9414 3670
rect 9448 3636 9483 3670
rect 9517 3636 9552 3670
rect 9586 3636 9602 3670
rect 9190 3620 9602 3636
rect 9782 3686 9882 3718
rect 9938 3686 10038 3718
rect 10094 3686 10194 3718
rect 10250 3686 10350 3718
rect 9782 3670 10350 3686
rect 9782 3636 9798 3670
rect 9832 3636 9869 3670
rect 9903 3636 9940 3670
rect 9974 3636 10012 3670
rect 10046 3636 10084 3670
rect 10118 3636 10156 3670
rect 10190 3636 10228 3670
rect 10262 3636 10300 3670
rect 10334 3636 10350 3670
rect 9782 3620 10350 3636
rect 10530 3669 10630 3718
rect 10530 3635 10580 3669
rect 10614 3635 10630 3669
rect 10530 3601 10630 3635
rect 10530 3567 10580 3601
rect 10614 3567 10630 3601
rect 9815 3538 9935 3564
rect 9991 3538 10111 3564
rect 10195 3538 10315 3564
rect 10530 3551 10630 3567
rect 10686 3669 10786 3718
rect 10686 3635 10719 3669
rect 10753 3635 10786 3669
rect 10686 3601 10786 3635
rect 11062 3693 11862 3747
rect 11062 3659 11078 3693
rect 11112 3659 11151 3693
rect 11185 3659 11224 3693
rect 11258 3659 11297 3693
rect 11331 3659 11370 3693
rect 11404 3659 11443 3693
rect 11477 3659 11516 3693
rect 11550 3659 11590 3693
rect 11624 3659 11664 3693
rect 11698 3659 11738 3693
rect 11772 3659 11812 3693
rect 11846 3659 11862 3693
rect 11062 3605 11862 3659
rect 10686 3567 10719 3601
rect 10753 3567 10786 3601
rect 10686 3551 10786 3567
rect 1159 3155 1433 3177
rect 1159 3121 1179 3155
rect 1213 3121 1247 3155
rect 1281 3121 1315 3155
rect 1349 3121 1383 3155
rect 1417 3121 1433 3155
rect 7513 3160 7861 3182
rect 1159 3105 1433 3121
rect 1737 3109 3337 3135
rect 7513 3126 7675 3160
rect 7709 3126 7743 3160
rect 7777 3126 7811 3160
rect 7845 3126 7861 3160
rect 7513 3110 7861 3126
rect -145 3013 -25 3039
rect 7587 3052 7721 3110
rect 1737 2977 3337 3025
rect 1737 2943 1767 2977
rect 1801 2943 1835 2977
rect 1869 2943 1903 2977
rect 1937 2943 1971 2977
rect 2005 2943 2039 2977
rect 2073 2943 2107 2977
rect 2141 2943 2175 2977
rect 2209 2943 2243 2977
rect 2277 2943 2311 2977
rect 2345 2943 2379 2977
rect 2413 2943 2447 2977
rect 2481 2943 2515 2977
rect 2549 2943 2583 2977
rect 2617 2943 2651 2977
rect 2685 2943 2719 2977
rect 2753 2943 2787 2977
rect 2821 2943 2855 2977
rect 2889 2943 2923 2977
rect 2957 2943 2991 2977
rect 3025 2943 3059 2977
rect 3093 2943 3127 2977
rect 3161 2943 3195 2977
rect 3229 2943 3263 2977
rect 3297 2943 3337 2977
rect 7587 3018 7603 3052
rect 7637 3018 7671 3052
rect 7705 3018 7721 3052
rect 7587 2996 7721 3018
rect 7925 3052 8059 3068
rect 7925 3018 7941 3052
rect 7975 3018 8009 3052
rect 8043 3018 8059 3052
rect 7925 2996 8059 3018
rect 8277 3052 8411 3068
rect 8277 3018 8293 3052
rect 8327 3018 8361 3052
rect 8395 3018 8411 3052
rect 8277 2996 8411 3018
rect 7587 2970 7707 2996
rect 7763 2970 7883 2996
rect 7939 2970 8059 2996
rect 8115 2970 8235 2996
rect 8291 2970 8411 2996
rect 8467 3052 9435 3068
rect 8467 3018 8628 3052
rect 8662 3018 8696 3052
rect 8730 3018 8764 3052
rect 8798 3018 8832 3052
rect 8866 3018 8900 3052
rect 8934 3018 8968 3052
rect 9002 3018 9036 3052
rect 9070 3018 9104 3052
rect 9138 3018 9172 3052
rect 9206 3018 9240 3052
rect 9274 3018 9308 3052
rect 9342 3018 9376 3052
rect 9410 3018 9435 3052
rect 8467 2996 9435 3018
rect 8467 2970 8667 2996
rect 8723 2970 8923 2996
rect 8979 2970 9179 2996
rect 9235 2970 9435 2996
rect 1737 2927 3337 2943
rect -425 2881 -325 2907
rect 12039 3539 12137 3600
rect 11062 3472 11862 3521
rect 11062 3438 11088 3472
rect 11122 3438 11157 3472
rect 11191 3438 11226 3472
rect 11260 3438 11294 3472
rect 11328 3438 11362 3472
rect 11396 3438 11430 3472
rect 11464 3438 11498 3472
rect 11532 3438 11566 3472
rect 11600 3438 11634 3472
rect 11668 3438 11702 3472
rect 11736 3438 11770 3472
rect 11804 3438 11862 3472
rect 11062 3389 11862 3438
rect 12039 3505 12055 3539
rect 12089 3505 12137 3539
rect 12039 3454 12137 3505
rect 12039 3420 12055 3454
rect 12089 3420 12137 3454
rect 12039 3400 12137 3420
rect 12221 3400 12253 3600
rect 11062 3273 11862 3305
rect 10881 3209 11025 3225
rect 10881 3175 10897 3209
rect 10931 3175 10975 3209
rect 11009 3175 11025 3209
rect 10881 3159 11025 3175
rect 10905 3127 11025 3159
rect 11081 3209 11377 3225
rect 11081 3175 11097 3209
rect 11131 3175 11174 3209
rect 11208 3175 11251 3209
rect 11285 3175 11327 3209
rect 11361 3175 11377 3209
rect 11081 3159 11377 3175
rect 11081 3127 11201 3159
rect 11257 3127 11377 3159
rect 11433 3209 11729 3273
rect 11433 3175 11449 3209
rect 11483 3175 11526 3209
rect 11560 3175 11603 3209
rect 11637 3175 11679 3209
rect 11713 3175 11729 3209
rect 11433 3159 11729 3175
rect 11433 3127 11553 3159
rect 11609 3127 11729 3159
rect 11785 3209 12081 3225
rect 11785 3175 11801 3209
rect 11835 3175 11877 3209
rect 11911 3175 11954 3209
rect 11988 3175 12031 3209
rect 12065 3175 12081 3209
rect 11785 3159 12081 3175
rect 11785 3127 11905 3159
rect 11961 3127 12081 3159
rect 9815 2890 9935 2938
rect 9815 2856 9858 2890
rect 9892 2856 9935 2890
rect 9815 2822 9935 2856
rect 9815 2788 9858 2822
rect 9892 2788 9935 2822
rect 7587 2744 7707 2770
rect 7763 2744 7883 2770
rect 7939 2744 8059 2770
rect 8115 2744 8235 2770
rect 8291 2744 8411 2770
rect 8467 2744 8667 2770
rect -408 2669 -288 2695
rect -232 2669 -112 2695
rect -56 2669 64 2695
rect 7760 2722 7894 2744
rect 7760 2688 7776 2722
rect 7810 2688 7844 2722
rect 7878 2688 7894 2722
rect 7760 2672 7894 2688
rect 8112 2722 8246 2744
rect 8112 2688 8128 2722
rect 8162 2688 8196 2722
rect 8230 2688 8246 2722
rect 8723 2734 8923 2770
rect 8979 2744 9179 2770
rect 9235 2744 9435 2770
rect 8723 2708 8843 2734
rect 8112 2672 8246 2688
rect 7512 2597 7584 2611
rect 7512 2595 7610 2597
rect 7512 2561 7528 2595
rect 7562 2561 7610 2595
rect 7512 2527 7610 2561
rect 7512 2493 7528 2527
rect 7562 2493 7610 2527
rect 7512 2477 7610 2493
rect 8610 2477 8636 2597
rect -408 2401 -288 2469
rect -232 2401 -112 2469
rect -56 2401 64 2469
rect 7599 2386 7743 2402
rect 7599 2352 7619 2386
rect 7653 2352 7687 2386
rect 7721 2352 7743 2386
rect 7599 2333 7743 2352
rect 7623 2307 7743 2333
rect 7799 2386 7941 2402
rect 7799 2352 7819 2386
rect 7853 2352 7887 2386
rect 7921 2352 7941 2386
rect 7799 2333 7941 2352
rect 7799 2307 7919 2333
rect -408 2153 -288 2201
rect -408 2119 -366 2153
rect -332 2119 -288 2153
rect -408 2085 -288 2119
rect -408 2051 -366 2085
rect -332 2051 -288 2085
rect -408 2003 -288 2051
rect -232 2153 -112 2201
rect -232 2119 -186 2153
rect -152 2119 -112 2153
rect -232 2085 -112 2119
rect -232 2051 -186 2085
rect -152 2051 -112 2085
rect -232 2003 -112 2051
rect -56 2153 64 2201
rect -56 2119 -15 2153
rect 19 2119 64 2153
rect -56 2085 64 2119
rect -56 2051 -15 2085
rect 19 2051 64 2085
rect -56 2003 64 2051
rect -408 1837 -288 1863
rect -232 1837 -112 1863
rect -56 1837 64 1863
rect 9815 2678 9935 2788
rect 9991 2890 10111 2938
rect 9991 2856 10034 2890
rect 10068 2856 10111 2890
rect 9991 2822 10111 2856
rect 9991 2788 10034 2822
rect 10068 2788 10111 2822
rect 9991 2678 10111 2788
rect 10195 2890 10315 2938
rect 10195 2856 10211 2890
rect 10245 2856 10315 2890
rect 10195 2822 10315 2856
rect 10195 2788 10211 2822
rect 10245 2788 10315 2822
rect 10195 2678 10315 2788
rect 9582 2613 9648 2629
rect 9582 2597 9598 2613
rect 8930 2497 8956 2597
rect 9556 2579 9598 2597
rect 9632 2579 9648 2613
rect 9556 2545 9648 2579
rect 9556 2511 9598 2545
rect 9632 2511 9648 2545
rect 9556 2497 9648 2511
rect 9582 2495 9648 2497
rect 10905 2495 11025 2527
rect 11081 2495 11201 2527
rect 11257 2495 11377 2527
rect 11433 2495 11553 2527
rect 11609 2495 11729 2527
rect 11785 2495 11905 2527
rect 11961 2495 12081 2527
rect 9815 2452 9935 2478
rect 9991 2452 10111 2478
rect 10195 2452 10315 2478
rect 8998 2390 9142 2410
rect 8998 2356 9018 2390
rect 9052 2356 9086 2390
rect 9120 2356 9142 2390
rect 8998 2334 9142 2356
rect 9022 2308 9142 2334
rect 9198 2390 9340 2410
rect 9198 2356 9218 2390
rect 9252 2356 9286 2390
rect 9320 2356 9340 2390
rect 9198 2334 9340 2356
rect 9709 2390 10005 2410
rect 9709 2356 9738 2390
rect 9772 2356 9806 2390
rect 9840 2356 9874 2390
rect 9908 2356 9942 2390
rect 9976 2356 10005 2390
rect 9709 2334 10005 2356
rect 9198 2308 9318 2334
rect 9709 2308 9829 2334
rect 9885 2308 10005 2334
rect 10061 2390 10357 2410
rect 10061 2356 10090 2390
rect 10124 2356 10158 2390
rect 10192 2356 10226 2390
rect 10260 2356 10294 2390
rect 10328 2356 10357 2390
rect 10829 2372 10949 2404
rect 11005 2372 11125 2404
rect 11181 2372 11301 2404
rect 11357 2372 11477 2404
rect 11533 2372 11653 2404
rect 11709 2372 11829 2404
rect 11885 2372 12005 2404
rect 10061 2334 10357 2356
rect 10061 2308 10181 2334
rect 10237 2308 10357 2334
rect 10829 1740 10949 1772
rect 11005 1740 11125 1772
rect 11181 1740 11301 1772
rect 11357 1740 11477 1772
rect 11533 1740 11653 1772
rect 10829 1724 11653 1740
rect 7623 1681 7743 1707
rect 7799 1681 7919 1707
rect 8723 1682 8843 1708
rect 9022 1682 9142 1708
rect 9198 1682 9318 1708
rect 9709 1682 9829 1708
rect 9885 1682 10005 1708
rect 7406 1636 7743 1681
rect 7406 1602 7426 1636
rect 7460 1602 7494 1636
rect 7528 1602 7743 1636
rect 7406 1570 7743 1602
rect 7819 1640 7964 1681
rect 7819 1606 7842 1640
rect 7876 1606 7910 1640
rect 7944 1606 7964 1640
rect 8723 1660 8857 1682
rect 8723 1626 8739 1660
rect 8773 1626 8807 1660
rect 8841 1626 8857 1660
rect 8723 1610 8857 1626
rect 8929 1659 9142 1682
rect 8929 1625 8952 1659
rect 8986 1625 9020 1659
rect 9054 1625 9088 1659
rect 9122 1625 9142 1659
rect 7819 1570 7964 1606
rect 8929 1570 9142 1625
rect 9241 1659 9558 1682
rect 9241 1625 9436 1659
rect 9470 1625 9504 1659
rect 9538 1625 9558 1659
rect 9241 1570 9558 1625
rect 9709 1659 10005 1682
rect 9709 1625 9738 1659
rect 9772 1625 9806 1659
rect 9840 1625 9874 1659
rect 9908 1625 9942 1659
rect 9976 1625 10005 1659
rect 9709 1570 10005 1625
rect 10061 1682 10181 1708
rect 10237 1682 10357 1708
rect 10829 1690 10845 1724
rect 10879 1690 10914 1724
rect 10948 1690 10983 1724
rect 11017 1690 11052 1724
rect 11086 1690 11121 1724
rect 11155 1690 11190 1724
rect 11224 1690 11259 1724
rect 11293 1690 11328 1724
rect 11362 1690 11397 1724
rect 11431 1690 11466 1724
rect 11500 1690 11535 1724
rect 11569 1690 11603 1724
rect 11637 1690 11653 1724
rect 10061 1666 10411 1682
rect 10829 1674 11653 1690
rect 11709 1740 11829 1772
rect 11885 1740 12005 1772
rect 11709 1724 12005 1740
rect 11709 1690 11725 1724
rect 11759 1690 11802 1724
rect 11836 1690 11879 1724
rect 11913 1690 11955 1724
rect 11989 1690 12005 1724
rect 11709 1674 12005 1690
rect 10061 1632 10152 1666
rect 10186 1662 10411 1666
rect 10186 1632 10289 1662
rect 10061 1628 10289 1632
rect 10323 1628 10357 1662
rect 10391 1628 10411 1662
rect 10061 1614 10411 1628
rect 10269 1570 10411 1614
rect 10929 1614 11029 1630
rect 10929 1580 10959 1614
rect 10993 1580 11029 1614
rect 7467 1544 7587 1570
rect 7643 1544 7763 1570
rect 7819 1544 7939 1570
rect 8929 1544 9029 1570
rect 9085 1544 9185 1570
rect 9241 1544 9341 1570
rect 9397 1544 9497 1570
rect 9801 1544 9901 1570
rect 9957 1544 10057 1570
rect 10113 1544 10213 1570
rect 10269 1544 10369 1570
rect 10617 1537 10873 1553
rect 10617 1503 10633 1537
rect 10667 1503 10728 1537
rect 10762 1503 10823 1537
rect 10857 1503 10873 1537
rect 10617 1487 10873 1503
rect 10617 1455 10717 1487
rect 10773 1455 10873 1487
rect 10929 1546 11029 1580
rect 10929 1512 10959 1546
rect 10993 1512 11029 1546
rect 10929 1455 11029 1512
rect 11085 1614 11185 1630
rect 11085 1580 11118 1614
rect 11152 1580 11185 1614
rect 11085 1546 11185 1580
rect 11085 1512 11118 1546
rect 11152 1512 11185 1546
rect 11085 1455 11185 1512
rect 11414 1431 12214 1447
rect 11414 1397 11430 1431
rect 11464 1397 11499 1431
rect 11533 1397 11568 1431
rect 11602 1397 11637 1431
rect 11671 1397 11706 1431
rect 11740 1397 11775 1431
rect 11809 1397 11844 1431
rect 11878 1397 11913 1431
rect 11947 1397 11982 1431
rect 12016 1397 12051 1431
rect 12085 1397 12120 1431
rect 12154 1397 12214 1431
rect 11414 1349 12214 1397
rect 11414 1217 12214 1265
rect 11414 1183 11430 1217
rect 11464 1183 11503 1217
rect 11537 1183 11576 1217
rect 11610 1183 11649 1217
rect 11683 1183 11722 1217
rect 11756 1183 11795 1217
rect 11829 1183 11868 1217
rect 11902 1183 11942 1217
rect 11976 1183 12016 1217
rect 12050 1183 12090 1217
rect 12124 1183 12164 1217
rect 12198 1183 12214 1217
rect 11414 1167 12214 1183
rect 10617 1123 10717 1155
rect 10773 1123 10873 1155
rect 10929 1123 11029 1155
rect 11085 1123 11185 1155
rect 11814 1115 12214 1167
rect 11814 1081 11843 1115
rect 11877 1081 11922 1115
rect 11956 1081 12000 1115
rect 12034 1081 12214 1115
rect 8929 918 9029 944
rect 9085 918 9185 944
rect 8929 896 9185 918
rect 8929 862 8979 896
rect 9013 862 9047 896
rect 9081 862 9115 896
rect 9149 862 9185 896
rect 8929 846 9185 862
rect 9241 918 9341 944
rect 9397 918 9497 944
rect 9241 896 9497 918
rect 9241 862 9272 896
rect 9306 862 9340 896
rect 9374 862 9408 896
rect 9442 862 9497 896
rect 9241 846 9497 862
rect 9801 918 9901 944
rect 9957 918 10057 944
rect 10113 918 10213 944
rect 10269 918 10369 944
rect 10902 1009 11758 1025
rect 10902 975 10943 1009
rect 10977 975 11012 1009
rect 11046 975 11081 1009
rect 11115 975 11150 1009
rect 11184 975 11219 1009
rect 11253 975 11288 1009
rect 11322 975 11358 1009
rect 11392 975 11428 1009
rect 11462 975 11498 1009
rect 11532 975 11568 1009
rect 11602 975 11638 1009
rect 11672 975 11708 1009
rect 11742 975 11758 1009
rect 10902 959 11758 975
rect 10902 927 11302 959
rect 11358 927 11758 959
rect 11814 1009 12214 1081
rect 11814 975 11830 1009
rect 11864 975 11914 1009
rect 11948 975 11998 1009
rect 12032 975 12081 1009
rect 12115 975 12164 1009
rect 12198 975 12214 1009
rect 11814 927 12214 975
rect 9801 896 10213 918
rect 9801 862 9855 896
rect 9889 862 9923 896
rect 9957 862 9991 896
rect 10025 862 10059 896
rect 10093 862 10127 896
rect 10161 862 10213 896
rect 9801 846 10213 862
rect 10902 811 11302 843
rect 11358 811 11758 843
rect 11814 811 12214 843
rect 10451 725 10707 741
rect 10451 691 10467 725
rect 10501 691 10562 725
rect 10596 691 10657 725
rect 10691 691 10707 725
rect 10451 675 10707 691
rect 10919 725 11053 741
rect 10919 691 10935 725
rect 10969 691 11003 725
rect 11037 691 11053 725
rect 10919 675 11053 691
rect 11108 725 11242 741
rect 11108 691 11124 725
rect 11158 691 11192 725
rect 11226 691 11242 725
rect 11108 675 11242 691
rect 11389 725 11801 741
rect 11389 691 11405 725
rect 11439 691 11475 725
rect 11509 691 11544 725
rect 11578 691 11613 725
rect 11647 691 11682 725
rect 11716 691 11751 725
rect 11785 691 11801 725
rect 11389 675 11801 691
rect 10451 643 10551 675
rect 10607 643 10707 675
rect 10953 643 11053 675
rect 11109 643 11209 675
rect 11389 643 11489 675
rect 11545 643 11645 675
rect 7467 518 7587 544
rect 7643 518 7763 544
rect 7819 518 7939 544
rect 7467 496 7763 518
rect 7467 462 7496 496
rect 7530 462 7564 496
rect 7598 462 7632 496
rect 7666 462 7700 496
rect 7734 462 7763 496
rect 7467 442 7763 462
rect 10953 527 11053 559
rect 11109 527 11209 559
rect 11389 527 11489 559
rect 11545 527 11645 559
rect 10451 411 10551 443
rect 10607 411 10707 443
<< polycont >>
rect 13351 4563 13385 4597
rect 13419 4563 13453 4597
rect -366 4283 -332 4317
rect -366 4215 -332 4249
rect -186 4283 -152 4317
rect -186 4215 -152 4249
rect -15 4283 19 4317
rect -15 4215 19 4249
rect 4505 4301 4539 4335
rect 4573 4301 4607 4335
rect 4641 4301 4675 4335
rect 4709 4301 4743 4335
rect 4777 4301 4811 4335
rect 4845 4301 4879 4335
rect 4913 4301 4947 4335
rect 4981 4301 5015 4335
rect 5049 4301 5083 4335
rect 5117 4301 5151 4335
rect 5185 4301 5219 4335
rect 5253 4301 5287 4335
rect 5321 4301 5355 4335
rect 5389 4301 5423 4335
rect 5457 4301 5491 4335
rect 5525 4301 5559 4335
rect 5593 4301 5627 4335
rect 1609 4251 1643 4285
rect 1677 4251 1711 4285
rect 1745 4251 1779 4285
rect 1813 4251 1847 4285
rect 1881 4251 1915 4285
rect 1949 4251 1983 4285
rect 2017 4251 2051 4285
rect 2085 4251 2119 4285
rect 2233 4251 2267 4285
rect 2301 4251 2335 4285
rect 2369 4251 2403 4285
rect 2437 4251 2471 4285
rect 2505 4251 2539 4285
rect 2573 4251 2607 4285
rect 2641 4251 2675 4285
rect 2709 4251 2743 4285
rect 3061 4251 3095 4285
rect 3129 4251 3163 4285
rect 3197 4251 3231 4285
rect 3265 4251 3299 4285
rect 3333 4251 3367 4285
rect 3401 4251 3435 4285
rect 3469 4251 3503 4285
rect 3537 4251 3571 4285
rect 3605 4251 3639 4285
rect 3673 4251 3707 4285
rect 3741 4251 3775 4285
rect 3809 4251 3843 4285
rect 3877 4251 3911 4285
rect 3945 4251 3979 4285
rect 4013 4251 4047 4285
rect 4081 4251 4115 4285
rect 4149 4251 4183 4285
rect -394 3666 -360 3700
rect -394 3598 -360 3632
rect -101 3623 -67 3657
rect -101 3555 -67 3589
rect 5950 4251 5984 4285
rect 6018 4251 6052 4285
rect 6086 4251 6120 4285
rect 6154 4251 6188 4285
rect 6222 4251 6256 4285
rect 6290 4251 6324 4285
rect 6358 4251 6392 4285
rect 6426 4251 6460 4285
rect 6494 4251 6528 4285
rect 6562 4251 6596 4285
rect 6630 4251 6664 4285
rect 6698 4251 6732 4285
rect 6766 4251 6800 4285
rect 6834 4251 6868 4285
rect 6902 4251 6936 4285
rect 6970 4251 7004 4285
rect 7038 4251 7072 4285
rect 7177 4251 7211 4285
rect 7245 4251 7279 4285
rect 7478 4251 7512 4285
rect 7546 4251 7580 4285
rect 7830 4251 7864 4285
rect 7898 4251 7932 4285
rect 7654 3492 7688 3526
rect 7722 3492 7756 3526
rect 7944 3476 7978 3510
rect 7944 3408 7978 3442
rect 7944 3340 7978 3374
rect 7944 3272 7978 3306
rect 8278 3983 8312 4017
rect 8278 3914 8312 3948
rect 8278 3845 8312 3879
rect 8278 3775 8312 3809
rect 8278 3705 8312 3739
rect 8278 3635 8312 3669
rect 8278 3565 8312 3599
rect 8278 3495 8312 3529
rect 8278 3425 8312 3459
rect 8278 3355 8312 3389
rect 8278 3285 8312 3319
rect 8630 3979 8664 4013
rect 8630 3911 8664 3945
rect 8630 3843 8664 3877
rect 8630 3775 8664 3809
rect 8630 3707 8664 3741
rect 8630 3639 8664 3673
rect 8630 3571 8664 3605
rect 8630 3503 8664 3537
rect 8630 3435 8664 3469
rect 8630 3367 8664 3401
rect 8630 3299 8664 3333
rect 12055 4186 12089 4220
rect 11078 4073 11112 4107
rect 11152 4073 11186 4107
rect 11226 4073 11260 4107
rect 11300 4073 11334 4107
rect 11374 4073 11408 4107
rect 11447 4073 11481 4107
rect 11520 4073 11554 4107
rect 11593 4073 11627 4107
rect 11666 4073 11700 4107
rect 11739 4073 11773 4107
rect 11812 4073 11846 4107
rect 12055 4114 12089 4148
rect 12055 4042 12089 4076
rect 12055 3969 12089 4003
rect 12055 3896 12089 3930
rect 12055 3823 12089 3857
rect 9206 3636 9240 3670
rect 9276 3636 9310 3670
rect 9345 3636 9379 3670
rect 9414 3636 9448 3670
rect 9483 3636 9517 3670
rect 9552 3636 9586 3670
rect 9798 3636 9832 3670
rect 9869 3636 9903 3670
rect 9940 3636 9974 3670
rect 10012 3636 10046 3670
rect 10084 3636 10118 3670
rect 10156 3636 10190 3670
rect 10228 3636 10262 3670
rect 10300 3636 10334 3670
rect 10580 3635 10614 3669
rect 10580 3567 10614 3601
rect 10719 3635 10753 3669
rect 11078 3659 11112 3693
rect 11151 3659 11185 3693
rect 11224 3659 11258 3693
rect 11297 3659 11331 3693
rect 11370 3659 11404 3693
rect 11443 3659 11477 3693
rect 11516 3659 11550 3693
rect 11590 3659 11624 3693
rect 11664 3659 11698 3693
rect 11738 3659 11772 3693
rect 11812 3659 11846 3693
rect 10719 3567 10753 3601
rect 1179 3121 1213 3155
rect 1247 3121 1281 3155
rect 1315 3121 1349 3155
rect 1383 3121 1417 3155
rect 7675 3126 7709 3160
rect 7743 3126 7777 3160
rect 7811 3126 7845 3160
rect 1767 2943 1801 2977
rect 1835 2943 1869 2977
rect 1903 2943 1937 2977
rect 1971 2943 2005 2977
rect 2039 2943 2073 2977
rect 2107 2943 2141 2977
rect 2175 2943 2209 2977
rect 2243 2943 2277 2977
rect 2311 2943 2345 2977
rect 2379 2943 2413 2977
rect 2447 2943 2481 2977
rect 2515 2943 2549 2977
rect 2583 2943 2617 2977
rect 2651 2943 2685 2977
rect 2719 2943 2753 2977
rect 2787 2943 2821 2977
rect 2855 2943 2889 2977
rect 2923 2943 2957 2977
rect 2991 2943 3025 2977
rect 3059 2943 3093 2977
rect 3127 2943 3161 2977
rect 3195 2943 3229 2977
rect 3263 2943 3297 2977
rect 7603 3018 7637 3052
rect 7671 3018 7705 3052
rect 7941 3018 7975 3052
rect 8009 3018 8043 3052
rect 8293 3018 8327 3052
rect 8361 3018 8395 3052
rect 8628 3018 8662 3052
rect 8696 3018 8730 3052
rect 8764 3018 8798 3052
rect 8832 3018 8866 3052
rect 8900 3018 8934 3052
rect 8968 3018 9002 3052
rect 9036 3018 9070 3052
rect 9104 3018 9138 3052
rect 9172 3018 9206 3052
rect 9240 3018 9274 3052
rect 9308 3018 9342 3052
rect 9376 3018 9410 3052
rect 11088 3438 11122 3472
rect 11157 3438 11191 3472
rect 11226 3438 11260 3472
rect 11294 3438 11328 3472
rect 11362 3438 11396 3472
rect 11430 3438 11464 3472
rect 11498 3438 11532 3472
rect 11566 3438 11600 3472
rect 11634 3438 11668 3472
rect 11702 3438 11736 3472
rect 11770 3438 11804 3472
rect 12055 3505 12089 3539
rect 12055 3420 12089 3454
rect 10897 3175 10931 3209
rect 10975 3175 11009 3209
rect 11097 3175 11131 3209
rect 11174 3175 11208 3209
rect 11251 3175 11285 3209
rect 11327 3175 11361 3209
rect 11449 3175 11483 3209
rect 11526 3175 11560 3209
rect 11603 3175 11637 3209
rect 11679 3175 11713 3209
rect 11801 3175 11835 3209
rect 11877 3175 11911 3209
rect 11954 3175 11988 3209
rect 12031 3175 12065 3209
rect 9858 2856 9892 2890
rect 9858 2788 9892 2822
rect 7776 2688 7810 2722
rect 7844 2688 7878 2722
rect 8128 2688 8162 2722
rect 8196 2688 8230 2722
rect 7528 2561 7562 2595
rect 7528 2493 7562 2527
rect 7619 2352 7653 2386
rect 7687 2352 7721 2386
rect 7819 2352 7853 2386
rect 7887 2352 7921 2386
rect -366 2119 -332 2153
rect -366 2051 -332 2085
rect -186 2119 -152 2153
rect -186 2051 -152 2085
rect -15 2119 19 2153
rect -15 2051 19 2085
rect 10034 2856 10068 2890
rect 10034 2788 10068 2822
rect 10211 2856 10245 2890
rect 10211 2788 10245 2822
rect 9598 2579 9632 2613
rect 9598 2511 9632 2545
rect 9018 2356 9052 2390
rect 9086 2356 9120 2390
rect 9218 2356 9252 2390
rect 9286 2356 9320 2390
rect 9738 2356 9772 2390
rect 9806 2356 9840 2390
rect 9874 2356 9908 2390
rect 9942 2356 9976 2390
rect 10090 2356 10124 2390
rect 10158 2356 10192 2390
rect 10226 2356 10260 2390
rect 10294 2356 10328 2390
rect 7426 1602 7460 1636
rect 7494 1602 7528 1636
rect 7842 1606 7876 1640
rect 7910 1606 7944 1640
rect 8739 1626 8773 1660
rect 8807 1626 8841 1660
rect 8952 1625 8986 1659
rect 9020 1625 9054 1659
rect 9088 1625 9122 1659
rect 9436 1625 9470 1659
rect 9504 1625 9538 1659
rect 9738 1625 9772 1659
rect 9806 1625 9840 1659
rect 9874 1625 9908 1659
rect 9942 1625 9976 1659
rect 10845 1690 10879 1724
rect 10914 1690 10948 1724
rect 10983 1690 11017 1724
rect 11052 1690 11086 1724
rect 11121 1690 11155 1724
rect 11190 1690 11224 1724
rect 11259 1690 11293 1724
rect 11328 1690 11362 1724
rect 11397 1690 11431 1724
rect 11466 1690 11500 1724
rect 11535 1690 11569 1724
rect 11603 1690 11637 1724
rect 11725 1690 11759 1724
rect 11802 1690 11836 1724
rect 11879 1690 11913 1724
rect 11955 1690 11989 1724
rect 10152 1632 10186 1666
rect 10289 1628 10323 1662
rect 10357 1628 10391 1662
rect 10959 1580 10993 1614
rect 10633 1503 10667 1537
rect 10728 1503 10762 1537
rect 10823 1503 10857 1537
rect 10959 1512 10993 1546
rect 11118 1580 11152 1614
rect 11118 1512 11152 1546
rect 11430 1397 11464 1431
rect 11499 1397 11533 1431
rect 11568 1397 11602 1431
rect 11637 1397 11671 1431
rect 11706 1397 11740 1431
rect 11775 1397 11809 1431
rect 11844 1397 11878 1431
rect 11913 1397 11947 1431
rect 11982 1397 12016 1431
rect 12051 1397 12085 1431
rect 12120 1397 12154 1431
rect 11430 1183 11464 1217
rect 11503 1183 11537 1217
rect 11576 1183 11610 1217
rect 11649 1183 11683 1217
rect 11722 1183 11756 1217
rect 11795 1183 11829 1217
rect 11868 1183 11902 1217
rect 11942 1183 11976 1217
rect 12016 1183 12050 1217
rect 12090 1183 12124 1217
rect 12164 1183 12198 1217
rect 11843 1081 11877 1115
rect 11922 1081 11956 1115
rect 12000 1081 12034 1115
rect 8979 862 9013 896
rect 9047 862 9081 896
rect 9115 862 9149 896
rect 9272 862 9306 896
rect 9340 862 9374 896
rect 9408 862 9442 896
rect 10943 975 10977 1009
rect 11012 975 11046 1009
rect 11081 975 11115 1009
rect 11150 975 11184 1009
rect 11219 975 11253 1009
rect 11288 975 11322 1009
rect 11358 975 11392 1009
rect 11428 975 11462 1009
rect 11498 975 11532 1009
rect 11568 975 11602 1009
rect 11638 975 11672 1009
rect 11708 975 11742 1009
rect 11830 975 11864 1009
rect 11914 975 11948 1009
rect 11998 975 12032 1009
rect 12081 975 12115 1009
rect 12164 975 12198 1009
rect 9855 862 9889 896
rect 9923 862 9957 896
rect 9991 862 10025 896
rect 10059 862 10093 896
rect 10127 862 10161 896
rect 10467 691 10501 725
rect 10562 691 10596 725
rect 10657 691 10691 725
rect 10935 691 10969 725
rect 11003 691 11037 725
rect 11124 691 11158 725
rect 11192 691 11226 725
rect 11405 691 11439 725
rect 11475 691 11509 725
rect 11544 691 11578 725
rect 11613 691 11647 725
rect 11682 691 11716 725
rect 11751 691 11785 725
rect 7496 462 7530 496
rect 7564 462 7598 496
rect 7632 462 7666 496
rect 7700 462 7734 496
<< locali >>
rect 1508 6962 1546 6996
rect 12782 5876 13062 5915
rect -502 4907 -478 4941
rect -444 4907 -406 4941
rect -372 4939 -334 4941
rect -300 4939 -262 4941
rect -228 4939 -190 4941
rect -366 4907 -334 4939
rect -281 4907 -262 4939
rect -196 4907 -190 4939
rect -156 4939 -119 4941
rect -85 4939 -48 4941
rect -156 4907 -145 4939
rect -85 4907 -60 4939
rect -14 4907 23 4941
rect 57 4939 94 4941
rect 59 4907 94 4939
rect 128 4907 152 4941
rect -366 4905 -315 4907
rect -281 4905 -230 4907
rect -196 4905 -145 4907
rect -111 4905 -60 4907
rect -26 4905 25 4907
rect 12941 4898 13062 5876
rect 12941 4864 13028 4898
rect -453 4815 -419 4833
rect -453 4747 -419 4781
rect -453 4682 -419 4713
rect -277 4815 -243 4827
rect -277 4747 -243 4755
rect -430 4679 -392 4682
rect -419 4648 -392 4679
rect -277 4679 -243 4713
rect -453 4553 -419 4645
rect -453 4485 -419 4519
rect -453 4417 -419 4451
rect -453 4155 -419 4383
rect -277 4553 -243 4645
rect -277 4485 -243 4519
rect -101 4815 -67 4833
rect -101 4747 -67 4781
rect -101 4679 -67 4713
rect -101 4553 -67 4645
rect -101 4518 -67 4519
rect 75 4815 109 4827
rect 75 4747 109 4755
rect 75 4679 109 4713
rect 12941 4826 13062 4864
rect 12941 4792 13028 4826
rect 12941 4754 13062 4792
rect 12941 4720 13028 4754
rect 12941 4662 13062 4720
rect 75 4553 109 4645
rect 12392 4642 13062 4662
rect -134 4485 -96 4518
rect -134 4484 -101 4485
rect 75 4485 109 4519
rect 10793 4584 13062 4642
rect 13332 4597 13901 4644
rect 10793 4580 12400 4584
rect 10793 4546 10909 4580
rect 10943 4546 10980 4580
rect 11014 4546 11051 4580
rect 11085 4546 11122 4580
rect 11156 4546 11193 4580
rect 11227 4546 11264 4580
rect 11298 4546 11335 4580
rect 11369 4546 11406 4580
rect 11440 4546 11477 4580
rect 11511 4546 11548 4580
rect 11582 4546 11619 4580
rect 11653 4546 11690 4580
rect 11724 4546 11761 4580
rect 11795 4546 11832 4580
rect 11866 4546 11903 4580
rect 11937 4546 11974 4580
rect 12008 4546 12045 4580
rect 12079 4546 12116 4580
rect 12150 4546 12187 4580
rect 12221 4546 12258 4580
rect 12292 4546 12329 4580
rect 12363 4546 12400 4580
rect 13332 4563 13351 4597
rect 13385 4563 13419 4597
rect 13453 4563 13901 4597
rect 10793 4506 12400 4546
rect 10793 4499 10839 4506
rect 10873 4499 12400 4506
rect 10793 4493 10807 4499
rect -277 4417 -243 4451
rect -277 4367 -243 4383
rect -202 4403 -177 4414
rect -101 4417 -67 4451
rect -143 4403 -136 4414
rect -202 4365 -136 4403
rect -202 4331 -177 4365
rect -143 4331 -136 4365
rect -202 4317 -136 4331
rect -382 4283 -367 4317
rect -332 4283 -316 4317
rect -382 4249 -316 4283
rect -382 4245 -366 4249
rect -382 4215 -367 4245
rect -332 4215 -316 4249
rect -202 4283 -186 4317
rect -152 4283 -136 4317
rect -202 4249 -136 4283
rect -202 4215 -186 4249
rect -152 4215 -136 4249
rect -644 4108 -532 4115
rect -644 4074 -638 4108
rect -604 4091 -566 4108
rect -581 4074 -566 4091
rect -644 4057 -615 4074
rect -581 4057 -532 4074
rect -644 4031 -532 4057
rect -453 4087 -419 4121
rect -453 4037 -419 4053
rect -277 4155 -243 4171
rect -277 4110 -243 4121
rect -101 4144 -67 4383
rect 75 4417 109 4451
rect 75 4367 109 4383
rect 271 4465 10807 4493
rect 10873 4472 10879 4499
rect 10841 4465 10879 4472
rect 10913 4465 10951 4499
rect 10985 4465 11023 4499
rect 11057 4465 11095 4499
rect 11129 4465 11167 4499
rect 11201 4465 11239 4499
rect 11273 4465 11311 4499
rect 11345 4465 11383 4499
rect 11417 4465 11455 4499
rect 11489 4465 11527 4499
rect 11561 4465 11599 4499
rect 11633 4465 11671 4499
rect 11705 4465 11743 4499
rect 11777 4465 11815 4499
rect 11849 4465 11887 4499
rect 11921 4496 12400 4499
rect 11921 4465 12366 4496
rect 271 4460 10893 4465
rect 271 4426 409 4460
rect 443 4426 477 4460
rect 515 4426 545 4460
rect 587 4426 613 4460
rect 659 4426 681 4460
rect 731 4426 749 4460
rect 803 4426 817 4460
rect 875 4426 885 4460
rect 947 4426 953 4460
rect 1019 4426 1021 4460
rect 1055 4426 1057 4460
rect 1123 4426 1129 4460
rect 1191 4426 1201 4460
rect 1259 4426 1273 4460
rect 1327 4426 1345 4460
rect 1395 4426 1417 4460
rect 1463 4426 1489 4460
rect 1531 4426 1561 4460
rect 1599 4426 1633 4460
rect 1667 4426 1701 4460
rect 1739 4426 1769 4460
rect 1811 4426 1837 4460
rect 1883 4426 1905 4460
rect 1955 4426 1973 4460
rect 2027 4426 2041 4460
rect 2099 4426 2109 4460
rect 2171 4426 2177 4460
rect 2243 4426 2245 4460
rect 2279 4426 2281 4460
rect 2347 4426 2353 4460
rect 2415 4426 2425 4460
rect 2483 4426 2497 4460
rect 2551 4426 2569 4460
rect 2619 4426 2641 4460
rect 2687 4426 2713 4460
rect 2755 4426 2785 4460
rect 2823 4426 2857 4460
rect 2891 4426 2925 4460
rect 2963 4426 2993 4460
rect 3035 4426 3061 4460
rect 3107 4426 3129 4460
rect 3179 4426 3197 4460
rect 3251 4426 3265 4460
rect 3323 4426 3333 4460
rect 3395 4426 3401 4460
rect 3467 4426 3469 4460
rect 3503 4426 3505 4460
rect 3571 4426 3577 4460
rect 3639 4426 3649 4460
rect 3707 4426 3721 4460
rect 3775 4426 3793 4460
rect 3843 4426 3865 4460
rect 3911 4426 3937 4460
rect 3979 4426 4009 4460
rect 4047 4426 4081 4460
rect 4115 4426 4149 4460
rect 4187 4426 4217 4460
rect 4259 4426 4285 4460
rect 4331 4426 4353 4460
rect 4403 4426 4421 4460
rect 4475 4426 4489 4460
rect 4547 4426 4557 4460
rect 4619 4426 4625 4460
rect 4691 4426 4693 4460
rect 4727 4426 4729 4460
rect 4795 4426 4801 4460
rect 4863 4426 4873 4460
rect 4931 4426 4945 4460
rect 4999 4426 5017 4460
rect 5067 4426 5089 4460
rect 5135 4426 5161 4460
rect 5203 4426 5233 4460
rect 5271 4426 5305 4460
rect 5339 4426 5373 4460
rect 5411 4426 5441 4460
rect 5483 4426 5509 4460
rect 5555 4426 5577 4460
rect 5627 4426 5645 4460
rect 5699 4426 5713 4460
rect 5771 4426 5781 4460
rect 5843 4426 5849 4460
rect 5915 4426 5917 4460
rect 5951 4426 5953 4460
rect 6019 4426 6025 4460
rect 6087 4426 6097 4460
rect 6155 4426 6169 4460
rect 6223 4426 6241 4460
rect 6291 4426 6313 4460
rect 6359 4426 6385 4460
rect 6427 4426 6457 4460
rect 6495 4426 6529 4460
rect 6563 4426 6597 4460
rect 6635 4426 6665 4460
rect 6707 4426 6733 4460
rect 6779 4426 6801 4460
rect 6851 4426 6869 4460
rect 6923 4426 6937 4460
rect 6995 4426 7005 4460
rect 7067 4426 7073 4460
rect 7139 4426 7141 4460
rect 7175 4426 7177 4460
rect 7243 4426 7249 4460
rect 7311 4426 7321 4460
rect 7379 4426 7393 4460
rect 7447 4426 7465 4460
rect 7515 4426 7537 4460
rect 7583 4426 7609 4460
rect 7651 4426 7681 4460
rect 7719 4426 7753 4460
rect 7787 4426 7821 4460
rect 7859 4426 7889 4460
rect 7931 4426 7957 4460
rect 8003 4426 8025 4460
rect 8075 4426 8093 4460
rect 8147 4426 8161 4460
rect 8219 4426 8229 4460
rect 8291 4426 8297 4460
rect 8363 4426 8365 4460
rect 8399 4426 8401 4460
rect 8467 4426 8473 4460
rect 8535 4426 8545 4460
rect 8603 4426 8617 4460
rect 8671 4426 8689 4460
rect 8739 4426 8761 4460
rect 8807 4426 8833 4460
rect 8875 4426 8905 4460
rect 8943 4426 8977 4460
rect 9011 4426 9045 4460
rect 9083 4426 9113 4460
rect 9155 4426 9181 4460
rect 9227 4426 9249 4460
rect 9299 4426 9317 4460
rect 9371 4426 9385 4460
rect 9443 4426 9453 4460
rect 9515 4426 9521 4460
rect 9587 4426 9589 4460
rect 9623 4426 9625 4460
rect 9691 4426 9697 4460
rect 9759 4426 9769 4460
rect 9827 4426 9841 4460
rect 9895 4426 9913 4460
rect 9963 4426 9985 4460
rect 10031 4426 10057 4460
rect 10099 4426 10129 4460
rect 10167 4426 10201 4460
rect 10235 4426 10269 4460
rect 10307 4426 10337 4460
rect 10379 4426 10405 4460
rect 10451 4426 10473 4460
rect 10523 4426 10541 4460
rect 10595 4426 10609 4460
rect 10643 4431 10893 4460
rect 10643 4426 10760 4431
rect 271 4409 10760 4426
rect 305 4397 10760 4409
rect 10794 4397 10893 4431
rect 11959 4462 12366 4465
rect 11959 4454 12400 4462
rect 11959 4420 12031 4454
rect 12065 4420 12112 4454
rect 12146 4420 12193 4454
rect 12227 4420 12274 4454
rect 12308 4428 12400 4454
rect 12308 4426 12366 4428
rect 305 4393 10893 4397
rect 305 4388 949 4393
rect 305 4375 371 4388
rect 271 4341 371 4375
rect -31 4283 -15 4317
rect 19 4283 35 4317
rect -31 4249 35 4283
rect -31 4240 -15 4249
rect 19 4240 35 4249
rect 305 4307 371 4341
rect 12366 4381 12368 4394
rect 12366 4360 12402 4381
rect 12400 4340 12402 4360
rect 271 4273 371 4307
rect 4489 4333 4505 4335
rect 4489 4299 4501 4333
rect 4539 4301 4573 4335
rect 4607 4301 4641 4335
rect 4675 4333 4709 4335
rect 4743 4333 4777 4335
rect 4811 4333 4845 4335
rect 4879 4333 4913 4335
rect 4947 4333 4981 4335
rect 5015 4333 5049 4335
rect 5083 4333 5117 4335
rect 5151 4333 5185 4335
rect 4679 4301 4709 4333
rect 4751 4301 4777 4333
rect 4823 4301 4845 4333
rect 4895 4301 4913 4333
rect 4967 4301 4981 4333
rect 5039 4301 5049 4333
rect 5111 4301 5117 4333
rect 5183 4301 5185 4333
rect 5219 4333 5253 4335
rect 5287 4333 5321 4335
rect 5355 4333 5389 4335
rect 5423 4333 5457 4335
rect 5491 4333 5525 4335
rect 5559 4333 5593 4335
rect 5219 4301 5221 4333
rect 5287 4301 5293 4333
rect 5355 4301 5365 4333
rect 5423 4301 5437 4333
rect 5491 4301 5509 4333
rect 5559 4301 5581 4333
rect 5627 4301 5643 4335
rect 4535 4299 4573 4301
rect 4607 4299 4645 4301
rect 4679 4299 4717 4301
rect 4751 4299 4789 4301
rect 4823 4299 4861 4301
rect 4895 4299 4933 4301
rect 4967 4299 5005 4301
rect 5039 4299 5077 4301
rect 5111 4299 5149 4301
rect 5183 4299 5221 4301
rect 5255 4299 5293 4301
rect 5327 4299 5365 4301
rect 5399 4299 5437 4301
rect 5471 4299 5509 4301
rect 5543 4299 5581 4301
rect 5615 4299 5643 4301
rect -31 4215 -26 4240
rect 19 4215 46 4240
rect 8 4206 46 4215
rect 305 4239 371 4273
rect 271 4205 371 4239
rect 305 4199 371 4205
rect 1536 4255 1609 4285
rect 1643 4255 1677 4285
rect 1711 4255 1745 4285
rect 1779 4255 1813 4285
rect 1847 4255 1881 4285
rect 1570 4251 1609 4255
rect 1647 4251 1677 4255
rect 1724 4251 1745 4255
rect 1801 4251 1813 4255
rect 1878 4251 1881 4255
rect 1915 4255 1949 4285
rect 1983 4255 2017 4285
rect 2051 4255 2085 4285
rect 2119 4255 2183 4285
rect 1915 4251 1921 4255
rect 1983 4251 1997 4255
rect 2051 4251 2073 4255
rect 2119 4251 2149 4255
rect 1570 4221 1613 4251
rect 1647 4221 1690 4251
rect 1724 4221 1767 4251
rect 1801 4221 1844 4251
rect 1878 4221 1921 4251
rect 1955 4221 1997 4251
rect 2031 4221 2073 4251
rect 2107 4221 2149 4251
rect 2217 4251 2233 4285
rect 2267 4255 2301 4285
rect 2300 4251 2301 4255
rect 2335 4255 2369 4285
rect 2403 4255 2437 4285
rect 2471 4255 2505 4285
rect 2335 4251 2343 4255
rect 2403 4251 2420 4255
rect 2471 4251 2497 4255
rect 2539 4251 2573 4285
rect 2607 4251 2641 4285
rect 2675 4251 2709 4285
rect 2743 4251 2761 4285
rect 2217 4221 2266 4251
rect 2300 4221 2343 4251
rect 2377 4221 2420 4251
rect 2454 4221 2497 4251
rect 2531 4221 2761 4251
rect 3045 4251 3061 4285
rect 3095 4255 3129 4285
rect 3163 4255 3197 4285
rect 3231 4255 3265 4285
rect 3299 4255 3333 4285
rect 3367 4255 3401 4285
rect 3435 4255 3469 4285
rect 3106 4251 3129 4255
rect 3178 4251 3197 4255
rect 3250 4251 3265 4255
rect 3322 4251 3333 4255
rect 3394 4251 3401 4255
rect 3466 4251 3469 4255
rect 3503 4255 3537 4285
rect 3571 4255 3605 4285
rect 3639 4255 3673 4285
rect 3707 4255 3741 4285
rect 3775 4255 3809 4285
rect 3843 4255 3877 4285
rect 3911 4255 3945 4285
rect 3979 4255 4013 4285
rect 4047 4255 4081 4285
rect 3503 4251 3504 4255
rect 3571 4251 3576 4255
rect 3639 4251 3648 4255
rect 3707 4251 3720 4255
rect 3775 4251 3792 4255
rect 3843 4251 3864 4255
rect 3911 4251 3936 4255
rect 3979 4251 4008 4255
rect 4047 4251 4080 4255
rect 4115 4251 4149 4285
rect 4183 4255 4199 4285
rect 4489 4265 5643 4299
rect 9145 4306 9179 4322
rect 3045 4221 3072 4251
rect 3106 4221 3144 4251
rect 3178 4221 3216 4251
rect 3250 4221 3288 4251
rect 3322 4221 3360 4251
rect 3394 4221 3432 4251
rect 3466 4221 3504 4251
rect 3538 4221 3576 4251
rect 3610 4221 3648 4251
rect 3682 4221 3720 4251
rect 3754 4221 3792 4251
rect 3826 4221 3864 4251
rect 3898 4221 3936 4251
rect 3970 4221 4008 4251
rect 4042 4221 4080 4251
rect 4114 4221 4152 4251
rect 4186 4221 4199 4255
rect 75 4155 109 4171
rect -101 4121 75 4144
rect -101 4110 109 4121
rect -277 4038 -243 4053
rect -644 3997 -638 4031
rect -604 4002 -566 4031
rect -581 3997 -566 4002
rect 70 4087 109 4110
rect 70 4053 75 4087
rect 70 4037 109 4053
rect 271 4137 305 4171
rect 271 4069 305 4100
rect -644 3968 -615 3997
rect -581 3968 -532 3997
rect -644 3954 -532 3968
rect -644 3920 -638 3954
rect -604 3920 -566 3954
rect -644 3912 -532 3920
rect -644 3878 -615 3912
rect -581 3878 -532 3912
rect -644 3876 -532 3878
rect -644 3842 -638 3876
rect -604 3842 -566 3876
rect 271 4001 305 4020
rect 271 3933 305 3940
rect 271 3893 305 3899
rect -644 3822 -532 3842
rect -644 3798 -615 3822
rect -581 3798 -532 3822
rect -644 3764 -638 3798
rect -581 3788 -566 3798
rect -604 3764 -566 3788
rect -470 3807 -436 3823
rect -470 3429 -436 3773
rect -314 3807 -280 3834
rect -314 3757 -280 3762
rect -190 3819 -156 3834
rect -190 3751 -156 3762
rect -394 3702 -360 3716
rect -190 3701 -156 3717
rect -14 3819 20 3835
rect -14 3751 20 3785
rect -394 3632 -360 3666
rect -394 3582 -360 3596
rect -117 3623 -101 3657
rect -67 3623 -51 3657
rect -117 3622 -51 3623
rect -117 3555 -101 3622
rect -67 3555 -51 3622
rect -101 3550 -67 3555
rect -190 3489 -156 3505
rect -470 3361 -436 3395
rect -470 3293 -436 3327
rect -470 3225 -436 3259
rect -470 3157 -436 3189
rect -470 3089 -436 3117
rect -470 3021 -436 3055
rect -470 2953 -436 2987
rect -470 2903 -436 2919
rect -314 3429 -280 3445
rect -314 3361 -280 3395
rect -314 3293 -280 3327
rect -314 3225 -280 3259
rect -314 3157 -280 3191
rect -314 3118 -280 3123
rect -314 3046 -280 3055
rect -190 3421 -156 3455
rect -190 3353 -156 3387
rect -190 3227 -156 3319
rect -190 3159 -156 3193
rect -190 3117 -156 3125
rect -190 3045 -156 3057
rect -14 3489 20 3717
rect -14 3421 20 3455
rect 271 3812 305 3831
rect 1016 4164 1050 4199
rect 1016 4096 1050 4130
rect 1016 4028 1050 4062
rect 1016 3960 1050 3994
rect 1016 3892 1050 3926
rect 1016 3824 1050 3858
rect 271 3729 305 3763
rect 271 3661 305 3695
rect 271 3593 305 3627
rect 271 3525 305 3559
rect 271 3457 305 3491
rect 20 3387 129 3395
rect -14 3361 129 3387
rect -14 3353 163 3361
rect 20 3323 163 3353
rect 20 3319 129 3323
rect -14 3289 129 3319
rect 271 3389 305 3423
rect 707 3719 813 3808
rect 741 3685 779 3719
rect 707 3414 813 3685
rect 1016 3756 1050 3790
rect 1016 3688 1050 3722
rect 1016 3643 1050 3654
rect 1016 3571 1050 3586
rect 1016 3499 1050 3518
rect 1016 3416 1050 3450
rect 271 3321 305 3355
rect -14 3227 20 3289
rect -14 3159 20 3193
rect -14 3091 20 3125
rect -14 3039 20 3057
rect 271 3253 305 3287
rect 271 3185 305 3219
rect 1016 3348 1050 3382
rect 1016 3280 1050 3314
rect 1016 3211 1050 3246
rect 1114 4133 1148 4149
rect 1114 4065 1148 4099
rect 1114 3997 1148 4031
rect 1114 3929 1148 3963
rect 1114 3861 1148 3895
rect 1114 3793 1148 3827
rect 1114 3725 1148 3759
rect 1114 3657 1148 3691
rect 1114 3589 1148 3623
rect 1114 3521 1148 3555
rect 1114 3453 1148 3487
rect 1270 4133 1304 4149
rect 1270 4065 1304 4099
rect 1270 3997 1304 4031
rect 1270 3929 1304 3963
rect 1426 4133 1460 4149
rect 1426 4065 1460 4099
rect 1426 3997 1460 4031
rect 1426 3945 1460 3963
rect 1388 3911 1426 3945
rect 1270 3861 1304 3895
rect 1270 3793 1304 3827
rect 1270 3725 1304 3759
rect 1270 3657 1304 3691
rect 1270 3589 1304 3609
rect 1270 3521 1304 3537
rect 1270 3453 1304 3465
rect 1148 3385 1186 3419
rect 1270 3385 1304 3419
rect 1114 3317 1148 3351
rect 1114 3249 1148 3283
rect 1114 3199 1148 3215
rect 1270 3317 1304 3351
rect 1270 3249 1304 3283
rect 1270 3199 1304 3215
rect 1426 3861 1460 3895
rect 1426 3793 1460 3827
rect 1426 3725 1460 3759
rect 1426 3657 1460 3691
rect 1426 3589 1460 3623
rect 1426 3521 1460 3555
rect 1426 3453 1460 3487
rect 1426 3385 1460 3419
rect 1426 3317 1460 3351
rect 1426 3249 1460 3283
rect 1426 3199 1460 3215
rect 1536 4133 1570 4221
rect 1536 4065 1570 4099
rect 1536 3997 1570 4031
rect 1536 3929 1570 3963
rect 1692 4133 1726 4149
rect 1692 4065 1726 4099
rect 1692 3997 1726 4031
rect 1692 3945 1726 3963
rect 1848 4133 1882 4221
rect 2149 4149 2183 4221
rect 1848 4065 1882 4099
rect 1848 3997 1882 4031
rect 1689 3929 1727 3945
rect 1689 3911 1692 3929
rect 1536 3861 1570 3895
rect 1536 3793 1570 3827
rect 1536 3725 1570 3759
rect 1726 3911 1727 3929
rect 1848 3929 1882 3963
rect 2004 4133 2038 4149
rect 2004 4065 2038 4099
rect 2004 3997 2038 4031
rect 2004 3945 2038 3963
rect 2149 4133 2194 4149
rect 2149 4099 2160 4133
rect 2149 4065 2194 4099
rect 2149 4031 2160 4065
rect 2149 3997 2194 4031
rect 2149 3963 2160 3997
rect 1692 3861 1726 3895
rect 1692 3793 1726 3827
rect 1692 3725 1726 3759
rect 1570 3689 1608 3723
rect 2000 3929 2038 3945
rect 2000 3911 2004 3929
rect 1848 3861 1882 3895
rect 1848 3793 1882 3827
rect 1848 3725 1882 3759
rect 1536 3657 1570 3689
rect 1536 3589 1570 3623
rect 1536 3521 1570 3555
rect 1536 3453 1570 3487
rect 1536 3385 1570 3419
rect 1536 3317 1570 3351
rect 1536 3249 1570 3283
rect 1536 3199 1570 3215
rect 1692 3657 1726 3691
rect 1844 3691 1848 3723
rect 2149 3929 2194 3963
rect 2004 3861 2038 3895
rect 2004 3793 2038 3827
rect 2004 3725 2038 3759
rect 1844 3689 1882 3691
rect 2149 3895 2160 3929
rect 2149 3861 2194 3895
rect 2149 3827 2160 3861
rect 2316 4133 2350 4221
rect 2316 4065 2350 4099
rect 2316 3997 2350 4031
rect 2316 3929 2350 3963
rect 2316 3861 2350 3895
rect 2149 3793 2194 3827
rect 2313 3827 2316 3859
rect 2472 4133 2506 4149
rect 2472 4065 2506 4099
rect 2472 3997 2506 4031
rect 2472 3929 2506 3963
rect 2472 3861 2506 3895
rect 2350 3827 2351 3859
rect 2313 3825 2351 3827
rect 2628 4133 2662 4221
rect 2882 4164 2916 4199
rect 2628 4065 2662 4099
rect 2628 3997 2662 4031
rect 2628 3929 2662 3963
rect 2628 3861 2662 3895
rect 2149 3759 2160 3793
rect 2149 3725 2194 3759
rect 2149 3723 2160 3725
rect 1692 3589 1726 3623
rect 1692 3521 1726 3555
rect 1692 3453 1726 3487
rect 1692 3385 1726 3419
rect 1692 3317 1726 3351
rect 1692 3249 1726 3283
rect 271 3117 305 3151
rect 1163 3126 1179 3155
rect 1163 3092 1175 3126
rect 1213 3121 1247 3155
rect 1281 3121 1315 3155
rect 1349 3126 1383 3155
rect 1417 3126 1433 3155
rect 1353 3121 1383 3126
rect 1209 3092 1247 3121
rect 1281 3092 1319 3121
rect 1353 3092 1391 3121
rect 1425 3092 1433 3126
rect 271 3049 305 3083
rect 1692 3071 1726 3215
rect 1848 3657 1882 3689
rect 1848 3589 1882 3623
rect 1848 3521 1882 3555
rect 1848 3453 1882 3487
rect 1848 3385 1882 3419
rect 1848 3317 1882 3351
rect 1848 3249 1882 3283
rect 1848 3199 1882 3215
rect 2004 3657 2038 3691
rect 2156 3691 2160 3723
rect 2316 3793 2350 3825
rect 2316 3725 2350 3759
rect 2156 3689 2194 3691
rect 2472 3793 2506 3827
rect 2624 3827 2628 3859
rect 2784 4133 2818 4149
rect 2784 4065 2818 4099
rect 2784 3997 2818 4031
rect 2784 3929 2818 3963
rect 2784 3861 2818 3895
rect 2624 3825 2662 3827
rect 2472 3725 2506 3759
rect 2004 3589 2038 3623
rect 2004 3521 2038 3555
rect 2004 3453 2038 3487
rect 2004 3385 2038 3419
rect 2004 3317 2038 3351
rect 2004 3249 2038 3283
rect 2149 3657 2194 3689
rect 2149 3623 2160 3657
rect 2149 3589 2194 3623
rect 2149 3555 2160 3589
rect 2149 3521 2194 3555
rect 2149 3487 2160 3521
rect 2149 3453 2194 3487
rect 2149 3419 2160 3453
rect 2149 3385 2194 3419
rect 2149 3351 2160 3385
rect 2149 3317 2194 3351
rect 2149 3283 2160 3317
rect 2149 3257 2194 3283
rect 2004 3199 2038 3215
rect 2160 3249 2194 3257
rect 2160 3199 2194 3215
rect 2316 3657 2350 3691
rect 2468 3691 2472 3723
rect 2628 3793 2662 3825
rect 2628 3725 2662 3759
rect 2468 3689 2506 3691
rect 2784 3793 2818 3827
rect 2784 3725 2818 3759
rect 2316 3589 2350 3623
rect 2316 3521 2350 3555
rect 2316 3453 2350 3487
rect 2316 3385 2350 3419
rect 2316 3317 2350 3351
rect 2316 3249 2350 3283
rect 2316 3199 2350 3215
rect 2472 3657 2506 3689
rect 2472 3589 2506 3623
rect 2472 3521 2506 3555
rect 2472 3453 2506 3487
rect 2472 3385 2506 3419
rect 2472 3317 2506 3351
rect 2472 3249 2506 3283
rect 2472 3199 2506 3215
rect 2628 3657 2662 3691
rect 2746 3689 2784 3723
rect 2628 3589 2662 3623
rect 2628 3521 2662 3555
rect 2628 3453 2662 3487
rect 2628 3385 2662 3419
rect 2628 3317 2662 3351
rect 2628 3249 2662 3283
rect 2628 3199 2662 3215
rect 2784 3657 2818 3689
rect 2784 3589 2818 3623
rect 2784 3521 2818 3555
rect 2784 3453 2818 3487
rect 2784 3385 2818 3419
rect 2784 3317 2818 3351
rect 2784 3249 2818 3283
rect 2784 3199 2818 3215
rect 4228 4164 4360 4199
rect 2882 4096 2916 4130
rect 2882 4028 2916 4062
rect 2882 3960 2916 3994
rect 2882 3892 2916 3926
rect 2882 3824 2916 3858
rect 2882 3756 2916 3790
rect 2882 3688 2916 3722
rect 2882 3643 2916 3654
rect 2980 4133 3014 4149
rect 2980 4065 3014 4099
rect 2980 3997 3014 4031
rect 2980 3929 3014 3963
rect 2980 3861 3014 3895
rect 2980 3793 3014 3827
rect 2980 3725 3014 3759
rect 3136 4133 3170 4149
rect 3136 4065 3170 4099
rect 3136 3997 3170 4031
rect 3136 3929 3170 3963
rect 3136 3861 3170 3895
rect 3136 3793 3170 3827
rect 3136 3725 3170 3759
rect 2980 3657 3014 3691
rect 3132 3691 3136 3723
rect 3292 4133 3382 4149
rect 3326 4099 3382 4133
rect 3292 4065 3382 4099
rect 3326 4031 3382 4065
rect 3292 3997 3382 4031
rect 3326 3963 3382 3997
rect 3292 3929 3382 3963
rect 3326 3895 3382 3929
rect 3292 3861 3382 3895
rect 3326 3827 3382 3861
rect 3292 3793 3382 3827
rect 3326 3759 3382 3793
rect 3292 3725 3382 3759
rect 3132 3689 3170 3691
rect 3326 3691 3382 3725
rect 3448 4133 3482 4149
rect 3448 4065 3482 4099
rect 3448 3997 3482 4031
rect 3448 3929 3482 3963
rect 3448 3861 3482 3895
rect 3448 3793 3482 3827
rect 3448 3725 3482 3759
rect 3604 4133 3638 4149
rect 3604 4065 3638 4099
rect 3604 3997 3638 4031
rect 3604 3929 3638 3963
rect 3604 3861 3638 3895
rect 3604 3793 3638 3827
rect 3604 3725 3638 3759
rect 3136 3657 3170 3689
rect 3292 3657 3382 3691
rect 3482 3691 3488 3723
rect 3450 3689 3488 3691
rect 3760 4133 3794 4149
rect 3760 4065 3794 4099
rect 3760 3997 3794 4031
rect 3760 3929 3794 3963
rect 3760 3861 3794 3895
rect 3760 3793 3794 3827
rect 3760 3725 3794 3759
rect 3326 3643 3382 3657
rect 3136 3589 3170 3623
rect 3136 3521 3170 3555
rect 2882 3416 2916 3450
rect 2882 3348 2916 3382
rect 2882 3280 2916 3314
rect 2882 3211 2916 3246
rect 2980 3453 3014 3465
rect 2980 3385 3014 3419
rect 2980 3317 3014 3351
rect 2980 3249 3014 3283
rect 2980 3199 3014 3215
rect 3136 3453 3170 3487
rect 3376 3465 3382 3643
rect 3136 3385 3170 3419
rect 3136 3317 3170 3351
rect 3136 3249 3170 3283
rect 3136 3199 3170 3215
rect 3292 3453 3382 3465
rect 3326 3419 3382 3453
rect 3292 3385 3382 3419
rect 3326 3351 3382 3385
rect 3292 3317 3382 3351
rect 3326 3283 3382 3317
rect 3292 3249 3382 3283
rect 3326 3215 3382 3249
rect 1692 3021 1726 3037
rect 3292 3071 3382 3215
rect 3448 3657 3482 3689
rect 3448 3589 3482 3623
rect 3448 3521 3482 3555
rect 3448 3453 3482 3487
rect 3448 3385 3482 3419
rect 3448 3317 3482 3351
rect 3448 3249 3482 3283
rect 3448 3199 3482 3215
rect 3604 3657 3638 3691
rect 3756 3691 3760 3723
rect 3916 4133 3950 4149
rect 3916 4065 3950 4099
rect 3916 3997 3950 4031
rect 3916 3929 3950 3963
rect 3916 3861 3950 3895
rect 3916 3793 3950 3827
rect 3916 3725 3950 3759
rect 3756 3689 3794 3691
rect 4072 4133 4106 4149
rect 4072 4065 4106 4099
rect 4072 3997 4106 4031
rect 4072 3929 4106 3963
rect 4072 3861 4106 3895
rect 4072 3793 4106 3827
rect 4072 3725 4106 3759
rect 4228 4133 4326 4164
rect 4262 4130 4326 4133
rect 4262 4099 4360 4130
rect 4228 4096 4360 4099
rect 4228 4065 4326 4096
rect 4262 4062 4326 4065
rect 4262 4031 4360 4062
rect 4228 4028 4360 4031
rect 4228 3997 4326 4028
rect 4262 3994 4326 3997
rect 4262 3963 4360 3994
rect 4228 3960 4360 3963
rect 4228 3929 4326 3960
rect 4262 3926 4326 3929
rect 4262 3895 4360 3926
rect 4228 3892 4360 3895
rect 4228 3861 4326 3892
rect 4262 3858 4326 3861
rect 4262 3827 4360 3858
rect 4228 3824 4360 3827
rect 4228 3793 4326 3824
rect 4262 3790 4326 3793
rect 4262 3759 4360 3790
rect 4228 3756 4360 3759
rect 4228 3725 4326 3756
rect 3604 3589 3638 3609
rect 3604 3521 3638 3537
rect 3604 3453 3638 3465
rect 3604 3385 3638 3419
rect 3604 3317 3638 3351
rect 3604 3249 3638 3283
rect 3604 3075 3638 3215
rect 3760 3657 3794 3689
rect 3760 3589 3794 3623
rect 3760 3521 3794 3555
rect 3760 3453 3794 3487
rect 3760 3385 3794 3419
rect 3760 3317 3794 3351
rect 3760 3249 3794 3283
rect 3760 3199 3794 3215
rect 3916 3657 3950 3691
rect 4067 3691 4072 3723
rect 4067 3689 4105 3691
rect 4262 3722 4326 3725
rect 4424 4183 4458 4199
rect 4424 4115 4458 4149
rect 4424 4047 4458 4081
rect 4424 3979 4458 4013
rect 4424 3911 4458 3945
rect 4424 3843 4458 3877
rect 4424 3775 4458 3809
rect 4424 3723 4458 3741
rect 4580 4183 4614 4265
rect 4580 4115 4614 4149
rect 4580 4047 4614 4081
rect 4580 3979 4614 4013
rect 4580 3911 4614 3945
rect 4580 3843 4614 3877
rect 4580 3775 4614 3809
rect 4262 3691 4360 3722
rect 3916 3589 3950 3609
rect 3916 3521 3950 3537
rect 3916 3453 3950 3465
rect 3916 3385 3950 3419
rect 3916 3317 3950 3351
rect 3916 3249 3950 3283
rect 3916 3075 3950 3215
rect 4072 3657 4106 3689
rect 4228 3688 4360 3691
rect 4457 3707 4495 3723
rect 4458 3689 4495 3707
rect 4580 3707 4614 3741
rect 4736 4183 4770 4199
rect 4736 4115 4770 4149
rect 4736 4047 4770 4081
rect 4736 3979 4770 4013
rect 4736 3911 4770 3945
rect 4736 3843 4770 3877
rect 4736 3775 4770 3809
rect 4736 3723 4770 3741
rect 4892 4183 4926 4265
rect 4892 4115 4926 4149
rect 4892 4047 4926 4081
rect 4892 3979 4926 4013
rect 4892 3911 4926 3945
rect 4892 3843 4926 3877
rect 4892 3775 4926 3809
rect 4228 3657 4326 3688
rect 4262 3654 4326 3657
rect 4262 3643 4360 3654
rect 4072 3589 4106 3623
rect 4072 3521 4106 3555
rect 4072 3453 4106 3487
rect 4359 3620 4360 3643
rect 4359 3552 4360 3586
rect 4359 3484 4360 3518
rect 4072 3385 4106 3419
rect 4072 3317 4106 3351
rect 4072 3249 4106 3283
rect 4072 3199 4106 3215
rect 4228 3453 4326 3465
rect 4262 3450 4326 3453
rect 4262 3419 4360 3450
rect 4228 3416 4360 3419
rect 4228 3385 4326 3416
rect 4262 3382 4326 3385
rect 4262 3351 4360 3382
rect 4228 3348 4360 3351
rect 4228 3317 4326 3348
rect 4262 3314 4326 3317
rect 4262 3283 4360 3314
rect 4228 3280 4360 3283
rect 4228 3249 4326 3280
rect 4262 3246 4326 3249
rect 4424 3639 4458 3673
rect 4424 3571 4458 3605
rect 4424 3503 4458 3537
rect 4424 3435 4458 3469
rect 4731 3707 4769 3723
rect 4731 3689 4736 3707
rect 4892 3707 4926 3741
rect 5048 4183 5082 4199
rect 5048 4115 5082 4149
rect 5048 4047 5082 4081
rect 5048 3979 5082 4013
rect 5048 3911 5082 3945
rect 5048 3843 5082 3877
rect 5048 3775 5082 3809
rect 5048 3723 5082 3741
rect 5204 4183 5238 4265
rect 5204 4115 5238 4149
rect 5204 4047 5238 4081
rect 5204 3979 5238 4013
rect 5204 3911 5238 3945
rect 5204 3843 5238 3877
rect 5204 3775 5238 3809
rect 4580 3639 4614 3673
rect 4580 3571 4614 3605
rect 4580 3503 4614 3537
rect 4580 3435 4614 3469
rect 4424 3367 4458 3401
rect 4576 3401 4580 3419
rect 4736 3639 4770 3673
rect 4736 3571 4770 3605
rect 4736 3503 4770 3537
rect 4736 3435 4770 3469
rect 4576 3385 4614 3401
rect 5043 3707 5081 3723
rect 5043 3689 5048 3707
rect 5204 3707 5238 3741
rect 5360 4183 5394 4199
rect 5360 4115 5394 4149
rect 5360 4047 5394 4081
rect 5360 3979 5394 4013
rect 5360 3911 5394 3945
rect 5360 3843 5394 3877
rect 5360 3775 5394 3809
rect 5360 3723 5394 3741
rect 5516 4183 5550 4265
rect 5677 4251 5950 4285
rect 5984 4251 6018 4285
rect 6052 4251 6086 4285
rect 6120 4251 6154 4285
rect 6188 4251 6222 4285
rect 6256 4251 6290 4285
rect 6324 4251 6358 4285
rect 6392 4251 6426 4285
rect 6460 4251 6494 4285
rect 6528 4251 6562 4285
rect 6596 4251 6630 4285
rect 6664 4251 6698 4285
rect 6732 4251 6766 4285
rect 6800 4251 6834 4285
rect 6868 4251 6902 4285
rect 6936 4251 6970 4285
rect 7004 4251 7038 4285
rect 7072 4251 7088 4285
rect 5677 4249 7088 4251
rect 5677 4199 5711 4249
rect 5934 4215 5951 4249
rect 5985 4215 6023 4249
rect 6057 4215 6095 4249
rect 6129 4215 6167 4249
rect 6201 4215 6239 4249
rect 6273 4215 6311 4249
rect 6345 4215 6383 4249
rect 6417 4215 6455 4249
rect 6489 4215 6527 4249
rect 6561 4215 6599 4249
rect 6633 4215 6671 4249
rect 6705 4215 6743 4249
rect 6777 4215 6815 4249
rect 6849 4215 6887 4249
rect 6921 4215 6959 4249
rect 6993 4215 7031 4249
rect 7065 4215 7088 4249
rect 7161 4251 7177 4285
rect 7211 4251 7245 4285
rect 7279 4251 7295 4285
rect 7161 4249 7295 4251
rect 7161 4215 7173 4249
rect 7207 4215 7245 4249
rect 7279 4215 7295 4249
rect 7462 4251 7478 4285
rect 7512 4251 7546 4285
rect 7580 4251 7596 4285
rect 7814 4251 7830 4285
rect 7864 4251 7898 4285
rect 7462 4217 7506 4251
rect 7540 4217 7578 4251
rect 7814 4217 7826 4251
rect 7860 4217 7898 4251
rect 7932 4217 7948 4285
rect 9145 4238 9179 4272
rect 9301 4306 9335 4322
rect 9301 4253 9335 4272
rect 9457 4306 9491 4322
rect 5516 4115 5550 4149
rect 5516 4047 5550 4081
rect 5516 3979 5550 4013
rect 5516 3911 5550 3945
rect 5516 3843 5550 3877
rect 5516 3775 5550 3809
rect 4892 3639 4926 3673
rect 4892 3571 4926 3605
rect 4892 3503 4926 3537
rect 4892 3435 4926 3469
rect 4424 3299 4458 3333
rect 4424 3249 4458 3265
rect 4580 3367 4614 3385
rect 4580 3299 4614 3333
rect 4580 3249 4614 3265
rect 4736 3367 4770 3401
rect 4888 3401 4892 3419
rect 5048 3639 5082 3673
rect 5048 3571 5082 3605
rect 5048 3503 5082 3537
rect 5048 3435 5082 3469
rect 4888 3385 4926 3401
rect 5355 3707 5393 3723
rect 5355 3689 5360 3707
rect 5516 3707 5550 3741
rect 5672 4183 5711 4199
rect 5706 4149 5711 4183
rect 5672 4115 5711 4149
rect 5706 4081 5711 4115
rect 5672 4047 5711 4081
rect 5706 4013 5711 4047
rect 5672 3979 5711 4013
rect 5706 3945 5711 3979
rect 5672 3911 5711 3945
rect 5706 3877 5711 3911
rect 5672 3843 5711 3877
rect 5706 3809 5711 3843
rect 5672 3775 5711 3809
rect 5706 3741 5711 3775
rect 5672 3723 5711 3741
rect 5204 3639 5238 3673
rect 5204 3571 5238 3605
rect 5204 3503 5238 3537
rect 5204 3435 5238 3469
rect 4736 3299 4770 3333
rect 4736 3249 4770 3265
rect 4892 3367 4926 3385
rect 4892 3299 4926 3333
rect 4892 3249 4926 3265
rect 5048 3367 5082 3401
rect 5200 3401 5204 3419
rect 5360 3639 5394 3673
rect 5360 3571 5394 3605
rect 5360 3503 5394 3537
rect 5360 3435 5394 3469
rect 5200 3385 5238 3401
rect 5633 3689 5671 3723
rect 5705 3707 5711 3723
rect 5516 3639 5550 3673
rect 5516 3571 5550 3605
rect 5516 3503 5550 3537
rect 5516 3435 5550 3469
rect 5048 3299 5082 3333
rect 5048 3249 5082 3265
rect 5204 3367 5238 3385
rect 5204 3299 5238 3333
rect 5204 3249 5238 3265
rect 5360 3367 5394 3401
rect 5512 3401 5516 3419
rect 5706 3673 5711 3707
rect 5672 3639 5711 3673
rect 5706 3605 5711 3639
rect 5672 3571 5711 3605
rect 5706 3537 5711 3571
rect 5672 3503 5711 3537
rect 5706 3469 5711 3503
rect 5672 3435 5711 3469
rect 5512 3385 5550 3401
rect 5706 3401 5711 3435
rect 5360 3299 5394 3333
rect 5360 3249 5394 3265
rect 5516 3367 5550 3385
rect 5516 3299 5550 3333
rect 5516 3249 5550 3265
rect 5672 3367 5711 3401
rect 5706 3333 5711 3367
rect 5672 3299 5711 3333
rect 5706 3265 5711 3299
rect 5672 3257 5711 3265
rect 5770 4164 5804 4199
rect 5770 4096 5804 4130
rect 5770 4028 5804 4062
rect 5770 3960 5804 3994
rect 5770 3892 5804 3926
rect 5770 3824 5804 3858
rect 5770 3756 5804 3790
rect 5770 3688 5804 3722
rect 5770 3643 5804 3654
rect 5868 4133 5902 4149
rect 5868 4065 5902 4099
rect 5868 3997 5902 4031
rect 5868 3929 5902 3963
rect 5868 3861 5902 3895
rect 5868 3793 5902 3827
rect 5868 3725 5902 3759
rect 5868 3657 5902 3691
rect 6024 4133 6058 4215
rect 6024 4065 6058 4099
rect 6024 3997 6058 4031
rect 6024 3929 6058 3963
rect 6024 3861 6058 3895
rect 6024 3793 6058 3827
rect 6024 3725 6058 3759
rect 6024 3657 6058 3691
rect 6024 3589 6058 3623
rect 6024 3521 6058 3555
rect 5770 3416 5804 3450
rect 5770 3348 5804 3382
rect 5770 3280 5804 3314
rect 5672 3249 5706 3257
rect 4262 3215 4360 3246
rect 4228 3075 4360 3215
rect 5770 3211 5804 3246
rect 5868 3453 5902 3465
rect 5868 3385 5902 3419
rect 5868 3317 5902 3351
rect 5868 3249 5902 3283
rect 5868 3199 5902 3215
rect 6024 3453 6058 3487
rect 6024 3385 6058 3419
rect 6024 3317 6058 3351
rect 6024 3249 6058 3283
rect 6024 3199 6058 3215
rect 6180 4133 6214 4149
rect 6180 4065 6214 4099
rect 6180 3997 6214 4031
rect 6180 3929 6214 3963
rect 6180 3861 6214 3895
rect 6180 3793 6214 3827
rect 6180 3725 6214 3759
rect 6180 3657 6214 3691
rect 6180 3589 6214 3609
rect 6180 3521 6214 3537
rect 6180 3453 6214 3465
rect 6180 3385 6214 3419
rect 6180 3317 6214 3351
rect 6180 3249 6214 3283
rect 6180 3199 6214 3215
rect 6336 4133 6370 4215
rect 6336 4065 6370 4099
rect 6336 3997 6370 4031
rect 6336 3929 6370 3963
rect 6336 3861 6370 3895
rect 6336 3793 6370 3827
rect 6336 3725 6370 3759
rect 6336 3657 6370 3691
rect 6336 3589 6370 3623
rect 6336 3521 6370 3555
rect 6336 3453 6370 3487
rect 6336 3385 6370 3419
rect 6336 3317 6370 3351
rect 6336 3249 6370 3283
rect 6336 3199 6370 3215
rect 6492 4133 6526 4149
rect 6492 4065 6526 4099
rect 6492 3997 6526 4031
rect 6492 3929 6526 3963
rect 6492 3861 6526 3895
rect 6492 3793 6526 3827
rect 6492 3725 6526 3759
rect 6492 3657 6526 3691
rect 6492 3589 6526 3609
rect 6492 3521 6526 3537
rect 6492 3453 6526 3465
rect 6492 3385 6526 3419
rect 6492 3317 6526 3351
rect 6492 3249 6526 3283
rect 6492 3199 6526 3215
rect 6648 4133 6682 4215
rect 6648 4065 6682 4099
rect 6648 3997 6682 4031
rect 6648 3929 6682 3963
rect 6648 3861 6682 3895
rect 6648 3793 6682 3827
rect 6648 3725 6682 3759
rect 6648 3657 6682 3691
rect 6648 3589 6682 3623
rect 6648 3521 6682 3555
rect 6648 3453 6682 3487
rect 6648 3385 6682 3419
rect 6648 3317 6682 3351
rect 6648 3249 6682 3283
rect 6648 3199 6682 3215
rect 6804 4133 6838 4149
rect 6804 4065 6838 4099
rect 6804 3997 6838 4031
rect 6804 3929 6838 3963
rect 6804 3861 6838 3895
rect 6804 3793 6838 3827
rect 6804 3725 6838 3759
rect 6804 3657 6838 3691
rect 6804 3589 6838 3609
rect 6804 3521 6838 3537
rect 6804 3453 6838 3465
rect 6804 3385 6838 3419
rect 6804 3317 6838 3351
rect 6804 3249 6838 3283
rect 6804 3199 6838 3215
rect 6960 4133 6994 4215
rect 9299 4238 9337 4253
rect 9299 4219 9301 4238
rect 7370 4164 7404 4199
rect 6960 4065 6994 4099
rect 6960 3997 6994 4031
rect 6960 3929 6994 3963
rect 6960 3861 6994 3895
rect 6960 3793 6994 3827
rect 6960 3725 6994 3759
rect 6960 3657 6994 3691
rect 6960 3589 6994 3623
rect 6960 3521 6994 3555
rect 6960 3453 6994 3487
rect 6960 3385 6994 3419
rect 6960 3317 6994 3351
rect 6960 3249 6994 3283
rect 6960 3199 6994 3215
rect 7116 4133 7150 4149
rect 7116 4065 7150 4099
rect 7116 3997 7150 4031
rect 7116 3929 7150 3963
rect 7116 3861 7150 3895
rect 7116 3793 7150 3827
rect 7116 3725 7150 3759
rect 7116 3657 7150 3691
rect 7116 3589 7150 3609
rect 7116 3521 7150 3537
rect 7116 3453 7150 3465
rect 7116 3385 7150 3419
rect 7116 3317 7150 3351
rect 7116 3249 7150 3283
rect 7116 3199 7150 3215
rect 7272 4133 7306 4149
rect 7272 4065 7306 4099
rect 7272 3997 7306 4031
rect 7272 3929 7306 3963
rect 7272 3861 7306 3895
rect 7272 3793 7306 3827
rect 7272 3725 7306 3759
rect 7272 3657 7306 3691
rect 8166 4164 8200 4199
rect 9145 4170 9179 4204
rect 7370 4096 7404 4130
rect 7370 4028 7404 4062
rect 7370 3960 7404 3994
rect 7370 3892 7404 3926
rect 7370 3824 7404 3858
rect 7370 3756 7404 3790
rect 7370 3688 7404 3722
rect 7370 3643 7404 3654
rect 7468 4125 7502 4141
rect 7468 4057 7502 4091
rect 7468 3989 7502 4023
rect 7468 3921 7502 3955
rect 7468 3853 7502 3887
rect 7468 3785 7502 3819
rect 7908 4125 7978 4141
rect 7942 4091 7978 4125
rect 7908 4057 7978 4091
rect 7942 4023 7978 4057
rect 7908 3989 7978 4023
rect 7942 3955 7978 3989
rect 7908 3921 7978 3955
rect 7942 3887 7978 3921
rect 7908 3853 7978 3887
rect 7942 3819 7978 3853
rect 7468 3717 7502 3751
rect 7468 3649 7502 3683
rect 7654 3761 7795 3795
rect 7654 3723 7829 3761
rect 7654 3689 7795 3723
rect 7908 3785 7978 3819
rect 7942 3751 7978 3785
rect 7908 3717 7978 3751
rect 7272 3589 7306 3623
rect 7272 3521 7306 3555
rect 7272 3453 7306 3487
rect 7654 3526 7756 3689
rect 7942 3683 7978 3717
rect 7688 3492 7722 3526
rect 7654 3476 7756 3492
rect 7790 3643 7824 3650
rect 7790 3571 7824 3609
rect 7790 3499 7824 3537
rect 7272 3413 7306 3419
rect 7272 3341 7306 3351
rect 7272 3249 7306 3283
rect 7370 3416 7404 3450
rect 7370 3348 7404 3382
rect 7370 3280 7404 3314
rect 7370 3230 7404 3246
rect 7468 3390 7502 3465
rect 7790 3406 7824 3465
rect 7468 3322 7502 3356
rect 7468 3254 7502 3288
rect 7272 3199 7306 3215
rect 7624 3390 7658 3406
rect 7624 3339 7658 3356
rect 7780 3390 7824 3406
rect 7814 3356 7824 3390
rect 7658 3305 7696 3339
rect 7780 3322 7824 3356
rect 7624 3254 7658 3288
rect 7468 3204 7502 3220
rect 7536 3220 7624 3228
rect 7536 3194 7658 3220
rect 7814 3288 7824 3322
rect 7780 3254 7824 3288
rect 7814 3220 7824 3254
rect 7780 3204 7824 3220
rect 7908 3649 7978 3683
rect 7942 3615 7978 3649
rect 7908 3510 7978 3615
rect 7908 3476 7944 3510
rect 7908 3442 7978 3476
rect 8022 4067 8038 4101
rect 8072 4067 8128 4101
rect 8022 3643 8128 4067
rect 8166 4096 8200 4130
rect 8350 4067 8366 4101
rect 8400 4067 8510 4101
rect 8544 4067 8560 4101
rect 8166 4028 8200 4062
rect 8166 3960 8200 3994
rect 8166 3892 8200 3926
rect 8166 3824 8200 3858
rect 8166 3756 8200 3790
rect 8166 3688 8200 3722
rect 8166 3643 8200 3654
rect 8022 3453 8128 3465
rect 7908 3408 7944 3442
rect 7908 3374 7978 3408
rect 7908 3340 7944 3374
rect 7908 3306 7978 3340
rect 7908 3272 7944 3306
rect 8166 3416 8200 3450
rect 8166 3348 8200 3382
rect 7536 3140 7570 3194
rect 7519 3126 7570 3140
rect 7469 3092 7507 3126
rect 7541 3092 7570 3126
rect 7519 3086 7570 3092
rect 7604 3126 7675 3160
rect 7709 3126 7743 3160
rect 7777 3126 7811 3160
rect 7845 3126 7868 3160
rect 7604 3092 7762 3126
rect 7796 3092 7834 3126
rect 7908 3126 7978 3272
rect 8060 3268 8098 3302
rect 8026 3245 8132 3268
rect 8022 3211 8038 3245
rect 8072 3211 8132 3245
rect 8166 3280 8200 3314
rect 8278 4017 8312 4033
rect 8278 3948 8312 3983
rect 8278 3888 8312 3914
rect 8630 4013 8664 4029
rect 8630 3945 8664 3979
rect 8630 3888 8664 3911
rect 8278 3886 8664 3888
rect 9145 4102 9179 4108
rect 9145 4046 9179 4068
rect 8751 3973 8985 3986
rect 8785 3939 8851 3973
rect 8885 3939 8951 3973
rect 8751 3900 8985 3939
rect 8278 3879 8611 3886
rect 8312 3852 8611 3879
rect 8645 3877 8683 3886
rect 8664 3852 8683 3877
rect 8785 3866 8851 3900
rect 8885 3866 8951 3900
rect 8312 3845 8630 3852
rect 8278 3843 8630 3845
rect 8278 3809 8664 3843
rect 8312 3775 8630 3809
rect 8278 3741 8664 3775
rect 8278 3739 8630 3741
rect 8312 3707 8630 3739
rect 8312 3705 8664 3707
rect 8278 3673 8664 3705
rect 8278 3669 8630 3673
rect 8312 3639 8630 3669
rect 8312 3635 8664 3639
rect 8278 3605 8664 3635
rect 8278 3599 8630 3605
rect 8312 3571 8630 3599
rect 8312 3565 8664 3571
rect 8278 3537 8664 3565
rect 8278 3529 8630 3537
rect 8312 3503 8630 3529
rect 8312 3495 8664 3503
rect 8278 3469 8664 3495
rect 8278 3459 8630 3469
rect 8312 3435 8630 3459
rect 8312 3425 8664 3435
rect 8278 3401 8664 3425
rect 8278 3389 8630 3401
rect 8312 3367 8630 3389
rect 8312 3355 8664 3367
rect 8278 3333 8664 3355
rect 8278 3329 8630 3333
rect 8278 3319 8312 3329
rect 8278 3269 8312 3285
rect 8630 3283 8664 3299
rect 8751 3827 8985 3866
rect 8785 3793 8851 3827
rect 8885 3793 8951 3827
rect 8751 3754 8985 3793
rect 9145 3966 9179 4000
rect 9145 3898 9179 3932
rect 9145 3830 9179 3864
rect 9145 3780 9179 3796
rect 9335 4219 9337 4238
rect 9457 4238 9491 4272
rect 9613 4306 9647 4322
rect 9613 4253 9647 4272
rect 9737 4306 9771 4322
rect 9301 4170 9335 4204
rect 9301 4102 9335 4136
rect 9301 4034 9335 4068
rect 9301 3966 9335 4000
rect 9301 3898 9335 3932
rect 9301 3830 9335 3864
rect 9301 3780 9335 3796
rect 9604 4238 9642 4253
rect 9604 4219 9613 4238
rect 9737 4238 9771 4272
rect 9457 4170 9491 4204
rect 9457 4102 9491 4108
rect 9457 4046 9491 4068
rect 9457 3966 9491 4000
rect 9457 3898 9491 3932
rect 9457 3830 9491 3864
rect 9457 3780 9491 3796
rect 9613 4170 9647 4204
rect 9737 4170 9771 4204
rect 9893 4306 9927 4322
rect 9893 4238 9927 4272
rect 9893 4170 9927 4204
rect 9613 4102 9647 4136
rect 9771 4136 9780 4167
rect 9742 4133 9780 4136
rect 10049 4306 10083 4322
rect 10049 4238 10083 4272
rect 10049 4170 10083 4204
rect 9613 4034 9647 4068
rect 9613 3966 9647 4000
rect 9613 3898 9647 3932
rect 9613 3830 9647 3864
rect 9613 3780 9647 3796
rect 9737 4102 9771 4133
rect 9893 4102 9927 4136
rect 10045 4136 10049 4167
rect 10205 4306 10239 4322
rect 10205 4238 10239 4272
rect 10205 4170 10239 4204
rect 10045 4133 10083 4136
rect 10361 4306 10395 4322
rect 10361 4238 10395 4272
rect 10361 4170 10395 4204
rect 9737 4034 9771 4068
rect 9891 4068 9893 4090
rect 10049 4102 10083 4133
rect 9927 4068 9929 4090
rect 9891 4056 9929 4068
rect 9737 3966 9771 4000
rect 9737 3898 9771 3932
rect 9737 3830 9771 3864
rect 9737 3780 9771 3796
rect 9893 4034 9927 4056
rect 9893 3966 9927 4000
rect 9893 3898 9927 3932
rect 9893 3830 9927 3864
rect 9893 3780 9927 3796
rect 10049 4034 10083 4068
rect 10205 4102 10239 4136
rect 10358 4136 10361 4167
rect 10485 4306 10519 4322
rect 10485 4238 10519 4272
rect 10641 4306 10675 4322
rect 10641 4253 10675 4272
rect 10797 4306 10831 4322
rect 10485 4170 10519 4204
rect 10395 4136 10396 4167
rect 10358 4133 10396 4136
rect 10205 4034 10239 4068
rect 10049 3966 10083 4000
rect 10204 4000 10205 4012
rect 10361 4102 10395 4133
rect 10485 4102 10519 4136
rect 10361 4034 10395 4068
rect 10484 4068 10485 4090
rect 10641 4238 10679 4253
rect 10607 4204 10641 4219
rect 10675 4219 10679 4238
rect 10675 4204 10713 4219
rect 10607 4170 10713 4204
rect 10607 4136 10641 4170
rect 10675 4136 10713 4170
rect 10607 4102 10713 4136
rect 10519 4068 10522 4090
rect 10484 4056 10522 4068
rect 10607 4068 10641 4102
rect 10675 4068 10713 4102
rect 10239 4000 10242 4012
rect 10204 3978 10242 4000
rect 10049 3898 10083 3932
rect 10205 3966 10239 3978
rect 10205 3898 10239 3932
rect 10049 3830 10083 3864
rect 10049 3780 10083 3796
rect 10125 3817 10159 3855
rect 8785 3720 8851 3754
rect 8885 3720 8951 3754
rect 8751 3681 8985 3720
rect 8785 3647 8851 3681
rect 8885 3647 8951 3681
rect 8751 3607 8985 3647
rect 9190 3723 9722 3746
rect 9190 3689 9599 3723
rect 9633 3689 9671 3723
rect 9705 3689 9722 3723
rect 9190 3670 9722 3689
rect 10125 3670 10159 3783
rect 10361 3966 10395 4000
rect 10361 3898 10395 3932
rect 10205 3830 10239 3864
rect 10205 3780 10239 3796
rect 10285 3817 10319 3855
rect 10285 3670 10319 3783
rect 10361 3830 10395 3864
rect 10361 3780 10395 3796
rect 10485 4034 10519 4056
rect 10485 3966 10519 4000
rect 10485 3898 10519 3932
rect 10485 3830 10519 3864
rect 10485 3780 10519 3796
rect 10607 4034 10713 4068
rect 10607 4000 10641 4034
rect 10675 4000 10713 4034
rect 10797 4238 10831 4272
rect 11873 4279 11874 4313
rect 11908 4279 11946 4313
rect 12366 4306 12368 4326
rect 12366 4292 12402 4306
rect 10970 4219 11008 4253
rect 11042 4219 11051 4253
rect 10797 4170 10831 4204
rect 11017 4201 11051 4219
rect 11017 4151 11051 4167
rect 11873 4201 11980 4279
rect 12133 4247 12149 4281
rect 12183 4247 12199 4281
rect 11907 4167 11980 4201
rect 11873 4151 11980 4167
rect 12055 4220 12089 4236
rect 10797 4102 10831 4136
rect 12055 4148 12089 4186
rect 10797 4034 10831 4068
rect 10944 4114 12055 4117
rect 12133 4220 12199 4247
rect 12133 4186 12145 4220
rect 12179 4186 12199 4220
rect 12133 4148 12199 4186
rect 12133 4114 12145 4148
rect 12179 4114 12199 4148
rect 12400 4265 12402 4292
rect 12366 4231 12368 4258
rect 12366 4224 12402 4231
rect 12400 4190 12402 4224
rect 12366 4156 12368 4190
rect 12400 4122 12402 4156
rect 12366 4115 12402 4122
rect 10944 4109 12089 4114
rect 10944 4075 10956 4109
rect 10990 4075 11028 4109
rect 11062 4107 12089 4109
rect 11062 4075 11078 4107
rect 10944 4073 11078 4075
rect 11112 4073 11152 4107
rect 11186 4073 11226 4107
rect 11260 4073 11300 4107
rect 11334 4073 11374 4107
rect 11408 4073 11447 4107
rect 11481 4073 11520 4107
rect 11554 4073 11593 4107
rect 11627 4073 11666 4107
rect 11700 4073 11739 4107
rect 11773 4073 11812 4107
rect 11846 4076 12089 4107
rect 11846 4073 12055 4076
rect 10944 4057 12055 4073
rect 10607 3966 10713 4000
rect 12366 4088 12368 4115
rect 10831 4000 10835 4012
rect 10797 3978 10835 4000
rect 12055 4003 12089 4042
rect 11017 3987 11051 4003
rect 10607 3932 10641 3966
rect 10675 3932 10713 3966
rect 10607 3898 10713 3932
rect 10607 3864 10641 3898
rect 10675 3864 10713 3898
rect 10607 3830 10713 3864
rect 10607 3799 10641 3830
rect 10675 3799 10713 3830
rect 10675 3796 10679 3799
rect 10641 3765 10679 3796
rect 10797 3966 10831 3978
rect 10797 3898 10831 3932
rect 10797 3830 10831 3864
rect 11017 3819 11051 3953
rect 11873 3987 12021 4003
rect 11907 3983 12021 3987
rect 11873 3949 11879 3953
rect 11913 3949 11951 3983
rect 11985 3949 12021 3983
rect 11873 3937 12021 3949
rect 10797 3780 10831 3796
rect 10908 3765 10946 3799
rect 10980 3765 10982 3799
rect 11017 3769 11051 3785
rect 11873 3834 11907 3835
rect 11873 3819 11945 3834
rect 11907 3785 11945 3819
rect 10550 3689 10588 3723
rect 10713 3689 10751 3723
rect 10785 3689 10786 3718
rect 9190 3636 9206 3670
rect 9240 3636 9276 3670
rect 9310 3636 9345 3670
rect 9379 3636 9414 3670
rect 9448 3636 9483 3670
rect 9517 3636 9552 3670
rect 9586 3636 9722 3670
rect 9782 3636 9798 3670
rect 9832 3636 9869 3670
rect 9903 3636 9940 3670
rect 9974 3636 10012 3670
rect 10046 3636 10084 3670
rect 10118 3636 10156 3670
rect 10190 3636 10228 3670
rect 10262 3636 10300 3670
rect 10334 3636 10350 3670
rect 10580 3669 10614 3689
rect 9190 3632 9722 3636
rect 8785 3573 8851 3607
rect 8885 3573 8951 3607
rect 8751 3533 8985 3573
rect 10483 3571 10517 3609
rect 8785 3499 8851 3533
rect 8885 3499 8951 3533
rect 8751 3459 8985 3499
rect 8785 3425 8851 3459
rect 8885 3425 8951 3459
rect 8751 3385 8985 3425
rect 8785 3351 8851 3385
rect 8885 3351 8951 3385
rect 8751 3311 8985 3351
rect 8785 3277 8851 3311
rect 8885 3277 8951 3311
rect 8751 3253 8985 3277
rect 9443 3518 9509 3537
rect 9477 3513 9515 3518
rect 9493 3484 9515 3513
rect 9640 3514 9674 3537
rect 9443 3479 9459 3484
rect 9493 3479 9509 3484
rect 9443 3412 9509 3479
rect 9443 3378 9459 3412
rect 9493 3378 9509 3412
rect 9443 3311 9509 3378
rect 9443 3277 9459 3311
rect 9493 3277 9509 3311
rect 9443 3253 9509 3277
rect 10136 3499 10170 3537
rect 9640 3440 9674 3465
rect 9640 3366 9674 3406
rect 9640 3292 9674 3332
rect 8166 3211 8200 3246
rect 8400 3211 8414 3245
rect 8486 3211 8510 3245
rect 8544 3211 8560 3245
rect 9640 3218 9674 3258
rect 7908 3092 7920 3126
rect 7954 3092 7992 3126
rect 3292 3037 3348 3071
rect 3292 3023 3382 3037
rect 3464 3067 4752 3075
rect 3464 3033 3488 3067
rect 3522 3033 3559 3067
rect 3593 3033 3630 3067
rect 3664 3033 3701 3067
rect 3735 3033 3772 3067
rect 3806 3033 3843 3067
rect 3877 3033 3914 3067
rect 3948 3033 3985 3067
rect 4019 3033 4056 3067
rect 4090 3033 4127 3067
rect 4161 3033 4198 3067
rect 4232 3033 4269 3067
rect 4303 3033 4340 3067
rect 4374 3033 4411 3067
rect 4445 3033 4482 3067
rect 4516 3033 4553 3067
rect 4587 3033 4624 3067
rect 4658 3033 4694 3067
rect 4728 3033 4752 3067
rect 3464 3025 4752 3033
rect 3348 3021 3382 3023
rect -314 2974 -280 2987
rect -314 2903 -280 2919
rect 271 2981 305 3015
rect 271 2913 305 2947
rect -135 2837 -111 2871
rect -77 2837 -50 2871
rect -16 2837 6 2871
rect 56 2837 64 2871
rect 271 2845 305 2879
rect 1801 2943 1823 2977
rect 1869 2943 1895 2977
rect 1937 2943 1967 2977
rect 2005 2943 2039 2977
rect 2073 2943 2107 2977
rect 2145 2943 2175 2977
rect 2217 2943 2243 2977
rect 2289 2943 2311 2977
rect 2361 2943 2379 2977
rect 2433 2943 2447 2977
rect 2505 2943 2515 2977
rect 2577 2943 2583 2977
rect 2649 2943 2651 2977
rect 2685 2943 2687 2977
rect 2753 2943 2759 2977
rect 2821 2943 2831 2977
rect 2889 2943 2903 2977
rect 2957 2943 2975 2977
rect 3025 2943 3047 2977
rect 3093 2943 3119 2977
rect 3161 2943 3191 2977
rect 3229 2943 3263 2977
rect 3297 2974 3313 2977
rect 7519 2974 7553 3086
rect 7604 3052 7868 3092
rect 7587 3018 7603 3052
rect 7637 3018 7671 3052
rect 7705 3018 7941 3052
rect 7975 3018 8009 3052
rect 8043 3018 8293 3052
rect 8327 3018 8361 3052
rect 8395 3018 8411 3052
rect 8486 2974 8552 3211
rect 9640 3144 9674 3184
rect 3297 2943 3358 2974
rect 1751 2940 3358 2943
rect 3392 2940 3432 2974
rect 3466 2940 3506 2974
rect 3540 2940 3580 2974
rect 3614 2940 3654 2974
rect 3688 2940 3728 2974
rect 3762 2940 3802 2974
rect 3836 2940 3876 2974
rect 3910 2940 3950 2974
rect 3984 2940 4024 2974
rect 4058 2940 4098 2974
rect 4132 2940 4172 2974
rect 4206 2940 4246 2974
rect 4280 2940 4320 2974
rect 4354 2940 4394 2974
rect 4428 2940 4468 2974
rect 4502 2940 4541 2974
rect 4575 2940 4614 2974
rect 4648 2940 4687 2974
rect 4721 2940 4760 2974
rect 4794 2940 4833 2974
rect 4867 2940 4906 2974
rect 7519 2958 7576 2974
rect 7718 2968 7752 2974
rect 1751 2871 4908 2940
rect 7519 2924 7542 2958
rect 7519 2890 7576 2924
rect 271 2777 305 2811
rect 7519 2856 7542 2890
rect 7519 2822 7576 2856
rect 7519 2788 7542 2822
rect 7519 2772 7576 2788
rect 7714 2958 7752 2968
rect 7714 2934 7718 2958
rect 7680 2924 7718 2934
rect 7752 2924 7786 2934
rect 7680 2890 7786 2924
rect 7680 2856 7718 2890
rect 7752 2856 7786 2890
rect 7680 2822 7786 2856
rect 7680 2788 7718 2822
rect 7752 2788 7786 2822
rect 7680 2772 7786 2788
rect 7894 2958 8036 2974
rect 7928 2924 8036 2958
rect 7894 2890 8036 2924
rect 7928 2856 8036 2890
rect 7894 2822 8036 2856
rect 7928 2788 8036 2822
rect 7894 2772 8036 2788
rect 8070 2968 8104 2974
rect 8104 2934 8142 2968
rect 8104 2924 8176 2934
rect 8070 2890 8176 2924
rect 8104 2856 8176 2890
rect 8070 2822 8176 2856
rect 8104 2788 8176 2822
rect 8070 2772 8176 2788
rect 8246 2958 8386 2974
rect 8280 2924 8386 2958
rect 8246 2890 8386 2924
rect 8280 2856 8386 2890
rect 8246 2822 8386 2856
rect 8280 2788 8386 2822
rect 8246 2772 8386 2788
rect 271 2709 305 2743
rect 7760 2713 7776 2722
rect 7810 2713 7844 2722
rect -453 2651 -419 2669
rect -453 2583 -419 2617
rect -453 2521 -419 2549
rect -453 2449 -419 2481
rect -453 2389 -419 2415
rect -453 2321 -419 2355
rect -453 2253 -419 2287
rect -453 1991 -419 2219
rect -277 2651 -243 2663
rect -277 2583 -243 2591
rect -277 2515 -243 2549
rect -277 2389 -243 2481
rect -277 2321 -243 2355
rect -277 2253 -243 2287
rect -277 2203 -243 2219
rect -101 2651 -67 2669
rect -101 2583 -67 2617
rect -101 2515 -67 2549
rect -101 2424 -67 2481
rect -101 2389 -67 2390
rect -101 2352 -67 2355
rect -101 2253 -67 2287
rect -382 2119 -366 2153
rect -329 2119 -316 2153
rect -382 2085 -316 2119
rect -382 2051 -366 2085
rect -332 2081 -316 2085
rect -329 2051 -316 2081
rect -202 2119 -186 2153
rect -149 2119 -136 2153
rect -202 2085 -136 2119
rect -202 2051 -186 2085
rect -152 2081 -136 2085
rect -149 2051 -136 2081
rect -453 1923 -419 1957
rect -453 1873 -419 1889
rect -277 1991 -243 2007
rect -277 1946 -243 1957
rect -101 1980 -67 2219
rect 75 2651 109 2663
rect 75 2583 109 2591
rect 75 2515 109 2549
rect 75 2389 109 2481
rect 75 2321 109 2355
rect 75 2253 109 2287
rect 75 2203 109 2219
rect 7718 2679 7756 2713
rect 7810 2688 7828 2713
rect 7878 2688 7894 2722
rect 7790 2679 7828 2688
rect 271 2641 305 2675
rect 7928 2642 8036 2772
rect 8112 2688 8122 2722
rect 8162 2688 8194 2722
rect 8230 2688 8246 2722
rect 8280 2710 8386 2772
rect 8456 2940 8494 2974
rect 8528 2940 8552 2974
rect 8586 3092 8639 3126
rect 8673 3092 8711 3126
rect 8745 3092 8783 3126
rect 8817 3092 8855 3126
rect 8889 3092 8927 3126
rect 8961 3092 8999 3126
rect 9033 3092 9071 3126
rect 9105 3092 9143 3126
rect 9177 3092 9215 3126
rect 9249 3092 9287 3126
rect 9321 3092 9359 3126
rect 9393 3092 9426 3126
rect 8586 3052 9426 3092
rect 8586 3018 8628 3052
rect 8662 3018 8696 3052
rect 8730 3018 8764 3052
rect 8798 3018 8832 3052
rect 8866 3018 8900 3052
rect 8934 3018 8968 3052
rect 9002 3018 9036 3052
rect 9070 3018 9104 3052
rect 9138 3018 9172 3052
rect 9206 3018 9240 3052
rect 9274 3018 9308 3052
rect 9342 3018 9376 3052
rect 9410 3018 9426 3052
rect 9756 3460 9790 3476
rect 9756 3392 9790 3426
rect 9756 3324 9790 3358
rect 9756 3256 9790 3290
rect 9756 3188 9790 3222
rect 9756 3126 9790 3154
rect 10580 3601 10614 3635
rect 10580 3551 10614 3567
rect 10679 3669 10786 3689
rect 10679 3635 10719 3669
rect 10753 3635 10786 3669
rect 10679 3601 10786 3635
rect 10679 3567 10719 3601
rect 10753 3567 10786 3601
rect 10483 3499 10517 3537
rect 10136 3460 10170 3465
rect 10136 3392 10170 3426
rect 10136 3324 10170 3358
rect 10136 3256 10170 3290
rect 10136 3188 10170 3222
rect 9640 3070 9674 3110
rect 9763 3120 9801 3126
rect 9790 3092 9801 3120
rect 10136 3120 10170 3154
rect 8456 2924 8528 2940
rect 8422 2890 8528 2924
rect 8456 2856 8528 2890
rect 8422 2822 8528 2856
rect 8456 2788 8528 2822
rect 8422 2771 8528 2788
rect 8314 2676 8352 2710
rect 8586 2642 8644 3018
rect 9640 2996 9674 3036
rect 8678 2958 8712 2974
rect 8678 2894 8712 2924
rect 8934 2968 9040 2975
rect 8968 2934 9006 2968
rect 8968 2924 9040 2934
rect 8712 2860 8750 2894
rect 8934 2890 9040 2924
rect 8678 2822 8712 2856
rect 8678 2772 8712 2788
rect 8968 2856 9040 2890
rect 8934 2822 9040 2856
rect 8968 2788 9040 2822
rect 8934 2771 9040 2788
rect 9190 2958 9224 2974
rect 9446 2968 9480 2974
rect 9396 2934 9434 2968
rect 9468 2958 9480 2968
rect 9640 2938 9674 2962
rect 9756 3052 9790 3086
rect 9756 2984 9790 3018
rect 9190 2890 9224 2924
rect 9446 2890 9480 2924
rect 9226 2856 9264 2890
rect 9190 2822 9224 2856
rect 9190 2772 9224 2788
rect 9446 2822 9480 2856
rect 9446 2772 9480 2788
rect 9756 2750 9790 2950
rect 10136 3052 10170 3086
rect 10136 2984 10170 3018
rect 10136 2934 10170 2950
rect 10326 3460 10360 3476
rect 10483 3428 10517 3465
rect 10326 3392 10360 3426
rect 10326 3324 10360 3358
rect 10326 3256 10360 3290
rect 10326 3188 10360 3222
rect 10326 3120 10360 3154
rect 10326 3052 10360 3086
rect 10326 2984 10360 3018
rect 9858 2890 9896 2894
rect 9842 2856 9858 2860
rect 9892 2860 9896 2890
rect 10031 2890 10069 2894
rect 10031 2860 10034 2890
rect 9892 2856 9908 2860
rect 9842 2822 9908 2856
rect 9842 2788 9858 2822
rect 9892 2788 9908 2822
rect 10018 2856 10034 2860
rect 10068 2860 10069 2890
rect 10068 2856 10084 2860
rect 10018 2822 10084 2856
rect 10018 2788 10034 2822
rect 10068 2788 10084 2822
rect 10195 2856 10211 2890
rect 10245 2856 10261 2890
rect 10195 2822 10261 2856
rect 10195 2788 10211 2822
rect 10245 2788 10261 2822
rect 10326 2812 10360 2950
rect 10442 3404 10517 3428
rect 10476 3370 10517 3404
rect 10442 3336 10517 3370
rect 10476 3302 10517 3336
rect 10442 3268 10517 3302
rect 10679 3326 10786 3567
rect 10874 3616 10982 3765
rect 11873 3737 11945 3785
rect 11062 3693 11862 3699
rect 11062 3659 11078 3693
rect 11112 3659 11151 3693
rect 11185 3659 11224 3693
rect 11258 3659 11297 3693
rect 11331 3659 11370 3693
rect 11404 3659 11443 3693
rect 11477 3659 11516 3693
rect 11550 3659 11590 3693
rect 11624 3659 11664 3693
rect 11698 3659 11738 3693
rect 11772 3659 11812 3693
rect 11846 3659 11862 3693
rect 11062 3653 11862 3659
rect 11904 3673 11945 3737
rect 11979 3769 12021 3937
rect 12055 3930 12089 3969
rect 12132 4025 12332 4070
rect 12132 3991 12149 4025
rect 12183 3991 12332 4025
rect 12132 3958 12332 3991
rect 12055 3857 12089 3896
rect 12055 3807 12089 3823
rect 12134 3892 12200 3897
rect 12134 3858 12145 3892
rect 12179 3858 12200 3892
rect 12134 3820 12200 3858
rect 12134 3786 12145 3820
rect 12179 3786 12200 3820
rect 12134 3769 12200 3786
rect 11979 3735 12149 3769
rect 12183 3735 12200 3769
rect 11979 3707 12200 3735
rect 10874 3567 11051 3616
rect 10874 3533 11017 3567
rect 10874 3516 11051 3533
rect 11433 3473 11728 3653
rect 11904 3645 12199 3673
rect 11904 3641 12149 3645
rect 12183 3641 12199 3645
rect 11904 3617 11937 3641
rect 11971 3607 12011 3641
rect 12045 3607 12084 3641
rect 12118 3611 12149 3641
rect 12118 3607 12157 3611
rect 12191 3607 12199 3641
rect 11873 3567 11911 3583
rect 11907 3533 11949 3567
rect 11072 3472 11820 3473
rect 11072 3438 11088 3472
rect 11122 3438 11157 3472
rect 11191 3438 11226 3472
rect 11260 3438 11294 3472
rect 11328 3438 11362 3472
rect 11396 3438 11430 3472
rect 11464 3438 11498 3472
rect 11532 3438 11566 3472
rect 11600 3438 11634 3472
rect 11668 3438 11702 3472
rect 11736 3438 11770 3472
rect 11804 3438 11820 3472
rect 11072 3437 11820 3438
rect 10679 3292 10680 3326
rect 10714 3292 10752 3326
rect 10679 3286 10786 3292
rect 10892 3379 10930 3413
rect 10964 3379 10983 3413
rect 10476 3234 10517 3268
rect 10442 3200 10517 3234
rect 10476 3166 10517 3200
rect 10858 3209 10983 3379
rect 11017 3351 11051 3367
rect 11051 3317 11256 3343
rect 11017 3316 11256 3317
rect 11017 3282 11149 3316
rect 11183 3282 11221 3316
rect 11255 3282 11256 3316
rect 11017 3277 11256 3282
rect 11138 3209 11180 3225
rect 11214 3209 11256 3225
rect 11290 3209 11331 3225
rect 11433 3209 11728 3437
rect 11873 3351 11949 3533
rect 11983 3539 12089 3573
rect 11983 3505 12055 3539
rect 11983 3454 12089 3505
rect 11983 3420 12055 3454
rect 11983 3419 12089 3420
rect 12017 3385 12055 3419
rect 12235 3389 12332 3958
rect 11907 3317 11949 3351
rect 11873 3301 11949 3317
rect 12133 3355 12149 3389
rect 12183 3355 12332 3389
rect 12133 3293 12332 3355
rect 12400 4054 12402 4081
rect 12366 4040 12402 4054
rect 12366 4020 12368 4040
rect 12400 3986 12402 4006
rect 12366 3965 12402 3986
rect 12366 3952 12368 3965
rect 12400 3918 12402 3931
rect 12366 3890 12402 3918
rect 12366 3884 12368 3890
rect 12400 3850 12402 3856
rect 12366 3816 12402 3850
rect 12400 3815 12402 3816
rect 12366 3781 12368 3782
rect 12366 3748 12400 3781
rect 12366 3680 12400 3714
rect 12366 3643 12400 3646
rect 13847 3585 13901 4563
rect 12366 3571 12400 3578
rect 12366 3499 12400 3510
rect 12366 3408 12400 3442
rect 12366 3340 12400 3356
rect 12366 3272 12400 3284
rect 11842 3209 11884 3225
rect 11918 3209 11960 3225
rect 11994 3209 12035 3225
rect 10858 3175 10897 3209
rect 10931 3175 10975 3209
rect 11009 3175 11025 3209
rect 11081 3175 11097 3209
rect 11138 3191 11174 3209
rect 11214 3191 11251 3209
rect 11290 3191 11327 3209
rect 11365 3191 11377 3209
rect 11131 3175 11174 3191
rect 11208 3175 11251 3191
rect 11285 3175 11327 3191
rect 11361 3175 11377 3191
rect 11433 3175 11449 3209
rect 11483 3175 11526 3209
rect 11560 3175 11603 3209
rect 11637 3175 11679 3209
rect 11713 3175 11729 3209
rect 11785 3175 11801 3209
rect 11842 3191 11877 3209
rect 11918 3191 11954 3209
rect 11994 3191 12031 3209
rect 12069 3191 12081 3209
rect 11835 3175 11877 3191
rect 11911 3175 11954 3191
rect 11988 3175 12031 3191
rect 12065 3175 12081 3191
rect 12366 3204 12400 3212
rect 10442 3132 10517 3166
rect 10476 3098 10517 3132
rect 11433 3145 11728 3175
rect 11433 3111 11493 3145
rect 11527 3111 11565 3145
rect 11599 3111 11728 3145
rect 11433 3109 11728 3111
rect 12366 3136 12400 3140
rect 10442 3064 10517 3098
rect 10476 3030 10517 3064
rect 10442 2996 10517 3030
rect 10476 2962 10517 2996
rect 10442 2938 10517 2962
rect 10744 3073 10894 3097
rect 10778 3049 10894 3073
rect 10778 3012 10860 3049
rect 10744 3005 10894 3012
rect 10778 2981 10894 3005
rect 10778 2940 10860 2981
rect 10744 2937 10894 2940
rect 10778 2913 10894 2937
rect 10778 2903 10860 2913
rect 10744 2879 10860 2903
rect 10744 2869 10894 2879
rect 10778 2845 10894 2869
rect 10778 2835 10860 2845
rect 10195 2750 10261 2788
rect 10345 2778 10383 2812
rect 10744 2811 10860 2835
rect 10744 2801 10894 2811
rect 271 2573 305 2607
rect 271 2505 305 2539
rect 7528 2595 7562 2611
rect 7664 2608 7680 2642
rect 7714 2608 7748 2642
rect 7782 2608 7816 2642
rect 7850 2608 7884 2642
rect 7918 2608 7952 2642
rect 7986 2608 8020 2642
rect 8054 2608 8088 2642
rect 8122 2608 8156 2642
rect 8190 2608 8224 2642
rect 8258 2608 8292 2642
rect 8326 2608 8360 2642
rect 8394 2608 8428 2642
rect 8462 2608 8496 2642
rect 8530 2608 8564 2642
rect 8598 2608 8644 2642
rect 8678 2696 8712 2712
rect 8678 2628 8712 2662
rect 7528 2527 7562 2561
rect 8678 2560 8712 2594
rect 7562 2493 7596 2510
rect 7558 2476 7596 2493
rect 8678 2492 8712 2526
rect 271 2437 305 2471
rect 7664 2432 7680 2466
rect 7714 2432 7748 2466
rect 7782 2432 7816 2466
rect 7850 2432 7884 2466
rect 7918 2432 7952 2466
rect 7986 2436 8020 2466
rect 8054 2436 8088 2466
rect 8122 2436 8156 2466
rect 7986 2432 7997 2436
rect 8054 2432 8069 2436
rect 8122 2432 8141 2436
rect 8190 2432 8224 2466
rect 8258 2432 8292 2466
rect 8326 2432 8360 2466
rect 8394 2432 8428 2466
rect 8462 2432 8496 2466
rect 8530 2432 8564 2466
rect 8598 2458 8678 2466
rect 8888 2694 8926 2728
rect 9756 2716 10261 2750
rect 8854 2628 8888 2662
rect 9756 2666 9790 2682
rect 9046 2642 9084 2652
rect 9118 2642 9156 2652
rect 9190 2642 9228 2652
rect 9262 2642 9300 2652
rect 9334 2642 9372 2652
rect 9406 2642 9444 2652
rect 8952 2608 8968 2642
rect 9002 2618 9012 2642
rect 9070 2618 9084 2642
rect 9138 2618 9156 2642
rect 9206 2618 9228 2642
rect 9274 2618 9300 2642
rect 9342 2618 9372 2642
rect 9002 2608 9036 2618
rect 9070 2608 9104 2618
rect 9138 2608 9172 2618
rect 9206 2608 9240 2618
rect 9274 2608 9308 2618
rect 9342 2608 9376 2618
rect 9410 2608 9444 2642
rect 9478 2613 9632 2642
rect 9478 2608 9598 2613
rect 8854 2560 8888 2594
rect 8854 2492 8888 2526
rect 9598 2545 9632 2579
rect 8712 2458 8720 2466
rect 8598 2432 8720 2458
rect 7664 2430 7997 2432
rect 271 2369 305 2403
rect 8031 2402 8069 2432
rect 8103 2402 8141 2432
rect 8175 2430 8720 2432
rect 271 2301 305 2335
rect 271 2233 305 2267
rect 271 2165 305 2199
rect -31 2119 -15 2153
rect 24 2119 35 2153
rect -31 2085 35 2119
rect -31 2051 -15 2085
rect 19 2081 35 2085
rect 24 2051 35 2081
rect 271 2097 305 2131
rect 271 2029 305 2063
rect 75 1991 109 2007
rect -101 1957 75 1980
rect -101 1946 109 1957
rect -277 1874 -243 1889
rect 70 1923 109 1946
rect 70 1889 75 1923
rect 70 1873 109 1889
rect 271 1961 305 1995
rect 271 1893 305 1927
rect 271 1825 305 1859
rect -433 1745 -423 1779
rect -375 1745 -344 1779
rect -297 1745 -265 1779
rect -219 1745 -187 1779
rect -141 1745 -109 1779
rect -63 1745 -31 1779
rect 14 1745 47 1779
rect 91 1745 115 1779
rect 271 1757 305 1791
rect 271 1689 305 1723
rect 7452 2386 7737 2390
rect 7452 2352 7619 2386
rect 7653 2352 7687 2386
rect 7721 2352 7737 2386
rect 7803 2352 7819 2386
rect 7853 2352 7887 2386
rect 7921 2352 7937 2386
rect 7452 2346 7737 2352
rect 7452 1678 7516 2346
rect 9046 2486 9084 2510
rect 9118 2486 9156 2510
rect 9190 2486 9228 2510
rect 9262 2486 9300 2510
rect 9334 2486 9372 2510
rect 9406 2486 9444 2510
rect 9598 2495 9632 2511
rect 9756 2598 9790 2632
rect 9756 2560 9790 2564
rect 9756 2488 9790 2496
rect 8854 2424 8888 2458
rect 8952 2452 8968 2486
rect 9002 2476 9012 2486
rect 9070 2476 9084 2486
rect 9138 2476 9156 2486
rect 9206 2476 9228 2486
rect 9274 2476 9300 2486
rect 9342 2476 9372 2486
rect 9002 2452 9036 2476
rect 9070 2452 9104 2476
rect 9138 2452 9172 2476
rect 9206 2452 9240 2476
rect 9274 2452 9308 2476
rect 9342 2452 9376 2476
rect 9410 2452 9444 2486
rect 9478 2452 9494 2486
rect 9946 2666 9980 2716
rect 9946 2598 9980 2632
rect 9946 2530 9980 2564
rect 9946 2480 9980 2496
rect 10136 2666 10170 2682
rect 10136 2598 10170 2632
rect 10136 2560 10170 2564
rect 10136 2488 10170 2496
rect 10326 2666 10360 2778
rect 10326 2598 10360 2632
rect 10326 2530 10360 2564
rect 10778 2777 10894 2801
rect 10778 2767 10860 2777
rect 10744 2743 10860 2767
rect 10744 2732 10894 2743
rect 10778 2709 10894 2732
rect 10778 2698 10860 2709
rect 10744 2675 10860 2698
rect 10744 2663 10894 2675
rect 10778 2641 10894 2663
rect 10778 2629 10860 2641
rect 10744 2607 10860 2629
rect 10744 2594 10894 2607
rect 10778 2573 10894 2594
rect 10778 2560 10860 2573
rect 10744 2539 10860 2560
rect 10744 2536 10894 2539
rect 10860 2523 10894 2536
rect 11036 3049 11070 3065
rect 11036 2981 11070 3015
rect 11036 2913 11070 2947
rect 11036 2845 11070 2879
rect 11036 2777 11070 2811
rect 11036 2709 11070 2743
rect 11036 2641 11070 2675
rect 11036 2573 11070 2607
rect 11036 2510 11070 2539
rect 11212 3049 11246 3065
rect 11212 2981 11246 3012
rect 11212 2913 11246 2940
rect 11212 2845 11246 2879
rect 11212 2777 11246 2811
rect 11212 2709 11246 2743
rect 11212 2641 11246 2675
rect 11212 2573 11246 2607
rect 11212 2523 11246 2539
rect 11388 3049 11422 3065
rect 11388 2981 11422 3015
rect 11388 2913 11422 2947
rect 11388 2845 11422 2879
rect 11388 2777 11422 2811
rect 11388 2709 11422 2743
rect 11388 2641 11422 2675
rect 11388 2573 11422 2607
rect 11388 2510 11422 2539
rect 11564 3049 11598 3065
rect 11564 2981 11598 3012
rect 11564 2913 11598 2940
rect 11564 2845 11598 2879
rect 11564 2777 11598 2811
rect 11564 2709 11598 2743
rect 11564 2641 11598 2675
rect 11564 2573 11598 2607
rect 11564 2523 11598 2539
rect 11740 3049 11774 3065
rect 11740 2981 11774 3015
rect 11740 2913 11774 2947
rect 11740 2845 11774 2879
rect 11740 2777 11774 2811
rect 11740 2709 11774 2743
rect 11740 2641 11774 2675
rect 11740 2573 11774 2607
rect 11740 2510 11774 2539
rect 11916 3049 11950 3065
rect 11916 2981 11950 3012
rect 11916 2913 11950 2940
rect 11916 2845 11950 2879
rect 11916 2777 11950 2811
rect 11916 2709 11950 2743
rect 11916 2641 11950 2675
rect 11916 2573 11950 2607
rect 11916 2523 11950 2539
rect 12092 3049 12126 3065
rect 12092 2981 12126 3015
rect 12092 2913 12126 2947
rect 12092 2845 12126 2879
rect 12092 2777 12126 2811
rect 12092 2709 12126 2743
rect 12092 2641 12126 2675
rect 12092 2573 12126 2607
rect 12092 2510 12126 2539
rect 12366 3030 12400 3034
rect 12366 2958 12400 2966
rect 12366 2886 12400 2898
rect 12366 2814 12400 2830
rect 12366 2742 12400 2762
rect 12366 2660 12400 2694
rect 12366 2592 12400 2626
rect 12366 2524 12400 2558
rect 10326 2480 10360 2496
rect 11045 2476 11083 2510
rect 11389 2476 11427 2510
rect 11743 2476 11781 2510
rect 12087 2476 12125 2510
rect 12366 2456 12400 2490
rect 12366 2413 12400 2422
rect 8854 2356 8888 2390
rect 9002 2356 9018 2390
rect 9052 2356 9086 2390
rect 9120 2356 9136 2390
rect 9202 2356 9218 2390
rect 9252 2356 9286 2390
rect 9320 2356 9628 2390
rect 9722 2356 9738 2390
rect 9772 2356 9806 2390
rect 9840 2356 9874 2390
rect 9908 2356 9942 2390
rect 9976 2356 9992 2390
rect 10074 2356 10090 2390
rect 10124 2356 10158 2390
rect 10192 2356 10226 2390
rect 10260 2356 10294 2390
rect 10328 2356 10344 2390
rect 10784 2360 10818 2376
rect 271 1621 305 1655
rect 7451 1636 7516 1678
rect 7578 2295 7612 2311
rect 7578 2227 7612 2261
rect 7578 2159 7612 2193
rect 7578 2091 7612 2125
rect 7578 2023 7612 2057
rect 7578 1955 7612 1989
rect 7578 1887 7612 1921
rect 7578 1819 7612 1853
rect 7578 1640 7612 1785
rect 7754 2295 7788 2311
rect 7754 2227 7788 2261
rect 7754 2159 7788 2193
rect 7754 2091 7788 2125
rect 7754 2023 7788 2057
rect 7754 1955 7788 1989
rect 7754 1887 7788 1921
rect 7754 1819 7788 1853
rect 7754 1769 7788 1785
rect 7930 2295 7964 2311
rect 7930 2227 7964 2261
rect 7930 2159 7964 2193
rect 7930 2091 7964 2125
rect 7930 2023 7964 2057
rect 7930 1955 7964 1985
rect 7930 1887 7964 1913
rect 7930 1819 7964 1841
rect 7930 1769 7964 1785
rect 8678 2288 8712 2322
rect 8678 2220 8712 2254
rect 8678 2152 8712 2186
rect 8678 2084 8712 2118
rect 8678 2018 8712 2050
rect 8678 1948 8712 1982
rect 8678 1880 8712 1912
rect 8678 1812 8712 1840
rect 8678 1762 8712 1778
rect 8854 2288 8888 2322
rect 8854 2220 8888 2254
rect 8854 2152 8888 2186
rect 8854 2084 8888 2118
rect 8854 2016 8888 2050
rect 8854 1948 8888 1982
rect 8854 1880 8888 1914
rect 8854 1812 8888 1846
rect 8854 1762 8888 1778
rect 8977 2296 9011 2312
rect 8977 2228 9011 2262
rect 8977 2160 9011 2194
rect 8977 2092 9011 2126
rect 8977 2024 9011 2058
rect 8977 1956 9011 1978
rect 8977 1888 9011 1906
rect 8977 1820 9011 1834
rect 8977 1770 9011 1786
rect 9045 1722 9119 2356
rect 8471 1686 8547 1720
rect 8581 1686 8619 1720
rect 8653 1686 8673 1720
rect 8471 1651 8673 1686
rect 8723 1686 8746 1720
rect 8780 1686 8818 1720
rect 8852 1686 8857 1720
rect 8723 1660 8857 1686
rect 271 1553 305 1587
rect 7410 1602 7426 1636
rect 7460 1602 7494 1636
rect 7528 1602 7544 1636
rect 7578 1606 7632 1640
rect 7826 1612 7840 1646
rect 7874 1640 7912 1646
rect 7826 1606 7842 1612
rect 7876 1606 7910 1640
rect 7946 1612 7960 1646
rect 8173 1612 8184 1627
rect 8218 1612 8256 1646
rect 8290 1612 8307 1627
rect 8723 1626 8739 1660
rect 8773 1626 8807 1660
rect 8841 1626 8857 1660
rect 8936 1688 8947 1722
rect 8981 1688 9019 1722
rect 9053 1688 9119 1722
rect 9153 2296 9258 2312
rect 9187 2262 9258 2296
rect 9153 2228 9258 2262
rect 9187 2194 9258 2228
rect 9153 2160 9258 2194
rect 9187 2126 9258 2160
rect 9153 2092 9258 2126
rect 9187 2058 9258 2092
rect 9153 2024 9258 2058
rect 9187 1990 9258 2024
rect 9153 1956 9258 1990
rect 9187 1922 9258 1956
rect 9153 1888 9258 1922
rect 9187 1854 9258 1888
rect 9153 1820 9258 1854
rect 9187 1786 9258 1820
rect 9153 1736 9258 1786
rect 9329 2296 9363 2312
rect 9329 2228 9363 2262
rect 9329 2160 9363 2194
rect 9329 2092 9363 2126
rect 9329 2024 9363 2058
rect 9445 2284 9547 2308
rect 9479 2250 9513 2284
rect 9445 2210 9547 2250
rect 9479 2176 9513 2210
rect 9445 2136 9547 2176
rect 9479 2102 9513 2136
rect 9445 2062 9547 2102
rect 9479 2028 9513 2062
rect 9445 2013 9547 2028
rect 9329 1956 9363 1978
rect 9329 1888 9363 1906
rect 9329 1820 9363 1834
rect 9329 1770 9363 1786
rect 9479 1806 9513 1835
rect 9445 1766 9547 1806
rect 9153 1702 9386 1736
rect 9479 1732 9513 1766
rect 9445 1708 9547 1732
rect 8936 1659 9119 1688
rect 8936 1625 8952 1659
rect 8986 1625 9020 1659
rect 9054 1625 9088 1659
rect 9122 1625 9138 1659
rect 7944 1606 7960 1612
rect 7410 1572 7544 1602
rect 7410 1538 7426 1572
rect 7460 1538 7498 1572
rect 7532 1538 7544 1572
rect 271 1485 305 1519
rect 271 1417 305 1451
rect 271 1349 305 1383
rect 271 1281 305 1315
rect 271 1213 305 1247
rect 271 1145 305 1179
rect 271 1077 305 1111
rect 271 1009 305 1043
rect 271 941 305 975
rect 271 873 305 907
rect 271 805 305 839
rect 7422 1486 7456 1490
rect 7422 1414 7456 1440
rect 7422 1342 7456 1372
rect 7422 1270 7456 1304
rect 7422 1202 7456 1236
rect 7422 1134 7456 1168
rect 7422 1066 7456 1100
rect 7422 998 7456 1032
rect 7422 930 7456 964
rect 7422 862 7456 896
rect 271 737 305 771
rect 271 669 305 703
rect 271 601 305 635
rect 609 770 633 796
rect 1075 770 1099 796
rect 609 664 621 770
rect 1087 664 1099 770
rect 609 626 633 664
rect 1075 626 1099 664
rect 7422 794 7456 828
rect 7422 726 7456 760
rect 7422 658 7456 692
rect 271 533 305 567
rect 7422 590 7456 624
rect 7422 540 7456 556
rect 271 465 305 499
rect 7496 496 7530 1538
rect 7598 1474 7632 1606
rect 9172 1516 9386 1702
rect 9581 1659 9628 2356
rect 9664 2296 9698 2312
rect 9664 2228 9698 2262
rect 9664 2160 9698 2194
rect 9664 2092 9698 2126
rect 9840 2296 9874 2312
rect 9840 2228 9874 2262
rect 9840 2160 9874 2194
rect 9732 2081 9770 2115
rect 9840 2092 9874 2126
rect 10016 2296 10050 2312
rect 10016 2228 10050 2262
rect 10016 2160 10050 2194
rect 10016 2115 10050 2126
rect 10192 2296 10226 2312
rect 10192 2228 10226 2262
rect 10192 2160 10226 2194
rect 9664 2024 9698 2058
rect 9664 1956 9698 1990
rect 9664 1888 9698 1922
rect 9664 1820 9698 1854
rect 9664 1770 9698 1786
rect 10016 2092 10054 2115
rect 9840 2024 9874 2058
rect 9840 1956 9874 1990
rect 9840 1888 9874 1922
rect 9840 1820 9874 1854
rect 9840 1736 9874 1786
rect 10050 2081 10054 2092
rect 10192 2092 10226 2126
rect 10368 2296 10402 2312
rect 10368 2228 10402 2262
rect 10368 2160 10402 2194
rect 10016 2024 10050 2058
rect 10016 1956 10050 1990
rect 10016 1888 10050 1922
rect 10016 1820 10050 1854
rect 10016 1770 10050 1786
rect 10296 2081 10334 2115
rect 10368 2092 10402 2126
rect 10192 2024 10226 2058
rect 10192 1956 10226 1978
rect 10192 1888 10226 1906
rect 10192 1820 10226 1834
rect 10192 1770 10226 1786
rect 10368 2024 10402 2058
rect 10368 1956 10402 1990
rect 10368 1888 10402 1922
rect 10368 1820 10402 1854
rect 10368 1770 10402 1786
rect 10486 2255 10520 2300
rect 10486 2187 10520 2221
rect 10486 2119 10520 2153
rect 10486 2051 10520 2085
rect 10486 2012 10520 2017
rect 10486 1940 10520 1949
rect 10486 1868 10520 1881
rect 10784 2292 10818 2326
rect 10784 2224 10818 2258
rect 10784 2156 10818 2190
rect 10784 2098 10818 2122
rect 10960 2360 10994 2376
rect 10960 2292 10994 2326
rect 10960 2224 10994 2258
rect 10960 2156 10994 2190
rect 10784 2088 10804 2098
rect 10838 2064 10876 2098
rect 10960 2088 10994 2122
rect 11136 2360 11170 2376
rect 11136 2292 11170 2326
rect 11136 2224 11170 2258
rect 11136 2156 11170 2190
rect 11136 2098 11170 2122
rect 11312 2360 11346 2376
rect 11312 2292 11346 2326
rect 11312 2224 11346 2258
rect 11312 2156 11346 2190
rect 10784 2020 10818 2054
rect 10784 1952 10818 1986
rect 10784 1884 10818 1918
rect 10784 1834 10818 1850
rect 11136 2088 11174 2098
rect 10960 2020 10994 2054
rect 10960 1952 10994 1984
rect 10960 1884 10994 1912
rect 10960 1834 10994 1840
rect 11170 2064 11174 2088
rect 11312 2088 11346 2122
rect 11136 2020 11170 2054
rect 11136 1952 11170 1986
rect 11136 1884 11170 1918
rect 11136 1834 11170 1850
rect 11312 2020 11346 2054
rect 11312 1952 11346 1984
rect 11312 1884 11346 1912
rect 11312 1834 11346 1840
rect 11459 2360 11571 2376
rect 11459 2326 11488 2360
rect 11522 2326 11571 2360
rect 11459 2292 11571 2326
rect 11459 2258 11488 2292
rect 11522 2258 11571 2292
rect 11459 2224 11571 2258
rect 11459 2190 11488 2224
rect 11522 2190 11571 2224
rect 11459 2156 11571 2190
rect 11459 2122 11488 2156
rect 11522 2122 11571 2156
rect 11459 2098 11571 2122
rect 11493 2088 11537 2098
rect 11522 2064 11537 2088
rect 11459 2054 11488 2064
rect 11522 2054 11571 2064
rect 11459 2020 11571 2054
rect 11459 1986 11488 2020
rect 11522 1986 11571 2020
rect 11459 1952 11571 1986
rect 11459 1918 11488 1952
rect 11522 1918 11571 1952
rect 11459 1884 11571 1918
rect 11459 1850 11488 1884
rect 11522 1850 11571 1884
rect 11459 1834 11571 1850
rect 11664 2360 11698 2376
rect 11664 2292 11698 2326
rect 11664 2224 11698 2258
rect 11664 2156 11698 2190
rect 11664 2088 11698 2122
rect 11664 2020 11698 2054
rect 11664 1952 11698 1984
rect 11664 1884 11698 1912
rect 11664 1834 11698 1840
rect 11806 2360 11918 2376
rect 11806 2326 11840 2360
rect 11874 2326 11918 2360
rect 11806 2292 11918 2326
rect 11806 2258 11840 2292
rect 11874 2258 11918 2292
rect 11806 2224 11918 2258
rect 11806 2190 11840 2224
rect 11874 2190 11918 2224
rect 11806 2156 11918 2190
rect 11806 2122 11840 2156
rect 11874 2122 11918 2156
rect 11806 2098 11918 2122
rect 11840 2088 11878 2098
rect 11806 2054 11840 2064
rect 11874 2064 11878 2088
rect 11912 2064 11918 2098
rect 11874 2054 11918 2064
rect 11806 2020 11918 2054
rect 11806 1986 11840 2020
rect 11874 1986 11918 2020
rect 11806 1952 11918 1986
rect 11806 1918 11840 1952
rect 11874 1918 11918 1952
rect 11806 1884 11918 1918
rect 11806 1850 11840 1884
rect 11874 1850 11918 1884
rect 11806 1834 11918 1850
rect 12016 2360 12050 2376
rect 12366 2337 12400 2354
rect 12050 2326 12167 2336
rect 12016 2312 12167 2326
rect 12016 2292 12133 2312
rect 12050 2278 12133 2292
rect 12050 2258 12167 2278
rect 12016 2237 12167 2258
rect 12016 2224 12133 2237
rect 12050 2203 12133 2224
rect 12050 2190 12167 2203
rect 12016 2162 12167 2190
rect 12016 2156 12133 2162
rect 12050 2128 12133 2156
rect 12050 2122 12167 2128
rect 12016 2088 12167 2122
rect 12050 2054 12133 2088
rect 12016 2020 12167 2054
rect 12050 2018 12167 2020
rect 12050 1984 12102 2018
rect 12136 2014 12167 2018
rect 12016 1980 12133 1984
rect 12016 1952 12167 1980
rect 12050 1946 12167 1952
rect 12050 1912 12102 1946
rect 12136 1940 12167 1946
rect 12016 1906 12133 1912
rect 12016 1884 12167 1906
rect 12050 1874 12167 1884
rect 12050 1840 12102 1874
rect 12136 1866 12167 1874
rect 12016 1834 12133 1840
rect 10486 1773 10520 1813
rect 12050 1832 12133 1834
rect 12050 1808 12167 1832
rect 12366 2261 12400 2286
rect 12366 2185 12400 2218
rect 12366 2116 12400 2150
rect 12366 2048 12400 2075
rect 12366 1980 12400 1999
rect 12366 1912 12400 1923
rect 12366 1844 12400 1847
rect 12366 1776 12400 1810
rect 9840 1693 10102 1736
rect 9420 1646 9436 1659
rect 9420 1612 9432 1646
rect 9470 1625 9504 1659
rect 9466 1612 9504 1625
rect 9538 1612 9628 1659
rect 9722 1625 9738 1659
rect 9772 1625 9806 1659
rect 9840 1625 9874 1659
rect 9908 1625 9942 1659
rect 9976 1625 9992 1659
rect 9722 1572 9992 1625
rect 9722 1565 9742 1572
rect 9728 1538 9742 1565
rect 9776 1538 9814 1572
rect 9848 1538 9886 1572
rect 9920 1538 9958 1572
rect 7598 1406 7632 1440
rect 7598 1338 7632 1372
rect 7598 1270 7632 1304
rect 7598 1202 7632 1236
rect 7774 1486 7808 1490
rect 7774 1414 7808 1440
rect 7774 1342 7808 1372
rect 7774 1270 7808 1304
rect 7774 1202 7808 1236
rect 7632 1168 7636 1188
rect 7598 1154 7636 1168
rect 7950 1474 7984 1490
rect 7950 1406 7984 1440
rect 7950 1338 7984 1372
rect 7950 1270 7984 1304
rect 7950 1202 7984 1236
rect 7598 1134 7632 1154
rect 7598 1066 7632 1100
rect 7598 998 7632 1032
rect 7598 930 7632 964
rect 7598 862 7632 896
rect 7598 794 7632 828
rect 7598 726 7632 760
rect 7598 658 7632 692
rect 7598 590 7632 624
rect 7598 540 7632 556
rect 7774 1134 7808 1168
rect 7912 1154 7950 1188
rect 7774 1066 7808 1100
rect 7774 998 7808 1032
rect 7774 930 7808 964
rect 7774 862 7808 896
rect 7774 794 7808 828
rect 7774 726 7808 760
rect 7774 658 7808 692
rect 7774 590 7808 624
rect 7774 540 7808 556
rect 7950 1134 7984 1154
rect 7950 1066 7984 1100
rect 7950 998 7984 1032
rect 7950 930 7984 964
rect 8884 1466 8918 1482
rect 8884 1398 8918 1432
rect 8884 1330 8918 1364
rect 8884 1268 8918 1296
rect 9040 1426 9074 1432
rect 9040 1354 9074 1364
rect 8918 1234 8956 1268
rect 9040 1262 9074 1296
rect 9196 1466 9230 1482
rect 9196 1398 9230 1432
rect 9196 1330 9230 1364
rect 9196 1268 9230 1296
rect 9352 1466 9386 1516
rect 9658 1514 9692 1536
rect 9352 1398 9386 1432
rect 9352 1330 9386 1364
rect 8884 1194 8918 1228
rect 8884 1126 8918 1160
rect 8884 1058 8918 1092
rect 8884 990 8918 1024
rect 8884 940 8918 956
rect 9194 1262 9232 1268
rect 9194 1234 9196 1262
rect 9040 1194 9074 1228
rect 9040 1126 9074 1160
rect 9040 1058 9074 1092
rect 9040 990 9074 1024
rect 9040 940 9074 956
rect 9230 1234 9232 1262
rect 9352 1262 9386 1296
rect 9196 1194 9230 1228
rect 9196 1126 9230 1160
rect 9196 1058 9230 1092
rect 9352 1194 9386 1228
rect 9352 1126 9386 1160
rect 9352 1070 9386 1092
rect 9508 1466 9542 1482
rect 9508 1398 9542 1432
rect 9508 1330 9542 1364
rect 9508 1268 9542 1296
rect 9658 1446 9692 1452
rect 9658 1378 9692 1380
rect 9658 1342 9692 1344
rect 9542 1234 9580 1268
rect 9658 1235 9692 1276
rect 9508 1194 9542 1228
rect 9508 1126 9542 1160
rect 9352 1058 9390 1070
rect 9196 990 9230 1024
rect 9196 940 9230 956
rect 9386 1036 9390 1058
rect 9508 1058 9542 1092
rect 9352 990 9386 1024
rect 9352 940 9386 956
rect 9508 990 9542 1024
rect 9658 1167 9692 1201
rect 9658 1099 9692 1133
rect 9658 1031 9692 1065
rect 9658 956 9692 997
rect 9756 1466 9790 1482
rect 9756 1398 9790 1432
rect 9756 1330 9790 1364
rect 9756 1262 9790 1296
rect 9756 1194 9790 1228
rect 9756 1126 9790 1160
rect 9912 1414 9946 1432
rect 9912 1342 9946 1364
rect 9912 1262 9946 1296
rect 9912 1194 9946 1228
rect 9912 1126 9946 1160
rect 9790 1078 9828 1112
rect 10068 1466 10102 1693
rect 10136 1666 10466 1707
rect 10136 1632 10152 1666
rect 10186 1662 10466 1666
rect 10186 1658 10289 1662
rect 10186 1632 10285 1658
rect 10136 1624 10285 1632
rect 10323 1628 10357 1662
rect 10391 1658 10466 1662
rect 10319 1624 10357 1628
rect 10391 1624 10429 1658
rect 10463 1624 10466 1658
rect 10136 1614 10466 1624
rect 10617 1690 10845 1724
rect 10879 1690 10914 1724
rect 10948 1690 10983 1724
rect 11017 1690 11052 1724
rect 11086 1690 11121 1724
rect 11155 1690 11190 1724
rect 11224 1690 11259 1724
rect 11293 1690 11328 1724
rect 11362 1690 11397 1724
rect 11431 1690 11466 1724
rect 11500 1690 11535 1724
rect 11569 1690 11603 1724
rect 11637 1690 11653 1724
rect 11709 1690 11725 1724
rect 11759 1690 11802 1724
rect 11836 1690 11879 1724
rect 11913 1690 11955 1724
rect 11989 1690 12005 1724
rect 10617 1572 10873 1690
rect 10617 1538 10639 1572
rect 10673 1538 10712 1572
rect 10746 1538 10785 1572
rect 10819 1538 10873 1572
rect 10617 1537 10873 1538
rect 10617 1503 10633 1537
rect 10667 1503 10728 1537
rect 10762 1503 10823 1537
rect 10857 1503 10873 1537
rect 10917 1614 11023 1630
rect 10917 1580 10959 1614
rect 10993 1580 11023 1614
rect 10917 1576 11023 1580
rect 10951 1546 10989 1576
rect 10951 1542 10959 1546
rect 11139 1616 11152 1630
rect 11105 1614 11152 1616
rect 11105 1580 11118 1614
rect 11105 1578 11152 1580
rect 11139 1546 11152 1578
rect 10917 1512 10959 1542
rect 10993 1512 11023 1542
rect 10917 1496 11023 1512
rect 11118 1496 11152 1512
rect 10068 1398 10102 1432
rect 10068 1330 10102 1364
rect 10068 1262 10102 1296
rect 10068 1194 10102 1228
rect 10068 1126 10102 1160
rect 10224 1414 10258 1432
rect 10224 1342 10258 1364
rect 10224 1262 10258 1296
rect 10224 1194 10258 1228
rect 10224 1126 10258 1160
rect 9756 1058 9790 1078
rect 9756 990 9790 1024
rect 9508 940 9542 956
rect 9756 940 9790 956
rect 9912 1058 9946 1092
rect 10056 1092 10068 1112
rect 10056 1078 10094 1092
rect 10380 1466 10414 1482
rect 10380 1398 10414 1432
rect 10380 1330 10414 1364
rect 10380 1262 10414 1296
rect 10380 1194 10414 1228
rect 10380 1126 10414 1160
rect 9912 990 9946 1024
rect 9912 940 9946 956
rect 10068 1058 10102 1078
rect 10068 990 10102 1024
rect 10068 940 10102 956
rect 10224 1058 10258 1092
rect 10330 1078 10368 1112
rect 10402 1078 10414 1092
rect 10224 990 10258 1024
rect 10224 940 10258 956
rect 10380 1058 10414 1078
rect 10380 990 10414 1024
rect 10380 940 10414 956
rect 10489 1458 10526 1492
rect 10455 1413 10526 1458
rect 10489 1379 10526 1413
rect 10455 1334 10526 1379
rect 10489 1300 10526 1334
rect 10455 1255 10526 1300
rect 10489 1221 10526 1255
rect 10455 1176 10526 1221
rect 10561 1443 10667 1459
rect 10561 1409 10572 1443
rect 10606 1409 10667 1443
rect 10561 1375 10667 1409
rect 10561 1341 10572 1375
rect 10606 1341 10667 1375
rect 10561 1307 10667 1341
rect 10561 1273 10572 1307
rect 10606 1273 10667 1307
rect 10561 1268 10667 1273
rect 10595 1239 10633 1268
rect 10606 1234 10633 1239
rect 10561 1205 10572 1234
rect 10606 1205 10667 1234
rect 10561 1189 10667 1205
rect 10702 1443 10762 1460
rect 10702 1409 10728 1443
rect 10702 1375 10762 1409
rect 10702 1341 10728 1375
rect 10702 1307 10762 1341
rect 10702 1273 10728 1307
rect 10702 1239 10762 1273
rect 10702 1205 10728 1239
rect 10489 1142 10526 1176
rect 10455 1078 10526 1142
rect 10455 1054 10530 1078
rect 10455 1020 10496 1054
rect 10455 986 10530 1020
rect 10455 952 10496 986
rect 10455 928 10530 952
rect 9572 896 10211 898
rect 7950 862 7984 896
rect 8963 862 8979 896
rect 9013 862 9025 896
rect 9081 862 9097 896
rect 9149 862 9165 896
rect 9256 862 9272 896
rect 9306 862 9340 896
rect 9386 862 9408 896
rect 9572 862 9855 896
rect 9889 862 9923 896
rect 9957 862 9991 896
rect 10025 862 10059 896
rect 10093 862 10127 896
rect 10161 862 10211 896
rect 7950 794 7984 828
rect 9572 851 10211 862
rect 9572 817 9578 851
rect 9612 817 9651 851
rect 9685 817 9724 851
rect 9758 817 9797 851
rect 9831 817 9870 851
rect 9904 817 9943 851
rect 9977 817 10016 851
rect 10050 817 10088 851
rect 10122 817 10160 851
rect 10194 817 10211 851
rect 10702 835 10762 1205
rect 10884 1443 10918 1459
rect 10884 1375 10918 1409
rect 10884 1307 10918 1341
rect 10884 1239 10918 1273
rect 10884 1189 10918 1205
rect 11040 1443 11074 1459
rect 11040 1375 11074 1388
rect 11040 1307 11074 1316
rect 11040 1239 11074 1273
rect 11040 1189 11074 1205
rect 11156 1443 11262 1459
rect 11156 1409 11196 1443
rect 11230 1409 11262 1443
rect 11709 1431 12005 1690
rect 12366 1708 12400 1742
rect 12366 1640 12400 1674
rect 12366 1572 12400 1606
rect 12366 1504 12400 1538
rect 12366 1436 12400 1458
rect 11156 1375 11262 1409
rect 11414 1397 11430 1431
rect 11464 1397 11499 1431
rect 11533 1397 11568 1431
rect 11602 1397 11637 1431
rect 11671 1397 11706 1431
rect 11740 1397 11775 1431
rect 11809 1397 11844 1431
rect 11878 1397 11913 1431
rect 11947 1397 11982 1431
rect 12016 1397 12051 1431
rect 12085 1397 12120 1431
rect 12154 1397 12170 1431
rect 11156 1341 11196 1375
rect 11230 1341 11262 1375
rect 11156 1307 11262 1341
rect 11156 1273 11196 1307
rect 11230 1273 11262 1307
rect 11156 1268 11262 1273
rect 11190 1239 11228 1268
rect 11190 1234 11196 1239
rect 11156 1205 11196 1234
rect 11230 1205 11262 1234
rect 11156 1189 11262 1205
rect 11311 1337 11403 1353
rect 11311 1303 11369 1337
rect 11311 1287 11403 1303
rect 11311 1100 11377 1287
rect 11709 1253 12081 1397
rect 12225 1349 12259 1387
rect 12225 1287 12259 1303
rect 12366 1368 12400 1386
rect 12366 1300 12400 1314
rect 11709 1219 11791 1253
rect 11825 1219 11872 1253
rect 11906 1219 11953 1253
rect 11987 1219 12034 1253
rect 12068 1219 12081 1253
rect 11709 1217 12081 1219
rect 12366 1232 12400 1266
rect 11414 1183 11430 1217
rect 11464 1183 11503 1217
rect 11537 1183 11576 1217
rect 11610 1183 11649 1217
rect 11683 1183 11722 1217
rect 11756 1183 11795 1217
rect 11829 1183 11868 1217
rect 11902 1183 11942 1217
rect 11976 1183 12016 1217
rect 12050 1183 12090 1217
rect 12124 1183 12164 1217
rect 12198 1183 12214 1217
rect 11709 1171 12081 1183
rect 11709 1156 11791 1171
rect 11825 1137 11872 1171
rect 11906 1137 11953 1171
rect 11987 1137 12034 1171
rect 12068 1137 12081 1171
rect 10827 1043 11377 1100
rect 11814 1115 12081 1137
rect 11814 1081 11843 1115
rect 11877 1081 11922 1115
rect 11956 1081 12000 1115
rect 12034 1081 12081 1115
rect 10827 915 10891 1043
rect 11814 1009 12081 1081
rect 12366 1164 12400 1198
rect 12366 1096 12400 1130
rect 12366 1028 12400 1047
rect 10927 975 10932 1009
rect 10977 975 11011 1009
rect 11046 975 11081 1009
rect 11124 975 11150 1009
rect 11203 975 11219 1009
rect 11282 975 11288 1009
rect 11322 975 11326 1009
rect 11392 975 11404 1009
rect 11462 975 11482 1009
rect 11532 975 11560 1009
rect 11602 975 11638 1009
rect 11672 975 11708 1009
rect 11750 975 11758 1009
rect 11814 975 11830 1009
rect 11864 975 11914 1009
rect 11948 975 11998 1009
rect 12032 975 12081 1009
rect 12115 975 12164 1009
rect 12198 975 12214 1009
rect 10827 881 10857 915
rect 10827 865 10891 881
rect 11313 915 11347 931
rect 11313 835 11347 881
rect 9572 805 10211 817
rect 10725 801 10763 835
rect 11343 801 11381 835
rect 7950 726 7984 760
rect 7950 658 7984 692
rect 10451 691 10467 725
rect 10506 696 10561 730
rect 10595 725 10651 730
rect 10596 696 10651 725
rect 10501 691 10562 696
rect 10596 691 10657 696
rect 10691 691 10707 725
rect 10900 725 10938 726
rect 11145 725 11220 730
rect 11497 725 11695 975
rect 12366 960 12400 974
rect 11769 915 11803 931
rect 11769 865 11803 881
rect 12183 915 12289 931
rect 12183 881 12225 915
rect 12259 881 12289 915
rect 12183 833 12289 881
rect 12217 799 12255 833
rect 12366 892 12400 901
rect 12366 824 12400 828
rect 12366 788 12400 790
rect 12700 1044 12734 1087
rect 12700 967 12734 1010
rect 12700 889 12734 933
rect 12700 811 12734 855
rect 12400 754 12427 763
rect 12366 729 12427 754
rect 10900 692 10935 725
rect 10972 692 11003 725
rect 10919 691 10935 692
rect 10969 691 11003 692
rect 11037 691 11053 725
rect 11108 696 11111 725
rect 11108 691 11124 696
rect 11158 691 11192 725
rect 11226 691 11242 696
rect 11389 691 11405 725
rect 11439 691 11475 725
rect 11509 691 11544 725
rect 11578 691 11613 725
rect 11647 691 11682 725
rect 11716 691 11751 725
rect 11785 691 11801 725
rect 12366 714 12393 729
rect 12700 733 12734 777
rect 12400 680 12427 695
rect 12393 661 12427 680
rect 7950 590 7984 624
rect 10286 618 10320 642
rect 10240 576 10278 610
rect 10312 576 10320 584
rect 7950 540 7984 556
rect 10286 550 10320 576
rect 10406 631 10440 647
rect 10562 631 10596 647
rect 10406 563 10440 597
rect 10560 597 10562 610
rect 10718 631 10752 647
rect 10596 597 10598 610
rect 10560 576 10598 597
rect 10406 520 10440 529
rect 10562 563 10596 576
rect 7480 462 7496 496
rect 7530 462 7564 496
rect 7598 462 7632 496
rect 7666 462 7700 496
rect 7734 462 7750 496
rect 10286 492 10320 516
rect 10404 495 10442 520
rect 10404 486 10406 495
rect 10440 486 10442 495
rect 10562 495 10596 529
rect 10718 563 10752 597
rect 10718 520 10752 529
rect 10908 631 10942 647
rect 11064 631 11098 647
rect 10908 520 10942 597
rect 11060 597 11064 610
rect 11220 631 11254 647
rect 11060 576 11098 597
rect 11344 631 11378 647
rect 11220 520 11254 597
rect 11342 597 11344 610
rect 11500 631 11534 647
rect 11378 597 11380 610
rect 11342 576 11380 597
rect 11656 631 11690 647
rect 11500 520 11534 597
rect 11654 597 11656 610
rect 11690 597 11692 610
rect 11654 576 11692 597
rect 12393 593 12427 627
rect 12393 525 12427 559
rect 10406 445 10440 461
rect 10716 495 10754 520
rect 10716 486 10718 495
rect 10562 445 10596 461
rect 10752 486 10754 495
rect 10909 486 10947 520
rect 11217 486 11255 520
rect 11497 486 11535 520
rect 10718 445 10752 461
rect 12393 457 12427 491
rect 271 349 305 431
rect 339 349 449 383
rect 483 349 517 383
rect 551 349 585 383
rect 619 349 653 383
rect 687 349 721 383
rect 755 349 789 383
rect 823 349 857 383
rect 891 349 925 383
rect 959 349 993 383
rect 1027 349 1061 383
rect 1095 349 1129 383
rect 1163 349 1197 383
rect 1231 349 1265 383
rect 1299 349 1333 383
rect 1367 349 1401 383
rect 1435 349 1469 383
rect 1503 349 1537 383
rect 1571 349 1605 383
rect 1639 349 1673 383
rect 1707 349 1741 383
rect 1775 349 1809 383
rect 1843 349 1877 383
rect 1911 349 1945 383
rect 1979 349 2013 383
rect 2047 349 2081 383
rect 2115 349 2149 383
rect 2183 349 2217 383
rect 2251 349 2285 383
rect 2319 349 2353 383
rect 2387 349 2421 383
rect 2455 349 2489 383
rect 2523 349 2557 383
rect 2591 349 2625 383
rect 2659 349 2693 383
rect 2727 349 2761 383
rect 2795 349 2829 383
rect 2863 349 2897 383
rect 2931 349 2965 383
rect 2999 349 3033 383
rect 3067 349 3101 383
rect 3135 349 3169 383
rect 3203 349 3237 383
rect 3271 349 3305 383
rect 3339 349 3373 383
rect 3407 349 3441 383
rect 3475 349 3509 383
rect 3543 349 3577 383
rect 3611 349 3645 383
rect 3679 349 3713 383
rect 3747 349 3781 383
rect 3815 349 3849 383
rect 3883 349 3917 383
rect 3951 349 3985 383
rect 4019 349 4053 383
rect 4087 349 4121 383
rect 4155 349 4189 383
rect 4223 349 4257 383
rect 4291 349 4325 383
rect 4359 349 4393 383
rect 4427 349 4461 383
rect 4495 349 4529 383
rect 4563 349 4597 383
rect 4631 349 4665 383
rect 4699 349 4733 383
rect 4767 349 4801 383
rect 4835 349 4869 383
rect 4903 349 4937 383
rect 4971 349 5005 383
rect 5039 349 5073 383
rect 5107 349 5141 383
rect 5175 349 5209 383
rect 5243 349 5277 383
rect 5311 349 5345 383
rect 5379 349 5413 383
rect 5447 349 5481 383
rect 5515 349 5549 383
rect 5583 349 5617 383
rect 5651 349 5685 383
rect 5719 349 5753 383
rect 5787 349 5821 383
rect 5855 349 5889 383
rect 5923 349 5957 383
rect 5991 349 6025 383
rect 6059 349 6093 383
rect 6127 349 6161 383
rect 6195 349 6229 383
rect 6263 349 6297 383
rect 6331 349 6365 383
rect 6399 349 6433 383
rect 6467 349 6501 383
rect 6535 349 6569 383
rect 6603 349 6637 383
rect 6671 349 6705 383
rect 6739 349 6773 383
rect 6807 349 6841 383
rect 6875 349 6909 383
rect 6943 349 6977 383
rect 7011 349 7045 383
rect 7079 349 7113 383
rect 7147 349 7181 383
rect 7215 349 7249 383
rect 7283 349 7317 383
rect 7351 349 7385 383
rect 7419 349 7453 383
rect 7487 349 7521 383
rect 7555 349 7589 383
rect 7623 349 7657 383
rect 7691 349 7725 383
rect 7759 349 7793 383
rect 7827 349 7861 383
rect 7895 349 7929 383
rect 7963 349 7997 383
rect 8031 349 8098 383
rect 8064 308 8098 349
rect 8132 308 8166 342
rect 8200 308 8234 342
rect 8268 308 8302 342
rect 8336 308 8370 342
rect 8404 308 8438 342
rect 8472 308 8506 342
rect 8540 308 8574 342
rect 8608 308 8642 342
rect 8676 308 8710 342
rect 8744 308 8778 342
rect 8812 308 8846 342
rect 8880 308 8914 342
rect 8948 308 8982 342
rect 9016 308 9050 342
rect 9084 308 9118 342
rect 9152 308 9186 342
rect 9220 308 9254 342
rect 9288 308 9322 342
rect 9356 308 9390 342
rect 9424 308 9458 342
rect 9492 308 9526 342
rect 9560 308 9594 342
rect 9628 308 9662 342
rect 9696 308 9730 342
rect 9764 308 9798 342
rect 9832 308 9866 342
rect 9900 308 9934 342
rect 9968 308 10002 342
rect 10036 308 10070 342
rect 10104 308 10138 342
rect 10172 308 10206 342
rect 10240 308 10274 342
rect 10308 308 10342 342
rect 10376 308 10410 342
rect 10444 308 10478 342
rect 10512 308 10546 342
rect 10580 308 10614 342
rect 10648 308 10682 342
rect 10716 308 10750 342
rect 10784 308 10818 342
rect 10852 308 10886 342
rect 10920 308 10954 342
rect 10988 308 11022 342
rect 11056 308 11090 342
rect 11124 308 11158 342
rect 11192 308 11226 342
rect 11260 308 11294 342
rect 11328 308 11362 342
rect 11396 308 11430 342
rect 11464 308 11498 342
rect 11532 308 11566 342
rect 11600 308 11634 342
rect 11668 308 11702 342
rect 11736 308 11770 342
rect 11804 308 11838 342
rect 11872 308 11906 342
rect 11940 308 11974 342
rect 12008 308 12042 342
rect 12076 308 12110 342
rect 12144 308 12178 342
rect 12212 308 12359 342
rect 12393 308 12427 423
<< viali >>
rect 1474 6962 1508 6996
rect 1546 6962 1580 6996
rect -400 4907 -372 4939
rect -372 4907 -366 4939
rect -315 4907 -300 4939
rect -300 4907 -281 4939
rect -230 4907 -228 4939
rect -228 4907 -196 4939
rect -145 4907 -119 4939
rect -119 4907 -111 4939
rect -60 4907 -48 4939
rect -48 4907 -26 4939
rect 25 4907 57 4939
rect 57 4907 59 4939
rect -400 4905 -366 4907
rect -315 4905 -281 4907
rect -230 4905 -196 4907
rect -145 4905 -111 4907
rect -60 4905 -26 4907
rect 25 4905 59 4907
rect 13028 4864 13062 4898
rect -277 4827 -243 4861
rect -277 4781 -243 4789
rect -277 4755 -243 4781
rect -464 4679 -430 4682
rect -464 4648 -453 4679
rect -453 4648 -430 4679
rect -392 4648 -358 4682
rect 75 4827 109 4861
rect 75 4781 109 4789
rect 75 4755 109 4781
rect 13028 4792 13062 4826
rect 13028 4720 13062 4754
rect -168 4484 -134 4518
rect -96 4485 -62 4518
rect -96 4484 -67 4485
rect -67 4484 -62 4485
rect -177 4403 -143 4437
rect -177 4331 -143 4365
rect -367 4283 -366 4317
rect -366 4283 -333 4317
rect -367 4215 -366 4245
rect -366 4215 -333 4245
rect -367 4211 -333 4215
rect -638 4091 -604 4108
rect -638 4074 -615 4091
rect -615 4074 -604 4091
rect -566 4074 -532 4108
rect 10807 4472 10839 4499
rect 10839 4472 10841 4499
rect 10807 4465 10841 4472
rect 10879 4465 10913 4499
rect 10951 4465 10985 4499
rect 11023 4465 11057 4499
rect 11095 4465 11129 4499
rect 11167 4465 11201 4499
rect 11239 4465 11273 4499
rect 11311 4465 11345 4499
rect 11383 4465 11417 4499
rect 11455 4465 11489 4499
rect 11527 4465 11561 4499
rect 11599 4465 11633 4499
rect 11671 4465 11705 4499
rect 11743 4465 11777 4499
rect 11815 4465 11849 4499
rect 11887 4465 11921 4499
rect 409 4426 443 4460
rect 481 4426 511 4460
rect 511 4426 515 4460
rect 553 4426 579 4460
rect 579 4426 587 4460
rect 625 4426 647 4460
rect 647 4426 659 4460
rect 697 4426 715 4460
rect 715 4426 731 4460
rect 769 4426 783 4460
rect 783 4426 803 4460
rect 841 4426 851 4460
rect 851 4426 875 4460
rect 913 4426 919 4460
rect 919 4426 947 4460
rect 985 4426 987 4460
rect 987 4426 1019 4460
rect 1057 4426 1089 4460
rect 1089 4426 1091 4460
rect 1129 4426 1157 4460
rect 1157 4426 1163 4460
rect 1201 4426 1225 4460
rect 1225 4426 1235 4460
rect 1273 4426 1293 4460
rect 1293 4426 1307 4460
rect 1345 4426 1361 4460
rect 1361 4426 1379 4460
rect 1417 4426 1429 4460
rect 1429 4426 1451 4460
rect 1489 4426 1497 4460
rect 1497 4426 1523 4460
rect 1561 4426 1565 4460
rect 1565 4426 1595 4460
rect 1633 4426 1667 4460
rect 1705 4426 1735 4460
rect 1735 4426 1739 4460
rect 1777 4426 1803 4460
rect 1803 4426 1811 4460
rect 1849 4426 1871 4460
rect 1871 4426 1883 4460
rect 1921 4426 1939 4460
rect 1939 4426 1955 4460
rect 1993 4426 2007 4460
rect 2007 4426 2027 4460
rect 2065 4426 2075 4460
rect 2075 4426 2099 4460
rect 2137 4426 2143 4460
rect 2143 4426 2171 4460
rect 2209 4426 2211 4460
rect 2211 4426 2243 4460
rect 2281 4426 2313 4460
rect 2313 4426 2315 4460
rect 2353 4426 2381 4460
rect 2381 4426 2387 4460
rect 2425 4426 2449 4460
rect 2449 4426 2459 4460
rect 2497 4426 2517 4460
rect 2517 4426 2531 4460
rect 2569 4426 2585 4460
rect 2585 4426 2603 4460
rect 2641 4426 2653 4460
rect 2653 4426 2675 4460
rect 2713 4426 2721 4460
rect 2721 4426 2747 4460
rect 2785 4426 2789 4460
rect 2789 4426 2819 4460
rect 2857 4426 2891 4460
rect 2929 4426 2959 4460
rect 2959 4426 2963 4460
rect 3001 4426 3027 4460
rect 3027 4426 3035 4460
rect 3073 4426 3095 4460
rect 3095 4426 3107 4460
rect 3145 4426 3163 4460
rect 3163 4426 3179 4460
rect 3217 4426 3231 4460
rect 3231 4426 3251 4460
rect 3289 4426 3299 4460
rect 3299 4426 3323 4460
rect 3361 4426 3367 4460
rect 3367 4426 3395 4460
rect 3433 4426 3435 4460
rect 3435 4426 3467 4460
rect 3505 4426 3537 4460
rect 3537 4426 3539 4460
rect 3577 4426 3605 4460
rect 3605 4426 3611 4460
rect 3649 4426 3673 4460
rect 3673 4426 3683 4460
rect 3721 4426 3741 4460
rect 3741 4426 3755 4460
rect 3793 4426 3809 4460
rect 3809 4426 3827 4460
rect 3865 4426 3877 4460
rect 3877 4426 3899 4460
rect 3937 4426 3945 4460
rect 3945 4426 3971 4460
rect 4009 4426 4013 4460
rect 4013 4426 4043 4460
rect 4081 4426 4115 4460
rect 4153 4426 4183 4460
rect 4183 4426 4187 4460
rect 4225 4426 4251 4460
rect 4251 4426 4259 4460
rect 4297 4426 4319 4460
rect 4319 4426 4331 4460
rect 4369 4426 4387 4460
rect 4387 4426 4403 4460
rect 4441 4426 4455 4460
rect 4455 4426 4475 4460
rect 4513 4426 4523 4460
rect 4523 4426 4547 4460
rect 4585 4426 4591 4460
rect 4591 4426 4619 4460
rect 4657 4426 4659 4460
rect 4659 4426 4691 4460
rect 4729 4426 4761 4460
rect 4761 4426 4763 4460
rect 4801 4426 4829 4460
rect 4829 4426 4835 4460
rect 4873 4426 4897 4460
rect 4897 4426 4907 4460
rect 4945 4426 4965 4460
rect 4965 4426 4979 4460
rect 5017 4426 5033 4460
rect 5033 4426 5051 4460
rect 5089 4426 5101 4460
rect 5101 4426 5123 4460
rect 5161 4426 5169 4460
rect 5169 4426 5195 4460
rect 5233 4426 5237 4460
rect 5237 4426 5267 4460
rect 5305 4426 5339 4460
rect 5377 4426 5407 4460
rect 5407 4426 5411 4460
rect 5449 4426 5475 4460
rect 5475 4426 5483 4460
rect 5521 4426 5543 4460
rect 5543 4426 5555 4460
rect 5593 4426 5611 4460
rect 5611 4426 5627 4460
rect 5665 4426 5679 4460
rect 5679 4426 5699 4460
rect 5737 4426 5747 4460
rect 5747 4426 5771 4460
rect 5809 4426 5815 4460
rect 5815 4426 5843 4460
rect 5881 4426 5883 4460
rect 5883 4426 5915 4460
rect 5953 4426 5985 4460
rect 5985 4426 5987 4460
rect 6025 4426 6053 4460
rect 6053 4426 6059 4460
rect 6097 4426 6121 4460
rect 6121 4426 6131 4460
rect 6169 4426 6189 4460
rect 6189 4426 6203 4460
rect 6241 4426 6257 4460
rect 6257 4426 6275 4460
rect 6313 4426 6325 4460
rect 6325 4426 6347 4460
rect 6385 4426 6393 4460
rect 6393 4426 6419 4460
rect 6457 4426 6461 4460
rect 6461 4426 6491 4460
rect 6529 4426 6563 4460
rect 6601 4426 6631 4460
rect 6631 4426 6635 4460
rect 6673 4426 6699 4460
rect 6699 4426 6707 4460
rect 6745 4426 6767 4460
rect 6767 4426 6779 4460
rect 6817 4426 6835 4460
rect 6835 4426 6851 4460
rect 6889 4426 6903 4460
rect 6903 4426 6923 4460
rect 6961 4426 6971 4460
rect 6971 4426 6995 4460
rect 7033 4426 7039 4460
rect 7039 4426 7067 4460
rect 7105 4426 7107 4460
rect 7107 4426 7139 4460
rect 7177 4426 7209 4460
rect 7209 4426 7211 4460
rect 7249 4426 7277 4460
rect 7277 4426 7283 4460
rect 7321 4426 7345 4460
rect 7345 4426 7355 4460
rect 7393 4426 7413 4460
rect 7413 4426 7427 4460
rect 7465 4426 7481 4460
rect 7481 4426 7499 4460
rect 7537 4426 7549 4460
rect 7549 4426 7571 4460
rect 7609 4426 7617 4460
rect 7617 4426 7643 4460
rect 7681 4426 7685 4460
rect 7685 4426 7715 4460
rect 7753 4426 7787 4460
rect 7825 4426 7855 4460
rect 7855 4426 7859 4460
rect 7897 4426 7923 4460
rect 7923 4426 7931 4460
rect 7969 4426 7991 4460
rect 7991 4426 8003 4460
rect 8041 4426 8059 4460
rect 8059 4426 8075 4460
rect 8113 4426 8127 4460
rect 8127 4426 8147 4460
rect 8185 4426 8195 4460
rect 8195 4426 8219 4460
rect 8257 4426 8263 4460
rect 8263 4426 8291 4460
rect 8329 4426 8331 4460
rect 8331 4426 8363 4460
rect 8401 4426 8433 4460
rect 8433 4426 8435 4460
rect 8473 4426 8501 4460
rect 8501 4426 8507 4460
rect 8545 4426 8569 4460
rect 8569 4426 8579 4460
rect 8617 4426 8637 4460
rect 8637 4426 8651 4460
rect 8689 4426 8705 4460
rect 8705 4426 8723 4460
rect 8761 4426 8773 4460
rect 8773 4426 8795 4460
rect 8833 4426 8841 4460
rect 8841 4426 8867 4460
rect 8905 4426 8909 4460
rect 8909 4426 8939 4460
rect 8977 4426 9011 4460
rect 9049 4426 9079 4460
rect 9079 4426 9083 4460
rect 9121 4426 9147 4460
rect 9147 4426 9155 4460
rect 9193 4426 9215 4460
rect 9215 4426 9227 4460
rect 9265 4426 9283 4460
rect 9283 4426 9299 4460
rect 9337 4426 9351 4460
rect 9351 4426 9371 4460
rect 9409 4426 9419 4460
rect 9419 4426 9443 4460
rect 9481 4426 9487 4460
rect 9487 4426 9515 4460
rect 9553 4426 9555 4460
rect 9555 4426 9587 4460
rect 9625 4426 9657 4460
rect 9657 4426 9659 4460
rect 9697 4426 9725 4460
rect 9725 4426 9731 4460
rect 9769 4426 9793 4460
rect 9793 4426 9803 4460
rect 9841 4426 9861 4460
rect 9861 4426 9875 4460
rect 9913 4426 9929 4460
rect 9929 4426 9947 4460
rect 9985 4426 9997 4460
rect 9997 4426 10019 4460
rect 10057 4426 10065 4460
rect 10065 4426 10091 4460
rect 10129 4426 10133 4460
rect 10133 4426 10163 4460
rect 10201 4426 10235 4460
rect 10273 4426 10303 4460
rect 10303 4426 10307 4460
rect 10345 4426 10371 4460
rect 10371 4426 10379 4460
rect 10417 4426 10439 4460
rect 10439 4426 10451 4460
rect 10489 4426 10507 4460
rect 10507 4426 10523 4460
rect 10561 4426 10575 4460
rect 10575 4426 10595 4460
rect 12031 4420 12065 4454
rect 12112 4420 12146 4454
rect 12193 4420 12227 4454
rect 12274 4420 12308 4454
rect 12368 4394 12400 4415
rect 12400 4394 12402 4415
rect 12368 4381 12402 4394
rect 4501 4301 4505 4333
rect 4505 4301 4535 4333
rect 4573 4301 4607 4333
rect 4645 4301 4675 4333
rect 4675 4301 4679 4333
rect 4717 4301 4743 4333
rect 4743 4301 4751 4333
rect 4789 4301 4811 4333
rect 4811 4301 4823 4333
rect 4861 4301 4879 4333
rect 4879 4301 4895 4333
rect 4933 4301 4947 4333
rect 4947 4301 4967 4333
rect 5005 4301 5015 4333
rect 5015 4301 5039 4333
rect 5077 4301 5083 4333
rect 5083 4301 5111 4333
rect 5149 4301 5151 4333
rect 5151 4301 5183 4333
rect 5221 4301 5253 4333
rect 5253 4301 5255 4333
rect 5293 4301 5321 4333
rect 5321 4301 5327 4333
rect 5365 4301 5389 4333
rect 5389 4301 5399 4333
rect 5437 4301 5457 4333
rect 5457 4301 5471 4333
rect 5509 4301 5525 4333
rect 5525 4301 5543 4333
rect 5581 4301 5593 4333
rect 5593 4301 5615 4333
rect 12368 4326 12400 4340
rect 12400 4326 12402 4340
rect 4501 4299 4535 4301
rect 4573 4299 4607 4301
rect 4645 4299 4679 4301
rect 4717 4299 4751 4301
rect 4789 4299 4823 4301
rect 4861 4299 4895 4301
rect 4933 4299 4967 4301
rect 5005 4299 5039 4301
rect 5077 4299 5111 4301
rect 5149 4299 5183 4301
rect 5221 4299 5255 4301
rect 5293 4299 5327 4301
rect 5365 4299 5399 4301
rect 5437 4299 5471 4301
rect 5509 4299 5543 4301
rect 5581 4299 5615 4301
rect -26 4215 -15 4240
rect -15 4215 8 4240
rect -26 4206 8 4215
rect 46 4206 80 4240
rect 1536 4221 1570 4255
rect 1613 4251 1643 4255
rect 1643 4251 1647 4255
rect 1690 4251 1711 4255
rect 1711 4251 1724 4255
rect 1767 4251 1779 4255
rect 1779 4251 1801 4255
rect 1844 4251 1847 4255
rect 1847 4251 1878 4255
rect 1921 4251 1949 4255
rect 1949 4251 1955 4255
rect 1997 4251 2017 4255
rect 2017 4251 2031 4255
rect 2073 4251 2085 4255
rect 2085 4251 2107 4255
rect 1613 4221 1647 4251
rect 1690 4221 1724 4251
rect 1767 4221 1801 4251
rect 1844 4221 1878 4251
rect 1921 4221 1955 4251
rect 1997 4221 2031 4251
rect 2073 4221 2107 4251
rect 2149 4221 2183 4255
rect 2266 4251 2267 4255
rect 2267 4251 2300 4255
rect 2343 4251 2369 4255
rect 2369 4251 2377 4255
rect 2420 4251 2437 4255
rect 2437 4251 2454 4255
rect 2497 4251 2505 4255
rect 2505 4251 2531 4255
rect 2266 4221 2300 4251
rect 2343 4221 2377 4251
rect 2420 4221 2454 4251
rect 2497 4221 2531 4251
rect 3072 4251 3095 4255
rect 3095 4251 3106 4255
rect 3144 4251 3163 4255
rect 3163 4251 3178 4255
rect 3216 4251 3231 4255
rect 3231 4251 3250 4255
rect 3288 4251 3299 4255
rect 3299 4251 3322 4255
rect 3360 4251 3367 4255
rect 3367 4251 3394 4255
rect 3432 4251 3435 4255
rect 3435 4251 3466 4255
rect 3504 4251 3537 4255
rect 3537 4251 3538 4255
rect 3576 4251 3605 4255
rect 3605 4251 3610 4255
rect 3648 4251 3673 4255
rect 3673 4251 3682 4255
rect 3720 4251 3741 4255
rect 3741 4251 3754 4255
rect 3792 4251 3809 4255
rect 3809 4251 3826 4255
rect 3864 4251 3877 4255
rect 3877 4251 3898 4255
rect 3936 4251 3945 4255
rect 3945 4251 3970 4255
rect 4008 4251 4013 4255
rect 4013 4251 4042 4255
rect 4080 4251 4081 4255
rect 4081 4251 4114 4255
rect 4152 4251 4183 4255
rect 4183 4251 4186 4255
rect 3072 4221 3106 4251
rect 3144 4221 3178 4251
rect 3216 4221 3250 4251
rect 3288 4221 3322 4251
rect 3360 4221 3394 4251
rect 3432 4221 3466 4251
rect 3504 4221 3538 4251
rect 3576 4221 3610 4251
rect 3648 4221 3682 4251
rect 3720 4221 3754 4251
rect 3792 4221 3826 4251
rect 3864 4221 3898 4251
rect 3936 4221 3970 4251
rect 4008 4221 4042 4251
rect 4080 4221 4114 4251
rect 4152 4221 4186 4251
rect -277 4087 -243 4110
rect -277 4076 -243 4087
rect -638 4002 -604 4031
rect -638 3997 -615 4002
rect -615 3997 -604 4002
rect -566 3997 -532 4031
rect -277 4004 -243 4038
rect 271 4103 305 4134
rect 271 4100 305 4103
rect 271 4035 305 4054
rect 271 4020 305 4035
rect -638 3920 -604 3954
rect -566 3920 -532 3954
rect -638 3842 -604 3876
rect -566 3842 -532 3876
rect 271 3967 305 3974
rect 271 3940 305 3967
rect -314 3834 -280 3868
rect -638 3788 -615 3798
rect -615 3788 -604 3798
rect -638 3764 -604 3788
rect -566 3764 -532 3798
rect -314 3773 -280 3796
rect -314 3762 -280 3773
rect -190 3834 -156 3868
rect 271 3865 305 3893
rect 271 3859 305 3865
rect -190 3785 -156 3796
rect -190 3762 -156 3785
rect -394 3700 -360 3702
rect -394 3668 -360 3700
rect -394 3598 -360 3630
rect -394 3596 -360 3598
rect -101 3589 -67 3622
rect -101 3588 -67 3589
rect -101 3516 -67 3550
rect -470 3191 -436 3223
rect -470 3189 -436 3191
rect -470 3123 -436 3151
rect -470 3117 -436 3123
rect -314 3089 -280 3118
rect -314 3084 -280 3089
rect -314 3021 -280 3046
rect -314 3012 -280 3021
rect -190 3091 -156 3117
rect -190 3083 -156 3091
rect -190 3011 -156 3045
rect 271 3797 305 3812
rect 271 3778 305 3797
rect 129 3361 163 3395
rect 129 3289 163 3323
rect 707 3685 741 3719
rect 779 3685 813 3719
rect 1016 3620 1050 3643
rect 1016 3609 1050 3620
rect 1016 3552 1050 3571
rect 1016 3537 1050 3552
rect 1016 3484 1050 3499
rect 1016 3465 1050 3484
rect 1354 3911 1388 3945
rect 1426 3929 1460 3945
rect 1426 3911 1460 3929
rect 1270 3623 1304 3643
rect 1270 3609 1304 3623
rect 1270 3555 1304 3571
rect 1270 3537 1304 3555
rect 1270 3487 1304 3499
rect 1270 3465 1304 3487
rect 1114 3385 1148 3419
rect 1186 3385 1220 3419
rect 1655 3911 1689 3945
rect 1727 3911 1761 3945
rect 1536 3691 1570 3723
rect 1536 3689 1570 3691
rect 1608 3689 1642 3723
rect 1966 3911 2000 3945
rect 1810 3689 1844 3723
rect 2038 3911 2072 3945
rect 1882 3689 1916 3723
rect 2279 3825 2313 3859
rect 2351 3825 2385 3859
rect 1175 3121 1179 3126
rect 1179 3121 1209 3126
rect 1247 3121 1281 3126
rect 1319 3121 1349 3126
rect 1349 3121 1353 3126
rect 1391 3121 1417 3126
rect 1417 3121 1425 3126
rect 1175 3092 1209 3121
rect 1247 3092 1281 3121
rect 1319 3092 1353 3121
rect 1391 3092 1425 3121
rect 2122 3689 2156 3723
rect 2194 3689 2228 3723
rect 2590 3825 2624 3859
rect 2662 3825 2696 3859
rect 2434 3689 2468 3723
rect 2506 3689 2540 3723
rect 2712 3689 2746 3723
rect 2784 3691 2818 3723
rect 2784 3689 2818 3691
rect 3098 3689 3132 3723
rect 3170 3689 3204 3723
rect 2882 3623 2980 3643
rect 2980 3623 3014 3643
rect 3014 3623 3060 3643
rect 2882 3620 3060 3623
rect 2882 3586 2916 3620
rect 2916 3589 3060 3620
rect 2916 3586 2980 3589
rect 2882 3555 2980 3586
rect 2980 3555 3014 3589
rect 3014 3555 3060 3589
rect 2882 3552 3060 3555
rect 2882 3518 2916 3552
rect 2916 3521 3060 3552
rect 2916 3518 2980 3521
rect 2882 3487 2980 3518
rect 2980 3487 3014 3521
rect 3014 3487 3060 3521
rect 2882 3484 3060 3487
rect 2882 3465 2916 3484
rect 2916 3465 3060 3484
rect 3416 3691 3448 3723
rect 3448 3691 3450 3723
rect 3416 3689 3450 3691
rect 3488 3689 3522 3723
rect 3270 3623 3292 3643
rect 3292 3623 3326 3643
rect 3326 3623 3376 3643
rect 3270 3589 3376 3623
rect 3270 3555 3292 3589
rect 3292 3555 3326 3589
rect 3326 3555 3376 3589
rect 3270 3521 3376 3555
rect 3270 3487 3292 3521
rect 3292 3487 3326 3521
rect 3326 3487 3376 3521
rect 3270 3465 3376 3487
rect 3722 3689 3756 3723
rect 3794 3689 3828 3723
rect 3604 3623 3638 3643
rect 3604 3609 3638 3623
rect 3604 3555 3638 3571
rect 3604 3537 3638 3555
rect 3604 3487 3638 3499
rect 3604 3465 3638 3487
rect 4033 3689 4067 3723
rect 4105 3691 4106 3723
rect 4106 3691 4139 3723
rect 4105 3689 4139 3691
rect 3916 3623 3950 3643
rect 3916 3609 3950 3623
rect 3916 3555 3950 3571
rect 3916 3537 3950 3555
rect 3916 3487 3950 3499
rect 3916 3465 3950 3487
rect 4423 3707 4457 3723
rect 4423 3689 4424 3707
rect 4424 3689 4457 3707
rect 4495 3689 4529 3723
rect 4181 3623 4228 3643
rect 4228 3623 4262 3643
rect 4262 3623 4359 3643
rect 4181 3620 4359 3623
rect 4181 3589 4326 3620
rect 4181 3555 4228 3589
rect 4228 3555 4262 3589
rect 4262 3586 4326 3589
rect 4326 3586 4359 3620
rect 4262 3555 4359 3586
rect 4181 3552 4359 3555
rect 4181 3521 4326 3552
rect 4181 3487 4228 3521
rect 4228 3487 4262 3521
rect 4262 3518 4326 3521
rect 4326 3518 4359 3552
rect 4262 3487 4359 3518
rect 4181 3484 4359 3487
rect 4181 3465 4326 3484
rect 4326 3465 4359 3484
rect 4697 3689 4731 3723
rect 4769 3707 4803 3723
rect 4769 3689 4770 3707
rect 4770 3689 4803 3707
rect 4542 3385 4576 3419
rect 4614 3385 4648 3419
rect 5009 3689 5043 3723
rect 5081 3707 5115 3723
rect 5081 3689 5082 3707
rect 5082 3689 5115 3707
rect 5951 4215 5985 4249
rect 6023 4215 6057 4249
rect 6095 4215 6129 4249
rect 6167 4215 6201 4249
rect 6239 4215 6273 4249
rect 6311 4215 6345 4249
rect 6383 4215 6417 4249
rect 6455 4215 6489 4249
rect 6527 4215 6561 4249
rect 6599 4215 6633 4249
rect 6671 4215 6705 4249
rect 6743 4215 6777 4249
rect 6815 4215 6849 4249
rect 6887 4215 6921 4249
rect 6959 4215 6993 4249
rect 7031 4215 7065 4249
rect 7173 4215 7207 4249
rect 7245 4215 7279 4249
rect 7506 4217 7540 4251
rect 7578 4217 7612 4251
rect 7826 4217 7860 4251
rect 7898 4217 7932 4251
rect 4854 3385 4888 3419
rect 4926 3385 4960 3419
rect 5321 3689 5355 3723
rect 5393 3707 5427 3723
rect 5393 3689 5394 3707
rect 5394 3689 5427 3707
rect 5166 3385 5200 3419
rect 5238 3385 5272 3419
rect 5599 3689 5633 3723
rect 5671 3707 5705 3723
rect 5671 3689 5672 3707
rect 5672 3689 5705 3707
rect 5478 3385 5512 3419
rect 5550 3385 5584 3419
rect 5770 3623 5868 3643
rect 5868 3623 5902 3643
rect 5902 3623 5948 3643
rect 5770 3620 5948 3623
rect 5770 3586 5804 3620
rect 5804 3589 5948 3620
rect 5804 3586 5868 3589
rect 5770 3555 5868 3586
rect 5868 3555 5902 3589
rect 5902 3555 5948 3589
rect 5770 3552 5948 3555
rect 5770 3518 5804 3552
rect 5804 3521 5948 3552
rect 5804 3518 5868 3521
rect 5770 3487 5868 3518
rect 5868 3487 5902 3521
rect 5902 3487 5948 3521
rect 5770 3484 5948 3487
rect 5770 3465 5804 3484
rect 5804 3465 5948 3484
rect 6180 3623 6214 3643
rect 6180 3609 6214 3623
rect 6180 3555 6214 3571
rect 6180 3537 6214 3555
rect 6180 3487 6214 3499
rect 6180 3465 6214 3487
rect 6492 3623 6526 3643
rect 6492 3609 6526 3623
rect 6492 3555 6526 3571
rect 6492 3537 6526 3555
rect 6492 3487 6526 3499
rect 6492 3465 6526 3487
rect 6804 3623 6838 3643
rect 6804 3609 6838 3623
rect 6804 3555 6838 3571
rect 6804 3537 6838 3555
rect 6804 3487 6838 3499
rect 6804 3465 6838 3487
rect 9265 4219 9299 4253
rect 7116 3623 7150 3643
rect 7116 3609 7150 3623
rect 7116 3555 7150 3571
rect 7116 3537 7150 3555
rect 7116 3487 7150 3499
rect 7116 3465 7150 3487
rect 7795 3761 7829 3795
rect 7795 3689 7829 3723
rect 7340 3620 7468 3643
rect 7340 3586 7370 3620
rect 7370 3586 7404 3620
rect 7404 3615 7468 3620
rect 7468 3615 7502 3643
rect 7502 3615 7518 3643
rect 7404 3586 7518 3615
rect 7340 3552 7518 3586
rect 7340 3518 7370 3552
rect 7370 3518 7404 3552
rect 7404 3518 7518 3552
rect 7340 3484 7518 3518
rect 7340 3465 7370 3484
rect 7370 3465 7404 3484
rect 7404 3465 7518 3484
rect 7790 3609 7824 3643
rect 7790 3537 7824 3571
rect 7790 3465 7824 3499
rect 7272 3385 7306 3413
rect 7272 3379 7306 3385
rect 7272 3317 7306 3341
rect 7272 3307 7306 3317
rect 7624 3322 7658 3339
rect 7624 3305 7658 3322
rect 7696 3305 7730 3339
rect 8751 4119 9001 4164
rect 8751 4085 8785 4119
rect 8785 4085 8851 4119
rect 8851 4085 8885 4119
rect 8885 4085 8951 4119
rect 8951 4085 8985 4119
rect 8985 4085 9001 4119
rect 8751 4046 9001 4085
rect 8022 3620 8200 3643
rect 8022 3586 8166 3620
rect 8166 3586 8200 3620
rect 8022 3552 8200 3586
rect 8022 3518 8166 3552
rect 8166 3518 8200 3552
rect 8022 3484 8200 3518
rect 8022 3465 8166 3484
rect 8166 3465 8200 3484
rect 7435 3092 7469 3126
rect 7507 3092 7541 3126
rect 7762 3092 7796 3126
rect 7834 3092 7868 3126
rect 8026 3268 8060 3302
rect 8098 3268 8132 3302
rect 8751 4012 8785 4046
rect 8785 4012 8851 4046
rect 8851 4012 8885 4046
rect 8885 4012 8951 4046
rect 8951 4012 8985 4046
rect 8985 4012 9001 4046
rect 8751 3986 9001 4012
rect 9145 4136 9179 4142
rect 9145 4108 9179 4136
rect 9145 4034 9179 4046
rect 9145 4012 9179 4034
rect 8611 3877 8645 3886
rect 8611 3852 8630 3877
rect 8630 3852 8645 3877
rect 8683 3852 8717 3886
rect 9337 4219 9371 4253
rect 9570 4219 9604 4253
rect 9642 4238 9676 4253
rect 9642 4219 9647 4238
rect 9647 4219 9676 4238
rect 9457 4136 9491 4142
rect 9457 4108 9491 4136
rect 9457 4034 9491 4046
rect 9457 4012 9491 4034
rect 9708 4136 9737 4167
rect 9737 4136 9742 4167
rect 9708 4133 9742 4136
rect 9780 4133 9814 4167
rect 10011 4133 10045 4167
rect 10083 4133 10117 4167
rect 9857 4056 9891 4090
rect 9929 4056 9963 4090
rect 10324 4133 10358 4167
rect 10396 4133 10430 4167
rect 10170 3978 10204 4012
rect 10450 4056 10484 4090
rect 10607 4219 10641 4253
rect 10679 4219 10713 4253
rect 10522 4056 10556 4090
rect 10242 3978 10276 4012
rect 10125 3855 10159 3889
rect 10125 3783 10159 3817
rect 9599 3689 9633 3723
rect 9671 3689 9705 3723
rect 10285 3855 10319 3889
rect 10285 3783 10319 3817
rect 11874 4279 11908 4313
rect 11946 4279 11980 4313
rect 12368 4306 12402 4326
rect 10936 4219 10970 4253
rect 11008 4219 11042 4253
rect 12145 4186 12179 4220
rect 12145 4114 12179 4148
rect 12368 4258 12400 4265
rect 12400 4258 12402 4265
rect 12368 4231 12402 4258
rect 12368 4156 12402 4190
rect 10956 4075 10990 4109
rect 11028 4075 11062 4109
rect 10763 3978 10797 4012
rect 12368 4088 12402 4115
rect 12368 4081 12400 4088
rect 12400 4081 12402 4088
rect 10835 3978 10869 4012
rect 10607 3765 10641 3799
rect 10679 3765 10713 3799
rect 11879 3953 11907 3983
rect 11907 3953 11913 3983
rect 11879 3949 11913 3953
rect 11951 3949 11985 3983
rect 10874 3765 10908 3799
rect 10946 3765 10980 3799
rect 10516 3689 10550 3723
rect 10588 3689 10622 3723
rect 10679 3689 10713 3723
rect 10751 3689 10785 3723
rect 10483 3609 10517 3643
rect 9640 3537 9674 3571
rect 9443 3513 9477 3518
rect 9443 3484 9459 3513
rect 9459 3484 9477 3513
rect 9515 3484 9549 3518
rect 9640 3480 9674 3499
rect 9640 3465 9674 3480
rect 10136 3537 10170 3571
rect 8342 3211 8366 3245
rect 8366 3211 8376 3245
rect 8414 3211 8448 3245
rect 7920 3092 7954 3126
rect 7992 3092 8026 3126
rect -314 2953 -280 2974
rect -314 2940 -280 2953
rect -50 2837 -16 2871
rect 22 2837 40 2871
rect 40 2837 56 2871
rect 1751 2943 1767 2977
rect 1767 2943 1785 2977
rect 1823 2943 1835 2977
rect 1835 2943 1857 2977
rect 1895 2943 1903 2977
rect 1903 2943 1929 2977
rect 1967 2943 1971 2977
rect 1971 2943 2001 2977
rect 2039 2943 2073 2977
rect 2111 2943 2141 2977
rect 2141 2943 2145 2977
rect 2183 2943 2209 2977
rect 2209 2943 2217 2977
rect 2255 2943 2277 2977
rect 2277 2943 2289 2977
rect 2327 2943 2345 2977
rect 2345 2943 2361 2977
rect 2399 2943 2413 2977
rect 2413 2943 2433 2977
rect 2471 2943 2481 2977
rect 2481 2943 2505 2977
rect 2543 2943 2549 2977
rect 2549 2943 2577 2977
rect 2615 2943 2617 2977
rect 2617 2943 2649 2977
rect 2687 2943 2719 2977
rect 2719 2943 2721 2977
rect 2759 2943 2787 2977
rect 2787 2943 2793 2977
rect 2831 2943 2855 2977
rect 2855 2943 2865 2977
rect 2903 2943 2923 2977
rect 2923 2943 2937 2977
rect 2975 2943 2991 2977
rect 2991 2943 3009 2977
rect 3047 2943 3059 2977
rect 3059 2943 3081 2977
rect 3119 2943 3127 2977
rect 3127 2943 3153 2977
rect 3191 2943 3195 2977
rect 3195 2943 3225 2977
rect 3263 2943 3297 2977
rect 3358 2940 3392 2974
rect 3432 2940 3466 2974
rect 3506 2940 3540 2974
rect 3580 2940 3614 2974
rect 3654 2940 3688 2974
rect 3728 2940 3762 2974
rect 3802 2940 3836 2974
rect 3876 2940 3910 2974
rect 3950 2940 3984 2974
rect 4024 2940 4058 2974
rect 4098 2940 4132 2974
rect 4172 2940 4206 2974
rect 4246 2940 4280 2974
rect 4320 2940 4354 2974
rect 4394 2940 4428 2974
rect 4468 2940 4502 2974
rect 4541 2940 4575 2974
rect 4614 2940 4648 2974
rect 4687 2940 4721 2974
rect 4760 2940 4794 2974
rect 4833 2940 4867 2974
rect 4906 2940 4940 2974
rect 7680 2934 7714 2968
rect 7752 2934 7786 2968
rect 8070 2958 8104 2968
rect 8070 2934 8104 2958
rect 8142 2934 8176 2968
rect -453 2515 -419 2521
rect -453 2487 -419 2515
rect -453 2415 -419 2449
rect -277 2663 -243 2697
rect -277 2617 -243 2625
rect -277 2591 -243 2617
rect -101 2390 -67 2424
rect -101 2321 -67 2352
rect -101 2318 -67 2321
rect -363 2119 -332 2153
rect -332 2119 -329 2153
rect -363 2051 -332 2081
rect -332 2051 -329 2081
rect -183 2119 -152 2153
rect -152 2119 -149 2153
rect -183 2051 -152 2081
rect -152 2051 -149 2081
rect -363 2047 -329 2051
rect -183 2047 -149 2051
rect 75 2663 109 2697
rect 75 2617 109 2625
rect 75 2591 109 2617
rect 7684 2679 7718 2713
rect 7756 2688 7776 2713
rect 7776 2688 7790 2713
rect 7828 2688 7844 2713
rect 7844 2688 7862 2713
rect 7756 2679 7790 2688
rect 7828 2679 7862 2688
rect 8122 2688 8128 2722
rect 8128 2688 8156 2722
rect 8194 2688 8196 2722
rect 8196 2688 8228 2722
rect 8422 2958 8456 2974
rect 8422 2940 8456 2958
rect 8494 2940 8528 2974
rect 8639 3092 8673 3126
rect 8711 3092 8745 3126
rect 8783 3092 8817 3126
rect 8855 3092 8889 3126
rect 8927 3092 8961 3126
rect 8999 3092 9033 3126
rect 9071 3092 9105 3126
rect 9143 3092 9177 3126
rect 9215 3092 9249 3126
rect 9287 3092 9321 3126
rect 9359 3092 9393 3126
rect 10136 3465 10170 3499
rect 10483 3537 10517 3571
rect 9729 3120 9763 3126
rect 9729 3092 9756 3120
rect 9756 3092 9763 3120
rect 9801 3092 9835 3126
rect 8280 2676 8314 2710
rect 8352 2676 8386 2710
rect 8934 2958 8968 2968
rect 8934 2934 8968 2958
rect 9006 2934 9040 2968
rect 8678 2890 8712 2894
rect 8678 2860 8712 2890
rect 8750 2860 8784 2894
rect 9362 2934 9396 2968
rect 9434 2958 9468 2968
rect 9434 2934 9446 2958
rect 9446 2934 9468 2958
rect 9192 2856 9224 2890
rect 9224 2856 9226 2890
rect 9264 2856 9298 2890
rect 10483 3465 10517 3499
rect 9824 2860 9858 2894
rect 9896 2860 9930 2894
rect 9997 2860 10031 2894
rect 10069 2860 10103 2894
rect 12145 3858 12179 3892
rect 12145 3786 12179 3820
rect 11937 3607 11971 3641
rect 12011 3607 12045 3641
rect 12084 3607 12118 3641
rect 12157 3611 12183 3641
rect 12183 3611 12191 3641
rect 12157 3607 12191 3611
rect 10680 3292 10714 3326
rect 10752 3292 10786 3326
rect 10858 3379 10892 3413
rect 10930 3379 10964 3413
rect 11149 3282 11183 3316
rect 11221 3282 11255 3316
rect 11104 3209 11138 3225
rect 11180 3209 11214 3225
rect 11256 3209 11290 3225
rect 11331 3209 11365 3225
rect 11983 3385 12017 3419
rect 12055 3385 12089 3419
rect 12368 4020 12402 4040
rect 12368 4006 12400 4020
rect 12400 4006 12402 4020
rect 12368 3952 12402 3965
rect 12368 3931 12400 3952
rect 12400 3931 12402 3952
rect 12368 3884 12402 3890
rect 12368 3856 12400 3884
rect 12400 3856 12402 3884
rect 12368 3782 12400 3815
rect 12400 3782 12402 3815
rect 12368 3781 12402 3782
rect 12366 3612 12400 3643
rect 12366 3609 12400 3612
rect 12366 3544 12400 3571
rect 12366 3537 12400 3544
rect 12366 3476 12400 3499
rect 12366 3465 12400 3476
rect 12366 3374 12400 3390
rect 12366 3356 12400 3374
rect 12366 3306 12400 3318
rect 12366 3284 12400 3306
rect 12366 3238 12400 3246
rect 11808 3209 11842 3225
rect 11884 3209 11918 3225
rect 11960 3209 11994 3225
rect 12035 3209 12069 3225
rect 12366 3212 12400 3238
rect 11104 3191 11131 3209
rect 11131 3191 11138 3209
rect 11180 3191 11208 3209
rect 11208 3191 11214 3209
rect 11256 3191 11285 3209
rect 11285 3191 11290 3209
rect 11331 3191 11361 3209
rect 11361 3191 11365 3209
rect 11808 3191 11835 3209
rect 11835 3191 11842 3209
rect 11884 3191 11911 3209
rect 11911 3191 11918 3209
rect 11960 3191 11988 3209
rect 11988 3191 11994 3209
rect 12035 3191 12065 3209
rect 12065 3191 12069 3209
rect 11493 3111 11527 3145
rect 11565 3111 11599 3145
rect 12366 3170 12400 3174
rect 12366 3140 12400 3170
rect 12366 3068 12400 3102
rect 10744 3039 10778 3046
rect 10744 3012 10778 3039
rect 10860 3015 10894 3046
rect 10860 3012 10894 3015
rect 10744 2971 10778 2974
rect 10744 2940 10778 2971
rect 10860 2947 10894 2974
rect 10860 2940 10894 2947
rect 10311 2778 10345 2812
rect 10383 2778 10417 2812
rect 7524 2493 7528 2510
rect 7528 2493 7558 2510
rect 7524 2476 7558 2493
rect 7596 2476 7630 2510
rect 7997 2432 8020 2436
rect 8020 2432 8031 2436
rect 8069 2432 8088 2436
rect 8088 2432 8103 2436
rect 8141 2432 8156 2436
rect 8156 2432 8175 2436
rect 8854 2696 8888 2728
rect 8854 2694 8888 2696
rect 8926 2694 8960 2728
rect 9012 2642 9046 2652
rect 9084 2642 9118 2652
rect 9156 2642 9190 2652
rect 9228 2642 9262 2652
rect 9300 2642 9334 2652
rect 9372 2642 9406 2652
rect 9444 2642 9478 2652
rect 9012 2618 9036 2642
rect 9036 2618 9046 2642
rect 9084 2618 9104 2642
rect 9104 2618 9118 2642
rect 9156 2618 9172 2642
rect 9172 2618 9190 2642
rect 9228 2618 9240 2642
rect 9240 2618 9262 2642
rect 9300 2618 9308 2642
rect 9308 2618 9334 2642
rect 9372 2618 9376 2642
rect 9376 2618 9406 2642
rect 9444 2618 9478 2642
rect 7997 2402 8031 2432
rect 8069 2402 8103 2432
rect 8141 2402 8175 2432
rect 8614 2424 8720 2430
rect 8614 2390 8678 2424
rect 8678 2390 8712 2424
rect 8712 2390 8720 2424
rect -10 2119 19 2153
rect 19 2119 24 2153
rect -10 2051 19 2081
rect 19 2051 24 2081
rect -10 2047 24 2051
rect -277 1923 -243 1946
rect -277 1912 -243 1923
rect -277 1840 -243 1874
rect -423 1745 -409 1779
rect -409 1745 -389 1779
rect -344 1745 -331 1779
rect -331 1745 -310 1779
rect -265 1745 -253 1779
rect -253 1745 -231 1779
rect -187 1745 -175 1779
rect -175 1745 -153 1779
rect -109 1745 -97 1779
rect -97 1745 -75 1779
rect -31 1745 -20 1779
rect -20 1745 3 1779
rect 47 1745 57 1779
rect 57 1745 81 1779
rect 8614 2356 8720 2390
rect 8614 2324 8678 2356
rect 8678 2324 8712 2356
rect 8712 2324 8720 2356
rect 9012 2486 9046 2510
rect 9084 2486 9118 2510
rect 9156 2486 9190 2510
rect 9228 2486 9262 2510
rect 9300 2486 9334 2510
rect 9372 2486 9406 2510
rect 9444 2486 9478 2510
rect 9756 2530 9790 2560
rect 9756 2526 9790 2530
rect 9012 2476 9036 2486
rect 9036 2476 9046 2486
rect 9084 2476 9104 2486
rect 9104 2476 9118 2486
rect 9156 2476 9172 2486
rect 9172 2476 9190 2486
rect 9228 2476 9240 2486
rect 9240 2476 9262 2486
rect 9300 2476 9308 2486
rect 9308 2476 9334 2486
rect 9372 2476 9376 2486
rect 9376 2476 9406 2486
rect 9444 2476 9478 2486
rect 9756 2454 9790 2488
rect 10136 2530 10170 2560
rect 10136 2526 10170 2530
rect 10136 2454 10170 2488
rect 11212 3015 11246 3046
rect 11212 3012 11246 3015
rect 11212 2947 11246 2974
rect 11212 2940 11246 2947
rect 11564 3015 11598 3046
rect 11564 3012 11598 3015
rect 11564 2947 11598 2974
rect 11564 2940 11598 2947
rect 11916 3015 11950 3046
rect 11916 3012 11950 3015
rect 11916 2947 11950 2974
rect 11916 2940 11950 2947
rect 12366 3000 12400 3030
rect 12366 2996 12400 3000
rect 12366 2932 12400 2958
rect 12366 2924 12400 2932
rect 12366 2864 12400 2886
rect 12366 2852 12400 2864
rect 12366 2796 12400 2814
rect 12366 2780 12400 2796
rect 12366 2728 12400 2742
rect 12366 2708 12400 2728
rect 11011 2476 11045 2510
rect 11083 2476 11117 2510
rect 11355 2476 11389 2510
rect 11427 2476 11461 2510
rect 11709 2476 11743 2510
rect 11781 2476 11815 2510
rect 12053 2476 12087 2510
rect 12125 2476 12159 2510
rect 12366 2388 12400 2413
rect 12366 2379 12400 2388
rect 7930 1989 7964 2019
rect 7930 1985 7964 1989
rect 7930 1921 7964 1947
rect 7930 1913 7964 1921
rect 7930 1853 7964 1875
rect 7930 1841 7964 1853
rect 8678 2016 8712 2018
rect 8678 1984 8712 2016
rect 8678 1914 8712 1946
rect 8678 1912 8712 1914
rect 8678 1846 8712 1874
rect 8678 1840 8712 1846
rect 8977 1990 9011 2012
rect 8977 1978 9011 1990
rect 8977 1922 9011 1940
rect 8977 1906 9011 1922
rect 8977 1854 9011 1868
rect 8977 1834 9011 1854
rect 8547 1686 8581 1720
rect 8619 1686 8653 1720
rect 8746 1686 8780 1720
rect 8818 1686 8852 1720
rect 7840 1640 7874 1646
rect 7912 1640 7946 1646
rect 7840 1612 7842 1640
rect 7842 1612 7874 1640
rect 7912 1612 7944 1640
rect 7944 1612 7946 1640
rect 8184 1612 8218 1646
rect 8256 1612 8290 1646
rect 8947 1688 8981 1722
rect 9019 1688 9053 1722
rect 9329 1990 9363 2012
rect 9329 1978 9363 1990
rect 9329 1922 9363 1940
rect 9329 1906 9363 1922
rect 9329 1854 9363 1868
rect 9329 1834 9363 1854
rect 9441 1988 9547 2013
rect 9441 1954 9445 1988
rect 9445 1954 9479 1988
rect 9479 1954 9513 1988
rect 9513 1954 9547 1988
rect 9441 1914 9547 1954
rect 9441 1880 9445 1914
rect 9445 1880 9479 1914
rect 9479 1880 9513 1914
rect 9513 1880 9547 1914
rect 9441 1840 9547 1880
rect 9441 1835 9445 1840
rect 9445 1835 9479 1840
rect 9479 1835 9513 1840
rect 9513 1835 9547 1840
rect 7426 1538 7460 1572
rect 7498 1538 7532 1572
rect 7422 1474 7456 1486
rect 7422 1452 7456 1474
rect 7422 1406 7456 1414
rect 7422 1380 7456 1406
rect 7422 1338 7456 1342
rect 7422 1308 7456 1338
rect 621 664 633 770
rect 633 664 1075 770
rect 1075 664 1087 770
rect 9698 2081 9732 2115
rect 9770 2081 9804 2115
rect 9982 2081 10016 2115
rect 10054 2081 10088 2115
rect 10262 2081 10296 2115
rect 10334 2081 10368 2115
rect 10192 1990 10226 2012
rect 10192 1978 10226 1990
rect 10192 1922 10226 1940
rect 10192 1906 10226 1922
rect 10192 1854 10226 1868
rect 10192 1834 10226 1854
rect 10486 1983 10520 2012
rect 10486 1978 10520 1983
rect 10486 1915 10520 1940
rect 10486 1906 10520 1915
rect 10486 1847 10520 1868
rect 10486 1834 10520 1847
rect 10804 2088 10838 2098
rect 10804 2064 10818 2088
rect 10818 2064 10838 2088
rect 10876 2064 10910 2098
rect 11102 2064 11136 2098
rect 10960 1986 10994 2018
rect 10960 1984 10994 1986
rect 10960 1918 10994 1946
rect 10960 1912 10994 1918
rect 10960 1850 10994 1874
rect 10960 1840 10994 1850
rect 11174 2064 11208 2098
rect 11312 1986 11346 2018
rect 11312 1984 11346 1986
rect 11312 1918 11346 1946
rect 11312 1912 11346 1918
rect 11312 1850 11346 1874
rect 11312 1840 11346 1850
rect 11459 2088 11493 2098
rect 11459 2064 11488 2088
rect 11488 2064 11493 2088
rect 11537 2064 11571 2098
rect 11664 1986 11698 2018
rect 11664 1984 11698 1986
rect 11664 1918 11698 1946
rect 11664 1912 11698 1918
rect 11664 1850 11698 1874
rect 11664 1840 11698 1850
rect 11806 2064 11840 2098
rect 11878 2064 11912 2098
rect 12016 1986 12050 2018
rect 12016 1984 12050 1986
rect 12102 2014 12136 2018
rect 12102 1984 12133 2014
rect 12133 1984 12136 2014
rect 12016 1918 12050 1946
rect 12016 1912 12050 1918
rect 12102 1940 12136 1946
rect 12102 1912 12133 1940
rect 12133 1912 12136 1940
rect 12016 1850 12050 1874
rect 12016 1840 12050 1850
rect 12102 1866 12136 1874
rect 12102 1840 12133 1866
rect 12133 1840 12136 1866
rect 12366 2320 12400 2337
rect 12366 2303 12400 2320
rect 12366 2252 12400 2261
rect 12366 2227 12400 2252
rect 12366 2184 12400 2185
rect 12366 2151 12400 2184
rect 12366 2082 12400 2109
rect 12366 2075 12400 2082
rect 12366 2014 12400 2033
rect 12366 1999 12400 2014
rect 12366 1946 12400 1957
rect 12366 1923 12400 1946
rect 12366 1878 12400 1881
rect 12366 1847 12400 1878
rect 9432 1625 9436 1646
rect 9436 1625 9466 1646
rect 9504 1625 9538 1646
rect 9432 1612 9466 1625
rect 9504 1612 9538 1625
rect 9742 1538 9776 1572
rect 9814 1538 9848 1572
rect 9886 1538 9920 1572
rect 9958 1538 9992 1572
rect 7564 1154 7598 1188
rect 7774 1474 7808 1486
rect 7774 1452 7808 1474
rect 7774 1406 7808 1414
rect 7774 1380 7808 1406
rect 7774 1338 7808 1342
rect 7774 1308 7808 1338
rect 7636 1154 7670 1188
rect 7878 1154 7912 1188
rect 7950 1168 7984 1188
rect 7950 1154 7984 1168
rect 9040 1466 9074 1498
rect 9040 1464 9074 1466
rect 9040 1398 9074 1426
rect 9040 1392 9074 1398
rect 9040 1330 9074 1354
rect 9040 1320 9074 1330
rect 8884 1262 8918 1268
rect 8884 1234 8918 1262
rect 8956 1234 8990 1268
rect 9160 1234 9194 1268
rect 9232 1234 9266 1268
rect 9658 1480 9692 1486
rect 9658 1452 9692 1480
rect 9658 1412 9692 1414
rect 9658 1380 9692 1412
rect 9658 1310 9692 1342
rect 9658 1308 9692 1310
rect 9508 1262 9542 1268
rect 9508 1234 9542 1262
rect 9580 1234 9614 1268
rect 9318 1036 9352 1070
rect 9390 1036 9424 1070
rect 9912 1466 9946 1486
rect 9912 1452 9946 1466
rect 9912 1398 9946 1414
rect 9912 1380 9946 1398
rect 9912 1330 9946 1342
rect 9912 1308 9946 1330
rect 9756 1092 9790 1112
rect 9756 1078 9790 1092
rect 9828 1078 9862 1112
rect 10285 1628 10289 1658
rect 10289 1628 10319 1658
rect 10357 1628 10391 1658
rect 10285 1624 10319 1628
rect 10357 1624 10391 1628
rect 10429 1624 10463 1658
rect 10639 1538 10673 1572
rect 10712 1538 10746 1572
rect 10785 1538 10819 1572
rect 10917 1542 10951 1576
rect 10989 1546 11023 1576
rect 10989 1542 10993 1546
rect 10993 1542 11023 1546
rect 11105 1616 11139 1650
rect 11105 1546 11139 1578
rect 11105 1544 11118 1546
rect 11118 1544 11139 1546
rect 10224 1466 10258 1486
rect 10224 1452 10258 1466
rect 10224 1398 10258 1414
rect 10224 1380 10258 1398
rect 10224 1330 10258 1342
rect 10224 1308 10258 1330
rect 10022 1078 10056 1112
rect 10094 1092 10102 1112
rect 10102 1092 10128 1112
rect 10094 1078 10128 1092
rect 10296 1078 10330 1112
rect 10368 1092 10380 1112
rect 10380 1092 10402 1112
rect 10368 1078 10402 1092
rect 10455 1458 10489 1492
rect 10455 1379 10489 1413
rect 10455 1300 10489 1334
rect 10455 1221 10489 1255
rect 10561 1239 10595 1268
rect 10561 1234 10572 1239
rect 10572 1234 10595 1239
rect 10633 1234 10667 1268
rect 10455 1142 10489 1176
rect 9025 862 9047 896
rect 9047 862 9059 896
rect 9097 862 9115 896
rect 9115 862 9131 896
rect 9352 862 9374 896
rect 9374 862 9386 896
rect 9424 862 9442 896
rect 9442 862 9458 896
rect 9578 817 9612 851
rect 9651 817 9685 851
rect 9724 817 9758 851
rect 9797 817 9831 851
rect 9870 817 9904 851
rect 9943 817 9977 851
rect 10016 817 10050 851
rect 10088 817 10122 851
rect 10160 817 10194 851
rect 11040 1409 11074 1422
rect 11040 1388 11074 1409
rect 11040 1341 11074 1350
rect 11040 1316 11074 1341
rect 12366 1470 12400 1492
rect 12366 1458 12400 1470
rect 11156 1234 11190 1268
rect 11228 1239 11262 1268
rect 11228 1234 11230 1239
rect 11230 1234 11262 1239
rect 12225 1387 12259 1421
rect 12225 1337 12259 1349
rect 12225 1315 12259 1337
rect 12366 1402 12400 1420
rect 12366 1386 12400 1402
rect 12366 1334 12400 1348
rect 12366 1314 12400 1334
rect 11791 1219 11825 1253
rect 11872 1219 11906 1253
rect 11953 1219 11987 1253
rect 12034 1219 12068 1253
rect 11791 1137 11825 1171
rect 11872 1137 11906 1171
rect 11953 1137 11987 1171
rect 12034 1137 12068 1171
rect 12366 1062 12400 1081
rect 12366 1047 12400 1062
rect 10932 975 10943 1009
rect 10943 975 10966 1009
rect 11011 975 11012 1009
rect 11012 975 11045 1009
rect 11090 975 11115 1009
rect 11115 975 11124 1009
rect 11169 975 11184 1009
rect 11184 975 11203 1009
rect 11248 975 11253 1009
rect 11253 975 11282 1009
rect 11326 975 11358 1009
rect 11358 975 11360 1009
rect 11404 975 11428 1009
rect 11428 975 11438 1009
rect 11482 975 11498 1009
rect 11498 975 11516 1009
rect 11560 975 11568 1009
rect 11568 975 11594 1009
rect 11638 975 11672 1009
rect 11716 975 11742 1009
rect 11742 975 11750 1009
rect 12366 994 12400 1008
rect 10691 801 10725 835
rect 10763 801 10797 835
rect 11309 801 11343 835
rect 11381 801 11415 835
rect 10472 725 10506 730
rect 10472 696 10501 725
rect 10501 696 10506 725
rect 10561 725 10595 730
rect 10651 725 10685 730
rect 10561 696 10562 725
rect 10562 696 10595 725
rect 10651 696 10657 725
rect 10657 696 10685 725
rect 10866 692 10900 726
rect 10938 725 10972 726
rect 11111 725 11145 730
rect 11220 725 11254 730
rect 12366 974 12400 994
rect 12183 799 12217 833
rect 12255 799 12289 833
rect 12366 926 12400 935
rect 12366 901 12400 926
rect 12366 858 12400 862
rect 12366 828 12400 858
rect 12366 754 12400 788
rect 12700 1087 12734 1121
rect 12700 1010 12734 1044
rect 12700 933 12734 967
rect 12700 855 12734 889
rect 12700 777 12734 811
rect 10938 692 10969 725
rect 10969 692 10972 725
rect 11111 696 11124 725
rect 11124 696 11145 725
rect 11220 696 11226 725
rect 11226 696 11254 725
rect 12366 695 12393 714
rect 12393 695 12400 714
rect 12700 699 12734 733
rect 12366 680 12400 695
rect 10206 576 10240 610
rect 10278 584 10286 610
rect 10286 584 10312 610
rect 10278 576 10312 584
rect 10526 576 10560 610
rect 10598 576 10632 610
rect 10370 486 10404 520
rect 10442 486 10476 520
rect 11026 576 11060 610
rect 11098 576 11132 610
rect 11308 576 11342 610
rect 11380 576 11414 610
rect 11620 576 11654 610
rect 11692 576 11726 610
rect 10682 486 10716 520
rect 10754 486 10788 520
rect 10875 486 10909 520
rect 10947 486 10981 520
rect 11183 486 11217 520
rect 11255 486 11289 520
rect 11463 486 11497 520
rect 11535 486 11569 520
<< metal1 >>
rect 1462 6953 1468 7005
rect 1520 6953 1534 7005
rect 1586 6953 1592 7005
rect 5095 6957 5128 6995
rect 5854 6502 5967 6850
rect 7271 6574 7277 6626
rect 7329 6574 7341 6626
rect 7393 6574 9428 6626
rect 9480 6574 9492 6626
rect 9544 6574 9550 6626
rect 14736 6434 14788 6440
rect 14854 6410 14989 6527
rect 14736 6370 14788 6382
rect 14736 6298 14788 6318
tri 14736 6297 14737 6298 ne
rect 14737 6297 14788 6298
tri 14788 6297 14803 6312 sw
tri 14737 6247 14787 6297 ne
rect 14787 6247 14803 6297
tri 14787 6231 14803 6247 ne
tri 14803 6231 14869 6297 sw
tri 14803 6211 14823 6231 ne
rect 14823 6141 14869 6231
rect 14824 6126 14868 6141
rect 288 5857 328 6059
tri 12592 5921 12598 5927 se
rect 12598 5875 12604 5927
rect 12656 5875 12668 5927
rect 12720 5875 12726 5927
tri 12726 5921 12732 5927 sw
rect 13102 5787 13142 5989
rect 13170 5809 13337 5965
tri 6699 5642 6713 5656 ne
rect 6713 5642 6735 5656
rect -370 5625 -318 5642
tri 6713 5631 6724 5642 ne
rect 6724 5631 6735 5642
tri 6724 5620 6735 5631 ne
tri 6831 5622 6865 5656 nw
rect 11679 5626 11685 5678
rect 11737 5626 11749 5678
rect 11801 5626 12949 5678
rect 13001 5626 13013 5678
rect 13065 5626 13071 5678
rect 13425 5630 13492 5674
rect -370 5561 -318 5573
rect 6870 5546 6876 5598
rect 6928 5546 6940 5598
rect 6992 5546 12200 5598
rect 12252 5546 12264 5598
rect 12316 5546 12322 5598
rect -370 5503 -318 5509
rect -18 5498 34 5504
rect -194 5492 -142 5498
rect -194 5406 -142 5440
tri 7432 5466 7449 5483 se
rect 7449 5480 8435 5483
tri 8435 5480 8438 5483 sw
rect 7449 5466 8438 5480
tri 8438 5466 8452 5480 sw
rect -18 5426 34 5446
tri 7395 5429 7432 5466 se
rect 7432 5445 8452 5466
rect 7432 5429 7449 5445
tri 7449 5429 7465 5445 nw
tri 8419 5429 8435 5445 ne
rect 8435 5429 8452 5445
tri 7378 5412 7395 5429 se
rect 7395 5412 7432 5429
tri 7432 5412 7449 5429 nw
tri 8435 5412 8452 5429 ne
tri 8452 5428 8490 5466 sw
rect 9422 5428 9428 5480
rect 9480 5428 9492 5480
rect 9544 5428 11573 5480
rect 11625 5428 11637 5480
rect 11689 5428 11695 5480
rect 12073 5443 12079 5495
rect 12131 5443 12143 5495
rect 12195 5443 12990 5495
tri 12910 5428 12925 5443 ne
rect 12925 5428 12990 5443
rect 8452 5412 8490 5428
tri 8490 5412 8506 5428 sw
tri 12925 5412 12941 5428 ne
rect 12941 5412 12990 5428
tri 7341 5375 7378 5412 se
rect 7378 5375 7395 5412
tri 7395 5375 7432 5412 nw
tri 8452 5375 8489 5412 ne
rect 8489 5409 8506 5412
tri 8506 5409 8509 5412 sw
tri 12941 5409 12944 5412 ne
rect 8489 5398 8509 5409
tri 8509 5398 8520 5409 sw
rect 8489 5375 8520 5398
rect -18 5368 34 5374
tri 7334 5368 7341 5375 se
rect 7341 5368 7378 5375
tri 7324 5358 7334 5368 se
rect 7334 5358 7378 5368
tri 7378 5358 7395 5375 nw
tri 8489 5358 8506 5375 ne
rect 8506 5368 8520 5375
tri 8520 5368 8550 5398 sw
rect 8506 5358 8550 5368
tri 8550 5358 8560 5368 sw
rect -194 5348 -142 5354
tri 7314 5348 7324 5358 se
rect 7324 5348 7341 5358
tri 7298 5332 7314 5348 se
rect 7314 5332 7341 5348
rect 715 5280 721 5332
rect 773 5280 785 5332
rect 837 5326 847 5332
tri 847 5326 853 5332 sw
tri 7292 5326 7298 5332 se
rect 7298 5326 7341 5332
rect 837 5280 6876 5326
rect 715 5274 6876 5280
rect 6928 5274 6940 5326
rect 6992 5274 6998 5326
tri 7287 5321 7292 5326 se
rect 7292 5321 7341 5326
tri 7341 5321 7378 5358 nw
tri 8506 5321 8543 5358 ne
rect 8543 5348 8560 5358
tri 8560 5348 8570 5358 sw
rect 8543 5346 8570 5348
tri 8570 5346 8572 5348 sw
rect 12194 5346 12200 5398
rect 12252 5346 12264 5398
rect 12316 5346 12863 5398
rect 8543 5332 8572 5346
tri 8572 5332 8586 5346 sw
tri 12777 5332 12791 5346 ne
rect 12791 5332 12863 5346
rect 8543 5326 8586 5332
tri 8586 5326 8592 5332 sw
tri 12791 5326 12797 5332 ne
rect 12797 5326 12863 5332
rect 8543 5321 8592 5326
tri 7270 5304 7287 5321 se
rect 7287 5304 7324 5321
tri 7324 5304 7341 5321 nw
tri 8543 5304 8560 5321 ne
rect 8560 5318 8592 5321
tri 8592 5318 8600 5326 sw
tri 12797 5318 12805 5326 ne
rect 12805 5318 12863 5326
rect 8560 5312 8600 5318
tri 8600 5312 8606 5318 sw
tri 9429 5312 9435 5318 se
rect 9435 5312 9441 5318
rect 8560 5304 8606 5312
tri 8606 5304 8614 5312 sw
tri 9421 5304 9429 5312 se
rect 9429 5304 9441 5312
tri 7240 5274 7270 5304 se
rect 7270 5274 7287 5304
tri 7233 5267 7240 5274 se
rect 7240 5267 7287 5274
tri 7287 5267 7324 5304 nw
tri 8560 5267 8597 5304 ne
rect 8597 5267 9441 5304
tri 7211 5245 7233 5267 se
rect 7233 5245 7265 5267
tri 7265 5245 7287 5267 nw
tri 8597 5266 8598 5267 ne
rect 8598 5266 9441 5267
rect 9493 5266 9505 5318
rect 9557 5266 9563 5318
tri 12805 5312 12811 5318 ne
rect 12811 5305 12863 5318
rect 12944 5351 12990 5412
tri 12990 5351 13024 5385 sw
tri 12863 5305 12869 5311 sw
rect 12944 5305 13136 5351
tri 13705 5305 13711 5311 se
rect 12811 5277 12869 5305
tri 12869 5277 12897 5305 sw
tri 13677 5277 13705 5305 se
rect 13705 5277 13711 5305
rect 14478 5304 14522 5348
rect 15042 5345 15116 5380
rect 5228 5239 7244 5245
rect 5280 5224 7244 5239
tri 7244 5224 7265 5245 nw
rect 5280 5207 7227 5224
tri 7227 5207 7244 5224 nw
rect 7411 5218 7463 5224
rect 12811 5219 13711 5277
rect 5228 5175 5280 5187
tri 5280 5134 5353 5207 nw
rect 7411 5154 7463 5166
rect 5228 5117 5280 5123
tri 7463 5148 7497 5182 sw
rect 7463 5102 8333 5148
rect 7411 5096 8333 5102
rect -508 4939 328 4945
rect -508 4905 -400 4939
rect -366 4905 -315 4939
rect -281 4905 -230 4939
rect -196 4905 -145 4939
rect -111 4905 -60 4939
rect -26 4905 25 4939
rect 59 4905 328 4939
rect 524 4938 564 5068
rect 12900 4938 12940 5068
rect 13335 4987 13341 4991
rect 13251 4939 13341 4987
rect 13393 4939 13413 4991
rect 13465 4939 13484 4991
rect 13536 4939 13555 4991
rect 13607 4939 13626 4991
rect 13678 4939 13684 4991
rect 13251 4916 13684 4939
rect -508 4861 328 4905
rect -508 4827 -277 4861
rect -243 4827 75 4861
rect 109 4827 328 4861
rect -508 4789 328 4827
rect -508 4755 -277 4789
rect -243 4755 75 4789
rect 109 4755 328 4789
rect -508 4743 328 4755
rect -508 4742 152 4743
rect 288 4708 328 4743
rect 823 4858 829 4910
rect 881 4858 894 4910
rect 946 4858 959 4910
rect 1011 4858 1024 4910
rect 1076 4858 1089 4910
rect 1141 4858 1153 4910
rect 1205 4858 1217 4910
rect 1269 4858 1281 4910
rect 1333 4858 1345 4910
rect 1397 4858 1409 4910
rect 1461 4858 1473 4910
rect 1525 4858 1531 4910
rect 823 4835 1531 4858
rect 823 4783 829 4835
rect 881 4783 894 4835
rect 946 4783 959 4835
rect 1011 4783 1024 4835
rect 1076 4783 1089 4835
rect 1141 4783 1153 4835
rect 1205 4783 1217 4835
rect 1269 4783 1281 4835
rect 1333 4783 1345 4835
rect 1397 4783 1409 4835
rect 1461 4783 1473 4835
rect 1525 4783 1531 4835
rect 823 4760 1531 4783
rect 823 4708 829 4760
rect 881 4708 894 4760
rect 946 4708 959 4760
rect 1011 4708 1024 4760
rect 1076 4708 1089 4760
rect 1141 4708 1153 4760
rect 1205 4708 1217 4760
rect 1269 4708 1281 4760
rect 1333 4708 1345 4760
rect 1397 4708 1409 4760
rect 1461 4708 1473 4760
rect 1525 4708 1531 4760
rect 12347 4904 12399 4910
rect 12347 4835 12399 4852
rect 12347 4766 12399 4783
rect 12347 4708 12399 4714
rect 12991 4898 13068 4910
rect 12991 4864 13028 4898
rect 13062 4864 13068 4898
rect 12991 4826 13068 4864
rect 12991 4792 13028 4826
rect 13062 4792 13068 4826
rect 13251 4864 13341 4916
rect 13393 4864 13413 4916
rect 13465 4864 13484 4916
rect 13536 4864 13555 4916
rect 13607 4864 13626 4916
rect 13678 4864 13684 4916
rect 13251 4841 13684 4864
rect 13251 4812 13341 4841
rect 12991 4754 13068 4792
rect 13335 4789 13341 4812
rect 13393 4789 13413 4841
rect 13465 4789 13484 4841
rect 13536 4789 13555 4841
rect 13607 4789 13626 4841
rect 13678 4789 13684 4841
rect 12991 4720 13028 4754
rect 13062 4720 13068 4754
rect 12991 4708 13068 4720
rect -476 4682 -282 4688
rect -476 4648 -464 4682
rect -430 4648 -392 4682
rect -358 4648 -282 4682
rect -476 4642 -282 4648
tri -352 4636 -346 4642 ne
rect -346 4636 -282 4642
rect -230 4636 -218 4688
rect -166 4636 -160 4688
rect 9930 4626 9936 4678
rect 9988 4626 10000 4678
rect 10052 4626 10190 4678
rect 10242 4626 10254 4678
rect 10306 4626 10312 4678
rect -463 4606 -406 4612
tri -406 4606 -400 4612 sw
rect -411 4596 219 4606
tri 219 4596 229 4606 sw
rect -411 4586 229 4596
tri 229 4586 239 4596 sw
rect -411 4554 3628 4586
rect -463 4544 -370 4554
tri -370 4544 -360 4554 nw
tri 197 4544 207 4554 ne
rect 207 4544 3628 4554
rect -463 4542 -380 4544
rect -411 4534 -380 4542
tri -380 4534 -370 4544 nw
tri 207 4534 217 4544 ne
rect 217 4534 3628 4544
rect 3680 4534 3692 4586
rect 3744 4534 3750 4586
rect 11615 4544 11621 4596
rect 11673 4544 11685 4596
rect 11737 4585 12071 4596
tri 12071 4585 12082 4596 sw
rect 12153 4585 12159 4637
rect 12211 4585 12224 4637
rect 12276 4585 14690 4637
rect 14742 4585 14754 4637
rect 14806 4585 14812 4637
rect 11737 4557 12082 4585
tri 12082 4557 12110 4585 sw
rect 11737 4544 14591 4557
tri 12049 4534 12059 4544 ne
rect 12059 4534 14591 4544
rect -411 4518 -396 4534
tri -396 4518 -380 4534 nw
tri 12059 4524 12069 4534 ne
rect 12069 4524 14591 4534
tri -251 4518 -245 4524 se
rect -245 4518 -50 4524
rect -411 4505 -409 4518
tri -409 4505 -396 4518 nw
tri -264 4505 -251 4518 se
rect -251 4505 -168 4518
tri -411 4503 -409 4505 nw
tri -266 4503 -264 4505 se
rect -264 4503 -168 4505
rect -463 4484 -411 4490
tri -285 4484 -266 4503 se
rect -266 4484 -168 4503
rect -134 4484 -96 4518
rect -62 4484 -50 4518
tri 12069 4505 12088 4524 ne
rect 12088 4505 14591 4524
rect 14643 4505 14655 4557
rect 14707 4505 14713 4557
tri -291 4478 -285 4484 se
rect -285 4478 -50 4484
tri -304 4465 -291 4478 se
rect -291 4465 -238 4478
tri -238 4465 -225 4478 nw
tri -307 4462 -304 4465 se
rect -304 4462 -241 4465
tri -241 4462 -238 4465 nw
tri -309 4460 -307 4462 se
rect -307 4460 -243 4462
tri -243 4460 -241 4462 nw
rect 369 4460 829 4505
tri -332 4437 -309 4460 se
rect -309 4458 -245 4460
tri -245 4458 -243 4460 nw
rect -309 4437 -266 4458
tri -266 4437 -245 4458 nw
rect -183 4443 -51 4449
rect -183 4437 -103 4443
tri -366 4403 -332 4437 se
rect -332 4403 -300 4437
tri -300 4403 -266 4437 nw
rect -183 4403 -177 4437
rect -143 4403 -103 4437
tri -373 4396 -366 4403 se
rect -366 4396 -307 4403
tri -307 4396 -300 4403 nw
rect -373 4381 -322 4396
tri -322 4381 -307 4396 nw
rect -183 4391 -103 4403
rect -373 4317 -327 4381
tri -327 4376 -322 4381 nw
rect -183 4377 -51 4391
rect 369 4426 409 4460
rect 443 4426 481 4460
rect 515 4426 553 4460
rect 587 4426 625 4460
rect 659 4426 697 4460
rect 731 4426 769 4460
rect 803 4453 829 4460
rect 881 4453 894 4505
rect 946 4460 959 4505
rect 1011 4460 1024 4505
rect 1076 4460 1089 4505
rect 1141 4460 1153 4505
rect 1205 4460 1217 4505
rect 1269 4460 1281 4505
rect 947 4453 959 4460
rect 1019 4453 1024 4460
rect 1269 4453 1273 4460
rect 1333 4453 1345 4505
rect 1397 4453 1409 4505
rect 1461 4453 1473 4505
rect 1525 4499 11999 4505
rect 1525 4465 10807 4499
rect 10841 4465 10879 4499
rect 10913 4465 10951 4499
rect 10985 4465 11023 4499
rect 11057 4465 11095 4499
rect 11129 4465 11167 4499
rect 11201 4465 11239 4499
rect 11273 4465 11311 4499
rect 11345 4465 11383 4499
rect 11417 4465 11455 4499
rect 11489 4465 11527 4499
rect 11561 4465 11599 4499
rect 11633 4465 11671 4499
rect 11705 4465 11743 4499
rect 11777 4465 11815 4499
rect 11849 4465 11887 4499
rect 11921 4473 11999 4499
tri 11999 4473 12031 4505 sw
rect 11921 4465 12408 4473
rect 1525 4460 12408 4465
rect 1525 4453 1561 4460
rect 803 4433 841 4453
rect 875 4433 913 4453
rect 947 4433 985 4453
rect 1019 4433 1057 4453
rect 1091 4433 1129 4453
rect 1163 4433 1201 4453
rect 1235 4433 1273 4453
rect 1307 4433 1345 4453
rect 1379 4433 1417 4453
rect 1451 4433 1489 4453
rect 1523 4433 1561 4453
rect 803 4426 829 4433
rect 369 4381 829 4426
rect 881 4381 894 4433
rect 947 4426 959 4433
rect 1019 4426 1024 4433
rect 1269 4426 1273 4433
rect 946 4381 959 4426
rect 1011 4381 1024 4426
rect 1076 4381 1089 4426
rect 1141 4381 1153 4426
rect 1205 4381 1217 4426
rect 1269 4381 1281 4426
rect 1333 4381 1345 4433
rect 1397 4381 1409 4433
rect 1461 4381 1473 4433
rect 1525 4426 1561 4433
rect 1595 4426 1633 4460
rect 1667 4426 1705 4460
rect 1739 4426 1777 4460
rect 1811 4426 1849 4460
rect 1883 4426 1921 4460
rect 1955 4426 1993 4460
rect 2027 4426 2065 4460
rect 2099 4426 2137 4460
rect 2171 4426 2209 4460
rect 2243 4426 2281 4460
rect 2315 4426 2353 4460
rect 2387 4426 2425 4460
rect 2459 4426 2497 4460
rect 2531 4426 2569 4460
rect 2603 4426 2641 4460
rect 2675 4426 2713 4460
rect 2747 4426 2785 4460
rect 2819 4426 2857 4460
rect 2891 4426 2929 4460
rect 2963 4426 3001 4460
rect 3035 4426 3073 4460
rect 3107 4426 3145 4460
rect 3179 4426 3217 4460
rect 3251 4426 3289 4460
rect 3323 4426 3361 4460
rect 3395 4426 3433 4460
rect 3467 4426 3505 4460
rect 3539 4426 3577 4460
rect 3611 4426 3649 4460
rect 3683 4426 3721 4460
rect 3755 4426 3793 4460
rect 3827 4426 3865 4460
rect 3899 4426 3937 4460
rect 3971 4426 4009 4460
rect 4043 4426 4081 4460
rect 4115 4426 4153 4460
rect 4187 4426 4225 4460
rect 4259 4426 4297 4460
rect 4331 4426 4369 4460
rect 4403 4426 4441 4460
rect 4475 4426 4513 4460
rect 4547 4426 4585 4460
rect 4619 4426 4657 4460
rect 4691 4426 4729 4460
rect 4763 4426 4801 4460
rect 4835 4426 4873 4460
rect 4907 4426 4945 4460
rect 4979 4426 5017 4460
rect 5051 4426 5089 4460
rect 5123 4426 5161 4460
rect 5195 4426 5233 4460
rect 5267 4426 5305 4460
rect 5339 4426 5377 4460
rect 5411 4426 5449 4460
rect 5483 4426 5521 4460
rect 5555 4426 5593 4460
rect 5627 4426 5665 4460
rect 5699 4426 5737 4460
rect 5771 4426 5809 4460
rect 5843 4426 5881 4460
rect 5915 4426 5953 4460
rect 5987 4426 6025 4460
rect 6059 4426 6097 4460
rect 6131 4426 6169 4460
rect 6203 4426 6241 4460
rect 6275 4426 6313 4460
rect 6347 4426 6385 4460
rect 6419 4426 6457 4460
rect 6491 4426 6529 4460
rect 6563 4426 6601 4460
rect 6635 4426 6673 4460
rect 6707 4426 6745 4460
rect 6779 4426 6817 4460
rect 6851 4426 6889 4460
rect 6923 4426 6961 4460
rect 6995 4426 7033 4460
rect 7067 4426 7105 4460
rect 7139 4426 7177 4460
rect 7211 4426 7249 4460
rect 7283 4426 7321 4460
rect 7355 4426 7393 4460
rect 7427 4426 7465 4460
rect 7499 4426 7537 4460
rect 7571 4426 7609 4460
rect 7643 4426 7681 4460
rect 7715 4426 7753 4460
rect 7787 4426 7825 4460
rect 7859 4426 7897 4460
rect 7931 4426 7969 4460
rect 8003 4426 8041 4460
rect 8075 4426 8113 4460
rect 8147 4426 8185 4460
rect 8219 4426 8257 4460
rect 8291 4426 8329 4460
rect 8363 4426 8401 4460
rect 8435 4426 8473 4460
rect 8507 4426 8545 4460
rect 8579 4426 8617 4460
rect 8651 4426 8689 4460
rect 8723 4426 8761 4460
rect 8795 4426 8833 4460
rect 8867 4426 8905 4460
rect 8939 4426 8977 4460
rect 9011 4426 9049 4460
rect 9083 4426 9121 4460
rect 9155 4426 9193 4460
rect 9227 4426 9265 4460
rect 9299 4426 9337 4460
rect 9371 4426 9409 4460
rect 9443 4426 9481 4460
rect 9515 4426 9553 4460
rect 9587 4426 9625 4460
rect 9659 4426 9697 4460
rect 9731 4426 9769 4460
rect 9803 4426 9841 4460
rect 9875 4426 9913 4460
rect 9947 4426 9985 4460
rect 10019 4426 10057 4460
rect 10091 4426 10129 4460
rect 10163 4426 10201 4460
rect 10235 4426 10273 4460
rect 10307 4426 10345 4460
rect 10379 4426 10417 4460
rect 10451 4426 10489 4460
rect 10523 4426 10561 4460
rect 10595 4454 12408 4460
rect 10595 4426 12031 4454
rect 1525 4420 12031 4426
rect 12065 4420 12112 4454
rect 12146 4420 12193 4454
rect 12227 4420 12274 4454
rect 12308 4420 12408 4454
rect 1525 4415 12408 4420
rect 1525 4381 12347 4415
rect 12402 4381 12408 4415
rect -183 4365 -103 4377
rect -183 4331 -177 4365
rect -143 4331 -103 4365
rect -183 4325 -103 4331
tri 11882 4349 11914 4381 ne
rect 11914 4363 12347 4381
rect 12399 4363 12408 4381
rect 11914 4350 12408 4363
rect 11914 4349 12347 4350
tri 12310 4342 12317 4349 ne
rect 12317 4342 12347 4349
tri 325 4340 327 4342 se
rect 327 4340 4286 4342
tri 4286 4340 4288 4342 sw
tri 12317 4340 12319 4342 ne
rect 12319 4340 12347 4342
rect 12399 4340 12408 4350
tri 323 4338 325 4340 se
rect 325 4338 4288 4340
tri 4288 4338 4290 4340 sw
tri 12319 4339 12320 4340 ne
rect 12320 4339 12347 4340
tri 318 4333 323 4338 se
rect 323 4333 4290 4338
tri 4290 4333 4295 4338 sw
rect 4489 4333 5636 4339
rect -183 4319 -51 4325
tri 304 4319 318 4333 se
rect 318 4319 4295 4333
rect -373 4283 -367 4317
rect -333 4283 -327 4317
tri 284 4299 304 4319 se
rect 304 4299 4295 4319
tri 4295 4299 4329 4333 sw
rect 4489 4299 4501 4333
rect 4535 4299 4573 4333
rect 4607 4299 4645 4333
rect 4679 4299 4717 4333
rect 4751 4299 4789 4333
rect 4823 4299 4861 4333
rect 4895 4299 4933 4333
rect 4967 4299 5005 4333
rect 5039 4299 5077 4333
rect 5111 4299 5149 4333
rect 5183 4299 5221 4333
rect 5255 4299 5293 4333
rect 5327 4299 5365 4333
rect 5399 4299 5437 4333
rect 5471 4299 5509 4333
rect 5543 4299 5581 4333
rect 5615 4321 5636 4333
tri 5636 4321 5654 4339 sw
tri 12320 4321 12338 4339 ne
rect 12338 4321 12347 4339
rect 5615 4319 5654 4321
tri 5654 4319 5656 4321 sw
tri 12338 4319 12340 4321 ne
rect 12340 4319 12347 4321
rect 5615 4313 5656 4319
tri 5656 4313 5662 4319 sw
rect 11862 4313 12285 4319
rect 5615 4312 5662 4313
tri 5662 4312 5663 4313 sw
rect 5615 4299 5663 4312
rect -373 4245 -327 4283
tri 265 4280 284 4299 se
rect 284 4290 4329 4299
rect 284 4280 338 4290
rect -373 4211 -367 4245
rect -333 4211 -327 4245
rect -373 4199 -327 4211
rect -187 4279 -135 4280
tri -135 4279 -134 4280 sw
tri 264 4279 265 4280 se
rect 265 4279 338 4280
tri 338 4279 349 4290 nw
tri 4264 4279 4275 4290 ne
rect 4275 4279 4329 4290
tri 4329 4279 4349 4299 sw
rect 4489 4293 5663 4299
tri 5616 4280 5629 4293 ne
rect 5629 4280 5663 4293
tri 5663 4280 5695 4312 sw
tri 5629 4279 5630 4280 ne
rect 5630 4279 5695 4280
tri 5695 4279 5696 4280 sw
rect 11862 4279 11874 4313
rect 11908 4279 11946 4313
rect 11980 4279 12233 4313
rect -187 4274 -134 4279
rect -135 4268 -134 4274
tri -134 4268 -123 4279 sw
tri 253 4268 264 4279 se
rect 264 4268 327 4279
tri 327 4268 338 4279 nw
tri 4275 4268 4286 4279 ne
rect 4286 4268 4349 4279
rect -135 4265 -123 4268
tri -123 4265 -120 4268 sw
tri 250 4265 253 4268 se
rect 253 4265 324 4268
tri 324 4265 327 4268 nw
tri 4286 4265 4289 4268 ne
rect 4289 4265 4349 4268
tri 4349 4265 4363 4279 sw
tri 5630 4265 5644 4279 ne
rect 5644 4273 5696 4279
tri 5696 4273 5702 4279 sw
rect 11862 4273 12233 4279
rect 5644 4265 5702 4273
tri 5702 4265 5710 4273 sw
tri 12186 4265 12194 4273 ne
rect 12194 4265 12233 4273
rect -135 4264 -120 4265
tri -120 4264 -119 4265 sw
tri 249 4264 250 4265 se
rect 250 4264 323 4265
tri 323 4264 324 4265 nw
tri 4289 4264 4290 4265 ne
rect 4290 4264 4363 4265
tri 4363 4264 4364 4265 sw
tri 5644 4264 5645 4265 ne
rect 5645 4264 5710 4265
rect -135 4261 -119 4264
tri -119 4261 -116 4264 sw
tri 246 4261 249 4264 se
rect 249 4261 314 4264
rect -135 4255 -116 4261
tri -116 4255 -110 4261 sw
tri 240 4255 246 4261 se
rect 246 4255 314 4261
tri 314 4255 323 4264 nw
tri 4290 4261 4293 4264 ne
rect 4293 4261 5178 4264
rect 1524 4255 2103 4261
rect 2155 4255 2167 4261
rect -135 4246 -110 4255
tri -110 4246 -101 4255 sw
tri 231 4246 240 4255 se
rect 240 4246 305 4255
tri 305 4246 314 4255 nw
rect -135 4240 280 4246
rect -135 4222 -26 4240
rect -187 4210 -26 4222
rect -135 4206 -26 4210
rect 8 4206 46 4240
rect 80 4221 280 4240
tri 280 4221 305 4246 nw
rect 1524 4221 1536 4255
rect 1570 4221 1613 4255
rect 1647 4221 1690 4255
rect 1724 4221 1767 4255
rect 1801 4221 1844 4255
rect 1878 4221 1921 4255
rect 1955 4221 1997 4255
rect 2031 4221 2073 4255
rect 80 4215 274 4221
tri 274 4215 280 4221 nw
rect 80 4206 259 4215
rect -135 4200 259 4206
tri 259 4200 274 4215 nw
rect 1524 4209 2103 4221
rect 2155 4209 2167 4221
rect 2219 4209 2225 4261
rect 2254 4255 2453 4261
rect 2505 4255 2517 4261
rect 2254 4221 2266 4255
rect 2300 4221 2343 4255
rect 2377 4221 2420 4255
rect 2254 4215 2453 4221
tri 2441 4212 2444 4215 ne
rect 2444 4212 2453 4215
tri 2444 4209 2447 4212 ne
rect 2447 4209 2453 4212
rect 2505 4209 2517 4221
rect 2569 4209 2575 4261
rect 2613 4209 2619 4261
rect 2671 4209 2683 4261
rect 2735 4255 4198 4261
rect 2735 4221 3072 4255
rect 3106 4221 3144 4255
rect 3178 4221 3216 4255
rect 3250 4221 3288 4255
rect 3322 4221 3360 4255
rect 3394 4221 3432 4255
rect 3466 4221 3504 4255
rect 3538 4221 3576 4255
rect 3610 4221 3648 4255
rect 3682 4221 3720 4255
rect 3754 4221 3792 4255
rect 3826 4221 3864 4255
rect 3898 4221 3936 4255
rect 3970 4221 4008 4255
rect 4042 4221 4080 4255
rect 4114 4221 4152 4255
rect 4186 4221 4198 4255
tri 4293 4253 4301 4261 ne
rect 4301 4253 5178 4261
tri 4301 4251 4303 4253 ne
rect 4303 4251 5178 4253
tri 4303 4249 4305 4251 ne
rect 4305 4249 5178 4251
tri 4305 4246 4308 4249 ne
rect 4308 4246 5178 4249
rect 2735 4209 4198 4221
tri 4308 4215 4339 4246 ne
rect 4339 4215 5178 4246
tri 4339 4212 4342 4215 ne
rect 4342 4212 5178 4215
rect 5230 4212 5242 4264
rect 5294 4212 5301 4264
tri 5645 4261 5648 4264 ne
rect 5648 4261 5710 4264
tri 5710 4261 5714 4265 sw
tri 12194 4261 12198 4265 ne
rect 12198 4261 12233 4265
tri 12340 4312 12347 4319 ne
tri 5648 4255 5654 4261 ne
rect 5654 4255 5714 4261
tri 5714 4255 5720 4261 sw
tri 5654 4253 5656 4255 ne
rect 5656 4253 5836 4255
tri 5656 4251 5658 4253 ne
rect 5658 4251 5836 4253
tri 5658 4249 5660 4251 ne
rect 5660 4249 5836 4251
tri 5660 4246 5663 4249 ne
rect 5663 4246 5836 4249
tri 5663 4215 5694 4246 ne
rect 5694 4215 5836 4246
tri 5694 4212 5697 4215 ne
rect 5697 4212 5836 4215
tri 5697 4209 5700 4212 ne
rect 5700 4209 5836 4212
rect 5837 4210 5838 4254
rect 5874 4210 5875 4254
rect 5876 4249 7077 4255
rect 5876 4215 5951 4249
rect 5985 4215 6023 4249
rect 6057 4215 6095 4249
rect 6129 4215 6167 4249
rect 6201 4215 6239 4249
rect 6273 4215 6311 4249
rect 6345 4215 6383 4249
rect 6417 4215 6455 4249
rect 6489 4215 6527 4249
rect 6561 4215 6599 4249
rect 6633 4215 6671 4249
rect 6705 4215 6743 4249
rect 6777 4215 6815 4249
rect 6849 4215 6887 4249
rect 6921 4215 6959 4249
rect 6993 4215 7031 4249
rect 7065 4215 7077 4249
rect 5876 4209 7077 4215
rect 7161 4249 7210 4261
rect 7262 4249 7274 4261
rect 7161 4215 7173 4249
rect 7207 4215 7210 4249
rect 7161 4209 7210 4215
rect 7262 4209 7274 4215
rect 7326 4209 7332 4261
rect 7462 4251 7602 4261
rect 7462 4217 7506 4251
rect 7540 4217 7578 4251
rect 7462 4209 7602 4217
rect 7654 4209 7666 4261
rect 7718 4209 7724 4261
rect 7752 4209 7758 4261
rect 7810 4209 7822 4261
rect 7874 4251 8837 4261
tri 12198 4259 12200 4261 ne
rect 12200 4259 12285 4261
rect 7874 4217 7898 4251
rect 7932 4217 8837 4251
rect 7874 4209 8837 4217
rect 9253 4253 10726 4259
rect 10837 4253 11054 4259
rect 9253 4219 9265 4253
rect 9299 4219 9337 4253
rect 9371 4219 9570 4253
rect 9604 4219 9642 4253
rect 9676 4219 10607 4253
rect 10641 4219 10679 4253
rect 10713 4219 10726 4253
tri 10803 4219 10837 4253 se
rect 9253 4213 10726 4219
tri 10797 4213 10803 4219 se
rect 10803 4213 10837 4219
tri 10793 4209 10797 4213 se
rect 10797 4209 10837 4213
tri 10784 4200 10793 4209 se
rect 10793 4201 10837 4209
rect 10889 4219 10936 4253
rect 10970 4219 11008 4253
rect 11042 4219 11054 4253
tri 12200 4232 12227 4259 ne
rect 12227 4249 12285 4259
rect 12227 4232 12233 4249
rect 10889 4213 11054 4219
rect 12139 4220 12185 4232
tri 12227 4231 12228 4232 ne
rect 12228 4231 12233 4232
tri 12228 4226 12233 4231 ne
rect 10889 4201 10902 4213
rect 10793 4200 10902 4201
rect -135 4186 -114 4200
tri -114 4186 -100 4200 nw
tri 10777 4193 10784 4200 se
rect 10784 4193 10902 4200
tri 10902 4193 10922 4213 nw
tri 10770 4186 10777 4193 se
rect 10777 4191 10900 4193
tri 10900 4191 10902 4193 nw
rect 10777 4189 10895 4191
rect 10777 4186 10837 4189
rect -135 4181 -119 4186
tri -119 4181 -114 4186 nw
tri 10765 4181 10770 4186 se
rect 10770 4181 10837 4186
rect -135 4167 -133 4181
tri -133 4167 -119 4181 nw
tri -135 4165 -133 4167 nw
rect -187 4152 -135 4158
rect 238 4140 311 4146
rect 290 4134 311 4140
rect -645 4116 152 4122
rect -593 4108 -545 4116
rect -493 4110 152 4116
rect -593 4074 -566 4108
rect -493 4076 -277 4110
rect -243 4076 152 4110
rect -593 4064 -545 4074
rect -493 4064 152 4076
rect -645 4039 152 4064
rect -593 4031 -545 4039
rect -493 4038 152 4039
rect -593 3997 -566 4031
rect -493 4004 -277 4038
rect -243 4004 152 4038
rect -593 3987 -545 3997
rect -493 3987 152 4004
rect -645 3962 152 3987
rect -593 3954 -545 3962
rect -593 3920 -566 3954
rect -593 3910 -545 3920
rect -493 3910 152 3962
rect -645 3885 152 3910
rect -593 3876 -545 3885
rect -593 3842 -566 3876
rect -493 3868 152 3885
rect -593 3833 -545 3842
rect -493 3834 -314 3868
rect -280 3834 -190 3868
rect -156 3834 152 3868
rect -493 3833 152 3834
rect -645 3808 152 3833
rect -593 3798 -545 3808
rect -593 3764 -566 3798
rect -493 3796 152 3808
rect -593 3756 -545 3764
rect -493 3762 -314 3796
rect -280 3762 -190 3796
rect -156 3762 152 3796
rect 305 4100 311 4134
rect 290 4088 311 4100
rect 238 4061 311 4088
rect 290 4054 311 4061
rect 305 4020 311 4054
rect 290 4009 311 4020
rect 238 3986 311 4009
rect 470 4129 1704 4181
rect 1756 4129 1773 4181
rect 1825 4129 1842 4181
rect 1894 4129 1911 4181
rect 1963 4129 1980 4181
rect 2032 4129 3156 4181
rect 3208 4129 3220 4181
rect 3272 4129 3284 4181
rect 3336 4129 3348 4181
rect 3400 4129 3412 4181
rect 3464 4129 3476 4181
rect 3528 4129 3540 4181
rect 3592 4164 9075 4181
tri 10757 4173 10765 4181 se
rect 10765 4173 10837 4181
rect 3592 4129 8751 4164
rect 470 4106 8751 4129
rect 470 4054 1704 4106
rect 1756 4054 1773 4106
rect 1825 4054 1842 4106
rect 1894 4054 1911 4106
rect 1963 4054 1980 4106
rect 2032 4054 3156 4106
rect 3208 4054 3220 4106
rect 3272 4054 3284 4106
rect 3336 4054 3348 4106
rect 3400 4054 3412 4106
rect 3464 4054 3476 4106
rect 3528 4054 3540 4106
rect 3592 4054 8751 4106
rect 470 4031 8751 4054
tri 311 3986 317 3992 sw
rect 238 3982 317 3986
rect 290 3979 317 3982
tri 317 3979 324 3986 sw
rect 470 3979 1704 4031
rect 1756 3979 1773 4031
rect 1825 3979 1842 4031
rect 1894 3979 1911 4031
rect 1963 3979 1980 4031
rect 2032 3979 3156 4031
rect 3208 3979 3220 4031
rect 3272 3979 3284 4031
rect 3336 3979 3348 4031
rect 3400 3979 3412 4031
rect 3464 3979 3476 4031
rect 3528 3979 3540 4031
rect 3592 3986 8751 4031
rect 9001 3986 9075 4164
rect 9696 4167 10837 4173
rect 9139 4152 9497 4154
rect 9139 4142 9147 4152
rect 9139 4108 9145 4142
rect 9139 4100 9147 4108
rect 9199 4100 9214 4152
rect 9266 4100 9280 4152
rect 9332 4142 9497 4152
rect 9332 4108 9457 4142
rect 9491 4108 9497 4142
rect 9696 4133 9708 4167
rect 9742 4133 9780 4167
rect 9814 4133 10011 4167
rect 10045 4133 10083 4167
rect 10117 4133 10324 4167
rect 10358 4133 10396 4167
rect 10430 4137 10837 4167
rect 10889 4186 10895 4189
tri 10895 4186 10900 4191 nw
rect 12139 4186 12145 4220
rect 12179 4186 12185 4220
rect 12233 4191 12285 4197
rect 12402 4306 12408 4340
rect 12399 4298 12408 4306
rect 12347 4285 12408 4298
rect 12399 4265 12408 4285
rect 12347 4231 12368 4233
rect 12402 4231 12408 4265
rect 14840 4258 15007 4414
rect 12347 4220 12408 4231
tri 10889 4180 10895 4186 nw
rect 10430 4133 10889 4137
rect 9696 4131 10889 4133
rect 12139 4148 12185 4186
rect 9696 4127 10777 4131
tri 10777 4127 10781 4131 nw
rect 9332 4100 9497 4108
rect 9139 4054 9497 4100
rect 10942 4109 11074 4115
rect 9139 4046 9147 4054
rect 9139 4012 9145 4046
rect 9139 4002 9147 4012
rect 9199 4002 9214 4054
rect 9266 4002 9280 4054
rect 9332 4046 9497 4054
rect 9845 4090 10568 4096
rect 9845 4056 9857 4090
rect 9891 4056 9929 4090
rect 9963 4056 10450 4090
rect 10484 4056 10522 4090
rect 10556 4056 10568 4090
rect 9845 4050 10568 4056
rect 10942 4075 10956 4109
rect 10990 4075 11000 4109
rect 11062 4075 11074 4109
rect 10942 4057 11000 4075
rect 11052 4057 11074 4075
rect 9332 4012 9457 4046
rect 9491 4012 9497 4046
rect 10942 4045 11074 4057
rect 9332 4002 9497 4012
rect 9139 4000 9497 4002
rect 10158 4012 10881 4018
rect 3592 3979 9075 3986
rect 290 3978 324 3979
tri 324 3978 325 3979 sw
rect 10158 3978 10170 4012
rect 10204 3978 10242 4012
rect 10276 3978 10763 4012
rect 10797 3978 10835 4012
rect 10869 3978 10881 4012
rect 290 3974 325 3978
rect 305 3951 325 3974
tri 325 3951 352 3978 sw
rect 10158 3972 10881 3978
rect 10942 3993 11000 4045
rect 11052 4009 11074 4045
rect 11052 4006 11071 4009
tri 11071 4006 11074 4009 nw
rect 12139 4114 12145 4148
rect 12179 4114 12185 4148
rect 10942 3987 11052 3993
tri 11052 3987 11071 4006 nw
rect 10942 3983 11048 3987
tri 11048 3983 11052 3987 nw
rect 11867 3986 11997 3992
rect 11867 3983 11886 3986
rect 11938 3983 11997 3986
rect 10942 3972 11037 3983
tri 11037 3972 11048 3983 nw
rect 305 3949 352 3951
tri 352 3949 354 3951 sw
rect 305 3945 354 3949
tri 354 3945 358 3949 sw
rect 1342 3945 2619 3951
rect 305 3940 358 3945
rect 290 3934 358 3940
tri 358 3934 369 3945 sw
rect 290 3930 1248 3934
rect 238 3923 1248 3930
rect 238 3903 829 3923
rect 290 3893 829 3903
rect 305 3871 829 3893
rect 881 3871 902 3923
rect 954 3871 974 3923
rect 1026 3871 1046 3923
rect 1098 3871 1118 3923
rect 1170 3871 1190 3923
rect 1242 3871 1248 3923
rect 1342 3911 1354 3945
rect 1388 3911 1426 3945
rect 1460 3911 1655 3945
rect 1689 3911 1727 3945
rect 1761 3911 1966 3945
rect 2000 3911 2038 3945
rect 2072 3911 2619 3945
rect 1342 3899 2619 3911
rect 2671 3899 2683 3951
rect 2735 3899 2741 3951
tri 3673 3899 3694 3920 se
rect 3694 3901 4087 3920
tri 4087 3901 4106 3920 sw
rect 3694 3899 4106 3901
tri 4106 3899 4108 3901 sw
rect 8031 3899 8037 3951
rect 8089 3899 8101 3951
rect 8153 3945 10053 3951
rect 8153 3923 10001 3945
rect 8153 3899 8522 3923
tri 8522 3899 8546 3923 nw
tri 9528 3899 9552 3923 ne
rect 9552 3899 10001 3923
tri 3666 3892 3673 3899 se
rect 3673 3895 4108 3899
tri 4108 3895 4112 3899 sw
tri 9552 3895 9556 3899 ne
rect 9556 3895 10001 3899
rect 3673 3892 4112 3895
tri 4112 3892 4115 3895 sw
tri 3663 3889 3666 3892 se
rect 3666 3891 4115 3892
tri 4115 3891 4116 3892 sw
rect 3666 3889 4116 3891
tri 4116 3889 4118 3891 sw
tri 7532 3889 7534 3891 se
rect 7534 3889 7870 3891
tri 7870 3889 7872 3891 sw
tri 3660 3886 3663 3889 se
rect 3663 3886 4118 3889
tri 4118 3886 4121 3889 sw
tri 7529 3886 7532 3889 se
rect 7532 3886 7872 3889
tri 7872 3886 7875 3889 sw
rect 8599 3886 9126 3895
tri 3653 3879 3660 3886 se
rect 3660 3879 4121 3886
tri 4121 3879 4128 3886 sw
tri 7522 3879 7529 3886 se
rect 7529 3879 7875 3886
tri 7875 3879 7882 3886 sw
tri 3645 3871 3653 3879 se
rect 3653 3871 4128 3879
tri 4128 3871 4136 3879 sw
tri 7514 3871 7522 3879 se
rect 7522 3871 7882 3879
rect 305 3861 1248 3871
rect 305 3859 379 3861
tri 379 3859 381 3861 nw
rect 2267 3859 2453 3871
rect 290 3851 345 3859
rect 238 3825 345 3851
tri 345 3825 379 3859 nw
rect 2267 3825 2279 3859
rect 2313 3825 2351 3859
rect 2385 3825 2453 3859
rect 238 3824 343 3825
rect 290 3823 343 3824
tri 343 3823 345 3825 nw
rect 290 3820 340 3823
tri 340 3820 343 3823 nw
rect 290 3817 337 3820
tri 337 3817 340 3820 nw
rect 2267 3819 2453 3825
rect 2505 3819 2517 3871
rect 2569 3868 7882 3871
tri 7882 3868 7893 3879 sw
rect 2569 3859 3700 3868
rect 2569 3825 2590 3859
rect 2624 3825 2662 3859
rect 2696 3852 3700 3859
tri 3700 3852 3716 3868 nw
tri 4065 3852 4081 3868 ne
rect 4081 3852 7893 3868
tri 7893 3852 7909 3868 sw
rect 8599 3852 8611 3886
rect 8645 3852 8683 3886
rect 8717 3852 9126 3886
rect 2696 3843 3691 3852
tri 3691 3843 3700 3852 nw
tri 4081 3843 4090 3852 ne
rect 4090 3843 7909 3852
tri 7909 3843 7918 3852 sw
rect 8599 3843 9126 3852
rect 9178 3843 9190 3895
rect 9242 3843 9296 3895
rect 9298 3894 9334 3895
rect 9297 3844 9335 3894
rect 9298 3843 9334 3844
rect 9336 3843 9371 3895
rect 9423 3843 9435 3895
rect 9487 3843 9493 3895
tri 9556 3892 9559 3895 ne
rect 9559 3893 10001 3895
rect 10942 3949 11014 3972
tri 11014 3949 11037 3972 nw
rect 11867 3949 11879 3983
rect 11938 3949 11951 3983
rect 11985 3949 11997 3983
rect 10942 3943 11008 3949
tri 11008 3943 11014 3949 nw
tri 10930 3931 10942 3943 se
rect 10942 3931 10996 3943
tri 10996 3931 11008 3943 nw
rect 11867 3934 11886 3949
rect 11938 3934 11997 3949
tri 10919 3920 10930 3931 se
rect 10930 3920 10966 3931
tri 10900 3901 10919 3920 se
rect 10919 3901 10966 3920
tri 10966 3901 10996 3931 nw
rect 11867 3922 11997 3934
rect 9559 3892 10053 3893
tri 9559 3889 9562 3892 ne
rect 9562 3889 10053 3892
tri 9562 3879 9572 3889 ne
rect 9572 3881 10053 3889
rect 9572 3879 10001 3881
tri 9945 3855 9969 3879 ne
rect 9969 3855 10001 3879
tri 9969 3843 9981 3855 ne
rect 9981 3843 10001 3855
rect 2696 3825 3671 3843
rect 2569 3823 3671 3825
tri 3671 3823 3691 3843 nw
tri 4090 3823 4110 3843 ne
rect 4110 3839 7918 3843
tri 7918 3839 7922 3843 sw
tri 9981 3839 9985 3843 ne
rect 9985 3839 10001 3843
rect 4110 3823 7540 3839
tri 7540 3823 7556 3839 nw
tri 7848 3823 7864 3839 ne
rect 7864 3823 7922 3839
tri 7922 3823 7938 3839 sw
tri 9985 3823 10001 3839 ne
rect 10001 3823 10053 3829
rect 10119 3892 10957 3901
tri 10957 3892 10966 3901 nw
rect 10119 3889 10923 3892
rect 10119 3855 10125 3889
rect 10159 3855 10285 3889
rect 10319 3858 10923 3889
tri 10923 3858 10957 3892 nw
rect 11867 3870 11886 3922
rect 11938 3870 11997 3922
rect 11867 3864 11997 3870
rect 12139 3892 12185 4114
rect 12139 3858 12145 3892
rect 12179 3858 12185 3892
rect 10319 3856 10921 3858
tri 10921 3856 10923 3858 nw
rect 10319 3855 10920 3856
tri 10920 3855 10921 3856 nw
rect 2569 3820 3668 3823
tri 3668 3820 3671 3823 nw
tri 4110 3820 4113 3823 ne
rect 4113 3820 7537 3823
tri 7537 3820 7540 3823 nw
tri 7864 3820 7867 3823 ne
rect 7867 3820 7938 3823
tri 7938 3820 7941 3823 sw
rect 10119 3820 10474 3855
tri 10474 3820 10509 3855 nw
rect 12139 3820 12185 3858
rect 2569 3819 3667 3820
tri 3667 3819 3668 3820 nw
tri 4113 3819 4114 3820 ne
rect 4114 3819 7536 3820
tri 7536 3819 7537 3820 nw
tri 7867 3819 7868 3820 ne
rect 7868 3819 7941 3820
tri 7868 3817 7870 3819 ne
rect 7870 3817 7941 3819
tri 7941 3817 7944 3820 sw
rect 10119 3817 10453 3820
rect 290 3812 315 3817
rect 305 3795 315 3812
tri 315 3795 337 3817 nw
tri 7870 3811 7876 3817 ne
rect 7876 3815 7944 3817
tri 7944 3815 7946 3817 sw
rect 7876 3811 9282 3815
tri 1973 3795 1985 3807 se
rect 1985 3795 2238 3807
tri 2238 3795 2250 3807 sw
rect 305 3778 311 3795
tri 311 3791 315 3795 nw
tri 1969 3791 1973 3795 se
rect 1973 3791 2250 3795
tri 2250 3791 2254 3795 sw
rect 290 3772 311 3778
tri 384 3773 402 3791 se
rect 402 3773 2871 3791
rect 238 3766 311 3772
tri 380 3769 384 3773 se
rect 384 3769 1995 3773
tri 1995 3769 1999 3773 nw
tri 2229 3769 2233 3773 ne
rect 2233 3769 2871 3773
tri 377 3766 380 3769 se
rect 380 3766 1987 3769
rect -493 3756 152 3762
tri 372 3761 377 3766 se
rect 377 3761 1987 3766
tri 1987 3761 1995 3769 nw
tri 2233 3761 2241 3769 ne
rect 2241 3761 2871 3769
tri 368 3757 372 3761 se
rect 372 3757 1983 3761
tri 1983 3757 1987 3761 nw
tri 2241 3757 2245 3761 ne
rect 2245 3757 2871 3761
rect -645 3750 152 3756
tri 361 3750 368 3757 se
rect 368 3750 409 3757
tri 409 3750 416 3757 nw
tri 2847 3750 2854 3757 ne
rect 2854 3750 2871 3757
tri 334 3723 361 3750 se
rect 361 3739 398 3750
tri 398 3739 409 3750 nw
tri 2854 3739 2865 3750 ne
rect 2865 3739 2871 3750
rect 2923 3739 2935 3791
rect 2987 3739 2993 3791
rect 3826 3757 3832 3809
rect 3884 3757 3896 3809
rect 3948 3795 3954 3809
tri 3954 3795 3968 3809 sw
rect 7672 3805 7726 3811
rect 3948 3791 3968 3795
tri 3968 3791 3972 3795 sw
rect 3948 3769 5956 3791
tri 5956 3769 5978 3791 sw
rect 3948 3766 5978 3769
tri 5978 3766 5981 3769 sw
rect 3948 3757 6753 3766
tri 5916 3739 5934 3757 ne
rect 5934 3739 6753 3757
rect 361 3725 384 3739
tri 384 3725 398 3739 nw
tri 5934 3735 5938 3739 ne
rect 5938 3735 6753 3739
tri 2091 3729 2097 3735 se
rect 2097 3729 2103 3735
rect 361 3723 382 3725
tri 382 3723 384 3725 nw
tri 430 3723 432 3725 se
rect 432 3723 825 3725
tri 330 3719 334 3723 se
rect 334 3719 378 3723
tri 378 3719 382 3723 nw
tri 426 3719 430 3723 se
rect 430 3719 825 3723
tri 325 3714 330 3719 se
rect 330 3714 372 3719
rect -463 3708 -354 3714
tri -243 3713 -242 3714 se
rect -242 3713 372 3714
tri 372 3713 378 3719 nw
tri 420 3713 426 3719 se
rect 426 3713 707 3719
tri -246 3710 -243 3713 se
rect -243 3710 369 3713
tri 369 3710 372 3713 nw
tri 417 3710 420 3713 se
rect 420 3710 707 3713
tri -247 3709 -246 3710 se
rect -246 3709 368 3710
tri 368 3709 369 3710 nw
tri 416 3709 417 3710 se
rect 417 3709 707 3710
rect -411 3702 -354 3708
rect -411 3668 -394 3702
rect -360 3668 -354 3702
tri -271 3685 -247 3709 se
rect -247 3685 344 3709
tri 344 3685 368 3709 nw
tri 392 3685 416 3709 se
rect 416 3685 707 3709
rect 741 3685 779 3719
rect 813 3685 825 3719
tri -276 3680 -271 3685 se
rect -271 3680 339 3685
tri 339 3680 344 3685 nw
tri 387 3680 392 3685 se
rect 392 3680 825 3685
rect 1524 3723 2103 3729
rect 2155 3723 2167 3735
rect 2219 3729 2225 3735
tri 2225 3729 2231 3735 sw
tri 5938 3729 5944 3735 ne
rect 5944 3729 6753 3735
rect 2219 3723 2830 3729
rect 1524 3689 1536 3723
rect 1570 3689 1608 3723
rect 1642 3689 1810 3723
rect 1844 3689 1882 3723
rect 1916 3689 2103 3723
rect 2156 3689 2167 3723
rect 2228 3689 2434 3723
rect 2468 3689 2506 3723
rect 2540 3689 2712 3723
rect 2746 3689 2784 3723
rect 2818 3689 2830 3723
rect 1524 3683 2103 3689
rect 2155 3683 2167 3689
rect 2219 3683 2830 3689
rect 3086 3723 4180 3729
rect 4182 3728 4218 3729
rect 3086 3689 3098 3723
rect 3132 3689 3170 3723
rect 3204 3689 3416 3723
rect 3450 3689 3488 3723
rect 3522 3689 3722 3723
rect 3756 3689 3794 3723
rect 3828 3689 4033 3723
rect 4067 3689 4105 3723
rect 4139 3689 4180 3723
rect 3086 3683 4180 3689
rect 4181 3684 4219 3728
rect 4220 3723 5717 3729
tri 5944 3723 5950 3729 ne
rect 5950 3723 6753 3729
rect 4220 3689 4423 3723
rect 4457 3689 4495 3723
rect 4529 3689 4697 3723
rect 4731 3689 4769 3723
rect 4803 3689 5009 3723
rect 5043 3689 5081 3723
rect 5115 3689 5321 3723
rect 5355 3689 5393 3723
rect 5427 3689 5599 3723
rect 5633 3689 5671 3723
rect 5705 3689 5717 3723
tri 5950 3714 5959 3723 ne
rect 5959 3714 6753 3723
rect 6805 3714 6817 3766
rect 6869 3714 6875 3766
rect 7724 3753 7726 3805
rect 7672 3741 7726 3753
rect 4182 3683 4218 3684
rect 4220 3683 5717 3689
rect 7724 3689 7726 3741
rect 7672 3683 7726 3689
rect 7727 3684 7728 3810
rect 7764 3684 7765 3810
rect 7766 3809 7836 3811
tri 7836 3809 7838 3811 sw
tri 7876 3809 7878 3811 ne
rect 7878 3809 9282 3811
rect 7766 3801 7838 3809
tri 7838 3801 7846 3809 sw
tri 7878 3801 7886 3809 ne
rect 7886 3801 9282 3809
rect 7766 3795 7846 3801
rect 7766 3761 7795 3795
rect 7829 3791 7846 3795
tri 7846 3791 7856 3801 sw
tri 7886 3791 7896 3801 ne
rect 7896 3791 9282 3801
rect 7829 3783 7856 3791
tri 7856 3783 7864 3791 sw
tri 7896 3783 7904 3791 ne
rect 7904 3783 9282 3791
rect 7829 3775 7864 3783
tri 7864 3775 7872 3783 sw
tri 7904 3775 7912 3783 ne
rect 7912 3775 9282 3783
rect 7829 3769 7872 3775
tri 7872 3769 7878 3775 sw
tri 7912 3769 7918 3775 ne
rect 7918 3769 9282 3775
rect 7829 3766 7878 3769
tri 7878 3766 7881 3769 sw
tri 7918 3766 7921 3769 ne
rect 7921 3766 9282 3769
rect 7829 3765 7881 3766
tri 7881 3765 7882 3766 sw
tri 7921 3765 7922 3766 ne
rect 7922 3765 9282 3766
rect 7829 3763 7882 3765
tri 7882 3763 7884 3765 sw
tri 7922 3763 7924 3765 ne
rect 7924 3763 9282 3765
rect 9334 3763 9346 3815
rect 9398 3763 9404 3815
rect 10119 3783 10125 3817
rect 10159 3783 10285 3817
rect 10319 3799 10453 3817
tri 10453 3799 10474 3820 nw
rect 10595 3799 10992 3805
rect 10319 3783 10425 3799
rect 10119 3771 10425 3783
tri 10425 3771 10453 3799 nw
rect 10595 3765 10607 3799
rect 10641 3765 10679 3799
rect 10713 3765 10874 3799
rect 10908 3765 10946 3799
rect 10980 3765 10992 3799
rect 12139 3786 12145 3820
rect 12179 3786 12185 3820
rect 12139 3774 12185 3786
rect 12399 4190 12408 4220
rect 12347 4156 12368 4168
rect 12402 4156 12408 4190
rect 12347 4155 12408 4156
rect 12399 4115 12408 4155
rect 12347 4090 12368 4103
rect 12402 4081 12408 4115
rect 12399 4040 12408 4081
rect 12347 4025 12368 4038
rect 12402 4006 12408 4040
rect 12399 3973 12408 4006
rect 12347 3965 12408 3973
rect 12347 3959 12368 3965
rect 12402 3931 12408 3965
rect 12399 3907 12408 3931
rect 12347 3893 12408 3907
rect 12399 3890 12408 3893
rect 12402 3856 12408 3890
rect 12399 3841 12408 3856
rect 12347 3827 12408 3841
rect 12399 3815 12408 3827
rect 12402 3781 12408 3815
rect 12399 3775 12408 3781
rect 12347 3769 12408 3775
rect 7829 3761 7884 3763
rect 7766 3759 7884 3761
tri 7884 3759 7888 3763 sw
rect 10595 3759 10992 3765
rect 7766 3735 7888 3759
tri 7888 3735 7912 3759 sw
rect 7766 3723 9371 3735
rect 7766 3689 7795 3723
rect 7829 3689 9371 3723
rect 7766 3683 9371 3689
rect 9423 3683 9435 3735
rect 9487 3683 9493 3735
rect 9587 3683 9593 3735
rect 9645 3683 9659 3735
rect 9711 3683 9717 3735
rect 10504 3723 10797 3729
rect 10504 3689 10516 3723
rect 10550 3689 10588 3723
rect 10622 3689 10679 3723
rect 10713 3689 10751 3723
rect 10785 3689 10797 3723
tri 12928 3710 12931 3713 se
rect 12931 3710 12965 3713
rect 10504 3683 10797 3689
tri 12901 3683 12928 3710 se
rect 12928 3683 12965 3710
rect -411 3656 -354 3668
rect -463 3642 -354 3656
tri -301 3655 -276 3680 se
rect -276 3655 -253 3680
tri -253 3655 -228 3680 nw
tri 386 3679 387 3680 se
rect 387 3679 825 3680
tri 12897 3679 12901 3683 se
rect 12901 3679 12965 3683
tri 362 3655 386 3679 se
rect 386 3655 428 3679
tri 428 3655 452 3679 nw
tri 12873 3655 12897 3679 se
rect 12897 3655 12965 3679
rect 13337 3704 13683 3710
tri -313 3643 -301 3655 se
rect -301 3643 -265 3655
tri -265 3643 -253 3655 nw
tri 356 3649 362 3655 se
rect 362 3651 424 3655
tri 424 3651 428 3655 nw
rect 938 3654 13026 3655
rect 362 3649 422 3651
tri 422 3649 424 3651 nw
tri 462 3649 464 3651 se
rect 464 3649 805 3651
rect 139 3643 191 3649
tri 191 3643 197 3649 sw
tri 350 3643 356 3649 se
rect 356 3643 416 3649
tri 416 3643 422 3649 nw
tri 456 3643 462 3649 se
rect 462 3643 805 3649
tri 805 3643 813 3651 sw
rect -411 3630 -354 3642
rect -411 3596 -394 3630
rect -360 3596 -354 3630
rect -411 3590 -354 3596
rect -463 3584 -354 3590
tri -324 3632 -313 3643 se
rect -313 3634 -274 3643
tri -274 3634 -265 3643 nw
rect -313 3632 -276 3634
tri -276 3632 -274 3634 nw
rect -324 3622 -286 3632
tri -286 3622 -276 3632 nw
rect -113 3622 -51 3634
tri -328 3535 -324 3539 se
rect -324 3535 -290 3622
tri -290 3618 -286 3622 nw
tri -339 3524 -328 3535 se
rect -328 3524 -290 3535
tri -347 3516 -339 3524 se
rect -339 3516 -298 3524
tri -298 3516 -290 3524 nw
rect -113 3570 -103 3622
rect -113 3558 -51 3570
tri -364 3499 -347 3516 se
rect -347 3499 -315 3516
tri -315 3499 -298 3516 nw
rect -113 3506 -103 3558
rect 191 3634 197 3643
tri 197 3634 206 3643 sw
tri 341 3634 350 3643 se
rect 350 3639 412 3643
tri 412 3639 416 3643 nw
tri 452 3639 456 3643 se
rect 456 3639 813 3643
rect 350 3634 407 3639
tri 407 3634 412 3639 nw
tri 447 3634 452 3639 se
rect 452 3634 813 3639
rect 191 3629 206 3634
tri 206 3629 211 3634 sw
tri 336 3629 341 3634 se
rect 341 3629 402 3634
tri 402 3629 407 3634 nw
tri 442 3629 447 3634 se
rect 447 3629 813 3634
rect 191 3613 386 3629
tri 386 3613 402 3629 nw
tri 426 3613 442 3629 se
rect 442 3613 813 3629
rect 191 3609 382 3613
tri 382 3609 386 3613 nw
tri 422 3609 426 3613 se
rect 426 3609 813 3613
tri 813 3609 847 3643 sw
rect 191 3605 378 3609
tri 378 3605 382 3609 nw
tri 418 3605 422 3609 se
rect 422 3605 847 3609
tri 847 3605 851 3609 sw
rect 191 3591 356 3605
rect 139 3583 356 3591
tri 356 3583 378 3605 nw
tri 396 3583 418 3605 se
rect 418 3583 462 3605
tri 462 3583 484 3605 nw
tri 785 3583 807 3605 ne
rect 807 3593 851 3605
tri 851 3593 863 3605 sw
rect 807 3583 863 3593
rect 139 3579 227 3583
rect 191 3571 227 3579
tri 227 3571 239 3583 nw
tri 384 3571 396 3583 se
rect 396 3573 452 3583
tri 452 3573 462 3583 nw
tri 807 3573 817 3583 ne
rect 396 3571 450 3573
tri 450 3571 452 3573 nw
rect 191 3537 193 3571
tri 193 3537 227 3571 nw
tri 352 3539 384 3571 se
rect 384 3569 448 3571
tri 448 3569 450 3571 nw
rect 384 3539 418 3569
tri 418 3539 448 3569 nw
tri 465 3539 495 3569 se
rect 495 3539 657 3569
tri 350 3537 352 3539 se
rect 352 3537 416 3539
tri 416 3537 418 3539 nw
tri 463 3537 465 3539 se
rect 465 3537 657 3539
tri 657 3537 689 3569 sw
tri 191 3535 193 3537 nw
tri 348 3535 350 3537 se
rect 350 3535 414 3537
tri 414 3535 416 3537 nw
tri 461 3535 463 3537 se
rect 463 3535 689 3537
tri 343 3530 348 3535 se
rect 348 3530 402 3535
rect 139 3521 191 3527
tri 334 3521 343 3530 se
rect 343 3523 402 3530
tri 402 3523 414 3535 nw
tri 449 3523 461 3535 se
rect 461 3523 689 3535
tri 689 3523 703 3537 sw
rect 343 3521 383 3523
tri 333 3520 334 3521 se
rect 334 3520 383 3521
rect -113 3504 -51 3506
tri -51 3504 -35 3520 sw
tri 317 3504 333 3520 se
rect 333 3504 383 3520
tri 383 3504 402 3523 nw
tri 430 3504 449 3523 se
rect 449 3504 496 3523
tri 496 3504 515 3523 nw
tri 631 3504 650 3523 ne
rect 650 3522 703 3523
tri 703 3522 704 3523 sw
rect 650 3504 704 3522
rect -113 3499 -35 3504
tri -35 3499 -30 3504 sw
tri 312 3499 317 3504 se
rect 317 3499 378 3504
tri 378 3499 383 3504 nw
tri 425 3499 430 3504 se
rect 430 3499 491 3504
tri 491 3499 496 3504 nw
tri 650 3499 655 3504 ne
rect 655 3499 704 3504
tri -388 3475 -364 3499 se
rect -364 3475 -339 3499
tri -339 3475 -315 3499 nw
rect -113 3491 -30 3499
tri -30 3491 -22 3499 sw
tri 304 3491 312 3499 se
rect 312 3491 354 3499
rect -113 3475 354 3491
tri 354 3475 378 3499 nw
tri 401 3475 425 3499 se
rect 425 3496 488 3499
tri 488 3496 491 3499 nw
tri 655 3496 658 3499 ne
rect 425 3475 467 3496
tri 467 3475 488 3496 nw
tri -398 3465 -388 3475 se
rect -388 3465 -349 3475
tri -349 3465 -339 3475 nw
rect -113 3473 352 3475
tri 352 3473 354 3475 nw
tri 399 3473 401 3475 se
rect 401 3473 465 3475
tri 465 3473 467 3475 nw
rect -113 3465 344 3473
tri 344 3465 352 3473 nw
tri 391 3465 399 3473 se
rect 399 3465 457 3473
tri 457 3465 465 3473 nw
tri -410 3453 -398 3465 se
rect -398 3453 -361 3465
tri -361 3453 -349 3465 nw
rect -113 3457 336 3465
tri 336 3457 344 3465 nw
tri 383 3457 391 3465 se
rect 391 3457 449 3465
tri 449 3457 457 3465 nw
rect -113 3454 333 3457
tri 333 3454 336 3457 nw
tri 380 3454 383 3457 se
rect 383 3454 445 3457
rect -113 3453 332 3454
tri 332 3453 333 3454 nw
tri 379 3453 380 3454 se
rect 380 3453 445 3454
tri 445 3453 449 3457 nw
tri -413 3450 -410 3453 se
rect -410 3450 -388 3453
rect -465 3444 -388 3450
rect -413 3426 -388 3444
tri -388 3426 -361 3453 nw
rect -113 3445 324 3453
tri 324 3445 332 3453 nw
tri 371 3445 379 3453 se
rect 379 3445 437 3453
tri 437 3445 445 3453 nw
tri 352 3426 371 3445 se
rect 371 3426 418 3445
tri 418 3426 437 3445 nw
rect -413 3419 -395 3426
tri -395 3419 -388 3426 nw
tri 345 3419 352 3426 se
rect 352 3419 411 3426
tri 411 3419 418 3426 nw
rect -413 3407 -407 3419
tri -407 3407 -395 3419 nw
tri 333 3407 345 3419 se
rect 345 3407 399 3419
tri 399 3407 411 3419 nw
rect -413 3402 -412 3407
tri -412 3402 -407 3407 nw
rect 121 3402 394 3407
tri 394 3402 399 3407 nw
tri -413 3401 -412 3402 nw
rect 121 3401 383 3402
rect -465 3380 -413 3392
rect -465 3322 -413 3328
rect 173 3391 383 3401
tri 383 3391 394 3402 nw
rect 173 3385 377 3391
tri 377 3385 383 3391 nw
rect 173 3379 371 3385
tri 371 3379 377 3385 nw
rect 173 3361 353 3379
tri 353 3361 371 3379 nw
rect 173 3356 225 3361
tri 225 3356 230 3361 nw
rect 173 3349 210 3356
rect 121 3341 210 3349
tri 210 3341 225 3356 nw
rect 121 3335 180 3341
rect 173 3311 180 3335
tri 180 3311 210 3341 nw
rect 173 3310 179 3311
tri 179 3310 180 3311 nw
rect 658 3310 704 3499
rect 817 3310 863 3583
rect 938 3602 947 3654
rect 999 3602 1013 3654
rect 1065 3602 1079 3654
rect 1131 3602 1145 3654
rect 1197 3602 1211 3654
rect 1263 3643 1277 3654
rect 1263 3609 1270 3643
rect 1263 3602 1277 3609
rect 1329 3602 1343 3654
rect 1395 3602 1408 3654
rect 1460 3602 1473 3654
rect 1525 3649 13026 3654
rect 1525 3643 8923 3649
rect 1525 3602 2882 3643
rect 938 3580 2882 3602
rect 938 3528 947 3580
rect 999 3528 1013 3580
rect 1065 3528 1079 3580
rect 1131 3528 1145 3580
rect 1197 3528 1211 3580
rect 1263 3571 1277 3580
rect 1263 3537 1270 3571
rect 1263 3528 1277 3537
rect 1329 3528 1343 3580
rect 1395 3528 1408 3580
rect 1460 3528 1473 3580
rect 1525 3528 2882 3580
rect 938 3506 2882 3528
rect 938 3454 947 3506
rect 999 3454 1013 3506
rect 1065 3454 1079 3506
rect 1131 3454 1145 3506
rect 1197 3454 1211 3506
rect 1263 3499 1277 3506
rect 1263 3465 1270 3499
rect 1263 3454 1277 3465
rect 1329 3454 1343 3506
rect 1395 3454 1408 3506
rect 1460 3454 1473 3506
rect 1525 3465 2882 3506
rect 3060 3465 3270 3643
rect 3376 3609 3604 3643
rect 3638 3609 3916 3643
rect 3950 3609 4181 3643
rect 3376 3571 4181 3609
rect 3376 3537 3604 3571
rect 3638 3537 3916 3571
rect 3950 3537 4181 3571
rect 3376 3499 4181 3537
rect 3376 3465 3604 3499
rect 3638 3465 3916 3499
rect 3950 3465 4181 3499
rect 4359 3465 5770 3643
rect 5948 3609 6180 3643
rect 6214 3609 6492 3643
rect 6526 3609 6804 3643
rect 6838 3609 7116 3643
rect 7150 3609 7340 3643
rect 5948 3571 7340 3609
rect 5948 3537 6180 3571
rect 6214 3537 6492 3571
rect 6526 3537 6804 3571
rect 6838 3537 7116 3571
rect 7150 3537 7340 3571
rect 5948 3499 7340 3537
rect 5948 3465 6180 3499
rect 6214 3465 6492 3499
rect 6526 3465 6804 3499
rect 6838 3465 7116 3499
rect 7150 3465 7340 3499
rect 7518 3609 7790 3643
rect 7824 3609 8022 3643
rect 7518 3571 8022 3609
rect 7518 3537 7790 3571
rect 7824 3537 8022 3571
rect 7518 3499 8022 3537
rect 7518 3465 7790 3499
rect 7824 3465 8022 3499
rect 8200 3597 8923 3643
rect 8975 3597 9027 3649
rect 9079 3643 12347 3649
rect 12399 3643 13026 3649
rect 9079 3609 10483 3643
rect 10517 3641 12347 3643
rect 10517 3609 11937 3641
rect 9079 3607 11937 3609
rect 11971 3607 12011 3641
rect 12045 3607 12084 3641
rect 12118 3607 12157 3641
rect 12191 3607 12347 3641
rect 12400 3609 13026 3643
rect 9079 3597 12347 3607
rect 12399 3597 13026 3609
rect 8200 3580 13026 3597
rect 8200 3528 8923 3580
rect 8975 3528 9027 3580
rect 9079 3571 12347 3580
rect 12399 3571 13026 3580
rect 9079 3537 9640 3571
rect 9674 3537 10136 3571
rect 10170 3537 10483 3571
rect 10517 3537 12347 3571
rect 12400 3566 13026 3571
rect 13337 3652 13338 3704
rect 13390 3652 13411 3704
rect 13463 3652 13484 3704
rect 13536 3652 13557 3704
rect 13609 3652 13630 3704
rect 13682 3652 13683 3704
rect 13337 3638 13683 3652
rect 13337 3586 13338 3638
rect 13390 3586 13411 3638
rect 13463 3586 13484 3638
rect 13536 3586 13557 3638
rect 13609 3586 13630 3638
rect 13682 3586 13683 3638
rect 13337 3572 13683 3586
rect 12400 3560 13216 3566
rect 12400 3537 12887 3560
rect 9079 3528 12347 3537
rect 12399 3528 12887 3537
rect 8200 3518 12887 3528
rect 8200 3511 9443 3518
rect 8200 3465 8923 3511
rect 1525 3459 8923 3465
rect 8975 3459 9027 3511
rect 9079 3484 9443 3511
rect 9477 3484 9515 3518
rect 9549 3511 12887 3518
rect 9549 3499 12347 3511
rect 12399 3508 12887 3511
rect 12939 3508 12956 3560
rect 13008 3508 13025 3560
rect 13077 3508 13094 3560
rect 13146 3508 13163 3560
rect 13215 3508 13216 3560
rect 12399 3499 13216 3508
rect 9549 3484 9640 3499
rect 9079 3465 9640 3484
rect 9674 3465 10136 3499
rect 10170 3465 10483 3499
rect 10517 3465 12347 3499
rect 12400 3490 13216 3499
rect 12400 3465 12887 3490
rect 9079 3459 12347 3465
rect 12399 3459 12887 3465
rect 1525 3454 12887 3459
rect 938 3453 12887 3454
tri 12547 3425 12575 3453 ne
rect 12575 3425 12749 3453
rect 1053 3419 8422 3425
rect 1053 3385 1114 3419
rect 1148 3385 1186 3419
rect 1220 3385 4542 3419
rect 4576 3385 4614 3419
rect 4648 3385 4854 3419
rect 4888 3385 4926 3419
rect 4960 3385 5166 3419
rect 5200 3385 5238 3419
rect 5272 3385 5478 3419
rect 5512 3385 5550 3419
rect 5584 3413 8422 3419
rect 5584 3385 7272 3413
rect 1053 3379 7272 3385
rect 7306 3379 8422 3413
rect 1053 3373 8422 3379
rect 8474 3373 8486 3425
rect 8538 3373 9582 3425
rect 9634 3373 9646 3425
rect 9698 3379 9704 3425
tri 11111 3424 11112 3425 se
rect 11112 3424 12101 3425
tri 11108 3421 11111 3424 se
rect 11111 3421 12101 3424
tri 9704 3379 9722 3397 sw
rect 9698 3378 9722 3379
tri 9722 3378 9723 3379 sw
rect 9698 3373 9723 3378
tri 7241 3356 7258 3373 ne
rect 7258 3356 7320 3373
tri 7320 3356 7337 3373 nw
tri 7989 3356 8006 3373 ne
rect 8006 3356 8152 3373
tri 8152 3356 8169 3373 nw
tri 9662 3356 9679 3373 ne
rect 9679 3356 9723 3373
tri 9723 3356 9745 3378 sw
rect 9812 3369 9818 3421
rect 9870 3369 9882 3421
rect 9934 3413 10976 3421
tri 11106 3419 11108 3421 se
rect 11108 3419 12101 3421
rect 9934 3379 10858 3413
rect 10892 3379 10930 3413
rect 10964 3379 10976 3413
tri 11089 3402 11106 3419 se
rect 11106 3402 11983 3419
tri 11072 3385 11089 3402 se
rect 11089 3385 11983 3402
rect 12017 3385 12055 3419
rect 12089 3385 12101 3419
tri 12575 3404 12596 3425 ne
rect 12596 3404 12749 3425
tri 12231 3402 12233 3404 se
rect 12233 3402 12285 3404
tri 12596 3402 12598 3404 ne
rect 12598 3402 12749 3404
tri 12219 3390 12231 3402 se
rect 12231 3398 12285 3402
rect 12231 3390 12233 3398
rect 9934 3369 10976 3379
tri 11056 3369 11072 3385 se
rect 11072 3379 12101 3385
tri 12208 3379 12219 3390 se
rect 12219 3379 12233 3390
rect 11072 3369 11112 3379
tri 11046 3359 11056 3369 se
rect 11056 3359 11112 3369
tri 11112 3359 11132 3379 nw
tri 12188 3359 12208 3379 se
rect 12208 3359 12233 3379
tri 11043 3356 11046 3359 se
rect 11046 3356 11109 3359
tri 11109 3356 11112 3359 nw
tri 12185 3356 12188 3359 se
rect 12188 3356 12233 3359
tri 7258 3348 7266 3356 ne
rect 7266 3341 7312 3356
tri 7312 3348 7320 3356 nw
tri 8006 3348 8014 3356 ne
rect 8014 3352 8148 3356
tri 8148 3352 8152 3356 nw
tri 9679 3352 9683 3356 ne
rect 9683 3352 9745 3356
tri 9745 3352 9749 3356 sw
tri 11039 3352 11043 3356 se
rect 11043 3352 11085 3356
rect 8014 3348 8144 3352
tri 8144 3348 8148 3352 nw
tri 9683 3348 9687 3352 ne
rect 9687 3348 9749 3352
tri 9687 3347 9688 3348 ne
rect 9688 3347 9749 3348
rect 8015 3346 8143 3347
tri 9688 3346 9689 3347 ne
rect 9689 3346 9749 3347
rect 173 3307 176 3310
tri 176 3307 179 3310 nw
rect 7266 3307 7272 3341
rect 7306 3307 7312 3341
rect 173 3305 174 3307
tri 174 3305 176 3307 nw
tri 173 3304 174 3305 nw
rect 7266 3295 7312 3307
rect 7612 3339 7742 3345
rect 7612 3305 7624 3339
rect 7658 3305 7696 3339
rect 7730 3305 7742 3339
rect 7612 3299 7742 3305
rect 8014 3310 8144 3346
tri 9689 3344 9691 3346 ne
rect 9691 3344 9749 3346
tri 8279 3326 8284 3331 se
rect 8284 3326 8775 3331
tri 8775 3326 8780 3331 sw
tri 8264 3311 8279 3326 se
rect 8279 3311 8780 3326
tri 8780 3311 8795 3326 sw
tri 8263 3310 8264 3311 se
rect 8264 3310 8795 3311
rect 8015 3309 8143 3310
tri 8262 3309 8263 3310 se
rect 8263 3309 8795 3310
tri 8261 3308 8262 3309 se
rect 8262 3308 8795 3309
rect 8014 3302 8144 3308
rect 121 3277 173 3283
rect 2367 3240 2373 3292
rect 2425 3240 2437 3292
rect 2489 3240 7005 3292
rect 7057 3240 7069 3292
rect 7121 3240 7127 3292
rect 8014 3268 8026 3302
rect 8060 3268 8098 3302
rect 8132 3268 8144 3302
tri 8245 3292 8261 3308 se
rect 8261 3292 8795 3308
tri 8795 3292 8814 3311 sw
rect 8983 3292 8989 3344
rect 9041 3292 9053 3344
rect 9105 3331 9542 3344
tri 9542 3331 9555 3344 sw
tri 9691 3331 9704 3344 ne
rect 9704 3332 9749 3344
tri 9749 3332 9769 3352 sw
tri 11019 3332 11039 3352 se
rect 11039 3332 11085 3352
tri 11085 3332 11109 3356 nw
tri 12161 3332 12185 3356 se
rect 12185 3346 12233 3356
rect 12185 3334 12285 3346
rect 12185 3332 12233 3334
rect 9704 3331 11071 3332
rect 9105 3326 9555 3331
tri 9555 3326 9560 3331 sw
tri 9704 3326 9709 3331 ne
rect 9709 3326 11071 3331
rect 9105 3311 9560 3326
tri 9560 3311 9575 3326 sw
tri 9709 3311 9724 3326 ne
rect 9724 3311 10680 3326
rect 9105 3292 9575 3311
tri 9575 3292 9594 3311 sw
tri 9724 3292 9743 3311 ne
rect 9743 3292 10680 3311
rect 10714 3292 10752 3326
rect 10786 3318 11071 3326
tri 11071 3318 11085 3332 nw
tri 12151 3322 12161 3332 se
rect 12161 3322 12233 3332
rect 10786 3316 11069 3318
tri 11069 3316 11071 3318 nw
rect 11137 3316 12233 3322
rect 10786 3311 11064 3316
tri 11064 3311 11069 3316 nw
rect 10786 3292 11039 3311
tri 8235 3282 8245 3292 se
rect 8245 3282 8814 3292
tri 8814 3282 8824 3292 sw
tri 9540 3282 9550 3292 ne
rect 9550 3282 9594 3292
tri 9594 3282 9604 3292 sw
tri 9743 3286 9749 3292 ne
rect 9749 3286 11039 3292
tri 11039 3286 11064 3311 nw
rect 11137 3282 11149 3316
rect 11183 3282 11221 3316
rect 11255 3282 12233 3316
tri 8232 3279 8235 3282 se
rect 8235 3279 8824 3282
tri 8824 3279 8827 3282 sw
tri 9550 3279 9553 3282 ne
rect 9553 3279 9604 3282
rect 8014 3256 8144 3268
tri 8209 3256 8232 3279 se
rect 8232 3256 8273 3279
tri 8199 3246 8209 3256 se
rect 8209 3246 8273 3256
tri 8273 3246 8306 3279 nw
tri 8765 3251 8793 3279 ne
rect 8793 3251 8827 3279
tri 8198 3245 8199 3246 se
rect 8199 3245 8272 3246
tri 8272 3245 8273 3246 nw
rect 8330 3245 8460 3251
tri 8793 3246 8798 3251 ne
rect 8798 3246 8827 3251
tri 8827 3246 8860 3279 sw
tri 9553 3252 9580 3279 ne
rect 9580 3252 9604 3279
tri 9604 3252 9634 3282 sw
rect 11137 3276 12285 3282
rect 12347 3396 12406 3402
rect 12399 3390 12406 3396
rect 12400 3356 12406 3390
rect 12399 3344 12406 3356
rect 12347 3332 12406 3344
rect 12399 3318 12406 3332
rect 12400 3284 12406 3318
tri 12598 3311 12689 3402 ne
rect 12689 3355 12749 3402
rect 12689 3311 12743 3355
tri 12743 3349 12749 3355 ne
rect 12886 3438 12887 3453
rect 12939 3438 12956 3490
rect 13008 3438 13025 3490
rect 13077 3438 13094 3490
rect 13146 3438 13163 3490
rect 13215 3438 13216 3490
rect 12886 3420 13216 3438
rect 12886 3368 12887 3420
rect 12939 3368 12956 3420
rect 13008 3368 13025 3420
rect 13077 3368 13094 3420
rect 13146 3368 13163 3420
rect 13215 3368 13216 3420
rect 12886 3349 13216 3368
rect 12399 3280 12406 3284
rect 12347 3268 12406 3280
tri 9580 3246 9586 3252 ne
rect 9586 3246 9634 3252
tri 9634 3246 9640 3252 sw
tri 9884 3246 9890 3252 se
rect 9890 3246 9942 3252
tri 8193 3240 8198 3245 se
rect 8198 3240 8249 3245
tri 8188 3235 8193 3240 se
rect 8193 3235 8249 3240
rect -476 3228 410 3235
tri 410 3228 417 3235 sw
tri 8181 3228 8188 3235 se
rect 8188 3228 8249 3235
rect -476 3223 417 3228
rect -476 3189 -470 3223
rect -436 3220 417 3223
tri 417 3220 425 3228 sw
rect -436 3212 425 3220
tri 425 3212 433 3220 sw
rect -436 3211 433 3212
tri 433 3211 434 3212 sw
rect -436 3199 434 3211
tri 434 3199 446 3211 sw
rect -436 3191 -397 3199
tri -397 3191 -389 3199 nw
tri 396 3191 404 3199 ne
rect 404 3191 446 3199
tri 446 3191 454 3199 sw
rect -436 3189 -414 3191
rect -476 3174 -414 3189
tri -414 3174 -397 3191 nw
tri 404 3174 421 3191 ne
rect 421 3174 454 3191
tri 454 3174 471 3191 sw
rect -476 3163 -425 3174
tri -425 3163 -414 3174 nw
tri 421 3163 432 3174 ne
rect 432 3163 471 3174
tri 471 3163 482 3174 sw
rect -476 3160 -428 3163
tri -428 3160 -425 3163 nw
tri 432 3160 435 3163 ne
rect 435 3160 482 3163
tri 482 3160 485 3163 sw
rect 2114 3160 2120 3212
rect 2172 3160 2184 3212
rect 2236 3160 6985 3212
rect 7037 3160 7049 3212
rect 7101 3160 7107 3212
rect 7204 3176 7210 3228
rect 7262 3176 7274 3228
rect 7326 3222 8249 3228
tri 8249 3222 8272 3245 nw
rect 7326 3220 8247 3222
tri 8247 3220 8249 3222 nw
rect 7326 3211 8238 3220
tri 8238 3211 8247 3220 nw
rect 8330 3211 8342 3245
rect 8376 3211 8414 3245
rect 8448 3211 8460 3245
tri 8798 3225 8819 3246 ne
rect 8819 3225 8860 3246
tri 8860 3225 8881 3246 sw
tri 9586 3225 9607 3246 ne
rect 9607 3230 9640 3246
tri 9640 3230 9656 3246 sw
tri 9868 3230 9884 3246 se
rect 9884 3230 9890 3246
rect 9607 3225 9890 3230
tri 8819 3222 8822 3225 ne
rect 8822 3222 8881 3225
tri 8881 3222 8884 3225 sw
tri 9607 3222 9610 3225 ne
rect 9610 3222 9890 3225
tri 8822 3220 8824 3222 ne
rect 8824 3220 8884 3222
tri 8884 3220 8886 3222 sw
tri 9610 3220 9612 3222 ne
rect 9612 3220 9890 3222
rect 7326 3205 8232 3211
tri 8232 3205 8238 3211 nw
rect 7326 3191 8218 3205
tri 8218 3191 8232 3205 nw
rect 8330 3197 8460 3211
tri 8824 3197 8847 3220 ne
rect 8847 3212 8886 3220
tri 8886 3212 8894 3220 sw
tri 9612 3212 9620 3220 ne
rect 9620 3212 9890 3220
rect 8847 3197 9450 3212
tri 8847 3196 8848 3197 ne
rect 8848 3196 9450 3197
rect 8331 3195 8459 3196
tri 8848 3195 8849 3196 ne
rect 8849 3195 9450 3196
rect 7326 3176 8203 3191
tri 8203 3176 8218 3191 nw
rect -476 3151 -430 3160
tri -430 3158 -428 3160 nw
tri 435 3158 437 3160 ne
rect 437 3158 485 3160
rect -476 3117 -470 3151
rect -436 3117 -430 3151
tri 437 3149 446 3158 ne
rect 446 3149 485 3158
tri 485 3149 496 3160 sw
rect 8330 3159 8460 3195
tri 8849 3191 8853 3195 ne
rect 8853 3191 9450 3195
tri 9450 3191 9471 3212 sw
tri 9620 3192 9640 3212 ne
rect 9640 3194 9890 3212
rect 12399 3246 12406 3268
rect 9640 3192 9942 3194
tri 9852 3191 9853 3192 ne
rect 9853 3191 9942 3192
tri 8853 3174 8870 3191 ne
rect 8870 3174 9471 3191
tri 9471 3174 9488 3191 sw
tri 9853 3174 9870 3191 ne
rect 9870 3182 9942 3191
rect 10619 3185 10625 3237
rect 10677 3185 10689 3237
rect 10741 3185 11006 3237
rect 11058 3185 11070 3237
rect 11122 3233 11128 3237
tri 11128 3233 11132 3237 sw
rect 11122 3231 11132 3233
tri 11132 3231 11134 3233 sw
rect 11122 3225 12081 3231
rect 11138 3191 11180 3225
rect 11214 3191 11256 3225
rect 11290 3191 11331 3225
rect 11365 3191 11808 3225
rect 11842 3191 11884 3225
rect 11918 3191 11960 3225
rect 11994 3191 12035 3225
rect 12069 3191 12081 3225
rect 12235 3227 12287 3233
tri 12234 3212 12235 3213 se
rect 11122 3185 12081 3191
tri 12207 3185 12234 3212 se
rect 12234 3185 12235 3212
rect 9870 3174 9890 3182
tri 8870 3160 8884 3174 ne
rect 8884 3160 9488 3174
tri 9488 3160 9502 3174 sw
tri 9870 3160 9884 3174 ne
rect 9884 3160 9890 3174
tri 9439 3159 9440 3160 ne
rect 9440 3159 9502 3160
rect 8331 3158 8459 3159
tri 9440 3158 9441 3159 ne
rect 9441 3158 9502 3159
tri 9441 3157 9442 3158 ne
rect 9442 3157 9502 3158
tri 8322 3149 8330 3157 se
rect 8330 3149 8460 3157
tri 8460 3149 8468 3157 sw
tri 9442 3149 9450 3157 ne
rect 9450 3149 9502 3157
tri 9502 3149 9513 3160 sw
tri 9884 3154 9890 3160 ne
tri 446 3145 450 3149 ne
rect 450 3145 496 3149
tri 496 3145 500 3149 sw
tri 8318 3145 8322 3149 se
rect 8322 3145 8468 3149
tri 8468 3145 8472 3149 sw
tri 9450 3145 9454 3149 ne
rect 9454 3145 9513 3149
tri 9513 3145 9517 3149 sw
tri 450 3132 463 3145 ne
rect 463 3132 500 3145
rect -476 3105 -430 3117
rect -389 3126 298 3132
tri 463 3130 465 3132 ne
rect 465 3130 500 3132
tri 500 3130 515 3145 sw
tri 8311 3138 8318 3145 se
rect 8318 3138 8472 3145
tri 8472 3138 8479 3145 sw
tri 9454 3138 9461 3145 ne
rect 9461 3138 9517 3145
tri 465 3126 469 3130 ne
rect 469 3127 515 3130
tri 515 3127 518 3130 sw
rect 469 3126 518 3127
rect -389 3118 238 3126
rect -389 3084 -314 3118
rect -280 3117 238 3118
rect -280 3084 -190 3117
rect -389 3083 -190 3084
rect -156 3083 238 3117
rect -389 3074 238 3083
rect 290 3074 298 3126
tri 469 3118 477 3126 ne
rect 477 3118 518 3126
tri 477 3113 482 3118 ne
rect -389 3054 298 3074
rect -389 3046 238 3054
rect -389 3012 -314 3046
rect -280 3045 238 3046
rect -280 3012 -190 3045
rect -389 3011 -190 3012
rect -156 3011 238 3045
rect -389 3002 238 3011
rect 290 3002 298 3054
rect -389 2982 298 3002
rect -389 2974 238 2982
rect -389 2940 -314 2974
rect -280 2940 238 2974
rect -389 2930 238 2940
rect 290 2930 298 2982
rect -389 2909 298 2930
tri -395 2894 -389 2900 se
rect -389 2894 238 2909
tri -418 2871 -395 2894 se
rect -395 2871 238 2894
tri -452 2837 -418 2871 se
rect -418 2837 -50 2871
rect -16 2837 22 2871
rect 56 2857 238 2871
rect 290 2857 298 2909
rect 56 2837 298 2857
tri -475 2814 -452 2837 se
rect -452 2836 298 2837
rect -452 2814 238 2836
tri -477 2812 -475 2814 se
rect -475 2812 238 2814
tri -508 2781 -477 2812 se
rect -477 2784 238 2812
rect 290 2784 298 2836
rect -477 2781 298 2784
rect -508 2778 298 2781
tri 298 2778 301 2781 sw
rect 482 2778 518 3118
rect 1162 3126 7553 3132
rect 1162 3092 1175 3126
rect 1209 3092 1247 3126
rect 1281 3092 1319 3126
rect 1353 3092 1391 3126
rect 1425 3092 7435 3126
rect 7469 3092 7507 3126
rect 7541 3092 7553 3126
rect 1162 3086 7553 3092
rect 7750 3086 7758 3138
rect 7810 3086 7822 3138
rect 7874 3086 7880 3138
tri 8305 3132 8311 3138 se
rect 8311 3132 8479 3138
tri 8479 3132 8485 3138 sw
tri 8667 3132 8673 3138 se
rect 8673 3132 8679 3138
rect 7908 3126 8679 3132
rect 8731 3126 8743 3138
rect 8795 3132 8801 3138
tri 8801 3132 8807 3138 sw
tri 9461 3132 9467 3138 ne
rect 9467 3132 9517 3138
tri 9517 3132 9530 3145 sw
rect 8795 3126 9427 3132
tri 9467 3130 9469 3132 ne
rect 9469 3130 9847 3132
tri 9469 3126 9473 3130 ne
rect 9473 3126 9847 3130
rect 7908 3092 7920 3126
rect 7954 3092 7992 3126
rect 8026 3092 8639 3126
rect 8673 3092 8679 3126
rect 8817 3092 8855 3126
rect 8889 3092 8927 3126
rect 8961 3092 8999 3126
rect 9033 3092 9071 3126
rect 9105 3092 9143 3126
rect 9177 3092 9215 3126
rect 9249 3092 9287 3126
rect 9321 3092 9359 3126
rect 9393 3092 9427 3126
tri 9473 3118 9481 3126 ne
rect 9481 3118 9729 3126
tri 9481 3092 9507 3118 ne
rect 9507 3092 9729 3118
rect 9763 3092 9801 3126
rect 9835 3092 9847 3126
tri 12196 3174 12207 3185 se
rect 12207 3175 12235 3185
rect 12207 3174 12287 3175
tri 12173 3151 12196 3174 se
rect 12196 3163 12287 3174
rect 12196 3151 12235 3163
rect 9890 3124 9942 3130
rect 11481 3145 12235 3151
rect 11481 3111 11493 3145
rect 11527 3111 11565 3145
rect 11599 3111 12235 3145
rect 11481 3105 12287 3111
rect 12347 3212 12366 3216
rect 12400 3212 12406 3246
rect 12886 3297 12887 3349
rect 12939 3297 12956 3349
rect 13008 3297 13025 3349
rect 13077 3297 13094 3349
rect 13146 3297 13163 3349
rect 13215 3297 13216 3349
rect 12886 3278 13216 3297
rect 12886 3226 12887 3278
rect 12939 3226 12956 3278
rect 13008 3226 13025 3278
rect 13077 3226 13094 3278
rect 13146 3226 13163 3278
rect 13215 3226 13216 3278
rect 12886 3220 13216 3226
rect 13337 3520 13338 3572
rect 13390 3520 13411 3572
rect 13463 3520 13484 3572
rect 13536 3520 13557 3572
rect 13609 3520 13630 3572
rect 13682 3520 13683 3572
rect 13337 3506 13683 3520
rect 13337 3454 13338 3506
rect 13390 3454 13411 3506
rect 13463 3454 13484 3506
rect 13536 3454 13557 3506
rect 13609 3454 13630 3506
rect 13682 3454 13683 3506
rect 13337 3440 13683 3454
rect 13337 3388 13338 3440
rect 13390 3388 13411 3440
rect 13463 3388 13484 3440
rect 13536 3388 13557 3440
rect 13609 3388 13630 3440
rect 13682 3388 13683 3440
rect 13337 3374 13683 3388
rect 13337 3322 13338 3374
rect 13390 3322 13411 3374
rect 13463 3322 13484 3374
rect 13536 3322 13557 3374
rect 13609 3322 13630 3374
rect 13682 3322 13683 3374
rect 13337 3308 13683 3322
rect 13337 3256 13338 3308
rect 13390 3256 13411 3308
rect 13463 3256 13484 3308
rect 13536 3256 13557 3308
rect 13609 3256 13630 3308
rect 13682 3256 13683 3308
rect 13337 3242 13683 3256
rect 14697 3248 15008 3480
rect 12347 3204 12406 3212
rect 12399 3174 12406 3204
rect 12347 3140 12366 3152
rect 12400 3140 12406 3174
rect 7908 3086 8679 3092
rect 8731 3086 8743 3092
rect 8795 3086 9427 3092
tri 9507 3086 9513 3092 ne
rect 9513 3086 9847 3092
rect 12399 3102 12406 3140
rect 13337 3190 13338 3242
rect 13390 3190 13411 3242
rect 13463 3190 13484 3242
rect 13536 3190 13557 3242
rect 13609 3190 13630 3242
rect 13682 3190 13683 3242
rect 13337 3176 13683 3190
rect 13337 3124 13338 3176
rect 13390 3124 13411 3176
rect 13463 3124 13484 3176
rect 13536 3124 13557 3176
rect 13609 3124 13630 3176
rect 13682 3124 13683 3176
rect 13337 3118 13683 3124
rect 12347 3076 12366 3088
rect 12400 3068 12406 3102
rect 1220 3057 12204 3058
rect 1220 3005 1704 3057
rect 1756 3005 1773 3057
rect 1825 3005 1842 3057
rect 1894 3005 1911 3057
rect 1963 3005 1980 3057
rect 2032 3005 3156 3057
rect 3208 3005 3220 3057
rect 3272 3005 3284 3057
rect 3336 3005 3348 3057
rect 3400 3005 3412 3057
rect 3464 3005 3476 3057
rect 3528 3005 3540 3057
rect 3592 3046 12204 3057
rect 3592 3012 10744 3046
rect 10778 3012 10860 3046
rect 10894 3012 11212 3046
rect 11246 3012 11564 3046
rect 11598 3012 11916 3046
rect 11950 3012 12204 3046
rect 3592 3005 12204 3012
rect 1220 2981 12204 3005
rect 1220 2929 1704 2981
rect 1756 2977 1773 2981
rect 1825 2977 1842 2981
rect 1894 2977 1911 2981
rect 1963 2977 1980 2981
rect 2032 2977 3156 2981
rect 3208 2977 3220 2981
rect 3272 2977 3284 2981
rect 1894 2943 1895 2977
rect 1963 2943 1967 2977
rect 2032 2943 2039 2977
rect 2073 2943 2111 2977
rect 2145 2943 2183 2977
rect 2217 2943 2255 2977
rect 2289 2943 2327 2977
rect 2361 2943 2399 2977
rect 2433 2943 2471 2977
rect 2505 2943 2543 2977
rect 2577 2943 2615 2977
rect 2649 2943 2687 2977
rect 2721 2943 2759 2977
rect 2793 2943 2831 2977
rect 2865 2943 2903 2977
rect 2937 2943 2975 2977
rect 3009 2943 3047 2977
rect 3081 2943 3119 2977
rect 3153 2943 3156 2977
rect 1756 2929 1773 2943
rect 1825 2929 1842 2943
rect 1894 2929 1911 2943
rect 1963 2929 1980 2943
rect 2032 2929 3156 2943
rect 3208 2929 3220 2943
rect 3272 2929 3284 2943
rect 3336 2929 3348 2981
rect 3400 2929 3412 2981
rect 3464 2974 3476 2981
rect 3528 2974 3540 2981
rect 3592 2974 12204 2981
rect 3466 2940 3476 2974
rect 3614 2940 3654 2974
rect 3688 2940 3728 2974
rect 3762 2940 3802 2974
rect 3836 2940 3876 2974
rect 3910 2940 3950 2974
rect 3984 2940 4024 2974
rect 4058 2940 4098 2974
rect 4132 2940 4172 2974
rect 4206 2940 4246 2974
rect 4280 2940 4320 2974
rect 4354 2940 4394 2974
rect 4428 2940 4468 2974
rect 4502 2940 4541 2974
rect 4575 2940 4614 2974
rect 4648 2940 4687 2974
rect 4721 2940 4760 2974
rect 4794 2940 4833 2974
rect 4867 2940 4906 2974
rect 4940 2968 8422 2974
rect 4940 2940 7680 2968
rect 3464 2929 3476 2940
rect 3528 2929 3540 2940
rect 3592 2934 7680 2940
rect 7714 2934 7752 2968
rect 7786 2934 8070 2968
rect 8104 2934 8142 2968
rect 8176 2940 8422 2968
rect 8456 2940 8494 2974
rect 8528 2968 10744 2974
rect 8528 2940 8934 2968
rect 8176 2934 8934 2940
rect 8968 2934 9006 2968
rect 9040 2934 9362 2968
rect 9396 2934 9434 2968
rect 9468 2940 10744 2968
rect 10778 2940 10860 2974
rect 10894 2940 11212 2974
rect 11246 2940 11564 2974
rect 11598 2940 11916 2974
rect 11950 2940 12204 2974
rect 9468 2934 12204 2940
rect 3592 2929 12204 2934
rect 1220 2928 12204 2929
rect 12399 3030 12406 3068
rect 12347 3012 12366 3024
rect 12400 2996 12406 3030
rect 12399 2960 12406 2996
rect 12347 2958 12406 2960
rect 12347 2948 12366 2958
rect 12400 2924 12406 2958
tri 1324 2894 1328 2898 se
rect 1328 2894 2120 2898
tri 1290 2860 1324 2894 se
rect 1324 2860 2120 2894
tri 1286 2856 1290 2860 se
rect 1290 2856 2120 2860
tri 1282 2852 1286 2856 se
rect 1286 2852 2120 2856
tri 1278 2848 1282 2852 se
rect 1282 2848 2120 2852
tri 1276 2846 1278 2848 se
rect 1278 2846 2120 2848
rect 2172 2846 2184 2898
rect 2236 2846 2242 2898
rect 6979 2848 6985 2900
rect 7037 2848 7049 2900
rect 7101 2894 8231 2900
rect 7101 2848 7758 2894
tri 7723 2846 7725 2848 ne
rect 7725 2846 7758 2848
tri 1250 2820 1276 2846 se
rect 1276 2820 1324 2846
tri 1324 2820 1350 2846 nw
tri 7725 2820 7751 2846 ne
rect 7751 2842 7758 2846
rect 7810 2848 8231 2894
rect 8283 2848 8295 2900
rect 8347 2848 8353 2900
rect 8416 2848 8422 2900
rect 8474 2848 8486 2900
rect 8538 2894 9137 2900
rect 9139 2899 9175 2900
rect 8538 2860 8678 2894
rect 8712 2860 8750 2894
rect 8784 2860 9137 2894
rect 8538 2848 9137 2860
rect 9138 2849 9176 2899
rect 9177 2890 9310 2900
rect 9177 2856 9192 2890
rect 9226 2856 9264 2890
rect 9298 2856 9310 2890
rect 9139 2848 9175 2849
rect 9177 2848 9310 2856
rect 9668 2848 9674 2900
rect 9726 2848 9738 2900
rect 9790 2894 9942 2900
rect 9790 2860 9824 2894
rect 9858 2860 9896 2894
rect 9930 2860 9942 2894
rect 9790 2848 9942 2860
rect 9982 2848 9988 2900
rect 10040 2848 10052 2900
rect 10104 2848 10115 2900
rect 10167 2848 10173 2900
rect 10225 2848 10237 2900
rect 10289 2894 12125 2900
rect 10289 2854 12073 2894
rect 10289 2852 10299 2854
tri 10299 2852 10301 2854 nw
tri 12039 2852 12041 2854 ne
rect 12041 2852 12073 2854
rect 10289 2848 10295 2852
tri 10295 2848 10299 2852 nw
tri 12041 2848 12045 2852 ne
rect 12045 2848 12073 2852
rect 7810 2842 7817 2848
rect 7751 2830 7817 2842
rect 7751 2820 7758 2830
tri 1244 2814 1250 2820 se
rect 1250 2814 1318 2820
tri 1318 2814 1324 2820 nw
tri 7751 2814 7757 2820 ne
rect 7757 2814 7758 2820
tri 1242 2812 1244 2814 se
rect 1244 2812 1316 2814
tri 1316 2812 1318 2814 nw
tri 7757 2813 7758 2814 ne
tri 1238 2808 1242 2812 se
rect 1242 2808 1282 2812
tri 1210 2780 1238 2808 se
rect 1238 2780 1282 2808
tri 518 2778 520 2780 sw
tri 1208 2778 1210 2780 se
rect 1210 2778 1282 2780
tri 1282 2778 1316 2812 nw
rect 7810 2820 7817 2830
tri 7817 2820 7845 2848 nw
tri 12045 2820 12073 2848 ne
rect 12073 2830 12125 2842
rect 7810 2814 7811 2820
tri 7811 2814 7817 2820 nw
tri 8025 2814 8031 2820 se
rect 8031 2814 10509 2820
tri 7810 2813 7811 2814 nw
tri 8024 2813 8025 2814 se
rect 8025 2813 10509 2814
tri 8023 2812 8024 2813 se
rect 8024 2812 10509 2813
tri 7989 2778 8023 2812 se
rect 8023 2778 10311 2812
rect 10345 2778 10383 2812
rect 10417 2778 10509 2812
rect -508 2772 301 2778
tri 301 2772 307 2778 sw
rect 482 2777 520 2778
tri 520 2777 521 2778 sw
tri 1207 2777 1208 2778 se
rect 1208 2777 1281 2778
tri 1281 2777 1282 2778 nw
rect 482 2772 521 2777
tri 521 2772 526 2777 sw
tri 1202 2772 1207 2777 se
rect 1207 2772 1276 2777
tri 1276 2772 1281 2777 nw
rect 7758 2772 7810 2778
tri 7988 2777 7989 2778 se
rect 7989 2777 10509 2778
tri 7983 2772 7988 2777 se
rect 7988 2772 10509 2777
rect -508 2763 307 2772
rect -508 2711 238 2763
rect 290 2742 307 2763
tri 307 2742 337 2772 sw
rect 482 2766 526 2772
tri 526 2766 532 2772 sw
tri 1196 2766 1202 2772 se
rect 1202 2770 1274 2772
tri 1274 2770 1276 2772 nw
tri 7981 2770 7983 2772 se
rect 7983 2770 10509 2772
rect 1202 2766 1246 2770
tri 482 2742 506 2766 ne
rect 506 2742 532 2766
tri 532 2742 556 2766 sw
tri 1192 2762 1196 2766 se
rect 1196 2762 1246 2766
rect 1192 2742 1246 2762
tri 1246 2742 1274 2770 nw
tri 4239 2742 4267 2770 se
rect 4267 2742 4504 2770
rect 290 2728 337 2742
tri 337 2728 351 2742 sw
tri 506 2741 507 2742 ne
rect 507 2741 556 2742
tri 556 2741 557 2742 sw
tri 507 2728 520 2741 ne
rect 520 2728 557 2741
tri 557 2728 570 2741 sw
rect 290 2722 351 2728
tri 351 2722 357 2728 sw
tri 520 2722 526 2728 ne
rect 526 2722 570 2728
tri 570 2722 576 2728 sw
rect 290 2713 357 2722
tri 357 2713 366 2722 sw
tri 526 2713 535 2722 ne
rect 535 2713 576 2722
tri 576 2713 585 2722 sw
rect 290 2711 366 2713
rect -508 2697 366 2711
rect -508 2663 -277 2697
rect -243 2663 75 2697
rect 109 2696 366 2697
tri 366 2696 383 2713 sw
tri 535 2696 552 2713 ne
rect 552 2696 585 2713
tri 585 2696 602 2713 sw
rect 109 2690 383 2696
rect 109 2663 238 2690
rect -508 2638 238 2663
rect 290 2679 383 2690
tri 383 2679 400 2696 sw
tri 552 2694 554 2696 ne
rect 554 2694 602 2696
tri 602 2694 604 2696 sw
rect 1192 2694 1238 2742
tri 1238 2734 1246 2742 nw
tri 4231 2734 4239 2742 se
rect 4239 2734 4504 2742
tri 4225 2728 4231 2734 se
rect 4231 2728 4504 2734
tri 4219 2722 4225 2728 se
rect 4225 2722 4504 2728
tri 4215 2718 4219 2722 se
rect 4219 2718 4504 2722
rect 4556 2718 4568 2770
rect 4620 2718 4626 2770
tri 7979 2768 7981 2770 se
rect 7981 2768 10509 2770
rect 10510 2769 10511 2819
rect 10547 2769 10548 2819
rect 10549 2768 10829 2820
rect 12073 2772 12125 2778
rect 12399 2896 12406 2924
rect 12347 2886 12406 2896
rect 12347 2884 12366 2886
rect 12400 2852 12406 2886
rect 12399 2832 12406 2852
rect 12347 2819 12406 2832
rect 12399 2814 12406 2819
rect 12400 2780 12406 2814
tri 7953 2742 7979 2768 se
rect 7979 2743 8028 2768
tri 8028 2743 8053 2768 nw
tri 10352 2743 10377 2768 ne
rect 10377 2743 10429 2768
tri 10429 2743 10454 2768 nw
tri 10752 2743 10777 2768 ne
rect 7979 2742 8027 2743
tri 8027 2742 8028 2743 nw
tri 7939 2728 7953 2742 se
rect 7953 2728 8013 2742
tri 8013 2728 8027 2742 nw
rect 10378 2741 10428 2742
rect 8842 2728 9282 2738
tri 7936 2725 7939 2728 se
rect 7939 2725 8007 2728
tri 4210 2713 4215 2718 se
rect 4215 2713 4284 2718
tri 4284 2713 4289 2718 nw
tri 4193 2696 4210 2713 se
rect 4210 2696 4267 2713
tri 4267 2696 4284 2713 nw
tri 4191 2694 4193 2696 se
rect 4193 2694 4250 2696
tri 554 2691 557 2694 ne
rect 557 2691 604 2694
tri 604 2691 607 2694 sw
tri 4188 2691 4191 2694 se
rect 4191 2691 4250 2694
tri 557 2679 569 2691 ne
rect 569 2679 607 2691
tri 607 2679 619 2691 sw
tri 4176 2679 4188 2691 se
rect 4188 2679 4250 2691
tri 4250 2679 4267 2696 nw
rect 290 2676 400 2679
tri 400 2676 403 2679 sw
tri 569 2676 572 2679 ne
rect 572 2676 619 2679
tri 619 2676 622 2679 sw
tri 4173 2676 4176 2679 se
rect 4176 2676 4247 2679
tri 4247 2676 4250 2679 nw
rect 290 2652 403 2676
tri 403 2652 427 2676 sw
tri 572 2652 596 2676 ne
rect 596 2652 622 2676
tri 622 2652 646 2676 sw
tri 4149 2652 4173 2676 se
rect 4173 2673 4244 2676
tri 4244 2673 4247 2676 nw
rect 7672 2673 7678 2725
rect 7730 2673 7742 2725
rect 7794 2722 8007 2725
tri 8007 2722 8013 2728 nw
rect 8110 2722 8240 2728
rect 7794 2713 7988 2722
rect 7794 2679 7828 2713
rect 7862 2703 7988 2713
tri 7988 2703 8007 2722 nw
rect 7862 2696 7981 2703
tri 7981 2696 7988 2703 nw
rect 7862 2694 7979 2696
tri 7979 2694 7981 2696 nw
rect 7862 2688 7973 2694
tri 7973 2688 7979 2694 nw
rect 8110 2688 8122 2722
rect 8156 2688 8194 2722
rect 8228 2688 8240 2722
rect 7862 2679 7963 2688
rect 7794 2678 7963 2679
tri 7963 2678 7973 2688 nw
rect 7794 2676 7961 2678
tri 7961 2676 7963 2678 nw
rect 7794 2673 7958 2676
tri 7958 2673 7961 2676 nw
rect 4173 2652 4223 2673
tri 4223 2652 4244 2673 nw
tri 8092 2652 8110 2670 se
rect 8110 2652 8240 2688
rect 290 2638 427 2652
rect -508 2625 427 2638
rect -508 2591 -277 2625
rect -243 2591 75 2625
rect 109 2619 427 2625
tri 427 2619 460 2652 sw
tri 596 2651 597 2652 ne
rect 597 2651 646 2652
tri 646 2651 647 2652 sw
tri 4148 2651 4149 2652 se
rect 4149 2651 4216 2652
tri 597 2644 604 2651 ne
rect 604 2644 647 2651
tri 647 2644 654 2651 sw
tri 4141 2644 4148 2651 se
rect 4148 2645 4216 2651
tri 4216 2645 4223 2652 nw
tri 8085 2645 8092 2652 se
rect 8092 2645 8240 2652
rect 4148 2644 4215 2645
tri 4215 2644 4216 2645 nw
tri 604 2641 607 2644 ne
rect 607 2641 654 2644
tri 654 2641 657 2644 sw
tri 4138 2641 4141 2644 se
rect 4141 2641 4189 2644
tri 607 2629 619 2641 ne
rect 619 2629 657 2641
tri 657 2629 669 2641 sw
tri 4126 2629 4138 2641 se
rect 4138 2629 4189 2641
rect 109 2617 460 2619
tri 619 2618 630 2629 ne
rect 630 2618 669 2629
tri 669 2618 680 2629 sw
rect 109 2591 238 2617
rect -508 2578 238 2591
tri 215 2560 233 2578 ne
rect 233 2565 238 2578
rect 290 2565 460 2617
tri 630 2591 657 2618 ne
rect 657 2591 680 2618
tri 680 2591 707 2618 sw
tri 657 2578 670 2591 ne
rect 670 2578 707 2591
tri 670 2577 671 2578 ne
rect 671 2577 707 2578
tri 707 2577 721 2591 sw
rect 2889 2577 2895 2629
rect 2947 2577 2959 2629
rect 3011 2618 4189 2629
tri 4189 2618 4215 2644 nw
rect 3011 2593 4164 2618
tri 4164 2593 4189 2618 nw
rect 7508 2593 7659 2645
rect 7711 2593 7723 2645
rect 7775 2593 8240 2645
rect 8268 2710 8398 2716
rect 8268 2676 8280 2710
rect 8314 2676 8352 2710
rect 8386 2676 8398 2710
rect 8842 2694 8854 2728
rect 8888 2694 8926 2728
rect 8960 2694 9282 2728
rect 3011 2577 4148 2593
tri 4148 2577 4164 2593 nw
rect 233 2560 460 2565
tri 671 2560 688 2577 ne
rect 688 2560 721 2577
tri 721 2560 738 2577 sw
tri 233 2559 234 2560 ne
rect 234 2559 460 2560
tri 234 2536 257 2559 ne
rect 257 2536 460 2559
tri 688 2545 703 2560 ne
rect 703 2545 738 2560
tri 738 2545 753 2560 sw
tri 703 2541 707 2545 ne
rect 707 2541 753 2545
tri 753 2541 757 2545 sw
tri 707 2536 712 2541 ne
rect 712 2536 757 2541
rect -187 2533 54 2536
tri 54 2533 57 2536 sw
tri 257 2533 260 2536 ne
rect 260 2533 460 2536
tri 712 2533 715 2536 ne
rect 715 2533 757 2536
rect -465 2527 -413 2533
rect -465 2461 -413 2475
rect -465 2403 -413 2409
rect -187 2531 57 2533
tri 57 2531 59 2533 sw
tri 260 2531 262 2533 ne
rect -187 2530 59 2531
rect -135 2526 59 2530
tri 59 2526 64 2531 sw
rect -135 2510 64 2526
tri 64 2510 80 2526 sw
rect -135 2491 80 2510
tri 80 2491 99 2510 sw
rect -135 2478 -120 2491
rect -187 2476 -120 2478
tri -120 2476 -105 2491 nw
tri 7 2476 22 2491 ne
rect 22 2476 99 2491
tri 99 2476 114 2491 sw
rect -187 2467 -129 2476
tri -129 2467 -120 2476 nw
tri 22 2467 31 2476 ne
rect 31 2467 114 2476
tri 114 2467 123 2476 sw
rect -187 2466 -135 2467
tri -135 2461 -129 2467 nw
tri 31 2461 37 2467 ne
rect 37 2461 123 2467
tri 37 2454 44 2461 ne
rect 44 2454 123 2461
tri 123 2454 136 2467 sw
tri 44 2442 56 2454 ne
rect 56 2452 136 2454
tri 136 2452 138 2454 sw
rect 56 2442 138 2452
tri 56 2436 62 2442 ne
rect 62 2436 138 2442
rect -187 2408 -135 2414
rect -107 2424 -61 2436
rect -107 2390 -101 2424
rect -67 2390 -61 2424
tri 62 2404 94 2436 ne
tri -132 2352 -107 2377 se
rect -107 2352 -61 2390
rect -369 2318 -101 2352
rect -67 2318 -61 2352
rect -369 2306 -61 2318
rect 3 2330 55 2336
rect -369 2303 -261 2306
tri -261 2303 -258 2306 nw
rect -369 2284 -280 2303
tri -280 2284 -261 2303 nw
tri -14 2284 3 2301 se
rect -369 2261 -303 2284
tri -303 2261 -280 2284 nw
tri -37 2261 -14 2284 se
rect -14 2278 3 2284
rect -14 2266 55 2278
rect -14 2261 3 2266
rect -369 2153 -323 2261
tri -323 2241 -303 2261 nw
tri -45 2253 -37 2261 se
rect -37 2253 3 2261
rect -369 2119 -363 2153
rect -329 2119 -323 2153
rect -369 2081 -323 2119
rect -369 2047 -363 2081
rect -329 2047 -323 2081
rect -369 2035 -323 2047
rect -189 2214 3 2253
rect -189 2207 55 2214
rect -189 2185 -107 2207
tri -107 2185 -85 2207 nw
tri 77 2185 94 2202 se
rect 94 2185 138 2436
rect -189 2165 -127 2185
tri -127 2165 -107 2185 nw
tri 58 2166 77 2185 se
rect 77 2166 138 2185
tri 57 2165 58 2166 se
rect 58 2165 137 2166
tri 137 2165 138 2166 nw
rect -189 2153 -139 2165
tri -139 2153 -127 2165 nw
rect -16 2154 126 2165
tri 126 2154 137 2165 nw
rect -16 2153 123 2154
rect -189 2119 -183 2153
rect -149 2119 -143 2153
tri -143 2149 -139 2153 nw
rect -189 2081 -143 2119
rect -189 2047 -183 2081
rect -149 2047 -143 2081
rect -189 2035 -143 2047
rect -16 2119 -10 2153
rect 24 2151 123 2153
tri 123 2151 126 2154 nw
rect 24 2119 87 2151
rect -16 2115 87 2119
tri 87 2115 123 2151 nw
rect -16 2086 58 2115
tri 58 2086 87 2115 nw
rect -16 2081 53 2086
tri 53 2081 58 2086 nw
rect -16 2047 -10 2081
rect 24 2064 36 2081
tri 36 2064 53 2081 nw
rect 24 2047 30 2064
tri 30 2058 36 2064 nw
rect -16 2035 30 2047
rect -508 1946 152 1958
rect -508 1912 -277 1946
rect -243 1912 152 1946
rect -508 1874 152 1912
rect -508 1840 -277 1874
rect -243 1840 152 1874
rect -508 1779 152 1840
rect -508 1745 -423 1779
rect -389 1745 -344 1779
rect -310 1745 -265 1779
rect -231 1745 -187 1779
rect -153 1745 -109 1779
rect -75 1745 -31 1779
rect 3 1745 47 1779
rect 81 1745 152 1779
rect -508 1743 152 1745
rect -435 1739 152 1743
rect 262 1612 460 2533
tri 715 2526 722 2533 ne
rect 722 2526 757 2533
tri 757 2526 772 2541 sw
tri 8253 2526 8268 2541 se
rect 8268 2526 8398 2676
rect 8445 2687 8500 2693
rect 8497 2645 8500 2687
rect 8842 2686 9282 2694
rect 9334 2686 9346 2738
rect 9398 2686 9404 2738
rect 10378 2704 10428 2705
tri 10370 2696 10377 2703 se
rect 10377 2696 10429 2703
tri 10429 2696 10436 2703 sw
tri 10360 2686 10370 2696 se
rect 10370 2689 10436 2696
tri 10436 2689 10443 2696 sw
rect 10370 2686 10443 2689
tri 10352 2678 10360 2686 se
rect 10360 2678 10443 2686
tri 10443 2678 10454 2689 sw
tri 10766 2678 10777 2689 se
rect 10777 2678 10829 2768
rect 12399 2767 12406 2780
rect 12347 2754 12406 2767
rect 12399 2742 12406 2754
rect 12400 2708 12406 2742
rect 12399 2702 12406 2708
rect 12347 2696 12406 2702
rect 8993 2652 9371 2658
tri 8500 2645 8503 2648 sw
rect 8497 2635 8503 2645
rect 8445 2626 8503 2635
tri 8503 2626 8522 2645 sw
rect 8445 2623 8522 2626
rect 8497 2618 8522 2623
tri 8522 2618 8530 2626 sw
rect 8993 2618 9012 2652
rect 9046 2618 9084 2652
rect 9118 2618 9156 2652
rect 9190 2618 9228 2652
rect 9262 2618 9300 2652
rect 9334 2618 9371 2652
rect 8497 2601 8530 2618
tri 8530 2601 8547 2618 sw
rect 8993 2606 9371 2618
rect 9423 2606 9435 2658
rect 9487 2606 9493 2658
rect 9576 2626 9582 2678
rect 9634 2626 9646 2678
rect 9698 2626 10311 2678
rect 10313 2677 10349 2678
rect 10312 2627 10350 2677
rect 10313 2626 10349 2627
rect 10351 2626 10457 2678
tri 10752 2664 10766 2678 se
rect 10766 2664 10829 2678
tri 10667 2626 10705 2664 se
rect 10705 2626 10829 2664
rect 8497 2597 8547 2601
tri 8547 2597 8551 2601 sw
rect 8497 2571 8823 2597
rect 8445 2545 8823 2571
rect 8875 2545 8887 2597
rect 8939 2545 8945 2597
rect 8993 2581 9493 2606
tri 10208 2601 10233 2626 ne
rect 8994 2579 9492 2580
rect 9750 2560 10176 2572
rect 8994 2542 9492 2543
tri 8398 2526 8413 2541 sw
tri 8978 2526 8993 2541 se
rect 8993 2526 9493 2541
tri 722 2510 738 2526 ne
rect 738 2510 772 2526
tri 772 2510 788 2526 sw
tri 8243 2516 8253 2526 se
rect 8253 2516 8413 2526
tri 8413 2516 8423 2526 sw
tri 8968 2516 8978 2526 se
rect 8978 2516 9493 2526
rect 7512 2510 9493 2516
tri 738 2491 757 2510 ne
rect 757 2491 788 2510
tri 788 2491 807 2510 sw
tri 757 2476 772 2491 ne
rect 772 2476 807 2491
tri 807 2476 822 2491 sw
rect 7512 2476 7524 2510
rect 7558 2476 7596 2510
rect 7630 2476 9012 2510
rect 9046 2476 9084 2510
rect 9118 2476 9156 2510
rect 9190 2476 9228 2510
rect 9262 2476 9300 2510
rect 9334 2476 9372 2510
rect 9406 2476 9444 2510
rect 9478 2476 9493 2510
tri 772 2467 781 2476 ne
rect 781 2467 822 2476
tri 822 2467 831 2476 sw
rect 7512 2470 9493 2476
rect 9750 2526 9756 2560
rect 9790 2526 10136 2560
rect 10170 2526 10176 2560
rect 9750 2488 10176 2526
tri 781 2454 794 2467 ne
rect 794 2454 831 2467
tri 831 2454 844 2467 sw
tri 9737 2454 9750 2467 se
rect 9750 2454 9756 2488
rect 9790 2454 10136 2488
rect 10170 2454 10176 2488
rect 10233 2522 10285 2626
tri 10285 2601 10310 2626 nw
tri 10642 2601 10667 2626 se
rect 10667 2612 10829 2626
rect 10667 2601 10711 2612
tri 10637 2596 10642 2601 se
rect 10642 2596 10711 2601
tri 10711 2596 10727 2612 nw
tri 10752 2596 10768 2612 ne
rect 10768 2596 10829 2612
tri 10588 2547 10637 2596 se
rect 10637 2590 10705 2596
tri 10705 2590 10711 2596 nw
tri 10768 2590 10774 2596 ne
rect 10774 2590 10829 2596
tri 10285 2522 10310 2547 sw
tri 10563 2522 10588 2547 se
rect 10588 2522 10637 2547
tri 10637 2522 10705 2590 nw
tri 10774 2587 10777 2590 ne
rect 10777 2587 10829 2590
rect 10778 2585 10828 2586
rect 10778 2548 10828 2549
tri 10752 2522 10777 2547 se
rect 10777 2522 10829 2547
rect 10233 2470 10374 2522
rect 10376 2521 10412 2522
rect 10375 2471 10413 2521
rect 10376 2470 10412 2471
rect 10414 2470 10462 2522
rect 10514 2470 10526 2522
rect 10578 2510 10625 2522
tri 10625 2510 10637 2522 nw
rect 10578 2476 10591 2510
tri 10591 2476 10625 2510 nw
rect 10578 2470 10585 2476
tri 10585 2470 10591 2476 nw
rect 10701 2470 10707 2522
rect 10759 2470 10771 2522
rect 10823 2470 10829 2522
rect 10889 2470 10895 2522
rect 10947 2470 10959 2522
rect 11011 2516 11017 2522
tri 11823 2516 11829 2522 se
rect 11829 2516 11835 2522
rect 11011 2510 11473 2516
rect 11045 2476 11083 2510
rect 11117 2476 11355 2510
rect 11389 2476 11427 2510
rect 11461 2476 11473 2510
rect 11011 2470 11473 2476
rect 11697 2510 11835 2516
rect 11697 2476 11709 2510
rect 11743 2476 11781 2510
rect 11815 2476 11835 2510
rect 11697 2470 11835 2476
rect 11887 2470 11899 2522
rect 11951 2516 11957 2522
tri 11957 2516 11963 2522 sw
rect 11951 2510 12492 2516
rect 11951 2476 12053 2510
rect 12087 2476 12125 2510
rect 12159 2476 12440 2510
rect 11951 2470 12440 2476
tri 12406 2467 12409 2470 ne
rect 12409 2467 12440 2470
tri 794 2443 805 2454 ne
rect 805 2443 844 2454
tri 844 2443 855 2454 sw
tri 9726 2443 9737 2454 se
rect 9737 2443 10176 2454
tri 805 2442 806 2443 ne
rect 806 2442 859 2443
tri 9725 2442 9726 2443 se
rect 9726 2442 10176 2443
tri 10176 2442 10201 2467 sw
tri 12409 2442 12434 2467 ne
rect 12434 2458 12440 2467
rect 12434 2446 12492 2458
rect 12434 2442 12440 2446
tri 806 2441 807 2442 ne
rect 807 2437 859 2442
rect 807 2373 859 2385
rect 807 2315 859 2321
rect 942 2390 1704 2442
rect 1756 2390 1773 2442
rect 1825 2390 1842 2442
rect 1894 2390 1911 2442
rect 1963 2390 1980 2442
rect 2032 2390 3156 2442
rect 3208 2390 3220 2442
rect 3272 2390 3284 2442
rect 3336 2390 3348 2442
rect 3400 2390 3412 2442
rect 3464 2390 3476 2442
rect 3528 2390 3540 2442
rect 3592 2436 12311 2442
tri 12434 2436 12440 2442 ne
rect 3592 2402 7997 2436
rect 8031 2402 8069 2436
rect 8103 2402 8141 2436
rect 8175 2430 12311 2436
rect 8175 2402 8614 2430
rect 3592 2390 8614 2402
rect 942 2364 8614 2390
rect 942 2312 1704 2364
rect 1756 2312 1773 2364
rect 1825 2312 1842 2364
rect 1894 2312 1911 2364
rect 1963 2312 1980 2364
rect 2032 2312 3156 2364
rect 3208 2312 3220 2364
rect 3272 2312 3284 2364
rect 3336 2312 3348 2364
rect 3400 2312 3412 2364
rect 3464 2312 3476 2364
rect 3528 2312 3540 2364
rect 3592 2324 8614 2364
rect 8720 2324 12311 2430
rect 3592 2312 12311 2324
rect 12347 2419 12406 2425
rect 12399 2413 12406 2419
rect 12400 2379 12406 2413
rect 12440 2388 12492 2394
rect 12399 2367 12406 2379
rect 12347 2354 12406 2367
rect 12399 2337 12406 2354
rect 12400 2303 12406 2337
rect 12399 2302 12406 2303
rect 12347 2289 12406 2302
tri 7420 2261 7443 2284 se
rect 7443 2261 9443 2284
tri 7391 2232 7420 2261 se
rect 7420 2232 9443 2261
rect 9495 2232 9507 2284
rect 9559 2278 11904 2284
rect 9559 2232 11852 2278
tri 7386 2227 7391 2232 se
rect 7391 2227 7460 2232
tri 7460 2227 7465 2232 nw
tri 11790 2227 11795 2232 ne
rect 11795 2227 11852 2232
tri 7366 2207 7386 2227 se
rect 7386 2207 7440 2227
tri 7440 2207 7460 2227 nw
tri 11795 2207 11815 2227 ne
rect 11815 2226 11852 2227
rect 11815 2214 11904 2226
rect 11815 2207 11852 2214
tri 7365 2206 7366 2207 se
rect 7366 2206 7418 2207
rect 6747 2154 6753 2206
rect 6805 2154 6817 2206
rect 6869 2185 7418 2206
tri 7418 2185 7440 2207 nw
tri 11815 2204 11818 2207 ne
rect 11818 2204 11852 2207
rect 6869 2170 7403 2185
tri 7403 2170 7418 2185 nw
rect 6869 2165 7398 2170
tri 7398 2165 7403 2170 nw
rect 6869 2158 7391 2165
tri 7391 2158 7398 2165 nw
rect 6869 2156 7389 2158
tri 7389 2156 7391 2158 nw
rect 6869 2154 7387 2156
tri 7387 2154 7389 2156 nw
rect 8891 2152 8898 2204
rect 8950 2152 8962 2204
rect 9014 2155 10566 2204
rect 9014 2154 9668 2155
tri 9668 2154 9669 2155 nw
tri 10397 2154 10398 2155 ne
rect 10398 2154 10566 2155
rect 9014 2152 9666 2154
tri 9666 2152 9668 2154 nw
tri 10398 2152 10400 2154 ne
rect 10400 2152 10566 2154
rect 10618 2152 10630 2204
rect 10682 2152 10688 2204
tri 11818 2203 11819 2204 ne
rect 11819 2203 11852 2204
tri 10770 2194 10779 2203 se
rect 10779 2194 10882 2203
tri 10761 2185 10770 2194 se
rect 10770 2185 10882 2194
tri 10746 2170 10761 2185 se
rect 10761 2170 10882 2185
tri 10732 2156 10746 2170 se
rect 10746 2156 10882 2170
tri 10728 2152 10732 2156 se
rect 10732 2152 10882 2156
tri 10727 2151 10728 2152 se
rect 10728 2151 10882 2152
rect 10934 2151 10946 2203
rect 10998 2151 11004 2203
tri 11819 2193 11829 2203 ne
rect 11829 2193 11852 2203
rect 11397 2187 11449 2193
tri 11392 2151 11397 2156 se
tri 10703 2127 10727 2151 se
rect 10727 2127 10770 2151
rect 9692 2115 10374 2127
tri 10700 2124 10703 2127 se
rect 10703 2124 10770 2127
tri 10770 2124 10797 2151 nw
tri 11365 2124 11392 2151 se
rect 11392 2135 11397 2151
tri 11829 2185 11837 2193 ne
rect 11837 2185 11852 2193
tri 11837 2170 11852 2185 ne
rect 11852 2156 11904 2162
rect 12399 2261 12406 2289
rect 12347 2227 12366 2237
rect 12400 2227 12406 2261
rect 12347 2223 12406 2227
rect 14840 2226 15007 2382
rect 12399 2185 12406 2223
rect 12347 2157 12366 2171
tri 11449 2151 11454 2156 sw
rect 12400 2151 12406 2185
rect 11449 2135 11454 2151
rect 11392 2124 11454 2135
tri 11454 2124 11481 2151 sw
rect 9692 2081 9698 2115
rect 9732 2081 9770 2115
rect 9804 2081 9982 2115
rect 10016 2081 10054 2115
rect 10088 2081 10262 2115
rect 10296 2081 10334 2115
rect 10368 2081 10374 2115
rect 9692 2069 10374 2081
rect 10462 2072 10468 2124
rect 10520 2072 10532 2124
rect 10584 2109 10755 2124
tri 10755 2109 10770 2124 nw
tri 11350 2109 11365 2124 se
rect 11365 2116 11481 2124
rect 11365 2109 11397 2116
rect 10584 2098 10744 2109
tri 10744 2098 10755 2109 nw
tri 11345 2104 11350 2109 se
rect 11350 2104 11397 2109
rect 10791 2098 11397 2104
rect 10584 2086 10732 2098
tri 10732 2086 10744 2098 nw
rect 10584 2072 10718 2086
tri 10718 2072 10732 2086 nw
rect 10791 2064 10804 2098
rect 10838 2064 10876 2098
rect 10910 2064 11102 2098
rect 11136 2064 11174 2098
rect 11208 2064 11397 2098
rect 11449 2109 11481 2116
tri 11481 2109 11496 2124 sw
rect 12399 2109 12406 2151
rect 11449 2104 11496 2109
tri 11496 2104 11501 2109 sw
rect 11449 2098 11936 2104
rect 11449 2064 11459 2098
rect 11493 2064 11537 2098
rect 11571 2064 11806 2098
rect 11840 2064 11878 2098
rect 11912 2064 11936 2098
rect 10791 2058 11936 2064
rect 12347 2091 12366 2105
rect 12400 2075 12406 2109
rect 12399 2039 12406 2075
rect 12347 2033 12406 2039
rect 948 2029 12211 2030
rect 948 1977 1704 2029
rect 1756 1977 1773 2029
rect 1825 1977 1842 2029
rect 1894 1977 1911 2029
rect 1963 1977 1980 2029
rect 2032 1977 3156 2029
rect 3208 1977 3220 2029
rect 3272 1977 3284 2029
rect 3336 1977 3348 2029
rect 3400 1977 3412 2029
rect 3464 1977 3476 2029
rect 3528 1977 3540 2029
rect 3592 2019 12211 2029
rect 3592 1985 7930 2019
rect 7964 2018 12211 2019
rect 7964 1985 8678 2018
rect 3592 1984 8678 1985
rect 8712 2013 10960 2018
rect 8712 2012 9441 2013
rect 8712 1984 8977 2012
rect 3592 1978 8977 1984
rect 9011 1978 9329 2012
rect 9363 1978 9441 2012
rect 3592 1977 9441 1978
rect 948 1955 9441 1977
rect 948 1903 1704 1955
rect 1756 1903 1773 1955
rect 1825 1903 1842 1955
rect 1894 1903 1911 1955
rect 1963 1903 1980 1955
rect 2032 1903 3156 1955
rect 3208 1903 3220 1955
rect 3272 1903 3284 1955
rect 3336 1903 3348 1955
rect 3400 1903 3412 1955
rect 3464 1903 3476 1955
rect 3528 1903 3540 1955
rect 3592 1947 9441 1955
rect 3592 1913 7930 1947
rect 7964 1946 9441 1947
rect 7964 1913 8678 1946
rect 3592 1912 8678 1913
rect 8712 1940 9441 1946
rect 8712 1912 8977 1940
rect 3592 1906 8977 1912
rect 9011 1906 9329 1940
rect 9363 1906 9441 1940
rect 3592 1903 9441 1906
rect 948 1881 9441 1903
rect 948 1829 1704 1881
rect 1756 1829 1773 1881
rect 1825 1829 1842 1881
rect 1894 1829 1911 1881
rect 1963 1829 1980 1881
rect 2032 1829 3156 1881
rect 3208 1829 3220 1881
rect 3272 1829 3284 1881
rect 3336 1829 3348 1881
rect 3400 1829 3412 1881
rect 3464 1829 3476 1881
rect 3528 1829 3540 1881
rect 3592 1875 9441 1881
rect 3592 1841 7930 1875
rect 7964 1874 9441 1875
rect 7964 1841 8678 1874
rect 3592 1840 8678 1841
rect 8712 1868 9441 1874
rect 8712 1840 8977 1868
rect 3592 1834 8977 1840
rect 9011 1834 9329 1868
rect 9363 1835 9441 1868
rect 9547 2012 10960 2013
rect 9547 1978 10192 2012
rect 10226 1978 10486 2012
rect 10520 1984 10960 2012
rect 10994 1984 11312 2018
rect 11346 1984 11664 2018
rect 11698 1984 12016 2018
rect 12050 1984 12102 2018
rect 12136 1984 12211 2018
rect 10520 1978 12211 1984
rect 9547 1946 12211 1978
rect 9547 1940 10960 1946
rect 9547 1906 10192 1940
rect 10226 1906 10486 1940
rect 10520 1912 10960 1940
rect 10994 1912 11312 1946
rect 11346 1912 11664 1946
rect 11698 1912 12016 1946
rect 12050 1912 12102 1946
rect 12136 1912 12211 1946
rect 10520 1906 12211 1912
rect 9547 1874 12211 1906
rect 9547 1873 10960 1874
rect 9547 1868 10560 1873
rect 9547 1835 10192 1868
rect 9363 1834 10192 1835
rect 10226 1834 10486 1868
rect 10520 1840 10560 1868
tri 10560 1840 10593 1873 nw
tri 10759 1840 10792 1873 ne
rect 10792 1840 10960 1873
rect 10994 1840 11312 1874
rect 11346 1840 11664 1874
rect 11698 1840 12016 1874
rect 12050 1840 12102 1874
rect 12136 1840 12211 1874
rect 10520 1834 10548 1840
rect 3592 1829 10548 1834
rect 948 1828 10548 1829
tri 10548 1828 10560 1840 nw
tri 10792 1828 10804 1840 ne
rect 10804 1828 12211 1840
rect 12347 2025 12366 2033
rect 12400 1999 12406 2033
rect 12399 1973 12406 1999
rect 12347 1959 12406 1973
rect 12399 1957 12406 1959
rect 12400 1923 12406 1957
rect 12399 1907 12406 1923
rect 12347 1893 12406 1907
rect 12399 1881 12406 1893
rect 12400 1847 12406 1881
rect 12399 1841 12406 1847
rect 12347 1835 12406 1841
rect 8535 1772 12799 1800
rect 7301 1765 7353 1771
tri 7353 1744 7380 1771 sw
rect 8535 1758 8685 1772
tri 8685 1758 8699 1772 nw
tri 12779 1758 12793 1772 ne
rect 12793 1758 12799 1772
tri 12799 1758 12841 1800 sw
rect 7353 1726 7380 1744
tri 7380 1726 7398 1744 sw
rect 7353 1722 7398 1726
tri 7398 1722 7402 1726 sw
rect 7353 1720 7402 1722
tri 7402 1720 7404 1722 sw
rect 8535 1720 8665 1758
tri 8665 1738 8685 1758 nw
tri 12793 1752 12799 1758 ne
rect 12799 1752 12841 1758
tri 12799 1744 12807 1752 ne
rect 12807 1744 12841 1752
tri 10232 1738 10238 1744 se
rect 10238 1738 10618 1744
tri 10226 1732 10232 1738 se
rect 10232 1732 10618 1738
rect 7353 1719 7404 1720
tri 7404 1719 7405 1720 sw
rect 7353 1713 8279 1719
rect 7301 1701 8279 1713
rect 706 1654 758 1660
tri 460 1612 480 1632 sw
rect 262 1578 480 1612
tri 480 1578 514 1612 sw
tri 672 1578 706 1612 se
rect 7163 1654 7215 1660
tri 758 1606 764 1612 sw
rect 758 1602 764 1606
rect 706 1590 764 1602
rect 262 1576 514 1578
tri 514 1576 516 1578 sw
rect 262 1572 516 1576
tri 516 1572 520 1576 sw
rect 262 1566 520 1572
tri 520 1566 526 1572 sw
rect 262 1538 526 1566
tri 526 1538 554 1566 sw
rect 686 1538 706 1578
rect 758 1578 764 1590
tri 764 1578 792 1606 sw
rect 7353 1692 8279 1701
tri 8279 1692 8306 1719 sw
rect 7353 1687 8306 1692
tri 8306 1687 8311 1692 sw
rect 7353 1686 7396 1687
tri 7396 1686 7397 1687 nw
tri 8137 1686 8138 1687 ne
rect 8138 1686 8311 1687
tri 8311 1686 8312 1687 sw
rect 8535 1686 8547 1720
rect 8581 1686 8619 1720
rect 8653 1686 8665 1720
rect 7353 1658 7368 1686
tri 7368 1658 7396 1686 nw
tri 8138 1658 8166 1686 ne
rect 8166 1658 8312 1686
tri 8312 1658 8340 1686 sw
rect 8535 1680 8665 1686
rect 8711 1680 8717 1732
rect 8769 1720 8806 1732
rect 8780 1686 8806 1720
rect 8769 1680 8806 1686
rect 8858 1680 8864 1732
rect 8935 1722 9019 1732
rect 8935 1688 8947 1722
rect 8981 1688 9019 1722
rect 8935 1680 9019 1688
rect 9071 1680 9083 1732
rect 9135 1680 9674 1732
rect 9726 1680 9738 1732
rect 9790 1680 9796 1732
tri 10186 1692 10226 1732 se
rect 10226 1692 10618 1732
rect 10670 1692 10682 1744
rect 10734 1692 10740 1744
tri 12807 1738 12813 1744 ne
tri 10174 1680 10186 1692 se
rect 10186 1680 10248 1692
tri 10248 1680 10260 1692 nw
tri 10152 1658 10174 1680 se
rect 10174 1658 10226 1680
tri 10226 1658 10248 1680 nw
rect 10273 1658 10373 1664
rect 10425 1658 10437 1664
rect 7353 1649 7356 1658
rect 7301 1646 7356 1649
tri 7356 1646 7368 1658 nw
rect 7828 1646 7997 1658
rect 7301 1643 7353 1646
tri 7353 1643 7356 1646 nw
rect 7828 1612 7840 1646
rect 7874 1612 7912 1646
rect 7946 1612 7997 1646
rect 7828 1606 7997 1612
rect 8049 1606 8061 1658
rect 8113 1606 8119 1658
tri 8166 1652 8172 1658 ne
rect 8172 1652 8340 1658
tri 8340 1652 8346 1658 sw
tri 10146 1652 10152 1658 se
rect 10152 1652 10220 1658
tri 10220 1652 10226 1658 nw
rect 8172 1646 9435 1652
rect 8172 1612 8184 1646
rect 8218 1612 8256 1646
rect 8290 1612 9432 1646
rect 8172 1606 9435 1612
tri 9423 1603 9426 1606 ne
rect 9426 1603 9435 1606
rect 7163 1590 7215 1602
rect 262 1532 554 1538
tri 554 1532 560 1538 sw
rect 686 1532 758 1538
tri 7215 1578 7240 1603 sw
tri 9426 1600 9429 1603 ne
rect 9429 1600 9435 1603
rect 9487 1600 9499 1652
rect 9551 1624 10192 1652
tri 10192 1624 10220 1652 nw
rect 10273 1624 10285 1658
rect 10319 1624 10357 1658
rect 10425 1624 10429 1658
rect 9551 1618 10186 1624
tri 10186 1618 10192 1624 nw
rect 9551 1616 10184 1618
tri 10184 1616 10186 1618 nw
rect 9551 1612 10180 1616
tri 10180 1612 10184 1616 nw
rect 10273 1612 10373 1624
rect 10425 1612 10437 1624
rect 10489 1612 10495 1664
rect 10523 1612 10707 1664
rect 10759 1612 10771 1664
rect 10823 1654 11150 1664
rect 10823 1612 11098 1654
rect 9551 1606 9563 1612
tri 9563 1606 9569 1612 nw
rect 9551 1603 9560 1606
tri 9560 1603 9563 1606 nw
rect 9551 1600 9557 1603
tri 9557 1600 9560 1603 nw
tri 9579 1578 9585 1584 se
rect 9585 1578 9591 1584
rect 7215 1576 9374 1578
tri 9374 1576 9376 1578 sw
tri 9577 1576 9579 1578 se
rect 9579 1576 9591 1578
rect 7215 1572 9376 1576
tri 9376 1572 9380 1576 sw
tri 9573 1572 9577 1576 se
rect 9577 1572 9591 1576
rect 7215 1538 7426 1572
rect 7460 1538 7498 1572
rect 7532 1538 9591 1572
rect 7163 1532 9591 1538
rect 9643 1532 9655 1584
rect 9707 1578 9713 1584
tri 9713 1578 9719 1584 sw
rect 9707 1572 10004 1578
rect 9707 1538 9742 1572
rect 9776 1538 9814 1572
rect 9848 1538 9886 1572
rect 9920 1538 9958 1572
rect 9992 1538 10004 1572
rect 9707 1532 10004 1538
rect 10523 1569 10575 1612
tri 10575 1587 10600 1612 nw
tri 11066 1587 11091 1612 ne
rect 11091 1602 11098 1612
rect 11091 1590 11150 1602
rect 11091 1587 11098 1590
tri 11091 1584 11094 1587 ne
rect 11094 1584 11098 1587
rect 10524 1567 10574 1568
rect 262 1504 560 1532
tri 560 1504 588 1532 sw
rect 10523 1531 10575 1567
rect 10627 1532 10633 1584
rect 10685 1532 10703 1584
rect 10755 1532 10773 1584
rect 10825 1532 10831 1584
rect 10903 1532 10909 1584
rect 10961 1532 10973 1584
rect 11025 1532 11035 1584
tri 11094 1580 11098 1584 ne
rect 11098 1532 11150 1538
rect 10524 1530 10574 1531
tri 10498 1504 10523 1529 se
rect 10523 1504 10575 1529
tri 10575 1504 10600 1529 sw
rect 262 1503 1799 1504
rect 262 1451 992 1503
rect 1044 1451 1061 1503
rect 1113 1451 1130 1503
rect 1182 1451 1199 1503
rect 1251 1451 1268 1503
rect 1320 1451 1337 1503
rect 1389 1451 1405 1503
rect 1457 1451 1473 1503
rect 1525 1500 1799 1503
tri 1799 1500 1803 1504 sw
tri 1981 1500 1985 1504 se
rect 1985 1500 12676 1504
rect 1525 1498 1803 1500
tri 1803 1498 1805 1500 sw
tri 1979 1498 1981 1500 se
rect 1981 1498 12676 1500
rect 1525 1486 1805 1498
tri 1805 1486 1817 1498 sw
tri 1967 1486 1979 1498 se
rect 1979 1486 9040 1498
rect 1525 1468 1817 1486
tri 1817 1468 1835 1486 sw
tri 1949 1468 1967 1486 se
rect 1967 1468 7422 1486
rect 1525 1452 7422 1468
rect 7456 1452 7774 1486
rect 7808 1464 9040 1486
rect 9074 1492 12347 1498
rect 12399 1492 12676 1498
rect 9074 1486 10455 1492
rect 9074 1464 9658 1486
rect 7808 1452 9658 1464
rect 9692 1452 9912 1486
rect 9946 1452 10224 1486
rect 10258 1458 10455 1486
rect 10489 1458 12347 1492
rect 12400 1489 12676 1492
tri 12676 1489 12691 1504 sw
rect 12813 1496 12841 1744
tri 12813 1489 12820 1496 ne
rect 12820 1489 12841 1496
tri 12841 1489 12875 1523 sw
tri 14792 1489 14826 1523 se
rect 12400 1468 12691 1489
tri 12691 1468 12712 1489 sw
tri 12820 1468 12841 1489 ne
rect 12841 1468 14872 1489
rect 12400 1461 12712 1468
tri 12712 1461 12719 1468 sw
tri 12841 1461 12848 1468 ne
rect 12848 1461 14872 1468
rect 12400 1458 12719 1461
rect 10258 1452 12347 1458
rect 1525 1451 12347 1452
rect 262 1446 12347 1451
rect 12399 1446 12719 1458
rect 262 1429 12719 1446
rect 262 1377 992 1429
rect 1044 1377 1061 1429
rect 1113 1377 1130 1429
rect 1182 1377 1199 1429
rect 1251 1377 1268 1429
rect 1320 1377 1337 1429
rect 1389 1377 1405 1429
rect 1457 1377 1473 1429
rect 1525 1426 12347 1429
rect 1525 1414 9040 1426
rect 1525 1380 7422 1414
rect 7456 1380 7774 1414
rect 7808 1392 9040 1414
rect 9074 1422 12347 1426
rect 9074 1414 11040 1422
rect 9074 1392 9658 1414
rect 7808 1380 9658 1392
rect 9692 1380 9912 1414
rect 9946 1380 10224 1414
rect 10258 1413 11040 1414
rect 10258 1380 10455 1413
rect 1525 1379 10455 1380
rect 10489 1388 11040 1413
rect 11074 1421 12347 1422
rect 11074 1388 12225 1421
rect 10489 1387 12225 1388
rect 12259 1387 12347 1421
rect 12399 1423 12719 1429
tri 12719 1423 12757 1461 sw
rect 12399 1420 12817 1423
rect 10489 1379 12347 1387
rect 12400 1386 12817 1420
rect 1525 1377 12347 1379
rect 12399 1377 12817 1386
rect 262 1360 12817 1377
rect 262 1355 12347 1360
rect 262 1303 992 1355
rect 1044 1303 1061 1355
rect 1113 1303 1130 1355
rect 1182 1303 1199 1355
rect 1251 1303 1268 1355
rect 1320 1303 1337 1355
rect 1389 1303 1405 1355
rect 1457 1303 1473 1355
rect 1525 1354 12347 1355
rect 1525 1342 9040 1354
rect 1525 1308 7422 1342
rect 7456 1308 7774 1342
rect 7808 1320 9040 1342
rect 9074 1350 12347 1354
rect 9074 1342 11040 1350
rect 9074 1320 9658 1342
rect 7808 1308 9658 1320
rect 9692 1308 9912 1342
rect 9946 1308 10224 1342
rect 10258 1334 11040 1342
rect 10258 1308 10455 1334
rect 1525 1303 10455 1308
rect 262 1302 10455 1303
rect 262 1300 337 1302
tri 337 1300 339 1302 nw
tri 10413 1300 10415 1302 ne
rect 10415 1300 10455 1302
rect 10489 1316 11040 1334
rect 11074 1349 12347 1350
rect 11074 1316 12225 1349
rect 10489 1315 12225 1316
rect 12259 1315 12347 1349
rect 12399 1348 12817 1360
rect 10489 1308 12347 1315
rect 12400 1314 12817 1348
rect 12399 1308 12817 1314
rect 10489 1302 12817 1308
rect 10489 1300 10506 1302
rect 262 801 314 1300
tri 314 1277 337 1300 nw
tri 10415 1277 10438 1300 ne
rect 10438 1277 10506 1300
tri 10506 1277 10531 1302 nw
tri 12599 1277 12624 1302 ne
rect 12624 1277 12817 1302
tri 10438 1274 10441 1277 ne
rect 10441 1274 10503 1277
tri 10503 1274 10506 1277 nw
tri 12624 1274 12627 1277 ne
rect 12627 1274 12817 1277
rect 6054 1228 6094 1274
rect 6190 1228 6231 1274
rect 7577 1222 7583 1274
rect 7635 1222 7647 1274
rect 7699 1268 8144 1274
tri 8144 1268 8150 1274 sw
rect 8872 1268 9626 1274
tri 10441 1268 10447 1274 ne
rect 10447 1268 10497 1274
tri 10497 1268 10503 1274 nw
rect 10549 1268 11274 1274
rect 7699 1237 8150 1268
tri 8150 1237 8181 1268 sw
rect 7699 1234 8181 1237
tri 8181 1234 8184 1237 sw
rect 8872 1234 8884 1268
rect 8918 1234 8956 1268
rect 8990 1234 9160 1268
rect 9194 1234 9232 1268
rect 9266 1234 9508 1268
rect 9542 1234 9580 1268
rect 9614 1234 9626 1268
tri 10447 1266 10449 1268 ne
rect 7699 1222 8184 1234
tri 8184 1222 8196 1234 sw
rect 8872 1228 9626 1234
rect 10449 1255 10495 1268
tri 10495 1266 10497 1268 nw
tri 8134 1221 8135 1222 ne
rect 8135 1221 8196 1222
tri 8196 1221 8197 1222 sw
rect 10449 1221 10455 1255
rect 10489 1221 10495 1255
rect 10549 1234 10561 1268
rect 10595 1234 10633 1268
rect 10667 1234 11156 1268
rect 11190 1234 11228 1268
rect 11262 1234 11274 1268
tri 12627 1259 12642 1274 ne
rect 12642 1259 12817 1274
tri 11773 1253 11779 1259 se
rect 11779 1253 12287 1259
tri 11757 1237 11773 1253 se
rect 11773 1237 11791 1253
rect 10549 1228 11274 1234
tri 11748 1228 11757 1237 se
rect 11757 1228 11791 1237
tri 11742 1222 11748 1228 se
rect 11748 1222 11791 1228
tri 8135 1219 8137 1221 ne
rect 8137 1219 8197 1221
tri 8197 1219 8199 1221 sw
tri 8137 1208 8148 1219 ne
rect 8148 1208 8199 1219
tri 8199 1208 8210 1219 sw
tri 8148 1194 8162 1208 ne
rect 8162 1198 8210 1208
tri 8210 1198 8220 1208 sw
rect 8162 1194 9674 1198
rect 7552 1188 7996 1194
rect 4498 1112 4504 1164
rect 4556 1112 4568 1164
rect 4620 1112 5478 1164
rect 5530 1112 5542 1164
rect 5594 1112 5600 1164
rect 7552 1154 7564 1188
rect 7598 1154 7636 1188
rect 7670 1154 7878 1188
rect 7912 1154 7950 1188
rect 7984 1154 7996 1188
tri 8162 1176 8180 1194 ne
rect 8180 1176 9674 1194
tri 8180 1164 8192 1176 ne
rect 8192 1164 9674 1176
rect 7552 1148 7996 1154
tri 8192 1148 8208 1164 ne
rect 8208 1148 9674 1164
tri 8208 1146 8210 1148 ne
rect 8210 1146 9674 1148
rect 9726 1146 9738 1198
rect 9790 1146 9796 1198
rect 10449 1176 10495 1221
tri 11739 1219 11742 1222 se
rect 11742 1219 11791 1222
rect 11825 1219 11872 1253
rect 11906 1219 11953 1253
rect 11987 1219 12034 1253
rect 12068 1219 12235 1253
tri 11728 1208 11739 1219 se
rect 11739 1208 12235 1219
tri 11718 1198 11728 1208 se
rect 11728 1201 12235 1208
tri 12642 1237 12664 1259 ne
rect 12664 1237 12817 1259
tri 12287 1203 12321 1237 sw
tri 12664 1203 12698 1237 ne
rect 12698 1203 12817 1237
rect 12287 1201 12499 1203
rect 11728 1198 12499 1201
tri 11713 1193 11718 1198 se
rect 11718 1193 12499 1198
tri 10657 1189 10661 1193 se
rect 10661 1189 12499 1193
rect 10449 1142 10455 1176
rect 10489 1142 10495 1176
tri 10639 1171 10657 1189 se
rect 10657 1171 12235 1189
tri 10617 1149 10639 1171 se
rect 10639 1149 11791 1171
tri 10614 1146 10617 1149 se
rect 10617 1146 10686 1149
tri 10686 1146 10689 1149 nw
tri 11761 1146 11764 1149 ne
rect 11764 1146 11791 1149
rect 10449 1130 10495 1142
tri 10605 1137 10614 1146 se
rect 10614 1137 10677 1146
tri 10677 1137 10686 1146 nw
tri 11764 1137 11773 1146 ne
rect 11773 1137 11791 1146
rect 11825 1137 11872 1171
rect 11906 1137 11953 1171
rect 11987 1137 12034 1171
rect 12068 1137 12235 1171
rect 12287 1179 12499 1189
tri 12499 1179 12523 1203 sw
tri 12698 1179 12722 1203 ne
rect 12722 1179 12817 1203
rect 12287 1151 12523 1179
tri 10604 1136 10605 1137 se
rect 10605 1136 10671 1137
tri 10599 1131 10604 1136 se
rect 10604 1131 10671 1136
tri 10671 1131 10677 1137 nw
tri 11773 1131 11779 1137 ne
rect 11779 1131 12287 1137
tri 12287 1131 12307 1151 nw
tri 12477 1131 12497 1151 ne
rect 12497 1131 12523 1151
tri 10598 1130 10599 1131 se
rect 10599 1130 10661 1131
tri 10589 1121 10598 1130 se
rect 10598 1121 10661 1130
tri 10661 1121 10671 1131 nw
tri 12497 1121 12507 1131 ne
rect 12507 1121 12523 1131
tri 12523 1121 12581 1179 sw
tri 12722 1133 12768 1179 ne
rect 12768 1133 12817 1179
rect 12694 1121 12740 1133
tri 10586 1118 10589 1121 se
rect 10589 1118 10657 1121
rect 9744 1112 10414 1118
tri 10585 1117 10586 1118 se
rect 10586 1117 10657 1118
tri 10657 1117 10661 1121 nw
tri 12507 1117 12511 1121 ne
rect 12511 1117 12581 1121
tri 10580 1112 10585 1117 se
rect 10585 1112 10657 1117
rect 9744 1078 9756 1112
rect 9790 1078 9828 1112
rect 9862 1078 10022 1112
rect 10056 1078 10094 1112
rect 10128 1078 10296 1112
rect 10330 1078 10368 1112
rect 10402 1078 10414 1112
tri 10573 1105 10580 1112 se
rect 10580 1105 10657 1112
tri 12511 1105 12523 1117 ne
rect 12523 1105 12581 1117
tri 12581 1105 12597 1121 sw
rect 409 1013 553 1044
rect 8148 1030 8194 1076
rect 9306 1070 9436 1076
rect 9744 1072 10414 1078
rect 10443 1091 10495 1097
rect 9306 1036 9318 1070
rect 9352 1036 9390 1070
rect 9424 1036 9436 1070
rect 9306 1030 9436 1036
rect 10529 1053 10535 1105
rect 10587 1053 10599 1105
rect 10651 1053 10657 1105
tri 12523 1096 12532 1105 ne
rect 12532 1096 12597 1105
rect 12153 1090 12205 1096
tri 12532 1093 12535 1096 ne
rect 12535 1093 12597 1096
rect 10443 1027 10495 1039
tri 10429 1013 10443 1027 se
tri 10426 1010 10429 1013 se
rect 10429 1010 10443 1013
tri 10425 1009 10426 1010 se
rect 10426 1009 10443 1010
tri 10418 1002 10425 1009 se
rect 10425 1002 10443 1009
rect 7426 975 10443 1002
rect 12153 1026 12205 1038
rect 7426 974 10495 975
tri 10438 969 10443 974 ne
rect 10443 969 10495 974
rect 10702 969 10708 1021
rect 10760 969 10773 1021
rect 10825 1015 10831 1021
tri 10831 1015 10837 1021 sw
rect 10825 1009 11762 1015
rect 10825 975 10932 1009
rect 10966 975 11011 1009
rect 11045 975 11090 1009
rect 11124 975 11169 1009
rect 11203 975 11248 1009
rect 11282 975 11326 1009
rect 11360 975 11404 1009
rect 11438 975 11482 1009
rect 11516 975 11560 1009
rect 11594 975 11638 1009
rect 11672 975 11716 1009
rect 11750 975 11762 1009
rect 10825 969 11762 975
tri 12148 969 12153 974 se
rect 12153 969 12205 974
tri 12147 968 12148 969 se
rect 12148 968 12205 969
tri 12146 967 12147 968 se
rect 12147 967 12205 968
tri 12124 945 12146 967 se
rect 12146 945 12205 967
tri 6887 940 6892 945 se
rect 6892 940 7834 945
tri 7834 940 7839 945 sw
tri 12119 940 12124 945 se
rect 12124 940 12205 945
tri 6882 935 6887 940 se
rect 6887 935 7839 940
tri 7839 935 7844 940 sw
tri 6873 926 6882 935 se
rect 6882 926 7844 935
rect 5472 874 5478 926
rect 5530 874 5542 926
rect 5594 920 5600 926
tri 5600 920 5606 926 sw
tri 6867 920 6873 926 se
rect 6873 920 7844 926
tri 7844 920 7859 935 sw
rect 5594 903 7859 920
tri 7859 903 7876 920 sw
rect 5594 901 7876 903
tri 7876 901 7878 903 sw
rect 5594 899 7878 901
tri 7878 899 7880 901 sw
rect 5594 896 6909 899
tri 6909 896 6912 899 nw
tri 7814 896 7817 899 ne
rect 7817 897 7880 899
tri 7880 897 7882 899 sw
rect 7817 896 8466 897
tri 8466 896 8467 897 sw
rect 5594 888 6901 896
tri 6901 888 6909 896 nw
tri 7817 888 7825 896 ne
rect 7825 888 8467 896
tri 8467 888 8475 896 sw
rect 5594 874 6887 888
tri 6887 874 6901 888 nw
tri 7825 874 7839 888 ne
rect 7839 874 8475 888
tri 7839 862 7851 874 ne
rect 7851 862 8475 874
tri 8475 862 8501 888 sw
tri 7851 851 7862 862 ne
rect 7862 851 8501 862
tri 8501 851 8512 862 sw
rect 9013 851 9019 903
rect 9071 851 9085 903
rect 9137 851 9143 903
tri 8446 822 8475 851 ne
rect 8475 822 8512 851
tri 8512 822 8541 851 sw
rect 9340 850 9346 902
rect 9398 896 9438 902
rect 9398 862 9424 896
rect 9398 850 9438 862
rect 9490 850 9496 902
rect 9668 887 9674 939
rect 9726 887 9738 939
rect 9790 887 10496 939
rect 10548 887 10560 939
rect 10612 887 10618 939
rect 10737 888 10743 940
rect 10795 888 10807 940
rect 10859 898 12205 940
rect 12347 1087 12406 1093
tri 12535 1087 12541 1093 ne
rect 12541 1087 12597 1093
rect 12399 1081 12406 1087
tri 12541 1084 12544 1087 ne
rect 12544 1084 12597 1087
tri 12544 1083 12545 1084 ne
rect 12400 1047 12406 1081
rect 12399 1035 12406 1047
rect 12347 1011 12406 1035
rect 12399 1008 12406 1011
rect 12400 974 12406 1008
rect 12399 959 12406 974
rect 12347 935 12406 959
rect 12347 934 12366 935
rect 12400 901 12406 935
rect 10859 889 10866 898
tri 10866 889 10875 898 nw
rect 10859 888 10865 889
tri 10865 888 10866 889 nw
rect 12399 882 12406 901
rect 12347 862 12406 882
rect 12347 857 12366 862
tri 8475 817 8480 822 ne
rect 8480 817 8541 822
tri 8541 817 8546 822 sw
tri 8480 815 8482 817 ne
rect 8482 815 8546 817
tri 314 801 328 815 sw
tri 8482 801 8496 815 ne
rect 8496 801 8546 815
tri 8546 801 8562 817 sw
rect 9554 805 9560 857
rect 9612 805 9624 857
rect 9676 851 10206 857
rect 9685 817 9724 851
rect 9758 817 9797 851
rect 9831 817 9870 851
rect 9904 817 9943 851
rect 9977 817 10016 851
rect 10050 817 10088 851
rect 10122 817 10160 851
rect 10194 817 10206 851
rect 9676 811 10206 817
rect 10679 835 11465 841
rect 9676 805 9682 811
tri 9682 805 9688 811 nw
rect 10679 801 10691 835
rect 10725 801 10763 835
rect 10797 801 11309 835
rect 11343 801 11381 835
rect 11415 801 11465 835
rect 262 799 328 801
tri 328 799 330 801 sw
tri 8496 799 8498 801 ne
rect 8498 799 8562 801
tri 8562 799 8564 801 sw
rect 262 790 330 799
tri 330 790 339 799 sw
tri 8498 790 8507 799 ne
rect 8507 790 8564 799
rect 262 770 992 790
rect 1044 770 1061 790
rect 262 664 621 770
rect 1113 738 1130 790
rect 1182 738 1199 790
rect 1251 738 1268 790
rect 1320 738 1337 790
rect 1389 738 1405 790
rect 1457 738 1473 790
rect 1525 788 8309 790
tri 8309 788 8311 790 sw
tri 8507 788 8509 790 ne
rect 8509 788 8564 790
tri 8564 788 8575 799 sw
rect 10679 795 11465 801
tri 11453 789 11459 795 ne
rect 11459 789 11465 795
rect 11517 789 11529 841
rect 11581 789 11587 841
rect 1525 754 8311 788
tri 8311 754 8345 788 sw
tri 8509 756 8541 788 ne
rect 8541 756 8575 788
tri 8575 756 8607 788 sw
rect 12111 787 12117 839
rect 12169 787 12181 839
rect 12233 833 12301 839
rect 12233 799 12255 833
rect 12289 799 12301 833
rect 12233 793 12301 799
rect 12400 828 12406 862
rect 12399 805 12406 828
rect 12233 788 12240 793
tri 12240 788 12245 793 nw
rect 12347 788 12406 805
rect 12233 787 12239 788
tri 12239 787 12240 788 nw
rect 12347 780 12366 788
tri 8541 754 8543 756 ne
rect 8543 754 8607 756
tri 8607 754 8609 756 sw
rect 12400 754 12406 788
rect 1525 738 8345 754
rect 1087 733 8345 738
tri 8345 733 8366 754 sw
tri 8543 736 8561 754 ne
rect 8561 736 8609 754
tri 8609 736 8627 754 sw
tri 10861 736 10863 738 se
rect 10863 736 10869 738
tri 8561 733 8564 736 ne
rect 8564 733 9812 736
rect 1087 730 8366 733
tri 8366 730 8369 733 sw
tri 8564 730 8567 733 ne
rect 8567 730 9812 733
rect 1087 727 8369 730
tri 8369 727 8372 730 sw
tri 8567 727 8570 730 ne
rect 8570 727 9812 730
rect 1087 696 8372 727
tri 8372 696 8403 727 sw
tri 8570 696 8601 727 ne
rect 8601 696 9812 727
rect 262 644 992 664
rect 1044 644 1061 664
rect 1113 644 1130 696
rect 1182 644 1199 696
rect 1251 644 1268 696
rect 1320 644 1337 696
rect 1389 644 1405 696
rect 1457 644 1473 696
rect 1525 692 8403 696
tri 8403 692 8407 696 sw
tri 8601 692 8605 696 ne
rect 8605 692 9812 696
rect 1525 680 8407 692
tri 8407 680 8419 692 sw
tri 8605 690 8607 692 ne
rect 8607 690 9812 692
tri 9800 684 9806 690 ne
rect 9806 684 9812 690
rect 9864 684 9876 736
rect 9928 730 10697 736
rect 9928 696 10472 730
rect 10506 696 10561 730
rect 10595 696 10651 730
rect 10685 696 10697 730
rect 9928 690 10697 696
rect 10854 726 10869 736
rect 10854 692 10866 726
rect 9928 686 9936 690
tri 9936 686 9940 690 nw
rect 10854 686 10869 692
rect 10921 686 10933 738
rect 10985 686 10991 738
rect 9928 684 9934 686
tri 9934 684 9936 686 nw
rect 11022 684 11028 736
rect 11080 684 11092 736
rect 11144 730 11266 736
rect 11145 696 11220 730
rect 11254 696 11266 730
rect 12399 728 12406 754
tri 12337 714 12347 724 se
rect 12347 714 12406 728
rect 11144 684 11266 696
tri 12307 684 12337 714 se
rect 12337 684 12366 714
tri 12303 680 12307 684 se
rect 12307 680 12366 684
rect 12400 680 12406 714
rect 1525 668 8419 680
tri 8419 668 8431 680 sw
tri 12291 668 12303 680 se
rect 12303 668 12406 680
rect 1525 656 8431 668
tri 8431 656 8443 668 sw
tri 12279 656 12291 668 se
rect 12291 656 12406 668
rect 1525 644 10644 656
rect 262 415 314 644
tri 314 619 339 644 nw
tri 8325 619 8350 644 ne
rect 8350 619 10644 644
tri 8350 610 8359 619 ne
rect 8359 610 10644 619
tri 12271 648 12279 656 se
rect 12279 648 12406 656
rect 12271 642 12406 648
tri 8359 576 8393 610 ne
rect 8393 576 10206 610
rect 10240 576 10278 610
rect 10312 576 10526 610
rect 10560 576 10598 610
rect 10632 576 10644 610
tri 8393 570 8399 576 ne
rect 8399 570 10644 576
rect 11014 610 11738 616
rect 11014 576 11026 610
rect 11060 576 11098 610
rect 11132 576 11308 610
rect 11342 576 11380 610
rect 11414 576 11620 610
rect 11654 576 11692 610
rect 11726 576 11738 610
rect 11014 570 11738 576
rect 12271 610 12323 642
tri 12323 610 12355 642 nw
rect 10358 520 11333 526
tri 11333 520 11339 526 sw
rect 11451 520 11465 532
rect 10358 486 10370 520
rect 10404 486 10442 520
rect 10476 486 10682 520
rect 10716 486 10754 520
rect 10788 486 10875 520
rect 10909 486 10947 520
rect 10981 486 11183 520
rect 11217 486 11255 520
rect 11289 490 11339 520
tri 11339 490 11369 520 sw
rect 11289 486 11369 490
tri 11369 486 11373 490 sw
rect 11451 486 11463 520
rect 10358 480 11373 486
tri 11373 480 11379 486 sw
rect 11451 480 11465 486
rect 11517 480 11529 532
rect 11581 480 11587 532
tri 11313 476 11317 480 ne
rect 11317 476 11379 480
tri 11379 476 11383 480 sw
tri 11317 424 11369 476 ne
rect 11369 452 11383 476
tri 11383 452 11407 476 sw
tri 12087 452 12111 476 se
rect 12111 452 12117 476
rect 11369 424 12117 452
rect 12169 424 12181 476
rect 12233 424 12239 476
tri 314 415 316 417 sw
rect 12271 415 12321 610
tri 12321 608 12323 610 nw
rect 12359 592 12427 598
rect 12359 540 12363 592
rect 12415 540 12427 592
rect 12545 571 12597 1084
rect 12694 1087 12700 1121
rect 12734 1087 12740 1121
tri 12768 1096 12805 1133 ne
rect 12805 1096 12817 1133
rect 12694 1074 12740 1087
tri 12805 1084 12817 1096 ne
rect 12886 1415 13216 1421
rect 12886 1363 12887 1415
rect 12939 1363 12956 1415
rect 13008 1363 13025 1415
rect 13077 1363 13094 1415
rect 13146 1363 13163 1415
rect 13215 1363 13216 1415
rect 12886 1345 13216 1363
rect 12886 1293 12887 1345
rect 12939 1293 12956 1345
rect 13008 1293 13025 1345
rect 13077 1293 13094 1345
rect 13146 1293 13163 1345
rect 13215 1293 13216 1345
rect 12886 1275 13216 1293
rect 12886 1223 12887 1275
rect 12939 1223 12956 1275
rect 13008 1223 13025 1275
rect 13077 1223 13094 1275
rect 13146 1223 13163 1275
rect 13215 1223 13216 1275
rect 12886 1204 13216 1223
rect 12886 1152 12887 1204
rect 12939 1152 12956 1204
rect 13008 1152 13025 1204
rect 13077 1152 13094 1204
rect 13146 1152 13163 1204
rect 13215 1152 13216 1204
rect 12886 1133 13216 1152
rect 14697 1137 15008 1369
rect 12886 1081 12887 1133
rect 12939 1081 12956 1133
rect 13008 1081 13025 1133
rect 13077 1081 13094 1133
rect 13146 1081 13163 1133
rect 13215 1081 13216 1133
rect 12886 1075 13216 1081
rect 12657 1044 12859 1074
rect 12657 1010 12700 1044
rect 12734 1010 12859 1044
rect 12657 1003 12859 1010
tri 12859 1003 12930 1074 nw
rect 12657 967 12832 1003
tri 12832 976 12859 1003 nw
rect 14823 997 14875 1003
rect 12657 933 12700 967
rect 12734 933 12832 967
rect 12657 889 12832 933
rect 12657 855 12700 889
rect 12734 855 12832 889
rect 14823 931 14875 945
rect 14823 873 14875 879
rect 12657 811 12832 855
tri 12636 790 12657 811 se
rect 12657 790 12700 811
rect 12636 777 12700 790
rect 12734 777 12832 811
rect 12636 733 12832 777
rect 12636 699 12700 733
rect 12734 699 12832 733
rect 12636 644 12832 699
tri 12752 610 12786 644 ne
tri 12545 540 12576 571 ne
rect 12576 540 12597 571
tri 12597 540 12650 593 sw
rect 12359 528 12427 540
rect 12359 476 12363 528
rect 12415 476 12427 528
tri 12576 519 12597 540 ne
rect 12597 519 12675 540
tri 12597 488 12628 519 ne
rect 12628 516 12675 519
tri 12675 516 12699 540 sw
tri 14711 516 14735 540 se
rect 14735 516 14753 540
rect 12628 488 14753 516
rect 14805 488 14817 540
rect 14869 488 14875 540
rect 12359 472 12427 476
tri 12427 472 12439 484 sw
rect 12359 470 12439 472
tri 12359 423 12406 470 ne
rect 12406 423 12439 470
tri 12439 423 12488 472 sw
tri 12321 415 12329 423 sw
tri 12406 415 12414 423 ne
rect 12414 415 12488 423
tri 12488 415 12496 423 sw
rect 262 392 316 415
tri 316 392 339 415 sw
tri 12248 392 12271 415 se
rect 12271 392 12329 415
rect 262 389 339 392
tri 339 389 342 392 sw
tri 12245 389 12248 392 se
rect 12248 389 12329 392
tri 12329 389 12355 415 sw
tri 12414 390 12439 415 ne
rect 12439 389 12496 415
tri 12496 389 12522 415 sw
rect 262 343 784 389
rect 12439 355 12522 389
tri 12522 355 12556 389 sw
rect 262 340 323 343
tri 323 340 326 343 nw
tri 12412 307 12439 334 se
rect 12439 307 12556 355
tri 12406 301 12412 307 se
rect 12412 301 12434 307
rect 12428 255 12434 301
rect 12486 255 12498 307
rect 12550 255 12556 307
rect 14840 260 15007 416
<< rmetal1 >>
rect 5836 4254 5838 4255
rect 5836 4210 5837 4254
rect 5836 4209 5838 4210
rect 5874 4254 5876 4255
rect 5875 4210 5876 4254
rect 5874 4209 5876 4210
rect 9296 3894 9298 3895
rect 9334 3894 9336 3895
rect 9296 3844 9297 3894
rect 9335 3844 9336 3894
rect 9296 3843 9298 3844
rect 9334 3843 9336 3844
rect 7726 3810 7728 3811
rect 4180 3728 4182 3729
rect 4218 3728 4220 3729
rect 4180 3684 4181 3728
rect 4219 3684 4220 3728
rect 4180 3683 4182 3684
rect 4218 3683 4220 3684
rect 7726 3684 7727 3810
rect 7726 3683 7728 3684
rect 7764 3810 7766 3811
rect 7765 3684 7766 3810
rect 7764 3683 7766 3684
rect 8014 3347 8144 3348
rect 8014 3346 8015 3347
rect 8143 3346 8144 3347
rect 8014 3309 8015 3310
rect 8143 3309 8144 3310
rect 8014 3308 8144 3309
rect 8330 3196 8460 3197
rect 8330 3195 8331 3196
rect 8459 3195 8460 3196
rect 8330 3158 8331 3159
rect 8459 3158 8460 3159
rect 8330 3157 8460 3158
rect 9137 2899 9139 2900
rect 9175 2899 9177 2900
rect 9137 2849 9138 2899
rect 9176 2849 9177 2899
rect 9137 2848 9139 2849
rect 9175 2848 9177 2849
rect 10509 2819 10511 2820
rect 10509 2769 10510 2819
rect 10509 2768 10511 2769
rect 10547 2819 10549 2820
rect 10548 2769 10549 2819
rect 10547 2768 10549 2769
rect 10377 2742 10429 2743
rect 10377 2741 10378 2742
rect 10428 2741 10429 2742
rect 10377 2704 10378 2705
rect 10428 2704 10429 2705
rect 10377 2703 10429 2704
rect 10311 2677 10313 2678
rect 10349 2677 10351 2678
rect 10311 2627 10312 2677
rect 10350 2627 10351 2677
rect 10311 2626 10313 2627
rect 10349 2626 10351 2627
rect 8993 2580 9493 2581
rect 8993 2579 8994 2580
rect 9492 2579 9493 2580
rect 8993 2542 8994 2543
rect 9492 2542 9493 2543
rect 8993 2541 9493 2542
rect 10777 2586 10829 2587
rect 10777 2585 10778 2586
rect 10828 2585 10829 2586
rect 10777 2548 10778 2549
rect 10828 2548 10829 2549
rect 10777 2547 10829 2548
rect 10374 2521 10376 2522
rect 10412 2521 10414 2522
rect 10374 2471 10375 2521
rect 10413 2471 10414 2521
rect 10374 2470 10376 2471
rect 10412 2470 10414 2471
rect 10523 1568 10575 1569
rect 10523 1567 10524 1568
rect 10574 1567 10575 1568
rect 10523 1530 10524 1531
rect 10574 1530 10575 1531
rect 10523 1529 10575 1530
<< via1 >>
rect 1468 6996 1520 7005
rect 1468 6962 1474 6996
rect 1474 6962 1508 6996
rect 1508 6962 1520 6996
rect 1468 6953 1520 6962
rect 1534 6996 1586 7005
rect 1534 6962 1546 6996
rect 1546 6962 1580 6996
rect 1580 6962 1586 6996
rect 1534 6953 1586 6962
rect 7277 6574 7329 6626
rect 7341 6574 7393 6626
rect 9428 6574 9480 6626
rect 9492 6574 9544 6626
rect 14736 6382 14788 6434
rect 14736 6318 14788 6370
rect 12604 5875 12656 5927
rect 12668 5875 12720 5927
rect -370 5573 -318 5625
rect 11685 5626 11737 5678
rect 11749 5626 11801 5678
rect 12949 5626 13001 5678
rect 13013 5626 13065 5678
rect -370 5509 -318 5561
rect 6876 5546 6928 5598
rect 6940 5546 6992 5598
rect 12200 5546 12252 5598
rect 12264 5546 12316 5598
rect -194 5440 -142 5492
rect -194 5354 -142 5406
rect -18 5446 34 5498
rect -18 5374 34 5426
rect 9428 5428 9480 5480
rect 9492 5428 9544 5480
rect 11573 5428 11625 5480
rect 11637 5428 11689 5480
rect 12079 5443 12131 5495
rect 12143 5443 12195 5495
rect 721 5280 773 5332
rect 785 5280 837 5332
rect 6876 5274 6928 5326
rect 6940 5274 6992 5326
rect 12200 5346 12252 5398
rect 12264 5346 12316 5398
rect 9441 5266 9493 5318
rect 9505 5266 9557 5318
rect 5228 5187 5280 5239
rect 5228 5123 5280 5175
rect 7411 5166 7463 5218
rect 7411 5102 7463 5154
rect 13341 4939 13393 4991
rect 13413 4939 13465 4991
rect 13484 4939 13536 4991
rect 13555 4939 13607 4991
rect 13626 4939 13678 4991
rect 829 4858 881 4910
rect 894 4858 946 4910
rect 959 4858 1011 4910
rect 1024 4858 1076 4910
rect 1089 4858 1141 4910
rect 1153 4858 1205 4910
rect 1217 4858 1269 4910
rect 1281 4858 1333 4910
rect 1345 4858 1397 4910
rect 1409 4858 1461 4910
rect 1473 4858 1525 4910
rect 829 4783 881 4835
rect 894 4783 946 4835
rect 959 4783 1011 4835
rect 1024 4783 1076 4835
rect 1089 4783 1141 4835
rect 1153 4783 1205 4835
rect 1217 4783 1269 4835
rect 1281 4783 1333 4835
rect 1345 4783 1397 4835
rect 1409 4783 1461 4835
rect 1473 4783 1525 4835
rect 829 4708 881 4760
rect 894 4708 946 4760
rect 959 4708 1011 4760
rect 1024 4708 1076 4760
rect 1089 4708 1141 4760
rect 1153 4708 1205 4760
rect 1217 4708 1269 4760
rect 1281 4708 1333 4760
rect 1345 4708 1397 4760
rect 1409 4708 1461 4760
rect 1473 4708 1525 4760
rect 12347 4852 12399 4904
rect 12347 4783 12399 4835
rect 12347 4714 12399 4766
rect 13341 4864 13393 4916
rect 13413 4864 13465 4916
rect 13484 4864 13536 4916
rect 13555 4864 13607 4916
rect 13626 4864 13678 4916
rect 13341 4789 13393 4841
rect 13413 4789 13465 4841
rect 13484 4789 13536 4841
rect 13555 4789 13607 4841
rect 13626 4789 13678 4841
rect -282 4636 -230 4688
rect -218 4636 -166 4688
rect 9936 4626 9988 4678
rect 10000 4626 10052 4678
rect 10190 4626 10242 4678
rect 10254 4626 10306 4678
rect -463 4554 -411 4606
rect -463 4490 -411 4542
rect 3628 4534 3680 4586
rect 3692 4534 3744 4586
rect 11621 4544 11673 4596
rect 11685 4544 11737 4596
rect 12159 4585 12211 4637
rect 12224 4585 12276 4637
rect 14690 4585 14742 4637
rect 14754 4585 14806 4637
rect 14591 4505 14643 4557
rect 14655 4505 14707 4557
rect 829 4460 881 4505
rect -103 4391 -51 4443
rect 829 4453 841 4460
rect 841 4453 875 4460
rect 875 4453 881 4460
rect 894 4460 946 4505
rect 959 4460 1011 4505
rect 1024 4460 1076 4505
rect 1089 4460 1141 4505
rect 1153 4460 1205 4505
rect 1217 4460 1269 4505
rect 1281 4460 1333 4505
rect 894 4453 913 4460
rect 913 4453 946 4460
rect 959 4453 985 4460
rect 985 4453 1011 4460
rect 1024 4453 1057 4460
rect 1057 4453 1076 4460
rect 1089 4453 1091 4460
rect 1091 4453 1129 4460
rect 1129 4453 1141 4460
rect 1153 4453 1163 4460
rect 1163 4453 1201 4460
rect 1201 4453 1205 4460
rect 1217 4453 1235 4460
rect 1235 4453 1269 4460
rect 1281 4453 1307 4460
rect 1307 4453 1333 4460
rect 1345 4460 1397 4505
rect 1345 4453 1379 4460
rect 1379 4453 1397 4460
rect 1409 4460 1461 4505
rect 1409 4453 1417 4460
rect 1417 4453 1451 4460
rect 1451 4453 1461 4460
rect 1473 4460 1525 4505
rect 1473 4453 1489 4460
rect 1489 4453 1523 4460
rect 1523 4453 1525 4460
rect 829 4426 841 4433
rect 841 4426 875 4433
rect 875 4426 881 4433
rect 829 4381 881 4426
rect 894 4426 913 4433
rect 913 4426 946 4433
rect 959 4426 985 4433
rect 985 4426 1011 4433
rect 1024 4426 1057 4433
rect 1057 4426 1076 4433
rect 1089 4426 1091 4433
rect 1091 4426 1129 4433
rect 1129 4426 1141 4433
rect 1153 4426 1163 4433
rect 1163 4426 1201 4433
rect 1201 4426 1205 4433
rect 1217 4426 1235 4433
rect 1235 4426 1269 4433
rect 1281 4426 1307 4433
rect 1307 4426 1333 4433
rect 894 4381 946 4426
rect 959 4381 1011 4426
rect 1024 4381 1076 4426
rect 1089 4381 1141 4426
rect 1153 4381 1205 4426
rect 1217 4381 1269 4426
rect 1281 4381 1333 4426
rect 1345 4426 1379 4433
rect 1379 4426 1397 4433
rect 1345 4381 1397 4426
rect 1409 4426 1417 4433
rect 1417 4426 1451 4433
rect 1451 4426 1461 4433
rect 1409 4381 1461 4426
rect 1473 4426 1489 4433
rect 1489 4426 1523 4433
rect 1523 4426 1525 4433
rect 1473 4381 1525 4426
rect 12347 4381 12368 4415
rect 12368 4381 12399 4415
rect -103 4325 -51 4377
rect 12347 4363 12399 4381
rect 12347 4340 12399 4350
rect -187 4222 -135 4274
rect 2103 4255 2155 4261
rect 2167 4255 2219 4261
rect -187 4158 -135 4210
rect 2103 4221 2107 4255
rect 2107 4221 2149 4255
rect 2149 4221 2155 4255
rect 2167 4221 2183 4255
rect 2183 4221 2219 4255
rect 2103 4209 2155 4221
rect 2167 4209 2219 4221
rect 2453 4255 2505 4261
rect 2517 4255 2569 4261
rect 2453 4221 2454 4255
rect 2454 4221 2497 4255
rect 2497 4221 2505 4255
rect 2517 4221 2531 4255
rect 2531 4221 2569 4255
rect 2453 4209 2505 4221
rect 2517 4209 2569 4221
rect 2619 4209 2671 4261
rect 2683 4209 2735 4261
rect 5178 4212 5230 4264
rect 5242 4212 5294 4264
rect 12233 4261 12285 4313
rect 7210 4249 7262 4261
rect 7274 4249 7326 4261
rect 7210 4215 7245 4249
rect 7245 4215 7262 4249
rect 7274 4215 7279 4249
rect 7279 4215 7326 4249
rect 7210 4209 7262 4215
rect 7274 4209 7326 4215
rect 7602 4251 7654 4261
rect 7602 4217 7612 4251
rect 7612 4217 7654 4251
rect 7602 4209 7654 4217
rect 7666 4209 7718 4261
rect 7758 4209 7810 4261
rect 7822 4251 7874 4261
rect 7822 4217 7826 4251
rect 7826 4217 7860 4251
rect 7860 4217 7874 4251
rect 7822 4209 7874 4217
rect 10837 4201 10889 4253
rect 238 4134 290 4140
rect -645 4108 -593 4116
rect -545 4108 -493 4116
rect -645 4074 -638 4108
rect -638 4074 -604 4108
rect -604 4074 -593 4108
rect -545 4074 -532 4108
rect -532 4074 -493 4108
rect -645 4064 -593 4074
rect -545 4064 -493 4074
rect -645 4031 -593 4039
rect -545 4031 -493 4039
rect -645 3997 -638 4031
rect -638 3997 -604 4031
rect -604 3997 -593 4031
rect -545 3997 -532 4031
rect -532 3997 -493 4031
rect -645 3987 -593 3997
rect -545 3987 -493 3997
rect -645 3954 -593 3962
rect -545 3954 -493 3962
rect -645 3920 -638 3954
rect -638 3920 -604 3954
rect -604 3920 -593 3954
rect -545 3920 -532 3954
rect -532 3920 -493 3954
rect -645 3910 -593 3920
rect -545 3910 -493 3920
rect -645 3876 -593 3885
rect -545 3876 -493 3885
rect -645 3842 -638 3876
rect -638 3842 -604 3876
rect -604 3842 -593 3876
rect -545 3842 -532 3876
rect -532 3842 -493 3876
rect -645 3833 -593 3842
rect -545 3833 -493 3842
rect -645 3798 -593 3808
rect -545 3798 -493 3808
rect -645 3764 -638 3798
rect -638 3764 -604 3798
rect -604 3764 -593 3798
rect -545 3764 -532 3798
rect -532 3764 -493 3798
rect -645 3756 -593 3764
rect -545 3756 -493 3764
rect 238 4100 271 4134
rect 271 4100 290 4134
rect 238 4088 290 4100
rect 238 4054 290 4061
rect 238 4020 271 4054
rect 271 4020 290 4054
rect 238 4009 290 4020
rect 1704 4129 1756 4181
rect 1773 4129 1825 4181
rect 1842 4129 1894 4181
rect 1911 4129 1963 4181
rect 1980 4129 2032 4181
rect 3156 4129 3208 4181
rect 3220 4129 3272 4181
rect 3284 4129 3336 4181
rect 3348 4129 3400 4181
rect 3412 4129 3464 4181
rect 3476 4129 3528 4181
rect 3540 4129 3592 4181
rect 1704 4054 1756 4106
rect 1773 4054 1825 4106
rect 1842 4054 1894 4106
rect 1911 4054 1963 4106
rect 1980 4054 2032 4106
rect 3156 4054 3208 4106
rect 3220 4054 3272 4106
rect 3284 4054 3336 4106
rect 3348 4054 3400 4106
rect 3412 4054 3464 4106
rect 3476 4054 3528 4106
rect 3540 4054 3592 4106
rect 238 3974 290 3982
rect 1704 3979 1756 4031
rect 1773 3979 1825 4031
rect 1842 3979 1894 4031
rect 1911 3979 1963 4031
rect 1980 3979 2032 4031
rect 3156 3979 3208 4031
rect 3220 3979 3272 4031
rect 3284 3979 3336 4031
rect 3348 3979 3400 4031
rect 3412 3979 3464 4031
rect 3476 3979 3528 4031
rect 3540 3979 3592 4031
rect 9147 4142 9199 4152
rect 9147 4108 9179 4142
rect 9179 4108 9199 4142
rect 9147 4100 9199 4108
rect 9214 4100 9266 4152
rect 9280 4100 9332 4152
rect 10837 4137 10889 4189
rect 12233 4197 12285 4249
rect 12347 4306 12368 4340
rect 12368 4306 12399 4340
rect 12347 4298 12399 4306
rect 12347 4265 12399 4285
rect 12347 4233 12368 4265
rect 12368 4233 12399 4265
rect 9147 4046 9199 4054
rect 9147 4012 9179 4046
rect 9179 4012 9199 4046
rect 9147 4002 9199 4012
rect 9214 4002 9266 4054
rect 9280 4002 9332 4054
rect 11000 4075 11028 4109
rect 11028 4075 11052 4109
rect 11000 4057 11052 4075
rect 238 3940 271 3974
rect 271 3940 290 3974
rect 11000 3993 11052 4045
rect 11886 3983 11938 3986
rect 238 3930 290 3940
rect 238 3893 290 3903
rect 238 3859 271 3893
rect 271 3859 290 3893
rect 829 3871 881 3923
rect 902 3871 954 3923
rect 974 3871 1026 3923
rect 1046 3871 1098 3923
rect 1118 3871 1170 3923
rect 1190 3871 1242 3923
rect 2619 3899 2671 3951
rect 2683 3899 2735 3951
rect 8037 3899 8089 3951
rect 8101 3899 8153 3951
rect 238 3851 290 3859
rect 238 3812 290 3824
rect 2453 3819 2505 3871
rect 2517 3819 2569 3871
rect 9126 3843 9178 3895
rect 9190 3843 9242 3895
rect 9371 3843 9423 3895
rect 9435 3843 9487 3895
rect 10001 3893 10053 3945
rect 11886 3949 11913 3983
rect 11913 3949 11938 3983
rect 11886 3934 11938 3949
rect 10001 3829 10053 3881
rect 11886 3870 11938 3922
rect 238 3778 271 3812
rect 271 3778 290 3812
rect 238 3772 290 3778
rect 2871 3739 2923 3791
rect 2935 3739 2987 3791
rect 3832 3757 3884 3809
rect 3896 3757 3948 3809
rect -463 3656 -411 3708
rect 2103 3723 2155 3735
rect 2167 3723 2219 3735
rect 2103 3689 2122 3723
rect 2122 3689 2155 3723
rect 2167 3689 2194 3723
rect 2194 3689 2219 3723
rect 2103 3683 2155 3689
rect 2167 3683 2219 3689
rect 6753 3714 6805 3766
rect 6817 3714 6869 3766
rect 7672 3753 7724 3805
rect 7672 3689 7724 3741
rect 9282 3763 9334 3815
rect 9346 3763 9398 3815
rect 12347 4190 12399 4220
rect 12347 4168 12368 4190
rect 12368 4168 12399 4190
rect 12347 4115 12399 4155
rect 12347 4103 12368 4115
rect 12368 4103 12399 4115
rect 12347 4081 12368 4090
rect 12368 4081 12399 4090
rect 12347 4040 12399 4081
rect 12347 4038 12368 4040
rect 12368 4038 12399 4040
rect 12347 4006 12368 4025
rect 12368 4006 12399 4025
rect 12347 3973 12399 4006
rect 12347 3931 12368 3959
rect 12368 3931 12399 3959
rect 12347 3907 12399 3931
rect 12347 3890 12399 3893
rect 12347 3856 12368 3890
rect 12368 3856 12399 3890
rect 12347 3841 12399 3856
rect 12347 3815 12399 3827
rect 12347 3781 12368 3815
rect 12368 3781 12399 3815
rect 12347 3775 12399 3781
rect 9371 3683 9423 3735
rect 9435 3683 9487 3735
rect 9593 3723 9645 3735
rect 9593 3689 9599 3723
rect 9599 3689 9633 3723
rect 9633 3689 9645 3723
rect 9593 3683 9645 3689
rect 9659 3723 9711 3735
rect 9659 3689 9671 3723
rect 9671 3689 9705 3723
rect 9705 3689 9711 3723
rect 9659 3683 9711 3689
rect -463 3590 -411 3642
rect -103 3588 -101 3622
rect -101 3588 -67 3622
rect -67 3588 -51 3622
rect -103 3570 -51 3588
rect -103 3550 -51 3558
rect -103 3516 -101 3550
rect -101 3516 -67 3550
rect -67 3516 -51 3550
rect 139 3591 191 3643
rect 139 3527 191 3579
rect -103 3506 -51 3516
rect -465 3392 -413 3444
rect -465 3328 -413 3380
rect 121 3395 173 3401
rect 121 3361 129 3395
rect 129 3361 163 3395
rect 163 3361 173 3395
rect 121 3349 173 3361
rect 121 3323 173 3335
rect 121 3289 129 3323
rect 129 3289 163 3323
rect 163 3289 173 3323
rect 947 3602 999 3654
rect 1013 3643 1065 3654
rect 1013 3609 1016 3643
rect 1016 3609 1050 3643
rect 1050 3609 1065 3643
rect 1013 3602 1065 3609
rect 1079 3602 1131 3654
rect 1145 3602 1197 3654
rect 1211 3602 1263 3654
rect 1277 3643 1329 3654
rect 1277 3609 1304 3643
rect 1304 3609 1329 3643
rect 1277 3602 1329 3609
rect 1343 3602 1395 3654
rect 1408 3602 1460 3654
rect 1473 3602 1525 3654
rect 947 3528 999 3580
rect 1013 3571 1065 3580
rect 1013 3537 1016 3571
rect 1016 3537 1050 3571
rect 1050 3537 1065 3571
rect 1013 3528 1065 3537
rect 1079 3528 1131 3580
rect 1145 3528 1197 3580
rect 1211 3528 1263 3580
rect 1277 3571 1329 3580
rect 1277 3537 1304 3571
rect 1304 3537 1329 3571
rect 1277 3528 1329 3537
rect 1343 3528 1395 3580
rect 1408 3528 1460 3580
rect 1473 3528 1525 3580
rect 947 3454 999 3506
rect 1013 3499 1065 3506
rect 1013 3465 1016 3499
rect 1016 3465 1050 3499
rect 1050 3465 1065 3499
rect 1013 3454 1065 3465
rect 1079 3454 1131 3506
rect 1145 3454 1197 3506
rect 1211 3454 1263 3506
rect 1277 3499 1329 3506
rect 1277 3465 1304 3499
rect 1304 3465 1329 3499
rect 1277 3454 1329 3465
rect 1343 3454 1395 3506
rect 1408 3454 1460 3506
rect 1473 3454 1525 3506
rect 8923 3597 8975 3649
rect 9027 3597 9079 3649
rect 12347 3643 12399 3649
rect 12347 3609 12366 3643
rect 12366 3609 12399 3643
rect 12347 3597 12399 3609
rect 8923 3528 8975 3580
rect 9027 3528 9079 3580
rect 12347 3571 12399 3580
rect 12347 3537 12366 3571
rect 12366 3537 12399 3571
rect 13338 3652 13390 3704
rect 13411 3652 13463 3704
rect 13484 3652 13536 3704
rect 13557 3652 13609 3704
rect 13630 3652 13682 3704
rect 13338 3586 13390 3638
rect 13411 3586 13463 3638
rect 13484 3586 13536 3638
rect 13557 3586 13609 3638
rect 13630 3586 13682 3638
rect 12347 3528 12399 3537
rect 8923 3459 8975 3511
rect 9027 3459 9079 3511
rect 12347 3499 12399 3511
rect 12887 3508 12939 3560
rect 12956 3508 13008 3560
rect 13025 3508 13077 3560
rect 13094 3508 13146 3560
rect 13163 3508 13215 3560
rect 12347 3465 12366 3499
rect 12366 3465 12399 3499
rect 12347 3459 12399 3465
rect 8422 3373 8474 3425
rect 8486 3373 8538 3425
rect 9582 3373 9634 3425
rect 9646 3373 9698 3425
rect 9818 3369 9870 3421
rect 9882 3369 9934 3421
rect 121 3283 173 3289
rect 2373 3240 2425 3292
rect 2437 3240 2489 3292
rect 7005 3240 7057 3292
rect 7069 3240 7121 3292
rect 8989 3292 9041 3344
rect 9053 3292 9105 3344
rect 12233 3346 12285 3398
rect 12233 3282 12285 3334
rect 12347 3390 12399 3396
rect 12347 3356 12366 3390
rect 12366 3356 12399 3390
rect 12347 3344 12399 3356
rect 12347 3318 12399 3332
rect 12347 3284 12366 3318
rect 12366 3284 12399 3318
rect 12887 3438 12939 3490
rect 12956 3438 13008 3490
rect 13025 3438 13077 3490
rect 13094 3438 13146 3490
rect 13163 3438 13215 3490
rect 12887 3368 12939 3420
rect 12956 3368 13008 3420
rect 13025 3368 13077 3420
rect 13094 3368 13146 3420
rect 13163 3368 13215 3420
rect 12347 3280 12399 3284
rect 2120 3160 2172 3212
rect 2184 3160 2236 3212
rect 6985 3160 7037 3212
rect 7049 3160 7101 3212
rect 7210 3176 7262 3228
rect 7274 3176 7326 3228
rect 9890 3194 9942 3246
rect 12347 3246 12399 3268
rect 10625 3185 10677 3237
rect 10689 3185 10741 3237
rect 11006 3185 11058 3237
rect 11070 3225 11122 3237
rect 11070 3191 11104 3225
rect 11104 3191 11122 3225
rect 11070 3185 11122 3191
rect 238 3074 290 3126
rect 238 3002 290 3054
rect 238 2930 290 2982
rect 238 2857 290 2909
rect 238 2784 290 2836
rect 7758 3126 7810 3138
rect 7758 3092 7762 3126
rect 7762 3092 7796 3126
rect 7796 3092 7810 3126
rect 7758 3086 7810 3092
rect 7822 3126 7874 3138
rect 7822 3092 7834 3126
rect 7834 3092 7868 3126
rect 7868 3092 7874 3126
rect 7822 3086 7874 3092
rect 8679 3126 8731 3138
rect 8743 3126 8795 3138
rect 8679 3092 8711 3126
rect 8711 3092 8731 3126
rect 8743 3092 8745 3126
rect 8745 3092 8783 3126
rect 8783 3092 8795 3126
rect 9890 3130 9942 3182
rect 12235 3175 12287 3227
rect 12235 3111 12287 3163
rect 12347 3216 12366 3246
rect 12366 3216 12399 3246
rect 12887 3297 12939 3349
rect 12956 3297 13008 3349
rect 13025 3297 13077 3349
rect 13094 3297 13146 3349
rect 13163 3297 13215 3349
rect 12887 3226 12939 3278
rect 12956 3226 13008 3278
rect 13025 3226 13077 3278
rect 13094 3226 13146 3278
rect 13163 3226 13215 3278
rect 13338 3520 13390 3572
rect 13411 3520 13463 3572
rect 13484 3520 13536 3572
rect 13557 3520 13609 3572
rect 13630 3520 13682 3572
rect 13338 3454 13390 3506
rect 13411 3454 13463 3506
rect 13484 3454 13536 3506
rect 13557 3454 13609 3506
rect 13630 3454 13682 3506
rect 13338 3388 13390 3440
rect 13411 3388 13463 3440
rect 13484 3388 13536 3440
rect 13557 3388 13609 3440
rect 13630 3388 13682 3440
rect 13338 3322 13390 3374
rect 13411 3322 13463 3374
rect 13484 3322 13536 3374
rect 13557 3322 13609 3374
rect 13630 3322 13682 3374
rect 13338 3256 13390 3308
rect 13411 3256 13463 3308
rect 13484 3256 13536 3308
rect 13557 3256 13609 3308
rect 13630 3256 13682 3308
rect 12347 3174 12399 3204
rect 12347 3152 12366 3174
rect 12366 3152 12399 3174
rect 8679 3086 8731 3092
rect 8743 3086 8795 3092
rect 12347 3102 12399 3140
rect 13338 3190 13390 3242
rect 13411 3190 13463 3242
rect 13484 3190 13536 3242
rect 13557 3190 13609 3242
rect 13630 3190 13682 3242
rect 13338 3124 13390 3176
rect 13411 3124 13463 3176
rect 13484 3124 13536 3176
rect 13557 3124 13609 3176
rect 13630 3124 13682 3176
rect 12347 3088 12366 3102
rect 12366 3088 12399 3102
rect 12347 3068 12366 3076
rect 12366 3068 12399 3076
rect 1704 3005 1756 3057
rect 1773 3005 1825 3057
rect 1842 3005 1894 3057
rect 1911 3005 1963 3057
rect 1980 3005 2032 3057
rect 3156 3005 3208 3057
rect 3220 3005 3272 3057
rect 3284 3005 3336 3057
rect 3348 3005 3400 3057
rect 3412 3005 3464 3057
rect 3476 3005 3528 3057
rect 3540 3005 3592 3057
rect 1704 2977 1756 2981
rect 1773 2977 1825 2981
rect 1842 2977 1894 2981
rect 1911 2977 1963 2981
rect 1980 2977 2032 2981
rect 3156 2977 3208 2981
rect 3220 2977 3272 2981
rect 3284 2977 3336 2981
rect 1704 2943 1751 2977
rect 1751 2943 1756 2977
rect 1773 2943 1785 2977
rect 1785 2943 1823 2977
rect 1823 2943 1825 2977
rect 1842 2943 1857 2977
rect 1857 2943 1894 2977
rect 1911 2943 1929 2977
rect 1929 2943 1963 2977
rect 1980 2943 2001 2977
rect 2001 2943 2032 2977
rect 3156 2943 3191 2977
rect 3191 2943 3208 2977
rect 3220 2943 3225 2977
rect 3225 2943 3263 2977
rect 3263 2943 3272 2977
rect 3284 2943 3297 2977
rect 3297 2943 3336 2977
rect 1704 2929 1756 2943
rect 1773 2929 1825 2943
rect 1842 2929 1894 2943
rect 1911 2929 1963 2943
rect 1980 2929 2032 2943
rect 3156 2929 3208 2943
rect 3220 2929 3272 2943
rect 3284 2929 3336 2943
rect 3348 2974 3400 2981
rect 3348 2940 3358 2974
rect 3358 2940 3392 2974
rect 3392 2940 3400 2974
rect 3348 2929 3400 2940
rect 3412 2974 3464 2981
rect 3476 2974 3528 2981
rect 3540 2974 3592 2981
rect 3412 2940 3432 2974
rect 3432 2940 3464 2974
rect 3476 2940 3506 2974
rect 3506 2940 3528 2974
rect 3540 2940 3580 2974
rect 3580 2940 3592 2974
rect 3412 2929 3464 2940
rect 3476 2929 3528 2940
rect 3540 2929 3592 2940
rect 12347 3030 12399 3068
rect 12347 3024 12366 3030
rect 12366 3024 12399 3030
rect 12347 2996 12366 3012
rect 12366 2996 12399 3012
rect 12347 2960 12399 2996
rect 12347 2924 12366 2948
rect 12366 2924 12399 2948
rect 2120 2846 2172 2898
rect 2184 2846 2236 2898
rect 6985 2848 7037 2900
rect 7049 2848 7101 2900
rect 7758 2842 7810 2894
rect 8231 2848 8283 2900
rect 8295 2848 8347 2900
rect 8422 2848 8474 2900
rect 8486 2848 8538 2900
rect 9674 2848 9726 2900
rect 9738 2848 9790 2900
rect 9988 2894 10040 2900
rect 9988 2860 9997 2894
rect 9997 2860 10031 2894
rect 10031 2860 10040 2894
rect 9988 2848 10040 2860
rect 10052 2894 10104 2900
rect 10052 2860 10069 2894
rect 10069 2860 10103 2894
rect 10103 2860 10104 2894
rect 10052 2848 10104 2860
rect 10173 2848 10225 2900
rect 10237 2848 10289 2900
rect 7758 2778 7810 2830
rect 12073 2842 12125 2894
rect 238 2711 290 2763
rect 238 2638 290 2690
rect 4504 2718 4556 2770
rect 4568 2718 4620 2770
rect 12073 2778 12125 2830
rect 12347 2896 12399 2924
rect 12347 2852 12366 2884
rect 12366 2852 12399 2884
rect 12347 2832 12399 2852
rect 12347 2814 12399 2819
rect 12347 2780 12366 2814
rect 12366 2780 12399 2814
rect 7678 2713 7730 2725
rect 7678 2679 7684 2713
rect 7684 2679 7718 2713
rect 7718 2679 7730 2713
rect 7678 2673 7730 2679
rect 7742 2713 7794 2725
rect 7742 2679 7756 2713
rect 7756 2679 7790 2713
rect 7790 2679 7794 2713
rect 7742 2673 7794 2679
rect 238 2565 290 2617
rect 2895 2577 2947 2629
rect 2959 2577 3011 2629
rect 7659 2593 7711 2645
rect 7723 2593 7775 2645
rect -465 2521 -413 2527
rect -465 2487 -453 2521
rect -453 2487 -419 2521
rect -419 2487 -413 2521
rect -465 2475 -413 2487
rect -465 2449 -413 2461
rect -465 2415 -453 2449
rect -453 2415 -419 2449
rect -419 2415 -413 2449
rect -465 2409 -413 2415
rect -187 2478 -135 2530
rect -187 2414 -135 2466
rect 3 2278 55 2330
rect 3 2214 55 2266
rect 8445 2635 8497 2687
rect 9282 2686 9334 2738
rect 9346 2686 9398 2738
rect 12347 2767 12399 2780
rect 12347 2742 12399 2754
rect 12347 2708 12366 2742
rect 12366 2708 12399 2742
rect 12347 2702 12399 2708
rect 9371 2652 9423 2658
rect 8445 2571 8497 2623
rect 9371 2618 9372 2652
rect 9372 2618 9406 2652
rect 9406 2618 9423 2652
rect 9371 2606 9423 2618
rect 9435 2652 9487 2658
rect 9435 2618 9444 2652
rect 9444 2618 9478 2652
rect 9478 2618 9487 2652
rect 9435 2606 9487 2618
rect 9582 2626 9634 2678
rect 9646 2626 9698 2678
rect 8823 2545 8875 2597
rect 8887 2545 8939 2597
rect 10462 2470 10514 2522
rect 10526 2470 10578 2522
rect 10707 2470 10759 2522
rect 10771 2470 10823 2522
rect 10895 2470 10947 2522
rect 10959 2470 11011 2522
rect 11835 2470 11887 2522
rect 11899 2470 11951 2522
rect 12440 2458 12492 2510
rect 807 2385 859 2437
rect 807 2321 859 2373
rect 1704 2390 1756 2442
rect 1773 2390 1825 2442
rect 1842 2390 1894 2442
rect 1911 2390 1963 2442
rect 1980 2390 2032 2442
rect 3156 2390 3208 2442
rect 3220 2390 3272 2442
rect 3284 2390 3336 2442
rect 3348 2390 3400 2442
rect 3412 2390 3464 2442
rect 3476 2390 3528 2442
rect 3540 2390 3592 2442
rect 1704 2312 1756 2364
rect 1773 2312 1825 2364
rect 1842 2312 1894 2364
rect 1911 2312 1963 2364
rect 1980 2312 2032 2364
rect 3156 2312 3208 2364
rect 3220 2312 3272 2364
rect 3284 2312 3336 2364
rect 3348 2312 3400 2364
rect 3412 2312 3464 2364
rect 3476 2312 3528 2364
rect 3540 2312 3592 2364
rect 12347 2413 12399 2419
rect 12347 2379 12366 2413
rect 12366 2379 12399 2413
rect 12440 2394 12492 2446
rect 12347 2367 12399 2379
rect 12347 2337 12399 2354
rect 12347 2303 12366 2337
rect 12366 2303 12399 2337
rect 12347 2302 12399 2303
rect 9443 2232 9495 2284
rect 9507 2232 9559 2284
rect 11852 2226 11904 2278
rect 6753 2154 6805 2206
rect 6817 2154 6869 2206
rect 8898 2152 8950 2204
rect 8962 2152 9014 2204
rect 10566 2152 10618 2204
rect 10630 2152 10682 2204
rect 10882 2151 10934 2203
rect 10946 2151 10998 2203
rect 11397 2135 11449 2187
rect 11852 2162 11904 2214
rect 12347 2261 12399 2289
rect 12347 2237 12366 2261
rect 12366 2237 12399 2261
rect 12347 2185 12399 2223
rect 12347 2171 12366 2185
rect 12366 2171 12399 2185
rect 12347 2151 12366 2157
rect 12366 2151 12399 2157
rect 10468 2072 10520 2124
rect 10532 2072 10584 2124
rect 11397 2064 11449 2116
rect 12347 2109 12399 2151
rect 12347 2105 12366 2109
rect 12366 2105 12399 2109
rect 12347 2075 12366 2091
rect 12366 2075 12399 2091
rect 12347 2039 12399 2075
rect 1704 1977 1756 2029
rect 1773 1977 1825 2029
rect 1842 1977 1894 2029
rect 1911 1977 1963 2029
rect 1980 1977 2032 2029
rect 3156 1977 3208 2029
rect 3220 1977 3272 2029
rect 3284 1977 3336 2029
rect 3348 1977 3400 2029
rect 3412 1977 3464 2029
rect 3476 1977 3528 2029
rect 3540 1977 3592 2029
rect 1704 1903 1756 1955
rect 1773 1903 1825 1955
rect 1842 1903 1894 1955
rect 1911 1903 1963 1955
rect 1980 1903 2032 1955
rect 3156 1903 3208 1955
rect 3220 1903 3272 1955
rect 3284 1903 3336 1955
rect 3348 1903 3400 1955
rect 3412 1903 3464 1955
rect 3476 1903 3528 1955
rect 3540 1903 3592 1955
rect 1704 1829 1756 1881
rect 1773 1829 1825 1881
rect 1842 1829 1894 1881
rect 1911 1829 1963 1881
rect 1980 1829 2032 1881
rect 3156 1829 3208 1881
rect 3220 1829 3272 1881
rect 3284 1829 3336 1881
rect 3348 1829 3400 1881
rect 3412 1829 3464 1881
rect 3476 1829 3528 1881
rect 3540 1829 3592 1881
rect 12347 1999 12366 2025
rect 12366 1999 12399 2025
rect 12347 1973 12399 1999
rect 12347 1957 12399 1959
rect 12347 1923 12366 1957
rect 12366 1923 12399 1957
rect 12347 1907 12399 1923
rect 12347 1881 12399 1893
rect 12347 1847 12366 1881
rect 12366 1847 12399 1881
rect 12347 1841 12399 1847
rect 7301 1713 7353 1765
rect 706 1602 758 1654
rect 706 1538 758 1590
rect 7163 1602 7215 1654
rect 7301 1649 7353 1701
rect 8717 1720 8769 1732
rect 8806 1720 8858 1732
rect 8717 1686 8746 1720
rect 8746 1686 8769 1720
rect 8806 1686 8818 1720
rect 8818 1686 8852 1720
rect 8852 1686 8858 1720
rect 8717 1680 8769 1686
rect 8806 1680 8858 1686
rect 9019 1722 9071 1732
rect 9019 1688 9053 1722
rect 9053 1688 9071 1722
rect 9019 1680 9071 1688
rect 9083 1680 9135 1732
rect 9674 1680 9726 1732
rect 9738 1680 9790 1732
rect 10618 1692 10670 1744
rect 10682 1692 10734 1744
rect 10373 1658 10425 1664
rect 10437 1658 10489 1664
rect 7997 1606 8049 1658
rect 8061 1606 8113 1658
rect 9435 1646 9487 1652
rect 9435 1612 9466 1646
rect 9466 1612 9487 1646
rect 7163 1538 7215 1590
rect 9435 1600 9487 1612
rect 9499 1646 9551 1652
rect 9499 1612 9504 1646
rect 9504 1612 9538 1646
rect 9538 1612 9551 1646
rect 10373 1624 10391 1658
rect 10391 1624 10425 1658
rect 10437 1624 10463 1658
rect 10463 1624 10489 1658
rect 10373 1612 10425 1624
rect 10437 1612 10489 1624
rect 10707 1612 10759 1664
rect 10771 1612 10823 1664
rect 11098 1650 11150 1654
rect 11098 1616 11105 1650
rect 11105 1616 11139 1650
rect 11139 1616 11150 1650
rect 9499 1600 9551 1612
rect 9591 1532 9643 1584
rect 9655 1532 9707 1584
rect 11098 1602 11150 1616
rect 10633 1572 10685 1584
rect 10633 1538 10639 1572
rect 10639 1538 10673 1572
rect 10673 1538 10685 1572
rect 10633 1532 10685 1538
rect 10703 1572 10755 1584
rect 10703 1538 10712 1572
rect 10712 1538 10746 1572
rect 10746 1538 10755 1572
rect 10703 1532 10755 1538
rect 10773 1572 10825 1584
rect 10773 1538 10785 1572
rect 10785 1538 10819 1572
rect 10819 1538 10825 1572
rect 10773 1532 10825 1538
rect 10909 1576 10961 1584
rect 10909 1542 10917 1576
rect 10917 1542 10951 1576
rect 10951 1542 10961 1576
rect 10909 1532 10961 1542
rect 10973 1576 11025 1584
rect 10973 1542 10989 1576
rect 10989 1542 11023 1576
rect 11023 1542 11025 1576
rect 10973 1532 11025 1542
rect 11098 1578 11150 1590
rect 11098 1544 11105 1578
rect 11105 1544 11139 1578
rect 11139 1544 11150 1578
rect 11098 1538 11150 1544
rect 992 1451 1044 1503
rect 1061 1451 1113 1503
rect 1130 1451 1182 1503
rect 1199 1451 1251 1503
rect 1268 1451 1320 1503
rect 1337 1451 1389 1503
rect 1405 1451 1457 1503
rect 1473 1451 1525 1503
rect 12347 1492 12399 1498
rect 12347 1458 12366 1492
rect 12366 1458 12399 1492
rect 12347 1446 12399 1458
rect 992 1377 1044 1429
rect 1061 1377 1113 1429
rect 1130 1377 1182 1429
rect 1199 1377 1251 1429
rect 1268 1377 1320 1429
rect 1337 1377 1389 1429
rect 1405 1377 1457 1429
rect 1473 1377 1525 1429
rect 12347 1420 12399 1429
rect 12347 1386 12366 1420
rect 12366 1386 12399 1420
rect 12347 1377 12399 1386
rect 992 1303 1044 1355
rect 1061 1303 1113 1355
rect 1130 1303 1182 1355
rect 1199 1303 1251 1355
rect 1268 1303 1320 1355
rect 1337 1303 1389 1355
rect 1405 1303 1457 1355
rect 1473 1303 1525 1355
rect 12347 1348 12399 1360
rect 12347 1314 12366 1348
rect 12366 1314 12399 1348
rect 12347 1308 12399 1314
rect 7583 1222 7635 1274
rect 7647 1222 7699 1274
rect 4504 1112 4556 1164
rect 4568 1112 4620 1164
rect 5478 1112 5530 1164
rect 5542 1112 5594 1164
rect 9674 1146 9726 1198
rect 9738 1146 9790 1198
rect 12235 1201 12287 1253
rect 12235 1137 12287 1189
rect 10443 1039 10495 1091
rect 10535 1053 10587 1105
rect 10599 1053 10651 1105
rect 10443 975 10495 1027
rect 12153 1038 12205 1090
rect 10708 969 10760 1021
rect 10773 969 10825 1021
rect 12153 974 12205 1026
rect 5478 874 5530 926
rect 5542 874 5594 926
rect 9019 896 9071 903
rect 9019 862 9025 896
rect 9025 862 9059 896
rect 9059 862 9071 896
rect 9019 851 9071 862
rect 9085 896 9137 903
rect 9085 862 9097 896
rect 9097 862 9131 896
rect 9131 862 9137 896
rect 9085 851 9137 862
rect 9346 896 9398 902
rect 9438 896 9490 902
rect 9346 862 9352 896
rect 9352 862 9386 896
rect 9386 862 9398 896
rect 9438 862 9458 896
rect 9458 862 9490 896
rect 9346 850 9398 862
rect 9438 850 9490 862
rect 9674 887 9726 939
rect 9738 887 9790 939
rect 10496 887 10548 939
rect 10560 887 10612 939
rect 10743 888 10795 940
rect 10807 888 10859 940
rect 12347 1081 12399 1087
rect 12347 1047 12366 1081
rect 12366 1047 12399 1081
rect 12347 1035 12399 1047
rect 12347 1008 12399 1011
rect 12347 974 12366 1008
rect 12366 974 12399 1008
rect 12347 959 12399 974
rect 12347 901 12366 934
rect 12366 901 12399 934
rect 12347 882 12399 901
rect 9560 851 9612 857
rect 9560 817 9578 851
rect 9578 817 9612 851
rect 9560 805 9612 817
rect 9624 851 9676 857
rect 9624 817 9651 851
rect 9651 817 9676 851
rect 9624 805 9676 817
rect 992 770 1044 790
rect 1061 770 1113 790
rect 992 738 1044 770
rect 1061 738 1087 770
rect 1087 738 1113 770
rect 1130 738 1182 790
rect 1199 738 1251 790
rect 1268 738 1320 790
rect 1337 738 1389 790
rect 1405 738 1457 790
rect 1473 738 1525 790
rect 11465 789 11517 841
rect 11529 789 11581 841
rect 12117 787 12169 839
rect 12181 833 12233 839
rect 12181 799 12183 833
rect 12183 799 12217 833
rect 12217 799 12233 833
rect 12181 787 12233 799
rect 12347 828 12366 857
rect 12366 828 12399 857
rect 12347 805 12399 828
rect 12347 754 12366 780
rect 12366 754 12399 780
rect 992 664 1044 696
rect 1061 664 1087 696
rect 1087 664 1113 696
rect 992 644 1044 664
rect 1061 644 1113 664
rect 1130 644 1182 696
rect 1199 644 1251 696
rect 1268 644 1320 696
rect 1337 644 1389 696
rect 1405 644 1457 696
rect 1473 644 1525 696
rect 9812 684 9864 736
rect 9876 684 9928 736
rect 10869 726 10921 738
rect 10869 692 10900 726
rect 10900 692 10921 726
rect 10869 686 10921 692
rect 10933 726 10985 738
rect 10933 692 10938 726
rect 10938 692 10972 726
rect 10972 692 10985 726
rect 10933 686 10985 692
rect 11028 684 11080 736
rect 11092 730 11144 736
rect 11092 696 11111 730
rect 11111 696 11144 730
rect 12347 728 12399 754
rect 11092 684 11144 696
rect 11465 520 11517 532
rect 11465 486 11497 520
rect 11497 486 11517 520
rect 11465 480 11517 486
rect 11529 520 11581 532
rect 11529 486 11535 520
rect 11535 486 11569 520
rect 11569 486 11581 520
rect 11529 480 11581 486
rect 12117 424 12169 476
rect 12181 424 12233 476
rect 12363 540 12415 592
rect 12887 1363 12939 1415
rect 12956 1363 13008 1415
rect 13025 1363 13077 1415
rect 13094 1363 13146 1415
rect 13163 1363 13215 1415
rect 12887 1293 12939 1345
rect 12956 1293 13008 1345
rect 13025 1293 13077 1345
rect 13094 1293 13146 1345
rect 13163 1293 13215 1345
rect 12887 1223 12939 1275
rect 12956 1223 13008 1275
rect 13025 1223 13077 1275
rect 13094 1223 13146 1275
rect 13163 1223 13215 1275
rect 12887 1152 12939 1204
rect 12956 1152 13008 1204
rect 13025 1152 13077 1204
rect 13094 1152 13146 1204
rect 13163 1152 13215 1204
rect 12887 1081 12939 1133
rect 12956 1081 13008 1133
rect 13025 1081 13077 1133
rect 13094 1081 13146 1133
rect 13163 1081 13215 1133
rect 14823 945 14875 997
rect 14823 879 14875 931
rect 12363 476 12415 528
rect 14753 488 14805 540
rect 14817 488 14869 540
rect 12434 255 12486 307
rect 12498 255 12550 307
<< metal2 >>
tri 1301 6953 1353 7005 se
rect 1353 6953 1468 7005
rect 1520 6953 1534 7005
rect 1586 6953 1592 7005
tri 1273 6925 1301 6953 se
rect 1301 6925 1347 6953
tri 1347 6925 1375 6953 nw
tri 1221 6873 1273 6925 se
rect 1221 5703 1273 6873
tri 1273 6851 1347 6925 nw
rect 3354 6878 3400 6924
rect 3827 6885 3879 6924
rect 7271 6574 7277 6626
rect 7329 6574 7341 6626
rect 7393 6574 7399 6626
tri 7271 6498 7347 6574 ne
tri 1221 5701 1223 5703 ne
rect 1223 5701 1273 5703
tri 1273 5701 1297 5725 sw
tri 1223 5678 1246 5701 ne
rect 1246 5678 1297 5701
tri 1297 5678 1320 5701 sw
tri 1246 5651 1273 5678 ne
rect 1273 5651 1320 5678
tri 1273 5631 1293 5651 ne
rect 1293 5631 1320 5651
rect -370 5625 -318 5631
tri 1293 5627 1297 5631 ne
rect 1297 5627 1320 5631
tri 1320 5627 1371 5678 sw
tri 1297 5626 1298 5627 ne
rect 1298 5626 1371 5627
tri 1371 5626 1372 5627 sw
tri 1298 5598 1326 5626 ne
rect 1326 5598 1372 5626
tri 1372 5598 1400 5626 sw
rect -370 5561 -318 5573
tri 1326 5553 1371 5598 ne
rect 1371 5553 1400 5598
tri 1400 5553 1445 5598 sw
tri 1371 5546 1378 5553 ne
rect 1378 5546 1445 5553
tri 1445 5546 1452 5553 sw
rect 6870 5546 6876 5598
rect 6928 5546 6940 5598
rect 6992 5546 6998 5598
rect -463 4606 -411 4612
rect -463 4542 -411 4554
rect -645 4116 -493 4122
rect -593 4064 -545 4116
rect -645 4039 -493 4064
rect -593 3987 -545 4039
rect -645 3962 -493 3987
rect -593 3910 -545 3962
rect -645 3885 -493 3910
rect -593 3833 -545 3885
rect -645 3808 -493 3833
rect -593 3756 -545 3808
rect -645 1977 -493 3756
rect -463 3708 -411 4490
rect -463 3642 -411 3656
rect -463 3584 -411 3590
rect -465 3444 -413 3450
rect -465 3380 -413 3392
rect -465 2527 -413 3328
rect -465 2461 -413 2475
rect -465 2403 -413 2409
tri -493 1977 -448 2022 sw
rect -645 1973 -448 1977
tri -448 1973 -444 1977 sw
rect -645 1959 -444 1973
tri -444 1959 -430 1973 sw
rect -645 1958 -430 1959
tri -430 1958 -429 1959 sw
rect -645 1854 -563 1958
tri -645 1829 -620 1854 ne
rect -620 1829 -563 1854
tri -620 1772 -563 1829 ne
tri -374 696 -370 700 se
rect -370 696 -318 5509
tri 1378 5504 1420 5546 ne
rect 1420 5512 1452 5546
tri 1452 5512 1486 5546 sw
tri 6874 5512 6908 5546 ne
rect 1420 5504 1486 5512
rect -18 5498 34 5504
rect -194 5492 -142 5498
rect -194 5406 -142 5440
rect -194 4885 -142 5354
tri 1420 5495 1429 5504 ne
rect 1429 5495 1486 5504
tri 1486 5495 1503 5512 sw
tri 1429 5480 1444 5495 ne
rect 1444 5480 1503 5495
tri 1503 5480 1518 5495 sw
tri 1444 5479 1445 5480 ne
rect 1445 5479 1518 5480
tri 1518 5479 1519 5480 sw
rect -18 5426 34 5446
tri 1445 5428 1496 5479 ne
rect 1496 5428 1519 5479
tri 1519 5428 1570 5479 sw
tri 1496 5405 1519 5428 ne
rect 1519 5405 1570 5428
tri 1570 5405 1593 5428 sw
tri 1519 5398 1526 5405 ne
rect 1526 5398 1593 5405
tri 1593 5398 1600 5405 sw
tri -142 4885 -136 4891 sw
rect -194 4869 -136 4885
tri -194 4858 -183 4869 ne
rect -183 4858 -136 4869
tri -136 4858 -109 4885 sw
tri -183 4852 -177 4858 ne
rect -177 4852 -109 4858
tri -109 4852 -103 4858 sw
tri -177 4841 -166 4852 ne
rect -166 4841 -103 4852
tri -103 4841 -92 4852 sw
tri -166 4835 -160 4841 ne
rect -160 4835 -92 4841
tri -92 4835 -86 4841 sw
tri -160 4827 -152 4835 ne
rect -152 4827 -86 4835
tri -86 4827 -78 4835 sw
tri -152 4817 -142 4827 ne
rect -142 4817 -78 4827
tri -142 4805 -130 4817 ne
rect -267 4709 -211 4718
tri -268 4708 -267 4709 se
tri -288 4688 -268 4708 se
rect -268 4688 -267 4708
tri -211 4708 -201 4718 sw
rect -211 4688 -201 4708
tri -201 4688 -181 4708 sw
rect -288 4636 -282 4688
rect -230 4636 -218 4653
rect -166 4636 -160 4688
tri -288 4626 -278 4636 ne
rect -278 4629 -191 4636
rect -278 4626 -267 4629
tri -278 4615 -267 4626 ne
rect -211 4626 -191 4629
tri -191 4626 -181 4636 nw
tri -211 4606 -191 4626 nw
rect -267 4564 -211 4573
tri -154 4534 -130 4558 se
rect -130 4534 -78 4817
rect -18 4708 34 5374
tri 1526 5346 1578 5398 ne
rect 1578 5360 1600 5398
tri 1600 5360 1638 5398 sw
rect 1578 5346 1638 5360
tri 1638 5346 1652 5360 sw
tri 6894 5346 6908 5360 se
rect 6908 5346 6960 5546
tri 6960 5512 6994 5546 nw
tri 6960 5346 6974 5360 sw
tri 1578 5332 1592 5346 ne
rect 1592 5332 1652 5346
tri 1652 5332 1666 5346 sw
tri 6880 5332 6894 5346 se
rect 6894 5332 6974 5346
rect 715 5280 721 5332
rect 773 5280 785 5332
rect 837 5280 843 5332
tri 1592 5331 1593 5332 ne
rect 1593 5331 1666 5332
tri 1666 5331 1667 5332 sw
tri 6879 5331 6880 5332 se
rect 6880 5331 6974 5332
tri 1593 5326 1598 5331 ne
rect 1598 5326 1667 5331
tri 1667 5326 1672 5331 sw
tri 6874 5326 6879 5331 se
rect 6879 5326 6974 5331
tri 6974 5326 6994 5346 sw
tri 7339 5326 7347 5334 se
rect 7347 5326 7399 6574
rect 9422 6574 9428 6626
rect 9480 6574 9492 6626
rect 9544 6574 9550 6626
tri 13110 6574 13136 6600 se
rect 13136 6574 14739 6600
tri 14739 6574 14765 6600 sw
tri 9422 6536 9460 6574 ne
tri 9437 5495 9460 5518 se
rect 9460 5512 9512 6574
tri 9512 6536 9550 6574 nw
tri 13087 6551 13110 6574 se
rect 13110 6551 14765 6574
tri 14765 6551 14788 6574 sw
tri 13072 6536 13087 6551 se
rect 13087 6548 14788 6551
rect 13087 6536 13136 6548
tri 13062 6526 13072 6536 se
rect 13072 6526 13136 6536
tri 13136 6526 13158 6548 nw
tri 14701 6526 14723 6548 ne
rect 14723 6526 14788 6548
tri 12988 6452 13062 6526 se
tri 13062 6452 13136 6526 nw
tri 14723 6513 14736 6526 ne
tri 12981 6445 12988 6452 se
rect 12988 6445 13055 6452
tri 13055 6445 13062 6452 nw
rect 12981 6434 13044 6445
tri 13044 6434 13055 6445 nw
rect 14736 6434 14788 6526
rect 12598 5875 12604 5927
rect 12656 5875 12668 5927
rect 12720 5875 12726 5927
tri 12618 5847 12646 5875 ne
rect 11679 5626 11685 5678
rect 11737 5626 11749 5678
rect 11801 5626 11807 5678
tri 11676 5598 11679 5601 se
rect 11679 5598 11774 5626
tri 11774 5598 11802 5626 nw
tri 12627 5598 12646 5617 se
rect 12646 5598 12698 5875
tri 12698 5847 12726 5875 nw
tri 12943 5678 12981 5716 se
rect 12981 5678 13033 6434
tri 13033 6423 13044 6434 nw
rect 14736 6370 14788 6382
rect 14736 6312 14788 6318
tri 13033 5678 13071 5716 sw
rect 12943 5626 12949 5678
rect 13001 5626 13013 5678
rect 13065 5626 13071 5678
tri 11624 5546 11676 5598 se
rect 11676 5546 11722 5598
tri 11722 5546 11774 5598 nw
rect 12194 5546 12200 5598
rect 12252 5546 12264 5598
rect 12316 5546 12322 5598
tri 12624 5595 12627 5598 se
rect 12627 5595 12698 5598
tri 12575 5546 12624 5595 se
tri 11597 5519 11624 5546 se
rect 11624 5519 11695 5546
tri 11695 5519 11722 5546 nw
tri 12198 5519 12225 5546 ne
rect 12225 5519 12284 5546
tri 11596 5518 11597 5519 se
rect 11597 5518 11695 5519
tri 9512 5512 9518 5518 sw
tri 11590 5512 11596 5518 se
rect 11596 5512 11695 5518
tri 12225 5512 12232 5519 ne
rect 9460 5495 9518 5512
tri 9518 5495 9535 5512 sw
tri 11573 5495 11590 5512 se
rect 11590 5495 11695 5512
tri 9422 5480 9437 5495 se
rect 9437 5480 9535 5495
tri 9535 5480 9550 5495 sw
rect 9422 5428 9428 5480
rect 9480 5428 9492 5480
rect 9544 5428 9550 5480
tri 11567 5489 11573 5495 se
rect 11573 5489 11695 5495
rect 11567 5480 11695 5489
rect 11567 5428 11573 5480
rect 11625 5428 11637 5480
rect 11689 5428 11695 5480
rect 12073 5443 12079 5495
rect 12131 5443 12143 5495
rect 12195 5443 12201 5495
tri 1598 5280 1644 5326 ne
rect 1644 5280 1672 5326
tri 1672 5280 1718 5326 sw
rect 715 5274 795 5280
tri 795 5274 801 5280 nw
tri 1644 5274 1650 5280 ne
rect 1650 5274 1718 5280
tri 1718 5274 1724 5280 sw
rect 6870 5274 6876 5326
rect 6928 5274 6940 5326
rect 6992 5274 6998 5326
tri 7331 5318 7339 5326 se
rect 7339 5318 7399 5326
tri 7287 5274 7331 5318 se
rect 7331 5312 7399 5318
rect 7331 5274 7353 5312
rect 715 5266 787 5274
tri 787 5266 795 5274 nw
tri 1650 5266 1658 5274 ne
rect 1658 5266 1724 5274
tri 1724 5266 1732 5274 sw
tri 7279 5266 7287 5274 se
rect 7287 5266 7353 5274
tri 7353 5266 7399 5312 nw
rect 9435 5266 9441 5318
rect 9493 5266 9505 5318
rect 9557 5266 9563 5318
tri 688 4858 715 4885 se
rect 715 4862 767 5266
tri 767 5246 787 5266 nw
tri 1658 5257 1667 5266 ne
rect 1667 5257 1732 5266
tri 1732 5257 1741 5266 sw
tri 7273 5260 7279 5266 se
rect 7279 5260 7347 5266
tri 7347 5260 7353 5266 nw
tri 9435 5260 9441 5266 ne
rect 9441 5260 9557 5266
tri 9557 5260 9563 5266 nw
tri 7270 5257 7273 5260 se
rect 7273 5257 7315 5260
tri 1667 5246 1678 5257 ne
rect 1678 5246 1741 5257
tri 1741 5246 1752 5257 sw
tri 7259 5246 7270 5257 se
rect 7270 5246 7315 5257
tri 1678 5239 1685 5246 ne
rect 1685 5239 1752 5246
tri 1752 5239 1759 5246 sw
tri 7258 5245 7259 5246 se
rect 7259 5245 7315 5246
rect 5228 5239 5280 5245
tri 1685 5187 1737 5239 ne
rect 1737 5187 1759 5239
tri 1759 5187 1811 5239 sw
tri 1737 5183 1741 5187 ne
rect 1741 5183 1811 5187
tri 1811 5183 1815 5187 sw
tri 1741 5175 1749 5183 ne
rect 1749 5175 1815 5183
tri 1815 5175 1823 5183 sw
rect 5228 5175 5280 5187
tri 1749 5123 1801 5175 ne
rect 1801 5123 1823 5175
tri 1823 5123 1875 5175 sw
tri 1801 5109 1815 5123 ne
rect 1815 5109 1875 5123
tri 1875 5109 1889 5123 sw
tri 1815 5102 1822 5109 ne
rect 1822 5102 1889 5109
tri 1889 5102 1896 5109 sw
tri 1822 5035 1889 5102 ne
rect 1889 5035 1896 5102
tri 1896 5035 1963 5102 sw
tri 1889 5013 1911 5035 ne
rect 715 4858 763 4862
tri 763 4858 767 4862 nw
rect 823 4858 829 4910
rect 881 4858 894 4910
rect 946 4858 959 4910
rect 1011 4858 1024 4910
rect 1076 4858 1089 4910
rect 1141 4858 1153 4910
rect 1205 4858 1217 4910
rect 1269 4858 1281 4910
rect 1333 4858 1345 4910
rect 1397 4858 1409 4910
rect 1461 4858 1473 4910
rect 1525 4858 1531 4910
tri 682 4852 688 4858 se
rect 688 4852 757 4858
tri 757 4852 763 4858 nw
tri 677 4847 682 4852 se
rect 682 4847 752 4852
tri 752 4847 757 4852 nw
rect 677 4841 746 4847
tri 746 4841 752 4847 nw
rect 677 4835 740 4841
tri 740 4835 746 4841 nw
rect 823 4835 1531 4858
tri 34 4708 45 4719 sw
rect -18 4697 45 4708
tri -18 4678 1 4697 ne
rect 1 4678 45 4697
tri 45 4678 75 4708 sw
tri 1 4649 30 4678 ne
rect 30 4649 75 4678
tri 75 4649 104 4678 sw
tri 30 4645 34 4649 ne
rect 34 4645 104 4649
tri 34 4627 52 4645 ne
tri -183 4505 -154 4534 se
rect -154 4518 -78 4534
rect -154 4505 -91 4518
tri -91 4505 -78 4518 nw
tri -193 4495 -183 4505 se
rect -183 4495 -101 4505
tri -101 4495 -91 4505 nw
tri -241 4391 -193 4439 se
rect -193 4417 -141 4495
tri -141 4455 -101 4495 nw
rect -193 4391 -167 4417
tri -167 4391 -141 4417 nw
rect -103 4443 -51 4449
tri -251 4381 -241 4391 se
rect -241 4381 -177 4391
tri -177 4381 -167 4391 nw
tri -255 4377 -251 4381 se
rect -251 4377 -181 4381
tri -181 4377 -177 4381 nw
rect -103 4377 -51 4391
tri -267 4365 -255 4377 se
rect -255 4365 -193 4377
tri -193 4365 -181 4377 nw
rect -374 687 -318 696
rect -374 607 -318 631
rect -374 541 -318 551
tri -277 4355 -267 4365 se
rect -267 4355 -203 4365
tri -203 4355 -193 4365 nw
tri -306 424 -277 453 se
rect -277 431 -225 4355
tri -225 4333 -203 4355 nw
rect -187 4274 -135 4280
rect -187 4210 -135 4222
rect -187 2530 -135 4158
rect -103 3622 -51 4325
rect -103 3558 -51 3570
rect -103 3500 -51 3506
tri 20 3454 52 3486 se
rect 52 3464 104 4645
rect 238 4140 290 4146
rect 238 4061 290 4088
rect 238 3982 290 4009
rect 238 3903 290 3930
rect 238 3824 290 3851
rect 136 3666 192 3675
rect 136 3591 139 3610
rect 191 3591 192 3610
rect 136 3586 192 3591
rect 136 3527 139 3530
rect 191 3527 192 3530
rect 136 3521 192 3527
rect 52 3454 94 3464
tri 94 3454 104 3464 nw
tri 4 3438 20 3454 se
rect 20 3438 78 3454
tri 78 3438 94 3454 nw
tri -9 3425 4 3438 se
rect 4 3425 65 3438
tri 65 3425 78 3438 nw
tri -22 3412 -9 3425 se
rect -9 3412 52 3425
tri 52 3412 65 3425 nw
tri -33 3401 -22 3412 se
rect -22 3401 41 3412
tri 41 3401 52 3412 nw
rect 121 3401 173 3407
tri -85 3349 -33 3401 se
rect -33 3349 -11 3401
tri -11 3349 41 3401 nw
tri -88 3346 -85 3349 se
rect -85 3346 -14 3349
tri -14 3346 -11 3349 nw
tri -90 3344 -88 3346 se
rect -88 3344 -16 3346
tri -16 3344 -14 3346 nw
tri -96 3338 -90 3344 se
rect -90 3338 -22 3344
tri -22 3338 -16 3344 nw
tri -99 3335 -96 3338 se
rect -96 3335 -25 3338
tri -25 3335 -22 3338 nw
rect 121 3335 173 3349
rect -187 2466 -135 2478
rect -187 2408 -135 2414
tri -105 3329 -99 3335 se
rect -99 3329 -31 3335
tri -31 3329 -25 3335 nw
rect -277 424 -232 431
tri -232 424 -225 431 nw
tri -126 2101 -105 2122 se
rect -105 2101 -53 3329
tri -53 3307 -31 3329 nw
tri 99 3103 121 3125 se
rect 121 3103 173 3283
tri 70 3074 99 3103 se
rect 99 3087 157 3103
tri 157 3087 173 3103 nw
rect 238 3126 290 3772
rect 99 3074 144 3087
tri 144 3074 157 3087 nw
tri 55 3059 70 3074 se
rect 70 3059 127 3074
tri 53 3057 55 3059 se
rect 55 3057 127 3059
tri 127 3057 144 3074 nw
tri 50 3054 53 3057 se
rect 53 3054 124 3057
tri 124 3054 127 3057 nw
rect 238 3054 290 3074
tri 25 3029 50 3054 se
rect 50 3029 99 3054
tri 99 3029 124 3054 nw
tri 3 3007 25 3029 se
rect 25 3007 72 3029
rect 3 3002 72 3007
tri 72 3002 99 3029 nw
rect 3 2330 55 3002
tri 55 2985 72 3002 nw
rect 238 2982 290 3002
rect 238 2909 290 2930
rect 677 2947 729 4835
tri 729 4824 740 4835 nw
rect 823 4783 829 4835
rect 881 4783 894 4835
rect 946 4783 959 4835
rect 1011 4783 1024 4835
rect 1076 4783 1089 4835
rect 1141 4783 1153 4835
rect 1205 4783 1217 4835
rect 1269 4783 1281 4835
rect 1333 4783 1345 4835
rect 1397 4783 1409 4835
rect 1461 4783 1473 4835
rect 1525 4783 1531 4835
rect 1911 4806 1963 5035
tri 1963 4806 1975 4818 sw
rect 1911 4796 1975 4806
tri 1911 4783 1924 4796 ne
rect 1924 4783 1975 4796
tri 1975 4783 1998 4806 sw
rect 823 4760 1531 4783
tri 1924 4766 1941 4783 ne
rect 1941 4766 1998 4783
tri 1998 4766 2015 4783 sw
rect 823 4708 829 4760
rect 881 4708 894 4760
rect 946 4708 959 4760
rect 1011 4708 1024 4760
rect 1076 4708 1089 4760
rect 1141 4708 1153 4760
rect 1205 4708 1217 4760
rect 1269 4708 1281 4760
rect 1333 4708 1345 4760
rect 1397 4708 1409 4760
rect 1461 4708 1473 4760
rect 1525 4708 1531 4760
tri 1941 4732 1975 4766 ne
rect 1975 4732 2015 4766
tri 2015 4732 2049 4766 sw
tri 1975 4714 1993 4732 ne
rect 1993 4714 2049 4732
tri 2049 4714 2067 4732 sw
rect 823 4505 1531 4708
tri 1993 4678 2029 4714 ne
rect 2029 4678 2067 4714
tri 2067 4678 2103 4714 sw
tri 2029 4658 2049 4678 ne
rect 2049 4658 2103 4678
tri 2103 4658 2123 4678 sw
tri 2049 4626 2081 4658 ne
rect 2081 4626 2123 4658
tri 2123 4626 2155 4658 sw
tri 2081 4596 2111 4626 ne
rect 2111 4596 2155 4626
tri 2155 4596 2185 4626 sw
tri 2111 4586 2121 4596 ne
rect 2121 4586 2185 4596
tri 2185 4586 2195 4596 sw
tri 2121 4584 2123 4586 ne
rect 2123 4584 2195 4586
tri 2195 4584 2197 4586 sw
tri 2123 4534 2173 4584 ne
rect 2173 4534 2197 4584
tri 2197 4534 2247 4584 sw
rect 3622 4534 3628 4586
rect 3680 4534 3692 4586
rect 3744 4544 3750 4586
tri 3750 4544 3792 4586 sw
rect 3744 4534 3792 4544
tri 3792 4534 3802 4544 sw
tri 2173 4510 2197 4534 ne
rect 2197 4510 2247 4534
tri 2247 4510 2271 4534 sw
tri 3732 4510 3756 4534 ne
rect 3756 4510 3802 4534
tri 2197 4505 2202 4510 ne
rect 2202 4505 2271 4510
tri 2271 4505 2276 4510 sw
tri 3756 4505 3761 4510 ne
rect 3761 4505 3802 4510
tri 3802 4505 3831 4534 sw
rect 823 4453 829 4505
rect 881 4453 894 4505
rect 946 4453 959 4505
rect 1011 4453 1024 4505
rect 1076 4453 1089 4505
rect 1141 4453 1153 4505
rect 1205 4453 1217 4505
rect 1269 4453 1281 4505
rect 1333 4453 1345 4505
rect 1397 4453 1409 4505
rect 1461 4453 1473 4505
rect 1525 4453 1531 4505
rect 823 4433 1531 4453
tri 2202 4436 2271 4505 ne
rect 2271 4436 2276 4505
tri 2276 4436 2345 4505 sw
tri 3761 4466 3800 4505 ne
rect 3800 4466 3831 4505
tri 3831 4466 3870 4505 sw
tri 3800 4449 3817 4466 ne
rect 3817 4449 3870 4466
tri 3817 4436 3830 4449 ne
rect 3830 4436 3870 4449
rect 823 4381 829 4433
rect 881 4381 894 4433
rect 946 4381 959 4433
rect 1011 4381 1024 4433
rect 1076 4381 1089 4433
rect 1141 4381 1153 4433
rect 1205 4381 1217 4433
rect 1269 4381 1281 4433
rect 1333 4381 1345 4433
rect 1397 4381 1409 4433
rect 1461 4381 1473 4433
rect 1525 4381 1531 4433
tri 2271 4415 2292 4436 ne
rect 2292 4415 2345 4436
tri 2345 4415 2366 4436 sw
tri 3830 4415 3851 4436 ne
rect 3851 4415 3870 4436
tri 3870 4415 3921 4466 sw
rect 823 3923 1531 4381
tri 2292 4363 2344 4415 ne
rect 2344 4363 2366 4415
tri 2366 4363 2418 4415 sw
tri 3851 4396 3870 4415 ne
rect 3870 4413 3921 4415
tri 3921 4413 3923 4415 sw
tri 2344 4362 2345 4363 ne
rect 2345 4362 2418 4363
tri 2418 4362 2419 4363 sw
tri 2345 4350 2357 4362 ne
rect 2357 4350 2419 4362
tri 2357 4340 2367 4350 ne
rect 2097 4209 2103 4261
rect 2155 4209 2167 4261
rect 2219 4209 2225 4261
rect 823 3871 829 3923
rect 881 3871 902 3923
rect 954 3871 974 3923
rect 1026 3871 1046 3923
rect 1098 3871 1118 3923
rect 1170 3871 1190 3923
rect 1242 3871 1531 3923
rect 823 3654 1531 3871
rect 823 3602 947 3654
rect 999 3602 1013 3654
rect 1065 3602 1079 3654
rect 1131 3602 1145 3654
rect 1197 3602 1211 3654
rect 1263 3602 1277 3654
rect 1329 3602 1343 3654
rect 1395 3602 1408 3654
rect 1460 3602 1473 3654
rect 1525 3602 1531 3654
rect 823 3580 1531 3602
rect 823 3528 947 3580
rect 999 3528 1013 3580
rect 1065 3528 1079 3580
rect 1131 3528 1145 3580
rect 1197 3528 1211 3580
rect 1263 3528 1277 3580
rect 1329 3528 1343 3580
rect 1395 3528 1408 3580
rect 1460 3528 1473 3580
rect 1525 3528 1531 3580
rect 823 3506 1531 3528
rect 823 3454 947 3506
rect 999 3454 1013 3506
rect 1065 3454 1079 3506
rect 1131 3454 1145 3506
rect 1197 3454 1211 3506
rect 1263 3454 1277 3506
rect 1329 3454 1343 3506
rect 1395 3454 1408 3506
rect 1460 3454 1473 3506
rect 1525 3454 1531 3506
rect 823 3445 1531 3454
tri 823 3438 830 3445 ne
rect 830 3438 1531 3445
tri 830 3425 843 3438 ne
rect 843 3425 1531 3438
tri 843 3373 895 3425 ne
rect 895 3373 1531 3425
tri 895 3369 899 3373 ne
rect 899 3369 1531 3373
tri 899 3346 922 3369 ne
rect 922 3346 1531 3369
tri 922 3344 924 3346 ne
rect 924 3344 1531 3346
tri 924 3292 976 3344 ne
rect 976 3292 1531 3344
tri 976 3282 986 3292 ne
tri 729 2947 751 2969 sw
tri 677 2929 695 2947 ne
rect 695 2940 751 2947
tri 751 2940 758 2947 sw
rect 695 2929 758 2940
tri 695 2918 706 2929 ne
rect 238 2836 290 2857
rect 238 2763 290 2784
rect 238 2690 290 2711
rect 238 2617 290 2638
rect 238 2559 290 2565
rect 3 2266 55 2278
rect 3 2208 55 2214
rect -126 2100 -53 2101
tri -351 379 -306 424 se
rect -306 379 -277 424
tri -277 379 -232 424 nw
tri -129 405 -126 408 se
rect -126 405 -74 2100
tri -74 2079 -53 2100 nw
rect 706 1654 758 2929
rect 986 2718 1531 3292
rect 1698 4129 1704 4181
rect 1756 4129 1773 4181
rect 1825 4129 1842 4181
rect 1894 4129 1911 4181
rect 1963 4129 1980 4181
rect 2032 4129 2038 4181
rect 1698 4106 2038 4129
rect 1698 4054 1704 4106
rect 1756 4054 1773 4106
rect 1825 4054 1842 4106
rect 1894 4054 1911 4106
rect 1963 4054 1980 4106
rect 2032 4054 2038 4106
rect 1698 4031 2038 4054
rect 1698 3979 1704 4031
rect 1756 3979 1773 4031
rect 1825 3979 1842 4031
rect 1894 3979 1911 4031
rect 1963 3979 1980 4031
rect 2032 3979 2038 4031
rect 1698 3057 2038 3979
rect 2097 3735 2225 4209
rect 2097 3683 2103 3735
rect 2155 3683 2167 3735
rect 2219 3683 2225 3735
rect 2367 3292 2419 4350
rect 2447 4209 2453 4261
rect 2505 4209 2517 4261
rect 2569 4209 2575 4261
rect 2447 3871 2575 4209
rect 2613 4209 2619 4261
rect 2671 4209 2683 4261
rect 2735 4209 2741 4261
rect 2613 3951 2741 4209
rect 2613 3899 2619 3951
rect 2671 3899 2683 3951
rect 2735 3899 2741 3951
rect 3150 4129 3156 4181
rect 3208 4129 3220 4181
rect 3272 4129 3284 4181
rect 3336 4129 3348 4181
rect 3400 4129 3412 4181
rect 3464 4129 3476 4181
rect 3528 4129 3540 4181
rect 3592 4129 3598 4181
rect 3150 4106 3598 4129
rect 3150 4054 3156 4106
rect 3208 4054 3220 4106
rect 3272 4054 3284 4106
rect 3336 4054 3348 4106
rect 3400 4054 3412 4106
rect 3464 4054 3476 4106
rect 3528 4054 3540 4106
rect 3592 4054 3598 4106
rect 3150 4031 3598 4054
rect 3150 3987 3156 4031
rect 3208 3987 3220 4031
rect 3272 3987 3284 4031
rect 3336 3987 3348 4031
rect 3400 3987 3412 4031
rect 3464 3987 3476 4031
rect 3528 3987 3540 4031
rect 3592 3987 3598 4031
rect 3150 3931 3154 3987
rect 3210 3979 3220 3987
rect 3336 3979 3346 3987
rect 3402 3979 3412 3987
rect 3528 3979 3538 3987
rect 3210 3931 3250 3979
rect 3306 3931 3346 3979
rect 3402 3931 3442 3979
rect 3498 3931 3538 3979
rect 3594 3931 3598 3987
rect 3150 3906 3598 3931
rect 2447 3819 2453 3871
rect 2505 3819 2517 3871
rect 2569 3819 2575 3871
rect 3150 3850 3154 3906
rect 3210 3850 3250 3906
rect 3306 3850 3346 3906
rect 3402 3850 3442 3906
rect 3498 3850 3538 3906
rect 3594 3850 3598 3906
rect 3150 3825 3598 3850
tri 3861 3843 3870 3852 se
rect 3870 3843 3923 4413
tri 5222 4313 5228 4319 se
rect 5228 4313 5280 5123
tri 7241 5228 7258 5245 se
rect 7258 5228 7315 5245
tri 7315 5228 7347 5260 nw
tri 9441 5244 9457 5260 ne
rect 9457 5244 9541 5260
tri 9541 5244 9557 5260 nw
tri 9457 5242 9459 5244 ne
rect 9459 5242 9541 5244
tri 9459 5228 9473 5242 ne
rect 9473 5228 9541 5242
tri 10508 5228 10522 5242 se
rect 10522 5228 11301 5242
tri 11301 5228 11315 5242 sw
rect 7241 5224 7311 5228
tri 7311 5224 7315 5228 nw
tri 9473 5224 9477 5228 ne
rect 9477 5224 9541 5228
tri 10504 5224 10508 5228 se
rect 10508 5224 11315 5228
tri 11315 5224 11319 5228 sw
rect 7241 5218 7305 5224
tri 7305 5218 7311 5224 nw
rect 7411 5218 7463 5224
tri 7212 4544 7241 4573 se
rect 7241 4551 7293 5218
tri 7293 5206 7305 5218 nw
rect 7241 4544 7286 4551
tri 7286 4544 7293 4551 nw
tri 9477 5208 9493 5224 ne
rect 7411 5154 7463 5166
tri 7178 4510 7212 4544 se
rect 7212 4510 7247 4544
tri 7173 4505 7178 4510 se
rect 7178 4505 7247 4510
tri 7247 4505 7286 4544 nw
tri 7389 4508 7411 4530 se
rect 7411 4508 7463 5102
rect 7960 5168 8051 5176
tri 8051 5168 8059 5176 nw
rect 7960 5133 8016 5168
tri 8016 5133 8051 5168 nw
tri 7957 4544 7960 4547 se
rect 7960 4544 8012 5133
tri 8012 5129 8016 5133 nw
tri 7386 4505 7389 4508 se
rect 7389 4505 7460 4508
tri 7460 4505 7463 4508 nw
tri 7918 4505 7957 4544 se
rect 7957 4525 8012 4544
rect 7957 4505 7992 4525
tri 7992 4505 8012 4525 nw
tri 7167 4499 7173 4505 se
rect 7173 4499 7241 4505
tri 7241 4499 7247 4505 nw
tri 7380 4499 7386 4505 se
rect 7386 4499 7454 4505
tri 7454 4499 7460 4505 nw
tri 7912 4499 7918 4505 se
rect 7918 4499 7986 4505
tri 7986 4499 7992 4505 nw
tri 7104 4436 7167 4499 se
tri 7093 4425 7104 4436 se
rect 7104 4425 7167 4436
tri 7167 4425 7241 4499 nw
tri 7360 4479 7380 4499 se
rect 7380 4479 7412 4499
tri 7083 4415 7093 4425 se
rect 7093 4415 7157 4425
tri 7157 4415 7167 4425 nw
tri 7082 4414 7083 4415 se
rect 7083 4414 7156 4415
tri 7156 4414 7157 4415 nw
tri 7031 4363 7082 4414 se
rect 7082 4363 7105 4414
tri 7105 4363 7156 4414 nw
tri 7019 4351 7031 4363 se
rect 7031 4351 7093 4363
tri 7093 4351 7105 4363 nw
tri 7018 4350 7019 4351 se
rect 7019 4350 7092 4351
tri 7092 4350 7093 4351 nw
tri 5193 4284 5222 4313 se
rect 5222 4284 5280 4313
tri 7010 4342 7018 4350 se
rect 7018 4342 7084 4350
tri 7084 4342 7092 4350 nw
tri 5173 4264 5193 4284 se
rect 5193 4264 5280 4284
tri 5280 4264 5300 4284 sw
rect 5172 4212 5178 4264
rect 5230 4212 5242 4264
rect 5294 4212 5300 4264
tri 3847 3829 3861 3843 se
rect 3861 3829 3923 3843
tri 3923 3829 3934 3840 sw
tri 3845 3827 3847 3829 se
rect 3847 3827 3934 3829
tri 3934 3827 3936 3829 sw
rect 2865 3739 2871 3791
rect 2923 3739 2935 3791
rect 2987 3739 2993 3791
tri 2865 3727 2877 3739 ne
rect 2877 3727 2981 3739
tri 2981 3727 2993 3739 nw
rect 3150 3769 3154 3825
rect 3210 3769 3250 3825
rect 3306 3769 3346 3825
rect 3402 3769 3442 3825
rect 3498 3769 3538 3825
rect 3594 3769 3598 3825
tri 3837 3819 3845 3827 se
rect 3845 3819 3936 3827
tri 3833 3815 3837 3819 se
rect 3837 3815 3936 3819
tri 3936 3815 3948 3827 sw
tri 3827 3809 3833 3815 se
rect 3833 3809 3948 3815
tri 3948 3809 3954 3815 sw
rect 3150 3744 3598 3769
rect 3826 3757 3832 3809
rect 3884 3757 3896 3809
rect 3948 3757 3954 3809
tri 2877 3714 2890 3727 ne
rect 2890 3714 2981 3727
tri 2890 3689 2915 3714 ne
rect 2915 3689 2981 3714
tri 2915 3686 2918 3689 ne
tri 2419 3292 2453 3326 sw
rect 2367 3240 2373 3292
rect 2425 3240 2437 3292
rect 2489 3240 2495 3292
rect 1698 3005 1704 3057
rect 1756 3005 1773 3057
rect 1825 3005 1842 3057
rect 1894 3005 1911 3057
rect 1963 3005 1980 3057
rect 2032 3005 2038 3057
rect 1698 2981 2038 3005
rect 1698 2929 1704 2981
rect 1756 2929 1773 2981
rect 1825 2929 1842 2981
rect 1894 2929 1911 2981
rect 1963 2929 1980 2981
rect 2032 2929 2038 2981
rect 986 2673 1397 2718
tri 1397 2673 1442 2718 nw
rect 986 2645 1369 2673
tri 1369 2645 1397 2673 nw
tri 886 2571 892 2577 se
rect 892 2571 944 2641
tri 881 2566 886 2571 se
rect 886 2566 944 2571
tri 860 2545 881 2566 se
rect 881 2555 944 2566
rect 881 2545 934 2555
tri 934 2545 944 2555 nw
rect 986 2629 1353 2645
tri 1353 2629 1369 2645 nw
rect 986 2577 1301 2629
tri 1301 2577 1353 2629 nw
rect 986 2571 1295 2577
tri 1295 2571 1301 2577 nw
tri 837 2522 860 2545 se
rect 860 2522 911 2545
tri 911 2522 934 2545 nw
tri 807 2492 837 2522 se
rect 837 2492 881 2522
tri 881 2492 911 2522 nw
rect 807 2437 859 2492
tri 859 2470 881 2492 nw
rect 807 2373 859 2385
rect 807 2315 859 2321
rect 706 1590 758 1602
rect 706 1532 758 1538
rect 986 2154 1279 2571
tri 1279 2555 1295 2571 nw
rect 1698 2442 2038 2929
rect 2114 3160 2120 3212
rect 2172 3160 2184 3212
rect 2236 3160 2242 3212
rect 2114 2898 2242 3160
rect 2114 2846 2120 2898
rect 2172 2846 2184 2898
rect 2236 2846 2242 2898
tri 2905 2645 2918 2658 se
rect 2918 2645 2981 3689
rect 3150 3688 3154 3744
rect 3210 3688 3250 3744
rect 3306 3688 3346 3744
rect 3402 3688 3442 3744
rect 3498 3688 3538 3744
rect 3594 3688 3598 3744
rect 6747 3714 6753 3766
rect 6805 3714 6817 3766
rect 6869 3714 6875 3766
tri 6747 3689 6772 3714 ne
rect 6772 3689 6850 3714
tri 6850 3689 6875 3714 nw
rect 3150 3663 3598 3688
tri 6772 3683 6778 3689 ne
rect 6778 3683 6844 3689
tri 6844 3683 6850 3689 nw
tri 6778 3681 6780 3683 ne
rect 6780 3681 6842 3683
tri 6842 3681 6844 3683 nw
tri 6780 3672 6789 3681 ne
rect 3150 3607 3154 3663
rect 3210 3607 3250 3663
rect 3306 3607 3346 3663
rect 3402 3607 3442 3663
rect 3498 3607 3538 3663
rect 3594 3607 3598 3663
rect 3150 3582 3598 3607
rect 3150 3526 3154 3582
rect 3210 3526 3250 3582
rect 3306 3526 3346 3582
rect 3402 3526 3442 3582
rect 3498 3526 3538 3582
rect 3594 3526 3598 3582
rect 3150 3501 3598 3526
rect 3150 3445 3154 3501
rect 3210 3445 3250 3501
rect 3306 3445 3346 3501
rect 3402 3445 3442 3501
rect 3498 3445 3538 3501
rect 3594 3445 3598 3501
rect 3150 3420 3598 3445
rect 3150 3364 3154 3420
rect 3210 3364 3250 3420
rect 3306 3364 3346 3420
rect 3402 3364 3442 3420
rect 3498 3364 3538 3420
rect 3594 3364 3598 3420
rect 3150 3339 3598 3364
rect 3150 3283 3154 3339
rect 3210 3283 3250 3339
rect 3306 3283 3346 3339
rect 3402 3283 3442 3339
rect 3498 3283 3538 3339
rect 3594 3283 3598 3339
rect 3150 3258 3598 3283
rect 3150 3202 3154 3258
rect 3210 3202 3250 3258
rect 3306 3202 3346 3258
rect 3402 3202 3442 3258
rect 3498 3202 3538 3258
rect 3594 3202 3598 3258
rect 3150 3177 3598 3202
rect 3150 3121 3154 3177
rect 3210 3121 3250 3177
rect 3306 3121 3346 3177
rect 3402 3121 3442 3177
rect 3498 3121 3538 3177
rect 3594 3121 3598 3177
rect 3150 3096 3598 3121
rect 3150 3040 3154 3096
rect 3210 3057 3250 3096
rect 3306 3057 3346 3096
rect 3402 3057 3442 3096
rect 3498 3057 3538 3096
rect 3210 3040 3220 3057
rect 3336 3040 3346 3057
rect 3402 3040 3412 3057
rect 3528 3040 3538 3057
rect 3594 3040 3598 3096
rect 3150 3015 3156 3040
rect 3208 3015 3220 3040
rect 3272 3015 3284 3040
rect 3336 3015 3348 3040
rect 3400 3015 3412 3040
rect 3464 3015 3476 3040
rect 3528 3015 3540 3040
rect 3592 3015 3598 3040
rect 3150 2959 3154 3015
rect 3210 3005 3220 3015
rect 3336 3005 3346 3015
rect 3402 3005 3412 3015
rect 3528 3005 3538 3015
rect 3210 2981 3250 3005
rect 3306 2981 3346 3005
rect 3402 2981 3442 3005
rect 3498 2981 3538 3005
rect 3210 2959 3220 2981
rect 3336 2959 3346 2981
rect 3402 2959 3412 2981
rect 3528 2959 3538 2981
rect 3594 2959 3598 3015
rect 3150 2934 3156 2959
rect 3208 2934 3220 2959
rect 3272 2934 3284 2959
rect 3336 2934 3348 2959
rect 3400 2934 3412 2959
rect 3464 2934 3476 2959
rect 3528 2934 3540 2959
rect 3592 2934 3598 2959
rect 3150 2878 3154 2934
rect 3210 2929 3220 2934
rect 3336 2929 3346 2934
rect 3402 2929 3412 2934
rect 3528 2929 3538 2934
rect 3210 2878 3250 2929
rect 3306 2878 3346 2929
rect 3402 2878 3442 2929
rect 3498 2878 3538 2929
rect 3594 2878 3598 2934
rect 3150 2853 3598 2878
rect 3150 2797 3154 2853
rect 3210 2797 3250 2853
rect 3306 2797 3346 2853
rect 3402 2797 3442 2853
rect 3498 2797 3538 2853
rect 3594 2797 3598 2853
rect 3150 2772 3598 2797
rect 3150 2716 3154 2772
rect 3210 2716 3250 2772
rect 3306 2716 3346 2772
rect 3402 2716 3442 2772
rect 3498 2716 3538 2772
rect 3594 2716 3598 2772
rect 3150 2691 3598 2716
tri 2981 2645 2994 2658 sw
tri 2901 2641 2905 2645 se
rect 2905 2641 2994 2645
tri 2889 2629 2901 2641 se
rect 2901 2629 2994 2641
tri 2994 2629 3010 2645 sw
rect 3150 2635 3154 2691
rect 3210 2635 3250 2691
rect 3306 2635 3346 2691
rect 3402 2635 3442 2691
rect 3498 2635 3538 2691
rect 3594 2635 3598 2691
rect 4498 2718 4504 2770
rect 4556 2718 4568 2770
rect 4620 2718 4626 2770
tri 4498 2690 4526 2718 ne
rect 4526 2690 4598 2718
tri 4598 2690 4626 2718 nw
tri 4526 2686 4530 2690 ne
rect 4530 2686 4594 2690
tri 4594 2686 4598 2690 nw
tri 4530 2673 4543 2686 ne
rect 4543 2673 4594 2686
tri 4543 2670 4546 2673 ne
rect 2889 2577 2895 2629
rect 2947 2577 2959 2629
rect 3011 2577 3017 2629
rect 3150 2610 3598 2635
rect 1698 2390 1704 2442
rect 1756 2390 1773 2442
rect 1825 2390 1842 2442
rect 1894 2390 1911 2442
rect 1963 2390 1980 2442
rect 2032 2390 2038 2442
rect 1698 2364 2038 2390
rect 1698 2312 1704 2364
rect 1756 2312 1773 2364
rect 1825 2312 1842 2364
rect 1894 2312 1911 2364
rect 1963 2312 1980 2364
rect 2032 2312 2038 2364
tri 1279 2154 1302 2177 sw
rect 986 2152 1302 2154
tri 1302 2152 1304 2154 sw
rect 986 2151 1304 2152
tri 1304 2151 1305 2152 sw
rect 986 2135 1305 2151
tri 1305 2135 1321 2151 sw
rect 986 2124 1321 2135
tri 1321 2124 1332 2135 sw
rect 986 2072 1332 2124
tri 1332 2072 1384 2124 sw
rect 986 2064 1384 2072
tri 1384 2064 1392 2072 sw
rect 986 2039 1392 2064
tri 1392 2039 1417 2064 sw
rect 986 2034 1417 2039
tri 1417 2034 1422 2039 sw
rect 986 1503 1531 2034
rect 1698 2029 2038 2312
rect 1698 1977 1704 2029
rect 1756 1977 1773 2029
rect 1825 1977 1842 2029
rect 1894 1977 1911 2029
rect 1963 1977 1980 2029
rect 2032 1977 2038 2029
rect 1698 1955 2038 1977
rect 1698 1903 1704 1955
rect 1756 1903 1773 1955
rect 1825 1903 1842 1955
rect 1894 1903 1911 1955
rect 1963 1903 1980 1955
rect 2032 1903 2038 1955
rect 1698 1881 2038 1903
rect 1698 1829 1704 1881
rect 1756 1829 1773 1881
rect 1825 1829 1842 1881
rect 1894 1829 1911 1881
rect 1963 1829 1980 1881
rect 2032 1829 2038 1881
rect 1698 1828 2038 1829
rect 3150 2554 3154 2610
rect 3210 2554 3250 2610
rect 3306 2554 3346 2610
rect 3402 2554 3442 2610
rect 3498 2554 3538 2610
rect 3594 2554 3598 2610
rect 3150 2529 3598 2554
rect 3150 2473 3154 2529
rect 3210 2473 3250 2529
rect 3306 2473 3346 2529
rect 3402 2473 3442 2529
rect 3498 2473 3538 2529
rect 3594 2473 3598 2529
rect 3150 2447 3598 2473
rect 3150 2391 3154 2447
rect 3210 2442 3250 2447
rect 3306 2442 3346 2447
rect 3402 2442 3442 2447
rect 3498 2442 3538 2447
rect 3210 2391 3220 2442
rect 3336 2391 3346 2442
rect 3402 2391 3412 2442
rect 3528 2391 3538 2442
rect 3594 2391 3598 2447
rect 3150 2390 3156 2391
rect 3208 2390 3220 2391
rect 3272 2390 3284 2391
rect 3336 2390 3348 2391
rect 3400 2390 3412 2391
rect 3464 2390 3476 2391
rect 3528 2390 3540 2391
rect 3592 2390 3598 2391
rect 3150 2365 3598 2390
rect 3150 2309 3154 2365
rect 3210 2364 3250 2365
rect 3306 2364 3346 2365
rect 3402 2364 3442 2365
rect 3498 2364 3538 2365
rect 3210 2312 3220 2364
rect 3336 2312 3346 2364
rect 3402 2312 3412 2364
rect 3528 2312 3538 2364
rect 3210 2309 3250 2312
rect 3306 2309 3346 2312
rect 3402 2309 3442 2312
rect 3498 2309 3538 2312
rect 3594 2309 3598 2365
rect 3150 2283 3598 2309
rect 3150 2227 3154 2283
rect 3210 2227 3250 2283
rect 3306 2227 3346 2283
rect 3402 2227 3442 2283
rect 3498 2227 3538 2283
rect 3594 2227 3598 2283
rect 3150 2201 3598 2227
rect 3150 2145 3154 2201
rect 3210 2145 3250 2201
rect 3306 2145 3346 2201
rect 3402 2145 3442 2201
rect 3498 2145 3538 2201
rect 3594 2145 3598 2201
rect 3150 2119 3598 2145
rect 3150 2063 3154 2119
rect 3210 2063 3250 2119
rect 3306 2063 3346 2119
rect 3402 2063 3442 2119
rect 3498 2063 3538 2119
rect 3594 2063 3598 2119
rect 3150 2037 3598 2063
rect 3150 1981 3154 2037
rect 3210 2029 3250 2037
rect 3306 2029 3346 2037
rect 3402 2029 3442 2037
rect 3498 2029 3538 2037
rect 3210 1981 3220 2029
rect 3336 1981 3346 2029
rect 3402 1981 3412 2029
rect 3528 1981 3538 2029
rect 3594 1981 3598 2037
rect 3150 1977 3156 1981
rect 3208 1977 3220 1981
rect 3272 1977 3284 1981
rect 3336 1977 3348 1981
rect 3400 1977 3412 1981
rect 3464 1977 3476 1981
rect 3528 1977 3540 1981
rect 3592 1977 3598 1981
rect 3150 1955 3598 1977
rect 3150 1899 3154 1955
rect 3210 1903 3220 1955
rect 3336 1903 3346 1955
rect 3402 1903 3412 1955
rect 3528 1903 3538 1955
rect 3210 1899 3250 1903
rect 3306 1899 3346 1903
rect 3402 1899 3442 1903
rect 3498 1899 3538 1903
rect 3594 1899 3598 1955
rect 3150 1881 3598 1899
rect 3150 1873 3156 1881
rect 3208 1873 3220 1881
rect 3272 1873 3284 1881
rect 3336 1873 3348 1881
rect 3400 1873 3412 1881
rect 3464 1873 3476 1881
rect 3528 1873 3540 1881
rect 3592 1873 3598 1881
rect 3150 1817 3154 1873
rect 3210 1829 3220 1873
rect 3336 1829 3346 1873
rect 3402 1829 3412 1873
rect 3528 1829 3538 1873
rect 3210 1817 3250 1829
rect 3306 1817 3346 1829
rect 3402 1817 3442 1829
rect 3498 1817 3538 1829
rect 3594 1817 3598 1873
rect 3150 1791 3598 1817
rect 3150 1735 3154 1791
rect 3210 1735 3250 1791
rect 3306 1735 3346 1791
rect 3402 1735 3442 1791
rect 3498 1735 3538 1791
rect 3594 1735 3598 1791
rect 3150 1709 3598 1735
rect 3150 1653 3154 1709
rect 3210 1653 3250 1709
rect 3306 1653 3346 1709
rect 3402 1653 3442 1709
rect 3498 1653 3538 1709
rect 3594 1653 3598 1709
rect 3150 1644 3598 1653
rect 986 1451 992 1503
rect 1044 1451 1061 1503
rect 1113 1451 1130 1503
rect 1182 1451 1199 1503
rect 1251 1451 1268 1503
rect 1320 1451 1337 1503
rect 1389 1451 1405 1503
rect 1457 1451 1473 1503
rect 1525 1451 1531 1503
rect 986 1429 1531 1451
rect 986 1377 992 1429
rect 1044 1377 1061 1429
rect 1113 1377 1130 1429
rect 1182 1377 1199 1429
rect 1251 1377 1268 1429
rect 1320 1377 1337 1429
rect 1389 1377 1405 1429
rect 1457 1377 1473 1429
rect 1525 1377 1531 1429
rect 986 1355 1531 1377
rect 986 1303 992 1355
rect 1044 1303 1061 1355
rect 1113 1303 1130 1355
rect 1182 1303 1199 1355
rect 1251 1303 1268 1355
rect 1320 1303 1337 1355
rect 1389 1303 1405 1355
rect 1457 1303 1473 1355
rect 1525 1303 1531 1355
rect 986 790 1531 1303
tri 4535 1201 4546 1212 se
rect 4546 1201 4594 2673
tri 6780 2239 6789 2248 se
rect 6789 2239 6842 3681
rect 7010 3346 7062 4342
tri 7062 4320 7084 4342 nw
rect 7204 4209 7210 4261
rect 7262 4209 7274 4261
rect 7326 4209 7332 4261
rect 7204 4201 7292 4209
tri 7292 4201 7300 4209 nw
rect 7204 4197 7288 4201
tri 7288 4197 7292 4201 nw
rect 7204 4189 7280 4197
tri 7280 4189 7288 4197 nw
tri 7062 3346 7073 3357 sw
rect 7010 3344 7073 3346
tri 7073 3344 7075 3346 sw
rect 7010 3303 7075 3344
tri 7075 3303 7116 3344 sw
tri 6999 3292 7010 3303 se
rect 7010 3292 7116 3303
tri 7116 3292 7127 3303 sw
rect 6999 3240 7005 3292
rect 7057 3240 7069 3292
rect 7121 3240 7127 3292
rect 7204 3246 7275 4189
tri 7275 4184 7280 4189 nw
tri 7275 3246 7282 3253 sw
rect 7204 3228 7282 3246
tri 7282 3228 7300 3246 sw
rect 6979 3160 6985 3212
rect 7037 3160 7049 3212
rect 7101 3160 7107 3212
rect 7204 3176 7210 3228
rect 7262 3176 7274 3228
rect 7326 3176 7332 3228
rect 6979 2900 7107 3160
tri 7359 2947 7360 2948 se
rect 7360 2947 7412 4479
tri 7412 4457 7454 4499 nw
tri 7886 4473 7912 4499 se
rect 7912 4473 7960 4499
tri 7960 4473 7986 4499 nw
tri 7871 4458 7886 4473 se
rect 7886 4458 7945 4473
tri 7945 4458 7960 4473 nw
tri 7870 4457 7871 4458 se
rect 7871 4457 7902 4458
tri 7828 4415 7870 4457 se
rect 7870 4415 7902 4457
tri 7902 4415 7945 4458 nw
tri 7794 4261 7828 4295 se
rect 7828 4261 7880 4415
tri 7880 4393 7902 4415 nw
rect 9493 4393 9541 5224
tri 10487 5207 10504 5224 se
rect 10504 5207 11319 5224
tri 11319 5207 11336 5224 sw
tri 10448 5168 10487 5207 se
rect 10487 5190 11336 5207
rect 10487 5168 10522 5190
tri 10522 5168 10544 5190 nw
tri 11279 5168 11301 5190 ne
rect 11301 5168 11336 5190
tri 10413 5133 10448 5168 se
rect 10448 5133 10487 5168
tri 10487 5133 10522 5168 nw
tri 11301 5133 11336 5168 ne
tri 11336 5133 11410 5207 sw
tri 10374 5094 10413 5133 se
rect 10413 5094 10448 5133
tri 10448 5094 10487 5133 nw
tri 11336 5094 11375 5133 ne
rect 11375 5094 11410 5133
tri 10339 5059 10374 5094 se
rect 10374 5059 10413 5094
tri 10413 5059 10448 5094 nw
tri 11375 5059 11410 5094 ne
tri 11410 5059 11484 5133 sw
tri 10300 5020 10339 5059 se
rect 10339 5020 10374 5059
tri 10374 5020 10413 5059 nw
tri 11410 5020 11449 5059 ne
rect 11449 5020 11484 5059
tri 10271 4991 10300 5020 se
rect 10300 4991 10345 5020
tri 10345 4991 10374 5020 nw
tri 11449 4991 11478 5020 ne
rect 11478 4991 11484 5020
tri 11484 4991 11552 5059 sw
tri 10265 4985 10271 4991 se
rect 10271 4985 10339 4991
tri 10339 4985 10345 4991 nw
tri 11478 4985 11484 4991 ne
rect 11484 4985 11552 4991
tri 11552 4985 11558 4991 sw
tri 10237 4957 10265 4985 se
rect 10265 4957 10311 4985
tri 10311 4957 10339 4985 nw
tri 11484 4957 11512 4985 ne
rect 11512 4957 11558 4985
rect 10237 4939 10293 4957
tri 10293 4939 10311 4957 nw
tri 11512 4939 11530 4957 ne
rect 11530 4939 11558 4957
tri 11558 4939 11604 4985 sw
tri 10220 4714 10237 4731 se
rect 10237 4714 10289 4939
tri 10289 4935 10293 4939 nw
tri 11530 4935 11534 4939 ne
rect 11534 4935 11604 4939
tri 11534 4916 11553 4935 ne
rect 11553 4916 11604 4935
tri 11604 4916 11627 4939 sw
tri 11553 4911 11558 4916 ne
rect 11558 4911 11627 4916
tri 11627 4911 11632 4916 sw
tri 11558 4904 11565 4911 ne
rect 11565 4904 11632 4911
tri 11565 4889 11580 4904 ne
tri 10184 4678 10220 4714 se
rect 10220 4678 10289 4714
tri 10289 4678 10312 4701 sw
rect 9930 4626 9936 4678
rect 9988 4626 10000 4678
rect 10052 4626 10058 4678
rect 10184 4626 10190 4678
rect 10242 4626 10254 4678
rect 10306 4626 10312 4678
rect 11580 4637 11632 4904
tri 11632 4637 11636 4641 sw
rect 11580 4626 11636 4637
tri 11636 4626 11647 4637 sw
rect 9930 4529 10058 4626
rect 11580 4596 11647 4626
tri 11647 4596 11677 4626 sw
rect 11580 4544 11621 4596
rect 11673 4544 11685 4596
rect 11737 4544 11743 4596
tri 9930 4505 9954 4529 ne
rect 9954 4505 10058 4529
tri 9954 4499 9960 4505 ne
rect 9960 4499 10058 4505
tri 9960 4458 10001 4499 ne
rect 10001 4426 10058 4499
tri 9541 4393 9543 4395 sw
rect 9493 4391 9543 4393
tri 9543 4391 9545 4393 sw
rect 9493 4375 9545 4391
tri 9493 4363 9505 4375 ne
rect 9505 4363 9545 4375
tri 9545 4363 9573 4391 sw
tri 9505 4350 9518 4363 ne
rect 9518 4350 9573 4363
tri 9573 4350 9586 4363 sw
tri 9518 4323 9545 4350 ne
rect 9545 4323 9586 4350
tri 9586 4323 9613 4350 sw
tri 9545 4313 9555 4323 ne
rect 9555 4313 9613 4323
tri 9613 4313 9623 4323 sw
tri 9555 4261 9607 4313 ne
rect 9607 4261 9623 4313
tri 9623 4261 9675 4313 sw
rect 7596 4209 7602 4261
rect 7654 4209 7666 4261
rect 7718 4209 7724 4261
rect 7752 4209 7758 4261
rect 7810 4209 7822 4261
rect 7874 4209 7880 4261
tri 9607 4255 9613 4261 ne
rect 9613 4255 9675 4261
tri 9675 4255 9681 4261 sw
tri 9613 4253 9615 4255 ne
rect 9615 4253 9681 4255
tri 9681 4253 9683 4255 sw
tri 7647 4201 7655 4209 ne
rect 7655 4201 7724 4209
tri 7803 4201 7811 4209 ne
rect 7811 4201 7880 4209
tri 9615 4201 9667 4253 ne
rect 9667 4201 9683 4253
tri 9683 4201 9735 4253 sw
tri 7655 4197 7659 4201 ne
rect 7659 4197 7724 4201
tri 7811 4197 7815 4201 ne
rect 7815 4197 7880 4201
tri 9667 4197 9671 4201 ne
rect 9671 4197 9735 4201
tri 9735 4197 9739 4201 sw
tri 7659 4189 7667 4197 ne
rect 7667 4189 7724 4197
tri 7815 4189 7823 4197 ne
rect 7823 4189 7880 4197
tri 9671 4189 9679 4197 ne
rect 9679 4189 9739 4197
tri 9739 4189 9747 4197 sw
tri 7667 4187 7669 4189 ne
rect 7669 4187 7724 4189
tri 7823 4187 7825 4189 ne
rect 7825 4187 7880 4189
tri 9679 4187 9681 4189 ne
rect 9681 4187 9747 4189
tri 9747 4187 9749 4189 sw
tri 7669 4184 7672 4187 ne
tri 7326 2914 7359 2947 se
rect 7359 2914 7412 2947
rect 6979 2848 6985 2900
rect 7037 2848 7049 2900
rect 7101 2848 7107 2900
rect 7163 2862 7412 2914
rect 7672 3805 7724 4187
tri 7825 4184 7828 4187 ne
rect 7672 3741 7724 3753
rect 7163 2842 7229 2862
tri 7229 2842 7249 2862 nw
rect 7163 2832 7219 2842
tri 7219 2832 7229 2842 nw
rect 7163 2830 7217 2832
tri 7217 2830 7219 2832 nw
tri 7146 2673 7163 2690 se
rect 7163 2673 7215 2830
tri 7215 2828 7217 2830 nw
rect 7672 2738 7724 3689
tri 7803 3138 7828 3163 se
rect 7828 3138 7880 4187
tri 9681 4156 9712 4187 ne
rect 9712 4156 9749 4187
tri 9016 4152 9020 4156 se
rect 9020 4152 9340 4156
tri 8983 4119 9016 4152 se
rect 9016 4119 9147 4152
tri 8964 4100 8983 4119 se
rect 8983 4100 9147 4119
rect 9199 4100 9214 4152
rect 9266 4100 9280 4152
rect 9332 4100 9340 4152
tri 9712 4137 9731 4156 ne
rect 9731 4137 9749 4156
tri 9749 4137 9799 4187 sw
tri 9731 4119 9749 4137 ne
rect 9749 4119 9799 4137
tri 9799 4119 9817 4137 sw
tri 9749 4109 9759 4119 ne
rect 9759 4109 9817 4119
tri 9817 4109 9827 4119 sw
tri 8921 4057 8964 4100 se
rect 8964 4057 9340 4100
tri 9759 4057 9811 4109 ne
rect 9811 4057 9827 4109
tri 9827 4057 9879 4109 sw
rect 8921 4054 9340 4057
rect 8921 4002 9147 4054
rect 9199 4002 9214 4054
rect 9266 4002 9280 4054
rect 9332 4002 9340 4054
tri 9811 4051 9817 4057 ne
rect 9817 4051 9879 4057
tri 9879 4051 9885 4057 sw
tri 9817 4045 9823 4051 ne
rect 9823 4045 9885 4051
tri 9823 4031 9837 4045 ne
rect 8921 3998 9340 4002
rect 8921 3993 9127 3998
tri 9127 3993 9132 3998 nw
rect 8921 3986 9120 3993
tri 9120 3986 9127 3993 nw
rect 8031 3899 8037 3951
rect 8089 3899 8101 3951
rect 8153 3899 8159 3951
tri 8031 3897 8033 3899 ne
rect 8033 3897 8157 3899
tri 8157 3897 8159 3899 nw
rect 7752 3086 7758 3138
rect 7810 3086 7822 3138
rect 7874 3086 7880 3138
rect 7752 3076 7870 3086
tri 7870 3076 7880 3086 nw
rect 8033 3895 8155 3897
tri 8155 3895 8157 3897 nw
rect 8033 3843 8103 3895
tri 8103 3843 8155 3895 nw
rect 8033 3829 8089 3843
tri 8089 3829 8103 3843 nw
rect 8033 3827 8087 3829
tri 8087 3827 8089 3829 nw
rect 7752 3024 7818 3076
tri 7818 3024 7870 3076 nw
rect 7752 2894 7813 3024
tri 7813 3019 7818 3024 nw
rect 7752 2842 7758 2894
rect 7810 2842 7813 2894
rect 7752 2830 7813 2842
rect 7752 2778 7758 2830
rect 7810 2778 7813 2830
rect 7752 2772 7813 2778
tri 7724 2738 7736 2750 sw
rect 7672 2725 7736 2738
tri 7736 2725 7749 2738 sw
rect 7672 2673 7678 2725
rect 7730 2673 7742 2725
rect 7794 2673 7800 2725
tri 7129 2656 7146 2673 se
rect 7146 2656 7215 2673
rect 7653 2593 7659 2645
rect 7711 2593 7723 2645
rect 7775 2593 7781 2645
rect 7653 2571 7708 2593
tri 7708 2571 7730 2593 nw
tri 6773 2232 6780 2239 se
rect 6780 2232 6842 2239
tri 6842 2232 6849 2239 sw
tri 6767 2226 6773 2232 se
rect 6773 2226 6849 2232
tri 6849 2226 6855 2232 sw
tri 6764 2223 6767 2226 se
rect 6767 2223 6855 2226
tri 6855 2223 6858 2226 sw
tri 6755 2214 6764 2223 se
rect 6764 2214 6858 2223
tri 6858 2214 6867 2223 sw
tri 6747 2206 6755 2214 se
rect 6755 2206 6867 2214
tri 6867 2206 6875 2214 sw
rect 6747 2154 6753 2206
rect 6805 2154 6817 2206
rect 6869 2154 6875 2206
rect 7301 1765 7353 1771
rect 7301 1701 7353 1713
rect 7163 1654 7215 1672
rect 7301 1643 7353 1649
rect 7163 1590 7215 1602
rect 7163 1532 7215 1538
tri 7647 1293 7653 1299 se
rect 7653 1293 7705 2571
tri 7705 2568 7708 2571 nw
tri 8013 1680 8033 1700 se
rect 8033 1680 8084 3827
tri 8084 3824 8087 3827 nw
rect 8921 3649 9079 3986
tri 9079 3945 9120 3986 nw
rect 9120 3843 9126 3895
rect 9178 3843 9190 3895
rect 9242 3843 9248 3895
rect 9365 3843 9371 3895
rect 9423 3843 9435 3895
rect 9487 3843 9493 3895
tri 9156 3829 9170 3843 ne
rect 9170 3829 9248 3843
tri 9416 3829 9430 3843 ne
rect 9430 3829 9493 3843
tri 9170 3827 9172 3829 ne
rect 9172 3827 9248 3829
tri 9430 3827 9432 3829 ne
rect 9432 3827 9493 3829
tri 9172 3818 9181 3827 ne
rect 8921 3597 8923 3649
rect 8975 3597 9027 3649
rect 8921 3580 9079 3597
rect 8921 3528 8923 3580
rect 8975 3528 9027 3580
rect 8921 3511 9079 3528
rect 8921 3459 8923 3511
rect 8975 3459 9027 3511
rect 8921 3453 9079 3459
rect 8416 3373 8422 3425
rect 8474 3373 8486 3425
rect 8538 3373 8544 3425
tri 8467 3369 8471 3373 ne
rect 8471 3369 8544 3373
tri 8471 3348 8492 3369 ne
tri 8467 2900 8492 2925 se
rect 8492 2900 8544 3369
rect 8983 3292 8989 3344
rect 9041 3292 9053 3344
rect 9105 3292 9111 3344
rect 8673 3086 8679 3138
rect 8731 3086 8743 3138
rect 8795 3086 8801 3138
rect 8983 3096 9111 3292
tri 9111 3096 9115 3100 sw
tri 8975 3088 8983 3096 se
rect 8983 3088 9115 3096
tri 9115 3088 9123 3096 sw
tri 8974 3087 8975 3088 se
rect 8975 3087 9123 3088
tri 8973 3086 8974 3087 se
rect 8974 3086 9123 3087
tri 8677 3076 8687 3086 ne
rect 8687 3076 8785 3086
tri 8785 3076 8795 3086 nw
tri 8972 3085 8973 3086 se
rect 8973 3085 9123 3086
tri 9123 3085 9126 3088 sw
tri 8687 3052 8711 3076 ne
rect 8225 2848 8231 2900
rect 8283 2848 8295 2900
rect 8347 2848 8353 2900
tri 8353 2848 8363 2858 sw
rect 8416 2848 8422 2900
rect 8474 2848 8486 2900
rect 8538 2848 8544 2900
tri 8289 2842 8295 2848 ne
rect 8295 2842 8363 2848
tri 8363 2842 8369 2848 sw
tri 8295 2832 8305 2842 ne
rect 8305 2832 8369 2842
tri 8369 2832 8379 2842 sw
tri 8305 2830 8307 2832 ne
rect 8307 2830 8379 2832
tri 8379 2830 8381 2832 sw
tri 8307 2826 8311 2830 ne
rect 8311 2826 8381 2830
tri 8381 2826 8385 2830 sw
tri 8311 2778 8359 2826 ne
rect 8359 2778 8385 2826
tri 8385 2778 8433 2826 sw
tri 8359 2772 8365 2778 ne
rect 8365 2772 8433 2778
tri 8433 2772 8439 2778 sw
tri 8365 2767 8370 2772 ne
rect 8370 2767 8439 2772
tri 8439 2767 8444 2772 sw
tri 8370 2754 8383 2767 ne
rect 8383 2754 8444 2767
tri 8444 2754 8457 2767 sw
tri 8383 2752 8385 2754 ne
rect 8385 2752 8457 2754
tri 8457 2752 8459 2754 sw
tri 8385 2750 8387 2752 ne
rect 8387 2750 8459 2752
tri 8387 2738 8399 2750 ne
rect 8399 2738 8459 2750
tri 8459 2738 8473 2752 sw
tri 8399 2725 8412 2738 ne
rect 8412 2725 8473 2738
tri 8412 2714 8423 2725 ne
rect 8423 2714 8473 2725
tri 8473 2714 8497 2738 sw
tri 8423 2693 8444 2714 ne
rect 8444 2693 8497 2714
tri 8444 2692 8445 2693 ne
rect 8445 2687 8497 2693
rect 8445 2623 8497 2635
rect 8445 2565 8497 2571
rect 8711 1757 8761 3076
tri 8761 3052 8785 3076 nw
rect 8972 3029 8981 3085
rect 9037 3029 9061 3085
rect 9117 3029 9126 3085
rect 9181 2658 9248 3827
tri 9432 3818 9441 3827 ne
rect 9276 3763 9282 3815
rect 9334 3763 9346 3815
rect 9398 3763 9404 3815
rect 9276 3760 9350 3763
tri 9350 3760 9353 3763 nw
rect 9276 3758 9348 3760
tri 9348 3758 9350 3760 nw
tri 9439 3758 9441 3760 se
rect 9441 3758 9493 3827
rect 9837 3775 9885 4045
rect 10001 3945 10053 4426
tri 10053 4421 10058 4426 nw
rect 10837 4253 10889 4259
rect 10837 4189 10889 4201
rect 10837 4131 10889 4137
tri 10837 4125 10843 4131 ne
rect 10001 3881 10053 3893
rect 10001 3823 10053 3829
tri 9885 3775 9892 3782 sw
rect 9837 3769 9892 3775
tri 9837 3758 9848 3769 ne
rect 9848 3758 9892 3769
tri 9892 3758 9909 3775 sw
rect 9276 2754 9328 3758
tri 9328 3738 9348 3758 nw
tri 9419 3738 9439 3758 se
rect 9439 3738 9493 3758
tri 9416 3735 9419 3738 se
rect 9419 3735 9493 3738
tri 9848 3735 9871 3758 ne
rect 9871 3735 9909 3758
rect 9365 3683 9371 3735
rect 9423 3683 9435 3735
rect 9487 3683 9493 3735
rect 9587 3683 9593 3735
rect 9645 3683 9659 3735
rect 9711 3721 9762 3735
tri 9762 3721 9776 3735 sw
tri 9871 3721 9885 3735 ne
rect 9885 3721 9909 3735
rect 9711 3704 9776 3721
tri 9776 3704 9793 3721 sw
tri 9885 3704 9902 3721 ne
rect 9902 3704 9909 3721
tri 9909 3704 9963 3758 sw
rect 9711 3697 9793 3704
tri 9793 3697 9800 3704 sw
tri 9902 3697 9909 3704 ne
rect 9909 3697 9963 3704
tri 9963 3697 9970 3704 sw
rect 9711 3683 9800 3697
tri 9800 3683 9814 3697 sw
tri 9909 3683 9923 3697 ne
rect 9923 3683 9970 3697
tri 9416 3658 9441 3683 ne
tri 9328 2754 9337 2763 sw
rect 9276 2738 9337 2754
tri 9337 2738 9353 2754 sw
rect 9276 2686 9282 2738
rect 9334 2686 9346 2738
rect 9398 2686 9404 2738
tri 9436 2678 9441 2683 se
rect 9441 2678 9493 3683
tri 9740 3680 9743 3683 ne
rect 9743 3680 9814 3683
tri 9814 3680 9817 3683 sw
tri 9923 3680 9926 3683 ne
rect 9926 3680 9970 3683
tri 9743 3661 9762 3680 ne
rect 9762 3661 9817 3680
tri 9762 3652 9771 3661 ne
rect 9771 3652 9817 3661
tri 9817 3652 9845 3680 sw
tri 9926 3652 9954 3680 ne
rect 9954 3652 9970 3680
tri 9970 3652 10015 3697 sw
tri 9771 3649 9774 3652 ne
rect 9774 3649 9845 3652
tri 9845 3649 9848 3652 sw
tri 9954 3649 9957 3652 ne
rect 9957 3649 10015 3652
tri 10015 3649 10018 3652 sw
tri 9774 3636 9787 3649 ne
rect 9787 3636 9848 3649
tri 9848 3636 9861 3649 sw
tri 9957 3636 9970 3649 ne
rect 9970 3636 10018 3649
tri 10018 3636 10031 3649 sw
tri 9787 3623 9800 3636 ne
rect 9800 3623 9861 3636
tri 9861 3623 9874 3636 sw
tri 9970 3623 9983 3636 ne
tri 9800 3606 9817 3623 ne
rect 9817 3606 9874 3623
tri 9874 3606 9891 3623 sw
tri 9817 3597 9826 3606 ne
rect 9826 3597 9891 3606
tri 9826 3586 9837 3597 ne
rect 9837 3586 9891 3597
tri 9837 3584 9839 3586 ne
tri 9829 3438 9839 3448 se
rect 9839 3438 9891 3586
tri 9891 3438 9901 3448 sw
tri 9816 3425 9829 3438 se
rect 9829 3425 9901 3438
tri 9431 2673 9436 2678 se
rect 9436 2673 9493 2678
tri 9422 2664 9431 2673 se
rect 9431 2664 9493 2673
tri 9248 2658 9254 2664 sw
tri 9416 2658 9422 2664 se
rect 9422 2658 9493 2664
rect 9181 2645 9254 2658
tri 9254 2645 9267 2658 sw
rect 9181 2637 9267 2645
tri 9267 2637 9275 2645 sw
tri 9181 2626 9192 2637 ne
rect 9192 2626 9275 2637
tri 9275 2626 9286 2637 sw
tri 9192 2606 9212 2626 ne
rect 9212 2606 9286 2626
tri 9286 2606 9306 2626 sw
rect 9365 2606 9371 2658
rect 9423 2606 9435 2658
rect 9487 2606 9493 2658
rect 9576 3373 9582 3425
rect 9634 3373 9646 3425
rect 9698 3373 9704 3425
tri 9812 3421 9816 3425 se
rect 9816 3421 9901 3425
tri 9901 3421 9918 3438 sw
rect 9576 3369 9661 3373
tri 9661 3369 9665 3373 nw
rect 9812 3369 9818 3421
rect 9870 3369 9882 3421
rect 9934 3369 9940 3421
rect 9576 2702 9640 3369
tri 9640 3348 9661 3369 nw
rect 9812 3348 9882 3369
tri 9882 3348 9903 3369 nw
rect 9812 3346 9880 3348
tri 9880 3346 9882 3348 nw
rect 9812 3344 9878 3346
tri 9878 3344 9880 3346 nw
rect 9812 3336 9870 3344
tri 9870 3336 9878 3344 nw
tri 9810 3334 9812 3336 se
rect 9812 3334 9868 3336
tri 9868 3334 9870 3336 nw
tri 9796 3320 9810 3334 se
rect 9810 3320 9854 3334
tri 9854 3320 9868 3334 nw
tri 9758 3282 9796 3320 se
rect 9796 3282 9816 3320
tri 9816 3282 9854 3320 nw
tri 9756 3280 9758 3282 se
rect 9758 3280 9814 3282
tri 9814 3280 9816 3282 nw
tri 9754 3278 9756 3280 se
rect 9756 3278 9812 3280
tri 9812 3278 9814 3280 nw
tri 9744 3268 9754 3278 se
rect 9754 3268 9802 3278
tri 9802 3268 9812 3278 nw
tri 9738 3262 9744 3268 se
rect 9744 3262 9796 3268
tri 9796 3262 9802 3268 nw
rect 9738 3252 9786 3262
tri 9786 3252 9796 3262 nw
rect 9738 3246 9780 3252
tri 9780 3246 9786 3252 nw
rect 9890 3246 9942 3252
rect 9738 3024 9778 3246
tri 9778 3244 9780 3246 nw
rect 9890 3182 9942 3194
tri 9778 3024 9779 3025 sw
rect 9738 3020 9779 3024
tri 9779 3020 9783 3024 sw
rect 9738 3012 9783 3020
tri 9783 3012 9791 3020 sw
rect 9738 3007 9791 3012
tri 9791 3007 9796 3012 sw
tri 9738 3000 9745 3007 ne
rect 9745 3000 9796 3007
tri 9796 3000 9803 3007 sw
tri 9745 2993 9752 3000 ne
rect 9752 2993 9803 3000
tri 9803 2993 9810 3000 sw
tri 9752 2972 9773 2993 ne
rect 9773 2972 9810 2993
tri 9810 2972 9831 2993 sw
rect 9890 2972 9942 3130
rect 9983 3048 10031 3636
rect 10619 3185 10625 3237
rect 10677 3185 10689 3237
rect 10741 3185 10747 3237
rect 10619 3175 10737 3185
tri 10737 3175 10747 3185 nw
rect 10619 3163 10725 3175
tri 10725 3163 10737 3175 nw
rect 10619 3111 10673 3163
tri 10673 3111 10725 3163 nw
tri 9983 3024 10007 3048 ne
rect 10007 3024 10031 3048
tri 10031 3024 10075 3068 sw
tri 10007 3020 10011 3024 ne
rect 10011 3020 10075 3024
tri 10075 3020 10079 3024 sw
tri 10011 3012 10019 3020 ne
rect 10019 3012 10140 3020
tri 10140 3012 10148 3020 sw
tri 10019 3000 10031 3012 ne
rect 10031 3000 10148 3012
tri 10031 2993 10038 3000 ne
rect 10038 2993 10148 3000
tri 10148 2993 10167 3012 sw
tri 10038 2990 10041 2993 ne
rect 10041 2990 10167 2993
tri 9942 2972 9960 2990 sw
tri 10041 2972 10059 2990 ne
rect 10059 2972 10167 2990
tri 9773 2966 9779 2972 ne
rect 9779 2966 9831 2972
tri 9831 2966 9837 2972 sw
rect 9890 2968 9960 2972
tri 9960 2968 9964 2972 sw
tri 10120 2968 10124 2972 ne
rect 10124 2968 10167 2972
tri 9890 2966 9892 2968 ne
rect 9892 2966 9964 2968
tri 9779 2960 9785 2966 ne
rect 9785 2960 9837 2966
tri 9837 2960 9843 2966 sw
tri 9892 2960 9898 2966 ne
rect 9898 2960 9964 2966
tri 9964 2960 9972 2968 sw
tri 10124 2960 10132 2968 ne
rect 10132 2960 10167 2968
tri 10167 2960 10200 2993 sw
tri 9785 2948 9797 2960 ne
rect 9797 2948 9843 2960
tri 9843 2948 9855 2960 sw
tri 9898 2948 9910 2960 ne
rect 9910 2948 9972 2960
tri 9972 2948 9984 2960 sw
tri 10132 2948 10144 2960 ne
rect 10144 2948 10200 2960
tri 10200 2948 10212 2960 sw
tri 9797 2925 9820 2948 ne
rect 9820 2926 9855 2948
tri 9855 2926 9877 2948 sw
rect 9820 2925 9877 2926
tri 9910 2925 9933 2948 ne
rect 9933 2925 9984 2948
tri 9984 2925 10007 2948 sw
tri 10144 2925 10167 2948 ne
rect 10167 2925 10212 2948
tri 10212 2925 10235 2948 sw
tri 9820 2922 9823 2925 ne
rect 9823 2922 9877 2925
tri 9933 2922 9936 2925 ne
rect 9936 2922 10007 2925
tri 10007 2922 10010 2925 sw
rect 10167 2922 10235 2925
tri 10235 2922 10238 2925 sw
tri 9823 2908 9837 2922 ne
rect 9668 2848 9674 2900
rect 9726 2848 9738 2900
rect 9790 2848 9796 2900
tri 9719 2842 9725 2848 ne
rect 9725 2842 9796 2848
tri 9725 2832 9735 2842 ne
rect 9735 2832 9796 2842
tri 9735 2830 9737 2832 ne
rect 9737 2830 9796 2832
tri 9737 2823 9744 2830 ne
tri 9640 2702 9641 2703 sw
rect 9576 2678 9641 2702
tri 9641 2678 9665 2702 sw
rect 9576 2626 9582 2678
rect 9634 2626 9646 2678
rect 9698 2626 9704 2678
tri 9212 2597 9221 2606 ne
rect 9221 2597 9306 2606
rect 8817 2545 8823 2597
rect 8875 2545 8887 2597
rect 8939 2545 8945 2597
tri 9221 2593 9225 2597 ne
rect 9225 2593 9306 2597
tri 9225 2569 9249 2593 ne
rect 9249 2569 9306 2593
tri 9306 2569 9343 2606 sw
tri 9249 2568 9250 2569 ne
rect 9250 2568 9343 2569
tri 8839 2522 8862 2545 ne
rect 8862 2522 8939 2545
tri 8939 2539 8945 2545 nw
tri 9250 2539 9279 2568 ne
rect 9279 2539 9343 2568
tri 9279 2522 9296 2539 ne
rect 9296 2522 9343 2539
tri 9343 2522 9390 2569 sw
tri 8862 2492 8892 2522 ne
rect 8892 2232 8939 2522
tri 9296 2475 9343 2522 ne
rect 9343 2475 9390 2522
tri 9390 2475 9437 2522 sw
tri 9343 2470 9348 2475 ne
rect 9348 2470 9437 2475
tri 9437 2470 9442 2475 sw
tri 9348 2458 9360 2470 ne
rect 9360 2458 9442 2470
tri 9442 2458 9454 2470 sw
tri 9360 2446 9372 2458 ne
rect 9372 2446 9454 2458
tri 9454 2446 9466 2458 sw
tri 9372 2419 9399 2446 ne
rect 9399 2419 9466 2446
tri 9466 2419 9493 2446 sw
tri 9399 2381 9437 2419 ne
rect 9437 2381 9493 2419
tri 9493 2381 9531 2419 sw
rect 9437 2367 9531 2381
tri 9531 2367 9545 2381 sw
rect 9437 2354 9545 2367
tri 9545 2354 9558 2367 sw
rect 9437 2347 9558 2354
tri 9558 2347 9565 2354 sw
rect 9437 2284 9565 2347
tri 8939 2232 8964 2257 sw
rect 9437 2232 9443 2284
rect 9495 2232 9507 2284
rect 9559 2232 9565 2284
rect 8892 2226 8964 2232
tri 8964 2226 8970 2232 sw
rect 8892 2223 8970 2226
tri 8970 2223 8973 2226 sw
rect 8892 2214 8973 2223
tri 8973 2214 8982 2223 sw
rect 8892 2204 8982 2214
tri 8982 2204 8992 2214 sw
rect 8892 2152 8898 2204
rect 8950 2152 8962 2204
rect 9014 2152 9020 2204
tri 8761 1757 8770 1766 sw
rect 8711 1744 8770 1757
tri 8770 1744 8783 1757 sw
tri 9731 1744 9744 1757 se
rect 9744 1744 9796 2830
rect 8711 1732 8783 1744
tri 8783 1732 8795 1744 sw
tri 9719 1732 9731 1744 se
rect 9731 1732 9796 1744
tri 8084 1680 8097 1693 sw
rect 8711 1680 8717 1732
rect 8769 1680 8806 1732
rect 8858 1680 8864 1732
rect 9013 1680 9019 1732
rect 9071 1680 9083 1732
rect 9135 1680 9141 1732
rect 9668 1680 9674 1732
rect 9726 1680 9738 1732
rect 9790 1680 9796 1732
tri 7997 1664 8013 1680 se
rect 8013 1664 8097 1680
tri 8097 1664 8113 1680 sw
tri 9013 1664 9029 1680 ne
rect 9029 1664 9125 1680
tri 9125 1664 9141 1680 nw
tri 9719 1664 9735 1680 ne
rect 9735 1664 9796 1680
tri 7991 1658 7997 1664 se
rect 7997 1658 8113 1664
tri 8113 1658 8119 1664 sw
rect 7991 1606 7997 1658
rect 8049 1606 8061 1658
rect 8113 1606 8119 1658
tri 9029 1652 9041 1664 ne
rect 9041 1652 9113 1664
tri 9113 1652 9125 1664 nw
tri 9735 1655 9744 1664 ne
tri 9041 1645 9048 1652 ne
tri 7629 1275 7647 1293 se
rect 7647 1275 7705 1293
tri 7628 1274 7629 1275 se
rect 7629 1274 7705 1275
rect 7577 1222 7583 1274
rect 7635 1222 7647 1274
rect 7699 1222 7705 1274
tri 4532 1198 4535 1201 se
rect 4535 1198 4594 1201
tri 4530 1196 4532 1198 se
rect 4532 1196 4594 1198
tri 4498 1164 4530 1196 se
rect 4530 1164 4594 1196
tri 4594 1164 4626 1196 sw
rect 4498 1112 4504 1164
rect 4556 1112 4568 1164
rect 4620 1112 4626 1164
rect 5472 1112 5478 1164
rect 5530 1112 5542 1164
rect 5594 1112 5600 1164
tri 5472 1105 5479 1112 ne
rect 5479 1105 5593 1112
tri 5593 1105 5600 1112 nw
tri 5479 1091 5493 1105 ne
rect 5493 1091 5579 1105
tri 5579 1091 5593 1105 nw
tri 5493 1087 5497 1091 ne
rect 5497 1087 5575 1091
tri 5575 1087 5579 1091 nw
tri 5497 1070 5514 1087 ne
rect 5514 1070 5575 1087
tri 5514 1065 5519 1070 ne
tri 5515 969 5519 973 se
rect 5519 969 5575 1070
tri 5514 968 5515 969 se
rect 5515 968 5575 969
tri 5505 959 5514 968 se
rect 5514 959 5575 968
tri 5497 951 5505 959 se
rect 5505 951 5575 959
tri 5491 945 5497 951 se
rect 5497 945 5575 951
tri 5575 945 5581 951 sw
tri 5486 940 5491 945 se
rect 5491 940 5581 945
tri 5581 940 5586 945 sw
rect 9048 940 9100 1652
tri 9100 1639 9113 1652 nw
rect 9429 1600 9435 1652
rect 9487 1600 9499 1652
rect 9551 1600 9557 1652
tri 9429 1590 9439 1600 ne
rect 9439 1590 9520 1600
tri 9520 1590 9530 1600 nw
tri 9439 1584 9445 1590 ne
rect 9445 1584 9514 1590
tri 9514 1584 9520 1590 nw
tri 9445 1565 9464 1584 ne
tri 9100 940 9104 944 sw
tri 5485 939 5486 940 se
rect 5486 939 5586 940
tri 5586 939 5587 940 sw
rect 9048 939 9104 940
tri 9104 939 9105 940 sw
tri 5484 938 5485 939 se
rect 5485 938 5587 939
tri 5587 938 5588 939 sw
tri 5472 926 5484 938 se
rect 5484 926 5588 938
tri 5588 926 5600 938 sw
rect 5472 874 5478 926
rect 5530 874 5542 926
rect 5594 874 5600 926
tri 9013 903 9048 938 se
rect 9048 903 9105 939
tri 9105 903 9141 939 sw
tri 9431 903 9464 936 se
rect 9464 903 9496 1584
tri 9496 1566 9514 1584 nw
rect 9585 1532 9591 1584
rect 9643 1532 9655 1584
rect 9707 1532 9713 1584
rect 9585 1498 9679 1532
tri 9679 1498 9713 1532 nw
tri 9560 1391 9585 1416 se
rect 9585 1391 9636 1498
tri 9636 1455 9679 1498 nw
rect 9013 851 9019 903
rect 9071 851 9085 903
rect 9137 851 9143 903
tri 9430 902 9431 903 se
rect 9431 902 9496 903
rect 9340 850 9346 902
rect 9398 850 9438 902
rect 9490 850 9496 902
tri 9554 1385 9560 1391 se
rect 9560 1385 9622 1391
rect 9554 1377 9622 1385
tri 9622 1377 9636 1391 nw
rect 9554 882 9608 1377
tri 9608 1363 9622 1377 nw
tri 9723 1253 9744 1274 se
rect 9744 1253 9796 1664
tri 9692 1222 9723 1253 se
rect 9723 1222 9796 1253
tri 9671 1201 9692 1222 se
rect 9692 1201 9796 1222
tri 9668 1198 9671 1201 se
rect 9671 1198 9796 1201
rect 9668 1146 9674 1198
rect 9726 1146 9738 1198
rect 9790 1146 9796 1198
tri 9668 1137 9677 1146 ne
rect 9677 1137 9796 1146
tri 9677 1133 9681 1137 ne
rect 9681 1133 9796 1137
tri 9681 1105 9709 1133 ne
rect 9709 1105 9796 1133
tri 9709 1091 9723 1105 ne
rect 9723 1091 9796 1105
tri 9723 1087 9727 1091 ne
rect 9727 1087 9796 1091
tri 9727 1070 9744 1087 ne
tri 9731 1002 9744 1015 se
rect 9744 1002 9796 1087
tri 9704 975 9731 1002 se
rect 9731 975 9796 1002
tri 9698 969 9704 975 se
rect 9704 969 9796 975
tri 9697 968 9698 969 se
rect 9698 968 9796 969
tri 9688 959 9697 968 se
rect 9697 959 9796 968
tri 9680 951 9688 959 se
rect 9688 951 9796 959
tri 9674 945 9680 951 se
rect 9680 945 9796 951
tri 9673 944 9674 945 se
rect 9674 944 9796 945
tri 9669 940 9673 944 se
rect 9673 940 9796 944
tri 9668 939 9669 940 se
rect 9669 939 9796 940
rect 9668 887 9674 939
rect 9726 887 9738 939
rect 9790 887 9796 939
tri 9608 882 9612 886 sw
rect 9554 879 9612 882
tri 9612 879 9615 882 sw
rect 9554 857 9615 879
tri 9615 857 9637 879 sw
rect 9554 805 9560 857
rect 9612 805 9624 857
rect 9676 805 9682 857
rect 986 738 992 790
rect 1044 738 1061 790
rect 1113 738 1130 790
rect 1182 738 1199 790
rect 1251 738 1268 790
rect 1320 738 1337 790
rect 1389 738 1405 790
rect 1457 738 1473 790
rect 1525 738 1531 790
rect 9837 767 9877 2922
tri 9936 2900 9958 2922 ne
rect 9958 2900 10010 2922
tri 10010 2900 10032 2922 sw
rect 10167 2900 10238 2922
tri 10238 2900 10260 2922 sw
tri 9958 2881 9977 2900 ne
rect 9977 2881 9988 2900
tri 9977 2876 9982 2881 ne
rect 9982 2848 9988 2881
rect 10040 2848 10052 2900
rect 10104 2848 10110 2900
rect 10167 2848 10173 2900
rect 10225 2848 10237 2900
rect 10289 2848 10295 2900
rect 10456 2470 10462 2522
rect 10514 2470 10526 2522
rect 10578 2470 10584 2522
tri 10507 2458 10519 2470 ne
rect 10519 2458 10584 2470
tri 10519 2446 10531 2458 ne
rect 10531 2446 10584 2458
tri 10531 2445 10532 2446 ne
tri 10530 2354 10532 2356 se
rect 10532 2354 10584 2446
tri 10522 2346 10530 2354 se
rect 10530 2346 10584 2354
tri 10510 2334 10522 2346 se
rect 10522 2334 10584 2346
tri 10478 2302 10510 2334 se
rect 10510 2302 10552 2334
tri 10552 2302 10584 2334 nw
tri 10470 2294 10478 2302 se
rect 10478 2294 10539 2302
rect 10470 2289 10539 2294
tri 10539 2289 10552 2302 nw
rect 10470 2278 10528 2289
tri 10528 2278 10539 2289 nw
rect 10470 2135 10522 2278
tri 10522 2272 10528 2278 nw
rect 10619 2234 10671 3111
tri 10671 3109 10673 3111 nw
rect 10843 2562 10889 4131
rect 11000 4109 11052 4115
rect 11000 4045 11052 4057
rect 11000 3987 11052 3993
rect 11000 3986 11051 3987
tri 11051 3986 11052 3987 nw
rect 11886 3986 11938 3992
rect 11000 3282 11046 3986
tri 11046 3981 11051 3986 nw
rect 11886 3922 11938 3934
rect 11886 3864 11938 3870
tri 11886 3845 11905 3864 ne
tri 11046 3282 11083 3319 sw
rect 11000 3280 11083 3282
tri 11083 3280 11085 3282 sw
rect 11000 3278 11085 3280
tri 11085 3278 11087 3280 sw
rect 11000 3268 11087 3278
tri 11087 3268 11097 3278 sw
rect 11000 3237 11097 3268
tri 11097 3237 11128 3268 sw
rect 11000 3185 11006 3237
rect 11058 3185 11070 3237
rect 11122 3185 11128 3237
tri 10889 2562 10898 2571 sw
rect 10843 2551 10898 2562
tri 10843 2522 10872 2551 ne
rect 10872 2522 10898 2551
tri 10898 2522 10938 2562 sw
tri 11865 2522 11905 2562 se
rect 11905 2522 11938 3864
rect 12073 2894 12125 5443
tri 12125 5409 12159 5443 nw
tri 12209 5409 12232 5432 se
rect 12232 5409 12284 5519
tri 12284 5512 12318 5546 nw
tri 12550 5521 12575 5546 se
rect 12575 5521 12624 5546
tri 12624 5521 12698 5595 nw
tri 12541 5512 12550 5521 se
tri 12476 5447 12541 5512 se
rect 12541 5447 12550 5512
tri 12550 5447 12624 5521 nw
tri 12461 5432 12476 5447 se
tri 12284 5409 12307 5432 sw
tri 12438 5409 12461 5432 se
rect 12461 5409 12476 5432
tri 12198 5398 12209 5409 se
rect 12209 5398 12307 5409
tri 12307 5398 12318 5409 sw
tri 12427 5398 12438 5409 se
rect 12438 5398 12476 5409
rect 12194 5346 12200 5398
rect 12252 5346 12264 5398
rect 12316 5346 12322 5398
tri 12402 5373 12427 5398 se
rect 12427 5373 12476 5398
tri 12476 5373 12550 5447 nw
tri 12375 5346 12402 5373 se
tri 12347 5318 12375 5346 se
rect 12375 5318 12402 5346
rect 12347 5299 12402 5318
tri 12402 5299 12476 5373 nw
rect 12347 4904 12399 5299
tri 12399 5296 12402 5299 nw
rect 12347 4835 12399 4852
rect 12347 4766 12399 4783
rect 12073 2830 12125 2842
rect 12073 2772 12125 2778
rect 12153 4585 12159 4637
rect 12211 4585 12224 4637
rect 12276 4585 12282 4637
rect 12153 4557 12214 4585
tri 12214 4557 12242 4585 nw
tri 11938 2522 11957 2541 sw
rect 10701 2470 10707 2522
rect 10759 2470 10771 2522
rect 10823 2470 10829 2522
tri 10872 2505 10889 2522 ne
rect 10889 2470 10895 2522
rect 10947 2470 10959 2522
rect 11011 2470 11017 2522
rect 11829 2470 11835 2522
rect 11887 2470 11899 2522
rect 11951 2470 11957 2522
tri 10752 2458 10764 2470 ne
rect 10764 2458 10829 2470
tri 11829 2458 11841 2470 ne
rect 11841 2458 11945 2470
tri 11945 2458 11957 2470 nw
tri 10764 2446 10776 2458 ne
rect 10776 2446 10829 2458
tri 11841 2447 11852 2458 ne
tri 10776 2445 10777 2446 ne
tri 10671 2234 10688 2251 sw
tri 10612 2226 10619 2233 se
rect 10619 2226 10688 2234
tri 10609 2223 10612 2226 se
rect 10612 2223 10688 2226
tri 10600 2214 10609 2223 se
rect 10609 2214 10688 2223
tri 10590 2204 10600 2214 se
rect 10600 2204 10688 2214
rect 10560 2152 10566 2204
rect 10618 2152 10630 2204
rect 10682 2152 10688 2204
tri 10603 2151 10604 2152 ne
rect 10604 2151 10688 2152
tri 10604 2150 10605 2151 ne
rect 10605 2150 10688 2151
tri 10522 2135 10537 2150 sw
tri 10605 2135 10620 2150 ne
rect 10620 2135 10688 2150
tri 10462 2124 10470 2132 se
rect 10470 2124 10537 2135
tri 10537 2124 10548 2135 sw
tri 10620 2124 10631 2135 ne
rect 10631 2124 10688 2135
rect 10462 2072 10468 2124
rect 10520 2072 10532 2124
rect 10584 2072 10590 2124
tri 10631 2118 10637 2124 ne
rect 10416 1794 10425 1850
rect 10481 1794 10505 1850
rect 10561 1794 10582 1850
tri 10500 1769 10525 1794 ne
rect 10525 1769 10582 1794
rect 10637 1769 10688 2124
tri 10688 1769 10693 1774 sw
tri 10525 1758 10536 1769 ne
rect 10367 1612 10373 1664
rect 10425 1612 10437 1664
rect 10489 1612 10495 1664
rect 10536 1626 10582 1769
tri 10612 1744 10637 1769 se
rect 10637 1744 10693 1769
tri 10693 1744 10718 1769 sw
rect 10612 1692 10618 1744
rect 10670 1692 10682 1744
rect 10734 1692 10740 1744
tri 10752 1664 10777 1689 se
rect 10777 1664 10829 2446
rect 11852 2446 11933 2458
tri 11933 2446 11945 2458 nw
rect 11852 2419 11906 2446
tri 11906 2419 11933 2446 nw
rect 11852 2278 11904 2419
tri 11904 2417 11906 2419 nw
rect 11852 2214 11904 2226
rect 10876 2151 10882 2203
rect 10934 2151 10946 2203
rect 10998 2151 11004 2203
tri 10876 2147 10880 2151 ne
rect 10880 2147 11000 2151
tri 11000 2147 11004 2151 nw
rect 11397 2187 11449 2193
tri 10880 2135 10892 2147 ne
rect 10892 2135 11000 2147
tri 10892 2116 10911 2135 ne
rect 10911 2116 11000 2135
tri 10911 2079 10948 2116 ne
tri 10582 1626 10602 1646 sw
tri 10536 1612 10550 1626 ne
rect 10550 1612 10602 1626
tri 10602 1612 10616 1626 sw
rect 10701 1612 10707 1664
rect 10759 1612 10771 1664
rect 10823 1612 10829 1664
tri 10943 1624 10948 1629 se
rect 10948 1624 11000 2116
rect 11852 2156 11904 2162
rect 11397 2116 11449 2135
rect 11397 1811 11449 2064
tri 11449 1811 11471 1833 sw
tri 11397 1737 11471 1811 ne
tri 11471 1744 11538 1811 sw
rect 11471 1737 11538 1744
tri 11538 1737 11545 1744 sw
tri 11471 1670 11538 1737 ne
rect 11538 1695 11545 1737
tri 11545 1695 11587 1737 sw
tri 10931 1612 10943 1624 se
rect 10943 1612 11000 1624
rect 11098 1654 11150 1660
tri 10418 1602 10428 1612 ne
rect 10428 1602 10495 1612
tri 10550 1602 10560 1612 ne
rect 10560 1602 10616 1612
tri 10616 1602 10626 1612 sw
tri 10921 1602 10931 1612 se
rect 10931 1602 11000 1612
tri 11000 1602 11013 1615 sw
tri 10428 1590 10440 1602 ne
rect 10440 1590 10495 1602
tri 10560 1598 10564 1602 ne
rect 10564 1598 10626 1602
tri 10626 1598 10630 1602 sw
tri 10917 1598 10921 1602 se
rect 10921 1598 11013 1602
tri 10564 1590 10572 1598 ne
rect 10572 1590 10630 1598
tri 10630 1590 10638 1598 sw
tri 10909 1590 10917 1598 se
rect 10917 1590 11013 1598
tri 11013 1590 11025 1602 sw
rect 11098 1590 11150 1602
tri 10440 1587 10443 1590 ne
rect 10443 1091 10495 1590
tri 10572 1584 10578 1590 ne
rect 10578 1584 10638 1590
tri 10638 1584 10644 1590 sw
tri 10903 1584 10909 1590 se
rect 10909 1584 11025 1590
tri 11025 1584 11031 1590 sw
tri 10578 1535 10627 1584 ne
rect 10627 1532 10633 1584
rect 10685 1532 10703 1584
rect 10755 1532 10773 1584
rect 10825 1532 10831 1584
tri 10721 1498 10755 1532 ne
rect 10755 1498 10831 1532
rect 10903 1532 10909 1584
rect 10961 1532 10973 1584
rect 11025 1532 11031 1584
tri 10903 1498 10937 1532 ne
rect 10937 1498 10997 1532
tri 10997 1498 11031 1532 nw
tri 10755 1496 10757 1498 ne
rect 10757 1496 10831 1498
tri 10937 1496 10939 1498 ne
tri 10757 1475 10778 1496 ne
tri 10429 1039 10443 1053 se
tri 10428 1038 10429 1039 se
rect 10429 1038 10495 1039
rect 10529 1053 10535 1105
rect 10587 1053 10599 1105
rect 10651 1053 10657 1105
tri 10529 1038 10544 1053 ne
rect 10544 1038 10642 1053
tri 10642 1038 10657 1053 nw
tri 10757 1038 10778 1059 se
rect 10778 1038 10831 1496
tri 10425 1035 10428 1038 se
rect 10428 1035 10495 1038
tri 10544 1035 10547 1038 ne
rect 10547 1035 10639 1038
tri 10639 1035 10642 1038 nw
tri 10754 1035 10757 1038 se
rect 10757 1035 10831 1038
tri 10420 1030 10425 1035 se
rect 10425 1030 10495 1035
tri 10547 1030 10552 1035 ne
tri 10417 1027 10420 1030 se
rect 10420 1027 10495 1030
tri 10404 1014 10417 1027 se
rect 10417 1014 10443 1027
tri 10314 1002 10326 1014 se
rect 10326 1002 10443 1014
tri 10294 982 10314 1002 se
rect 10314 982 10443 1002
rect 10294 975 10443 982
rect 10294 969 10495 975
rect 10552 1026 10630 1035
tri 10630 1026 10639 1035 nw
tri 10745 1026 10754 1035 se
rect 10754 1026 10831 1035
rect 10552 1021 10625 1026
tri 10625 1021 10630 1026 nw
tri 10740 1021 10745 1026 se
rect 10745 1021 10831 1026
rect 10294 968 10399 969
tri 10399 968 10400 969 nw
tri 10551 968 10552 969 se
rect 10552 968 10618 1021
tri 10618 1014 10625 1021 nw
rect 10702 969 10708 1021
rect 10760 969 10773 1021
rect 10825 969 10831 1021
rect 10294 959 10390 968
tri 10390 959 10399 968 nw
tri 10542 959 10551 968 se
rect 10551 959 10618 968
rect 10294 945 10376 959
tri 10376 945 10390 959 nw
tri 10528 945 10542 959 se
rect 10542 945 10618 959
rect 10294 940 10371 945
tri 10371 940 10376 945 nw
tri 10523 940 10528 945 se
rect 10528 940 10618 945
rect 10294 939 10370 940
tri 10370 939 10371 940 nw
tri 10522 939 10523 940 se
rect 10523 939 10618 940
rect 10294 802 10338 939
tri 10338 907 10370 939 nw
rect 10490 887 10496 939
rect 10548 887 10560 939
rect 10612 887 10618 939
rect 10737 888 10743 940
rect 10795 888 10807 940
rect 10859 888 10865 940
rect 10737 887 10842 888
tri 10842 887 10843 888 nw
rect 10737 882 10837 887
tri 10837 882 10842 887 nw
rect 10737 879 10834 882
tri 10834 879 10837 882 nw
rect 10737 857 10812 879
tri 10812 857 10834 879 nw
rect 10737 844 10799 857
tri 10799 844 10812 857 nw
tri 10734 841 10737 844 se
rect 10737 841 10796 844
tri 10796 841 10799 844 nw
tri 10713 820 10734 841 se
rect 10734 820 10744 841
tri 10338 802 10356 820 sw
tri 10695 802 10713 820 se
rect 10713 802 10744 820
tri 10294 789 10307 802 ne
rect 10307 791 10356 802
tri 10356 791 10367 802 sw
tri 10684 791 10695 802 se
rect 10695 791 10744 802
rect 10307 789 10744 791
tri 10744 789 10796 841 nw
tri 10934 789 10939 794 se
rect 10939 789 10991 1498
tri 10991 1492 10997 1498 nw
tri 10307 787 10309 789 ne
rect 10309 787 10742 789
tri 10742 787 10744 789 nw
tri 10932 787 10934 789 se
rect 10934 787 10991 789
tri 10309 782 10314 787 ne
rect 10314 782 10737 787
tri 10737 782 10742 787 nw
tri 10927 782 10932 787 se
rect 10932 782 10991 787
tri 10314 780 10316 782 ne
rect 10316 780 10735 782
tri 10735 780 10737 782 nw
tri 10925 780 10927 782 se
rect 10927 780 10991 782
tri 10316 768 10328 780 ne
rect 10328 768 10723 780
tri 10723 768 10735 780 nw
tri 10913 768 10925 780 se
rect 10925 768 10991 780
tri 11093 768 11098 773 se
rect 11098 768 11150 1538
tri 11506 888 11538 920 se
rect 11538 888 11587 1695
rect 12153 1090 12205 4557
tri 12205 4548 12214 4557 nw
rect 12347 4415 12399 4714
rect 12347 4350 12399 4363
rect 12233 4313 12285 4319
rect 12233 4249 12285 4261
rect 12233 3398 12285 4197
rect 12233 3334 12285 3346
rect 12233 3276 12285 3282
rect 12347 4285 12399 4298
rect 12347 4220 12399 4233
rect 12347 4155 12399 4168
rect 12347 4090 12399 4103
rect 12347 4025 12399 4038
rect 12347 3959 12399 3973
rect 12347 3893 12399 3907
rect 12347 3827 12399 3841
rect 12347 3649 12399 3775
rect 12347 3580 12399 3597
rect 13335 4939 13341 4991
rect 13393 4939 13413 4991
rect 13465 4939 13484 4991
rect 13536 4939 13555 4991
rect 13607 4939 13626 4991
rect 13678 4939 13684 4991
rect 13335 4916 13684 4939
rect 13335 4864 13341 4916
rect 13393 4864 13413 4916
rect 13465 4864 13484 4916
rect 13536 4864 13555 4916
rect 13607 4864 13626 4916
rect 13678 4864 13684 4916
rect 13335 4841 13684 4864
rect 13335 4789 13341 4841
rect 13393 4789 13413 4841
rect 13465 4789 13484 4841
rect 13536 4789 13555 4841
rect 13607 4789 13626 4841
rect 13678 4789 13684 4841
rect 13335 3704 13684 4789
rect 14684 4585 14690 4637
rect 14742 4585 14754 4637
rect 14806 4585 14812 4637
tri 14726 4557 14754 4585 ne
rect 14754 4557 14812 4585
rect 14585 4505 14591 4557
rect 14643 4505 14655 4557
rect 14707 4505 14713 4557
tri 14754 4551 14760 4557 ne
tri 14604 4474 14635 4505 ne
rect 14635 4100 14687 4505
tri 14687 4479 14713 4505 nw
tri 14726 3866 14760 3900 se
rect 14760 3866 14812 4557
rect 13335 3652 13338 3704
rect 13390 3652 13411 3704
rect 13463 3652 13484 3704
rect 13536 3652 13557 3704
rect 13609 3652 13630 3704
rect 13682 3652 13684 3704
rect 13335 3638 13684 3652
rect 13335 3586 13338 3638
rect 13390 3586 13411 3638
rect 13463 3586 13484 3638
rect 13536 3586 13557 3638
rect 13609 3586 13630 3638
rect 13682 3586 13684 3638
rect 13335 3572 13684 3586
rect 12347 3511 12399 3528
rect 12347 3396 12399 3459
rect 12347 3332 12399 3344
rect 12347 3268 12399 3280
rect 12235 3227 12287 3233
rect 12235 3163 12287 3175
rect 12235 1253 12287 3111
rect 12235 1189 12287 1201
rect 12235 1123 12287 1137
rect 12347 3204 12399 3216
rect 12347 3140 12399 3152
rect 12347 3076 12399 3088
rect 12347 3012 12399 3024
rect 12347 2948 12399 2960
rect 12347 2884 12399 2896
rect 12347 2819 12399 2832
rect 12347 2754 12399 2767
rect 12347 2419 12399 2702
rect 12886 3560 13216 3566
rect 12886 3508 12887 3560
rect 12939 3508 12956 3560
rect 13008 3508 13025 3560
rect 13077 3508 13094 3560
rect 13146 3508 13163 3560
rect 13215 3508 13216 3560
rect 12886 3490 13216 3508
rect 12886 3438 12887 3490
rect 12939 3438 12956 3490
rect 13008 3438 13025 3490
rect 13077 3438 13094 3490
rect 13146 3438 13163 3490
rect 13215 3438 13216 3490
rect 12886 3420 13216 3438
rect 12886 3368 12887 3420
rect 12939 3368 12956 3420
rect 13008 3368 13025 3420
rect 13077 3368 13094 3420
rect 13146 3368 13163 3420
rect 13215 3368 13216 3420
rect 12886 3349 13216 3368
rect 12886 3297 12887 3349
rect 12939 3297 12956 3349
rect 13008 3297 13025 3349
rect 13077 3297 13094 3349
rect 13146 3297 13163 3349
rect 13215 3297 13216 3349
rect 12886 3278 13216 3297
rect 12886 3226 12887 3278
rect 12939 3226 12956 3278
rect 13008 3226 13025 3278
rect 13077 3226 13094 3278
rect 13146 3226 13163 3278
rect 13215 3226 13216 3278
rect 12440 2510 12492 2516
rect 12440 2446 12492 2458
rect 12440 2388 12492 2394
rect 12347 2354 12399 2367
rect 12347 2289 12399 2302
rect 12347 2223 12399 2237
rect 12347 2157 12399 2171
rect 12347 2091 12399 2105
rect 12347 2025 12399 2039
rect 12347 1959 12399 1973
rect 12347 1893 12399 1907
rect 12347 1498 12399 1841
rect 12347 1429 12399 1446
rect 12347 1360 12399 1377
rect 12153 1026 12205 1038
rect 12153 968 12205 974
rect 12347 1087 12399 1308
rect 12886 1415 13216 3226
rect 13335 3520 13338 3572
rect 13390 3520 13411 3572
rect 13463 3520 13484 3572
rect 13536 3520 13557 3572
rect 13609 3520 13630 3572
rect 13682 3520 13684 3572
rect 13335 3506 13684 3520
rect 13335 3454 13338 3506
rect 13390 3454 13411 3506
rect 13463 3454 13484 3506
rect 13536 3454 13557 3506
rect 13609 3454 13630 3506
rect 13682 3454 13684 3506
rect 13335 3440 13684 3454
rect 13335 3388 13338 3440
rect 13390 3388 13411 3440
rect 13463 3388 13484 3440
rect 13536 3388 13557 3440
rect 13609 3388 13630 3440
rect 13682 3388 13684 3440
rect 13335 3374 13684 3388
rect 13335 3322 13338 3374
rect 13390 3322 13411 3374
rect 13463 3322 13484 3374
rect 13536 3322 13557 3374
rect 13609 3322 13630 3374
rect 13682 3322 13684 3374
rect 13335 3308 13684 3322
rect 13335 3256 13338 3308
rect 13390 3256 13411 3308
rect 13463 3256 13484 3308
rect 13536 3256 13557 3308
rect 13609 3256 13630 3308
rect 13682 3256 13684 3308
rect 13335 3242 13684 3256
rect 13335 3190 13338 3242
rect 13390 3190 13411 3242
rect 13463 3190 13484 3242
rect 13536 3190 13557 3242
rect 13609 3190 13630 3242
rect 13682 3190 13684 3242
rect 13335 3176 13684 3190
rect 13335 3124 13338 3176
rect 13390 3124 13411 3176
rect 13463 3124 13484 3176
rect 13536 3124 13557 3176
rect 13609 3124 13630 3176
rect 13682 3124 13684 3176
rect 13335 3118 13684 3124
rect 14554 3814 14812 3866
rect 14554 3038 14606 3814
tri 14606 3780 14640 3814 nw
rect 12886 1363 12887 1415
rect 12939 1363 12956 1415
rect 13008 1363 13025 1415
rect 13077 1363 13094 1415
rect 13146 1363 13163 1415
rect 13215 1363 13216 1415
rect 12886 1345 13216 1363
rect 12886 1293 12887 1345
rect 12939 1293 12956 1345
rect 13008 1293 13025 1345
rect 13077 1293 13094 1345
rect 13146 1293 13163 1345
rect 13215 1293 13216 1345
rect 12886 1275 13216 1293
rect 12886 1223 12887 1275
rect 12939 1223 12956 1275
rect 13008 1223 13025 1275
rect 13077 1223 13094 1275
rect 13146 1223 13163 1275
rect 13215 1223 13216 1275
rect 12886 1204 13216 1223
rect 12886 1152 12887 1204
rect 12939 1152 12956 1204
rect 13008 1152 13025 1204
rect 13077 1152 13094 1204
rect 13146 1152 13163 1204
rect 13215 1152 13216 1204
rect 12886 1133 13216 1152
rect 12886 1081 12887 1133
rect 12939 1081 12956 1133
rect 13008 1081 13025 1133
rect 13077 1081 13094 1133
rect 13146 1081 13163 1133
rect 13215 1081 13216 1133
rect 12886 1075 13216 1081
rect 12347 1011 12399 1035
tri 11505 887 11506 888 se
rect 11506 887 11587 888
tri 11500 882 11505 887 se
rect 11505 882 11587 887
tri 11497 879 11500 882 se
rect 11500 879 11587 882
tri 11475 857 11497 879 se
rect 11497 857 11587 879
tri 9877 767 9878 768 sw
tri 10328 767 10329 768 ne
rect 10329 767 10722 768
tri 10722 767 10723 768 nw
tri 10912 767 10913 768 se
rect 10913 767 10991 768
tri 11092 767 11093 768 se
rect 11093 767 11150 768
tri 9808 738 9837 767 se
rect 9837 738 9878 767
tri 9878 738 9907 767 sw
tri 10329 747 10349 767 ne
rect 10349 747 10702 767
tri 10702 747 10722 767 nw
tri 10892 747 10912 767 se
rect 10912 747 10991 767
tri 11072 747 11092 767 se
rect 11092 747 11150 767
tri 10883 738 10892 747 se
rect 10892 738 10991 747
rect 986 696 1531 738
rect 986 644 992 696
rect 1044 644 1061 696
rect 1113 644 1130 696
rect 1182 644 1199 696
rect 1251 644 1268 696
rect 1320 644 1337 696
rect 1389 644 1405 696
rect 1457 644 1473 696
rect 1525 644 1531 696
tri 9806 736 9808 738 se
rect 9808 736 9907 738
tri 9907 736 9909 738 sw
rect 9806 684 9812 736
rect 9864 684 9876 736
rect 9928 684 9934 736
rect 10863 686 10869 738
rect 10921 686 10933 738
rect 10985 686 10991 738
tri 11061 736 11072 747 se
rect 11072 736 11150 747
rect 11022 684 11028 736
rect 11080 684 11092 736
rect 11144 684 11150 736
tri 11459 841 11475 857 se
rect 11475 841 11587 857
rect 11459 789 11465 841
rect 11517 789 11529 841
rect 11581 789 11587 841
rect 12347 934 12399 959
rect 12347 857 12399 882
rect 986 643 1531 644
rect 11459 532 11587 789
rect 11459 480 11465 532
rect 11517 480 11529 532
rect 11581 480 11587 532
rect 12111 787 12117 839
rect 12169 787 12181 839
rect 12233 787 12239 839
rect 12111 782 12218 787
tri 12218 782 12223 787 nw
rect 12111 780 12216 782
tri 12216 780 12218 782 nw
rect 12347 780 12399 805
rect 12111 768 12204 780
tri 12204 768 12216 780 nw
rect 12111 767 12203 768
tri 12203 767 12204 768 nw
rect 12111 747 12183 767
tri 12183 747 12203 767 nw
rect 12111 736 12172 747
tri 12172 736 12183 747 nw
rect 12111 728 12164 736
tri 12164 728 12172 736 nw
rect 12111 722 12158 728
tri 12158 722 12164 728 nw
rect 12347 722 12399 728
rect 14823 997 14875 1003
rect 14823 931 14875 945
rect 12111 476 12157 722
tri 12157 721 12158 722 nw
rect 12255 591 12264 647
rect 12320 591 12344 647
rect 12400 592 12423 647
rect 12255 540 12363 591
rect 12415 540 12423 592
tri 14812 563 14823 574 se
rect 14823 563 14875 879
rect 12255 528 12423 540
tri 12157 476 12195 514 sw
rect 12255 504 12363 528
tri 12255 476 12283 504 ne
rect 12283 476 12363 504
rect 12415 476 12423 528
rect 12786 514 12812 563
tri 14789 540 14812 563 se
rect 14812 540 14875 563
rect 12111 424 12117 476
rect 12169 424 12181 476
rect 12233 424 12239 476
tri 12283 466 12293 476 ne
rect 12293 466 12423 476
tri 12764 424 12773 433 se
rect 12773 424 12825 505
rect 13257 485 13306 500
tri 12745 405 12764 424 se
rect 12764 411 12825 424
rect 12764 405 12819 411
tri 12819 405 12825 411 nw
tri -155 379 -129 405 se
rect -129 386 -74 405
rect -129 379 -123 386
tri -389 341 -351 379 se
rect -351 341 -315 379
tri -315 341 -277 379 nw
tri -193 341 -155 379 se
rect -155 341 -123 379
rect -389 340 -316 341
tri -316 340 -315 341 nw
tri -194 340 -193 341 se
rect -193 340 -123 341
rect -389 50 -333 340
tri -333 323 -316 340 nw
tri -197 337 -194 340 se
rect -194 337 -123 340
tri -123 337 -74 386 nw
rect 12334 379 12793 405
tri 12793 379 12819 405 nw
rect 12334 362 12767 379
rect -197 323 -137 337
tri -137 323 -123 337 nw
rect -389 -30 -333 -6
rect -389 -95 -333 -86
rect -197 -95 -145 323
tri -145 315 -137 323 nw
rect 12390 353 12767 362
tri 12767 353 12793 379 nw
rect 12390 341 12420 353
tri 12420 341 12432 353 nw
rect 12390 340 12419 341
tri 12419 340 12420 341 nw
rect 12390 323 12402 340
tri 12402 323 12419 340 nw
tri 13238 323 13255 340 se
rect 13255 323 13307 485
rect 13425 445 13474 498
rect 14747 488 14753 540
rect 14805 488 14817 540
rect 14869 488 14875 540
rect 13617 397 13652 442
rect 13789 394 13823 443
rect 14263 399 14307 448
tri 12390 311 12402 323 nw
tri 13226 311 13238 323 se
rect 13238 318 13307 323
rect 13238 311 13296 318
tri 13222 307 13226 311 se
rect 13226 307 13296 311
tri 13296 307 13307 318 nw
rect 12334 282 12390 306
rect 12428 255 12434 307
rect 12486 255 12498 307
rect 12550 255 13244 307
tri 13244 255 13296 307 nw
rect 12334 217 12390 226
tri -145 -95 -124 -74 sw
rect -197 -96 -124 -95
tri -124 -96 -123 -95 sw
tri -197 -170 -123 -96 ne
tri -123 -155 -64 -96 sw
rect -123 -170 -64 -155
tri -64 -170 -49 -155 sw
tri -123 -213 -80 -170 ne
rect -80 -207 -49 -170
tri -49 -207 -12 -170 sw
rect -80 -213 -12 -207
tri -80 -229 -64 -213 ne
tri -138 -1219 -64 -1145 se
rect -64 -1167 -12 -213
tri 11400 -315 11502 -213 sw
rect 11348 -371 11357 -315
rect 11413 -371 11437 -315
rect 11493 -371 11502 -315
tri 11400 -473 11502 -371 nw
tri -64 -1219 -12 -1167 nw
tri -197 -1278 -138 -1219 se
rect -138 -1278 -123 -1219
tri -123 -1278 -64 -1219 nw
rect -197 -1529 -145 -1278
tri -145 -1300 -123 -1278 nw
tri -145 -1529 -99 -1483 sw
tri -200 -1532 -197 -1529 se
rect -197 -1532 -99 -1529
tri -99 -1532 -96 -1529 sw
rect -200 -1588 -191 -1532
rect -135 -1588 -111 -1532
rect -55 -1588 -46 -1532
<< via2 >>
rect -267 4688 -211 4709
rect -267 4653 -230 4688
rect -230 4653 -218 4688
rect -218 4653 -211 4688
rect -267 4573 -211 4629
rect -374 631 -318 687
rect -374 551 -318 607
rect 136 3643 192 3666
rect 136 3610 139 3643
rect 139 3610 191 3643
rect 191 3610 192 3643
rect 136 3579 192 3586
rect 136 3530 139 3579
rect 139 3530 191 3579
rect 191 3530 192 3579
rect 3154 3979 3156 3987
rect 3156 3979 3208 3987
rect 3208 3979 3210 3987
rect 3250 3979 3272 3987
rect 3272 3979 3284 3987
rect 3284 3979 3306 3987
rect 3346 3979 3348 3987
rect 3348 3979 3400 3987
rect 3400 3979 3402 3987
rect 3442 3979 3464 3987
rect 3464 3979 3476 3987
rect 3476 3979 3498 3987
rect 3538 3979 3540 3987
rect 3540 3979 3592 3987
rect 3592 3979 3594 3987
rect 3154 3931 3210 3979
rect 3250 3931 3306 3979
rect 3346 3931 3402 3979
rect 3442 3931 3498 3979
rect 3538 3931 3594 3979
rect 3154 3850 3210 3906
rect 3250 3850 3306 3906
rect 3346 3850 3402 3906
rect 3442 3850 3498 3906
rect 3538 3850 3594 3906
rect 3154 3769 3210 3825
rect 3250 3769 3306 3825
rect 3346 3769 3402 3825
rect 3442 3769 3498 3825
rect 3538 3769 3594 3825
rect 3154 3688 3210 3744
rect 3250 3688 3306 3744
rect 3346 3688 3402 3744
rect 3442 3688 3498 3744
rect 3538 3688 3594 3744
rect 3154 3607 3210 3663
rect 3250 3607 3306 3663
rect 3346 3607 3402 3663
rect 3442 3607 3498 3663
rect 3538 3607 3594 3663
rect 3154 3526 3210 3582
rect 3250 3526 3306 3582
rect 3346 3526 3402 3582
rect 3442 3526 3498 3582
rect 3538 3526 3594 3582
rect 3154 3445 3210 3501
rect 3250 3445 3306 3501
rect 3346 3445 3402 3501
rect 3442 3445 3498 3501
rect 3538 3445 3594 3501
rect 3154 3364 3210 3420
rect 3250 3364 3306 3420
rect 3346 3364 3402 3420
rect 3442 3364 3498 3420
rect 3538 3364 3594 3420
rect 3154 3283 3210 3339
rect 3250 3283 3306 3339
rect 3346 3283 3402 3339
rect 3442 3283 3498 3339
rect 3538 3283 3594 3339
rect 3154 3202 3210 3258
rect 3250 3202 3306 3258
rect 3346 3202 3402 3258
rect 3442 3202 3498 3258
rect 3538 3202 3594 3258
rect 3154 3121 3210 3177
rect 3250 3121 3306 3177
rect 3346 3121 3402 3177
rect 3442 3121 3498 3177
rect 3538 3121 3594 3177
rect 3154 3057 3210 3096
rect 3250 3057 3306 3096
rect 3346 3057 3402 3096
rect 3442 3057 3498 3096
rect 3538 3057 3594 3096
rect 3154 3040 3156 3057
rect 3156 3040 3208 3057
rect 3208 3040 3210 3057
rect 3250 3040 3272 3057
rect 3272 3040 3284 3057
rect 3284 3040 3306 3057
rect 3346 3040 3348 3057
rect 3348 3040 3400 3057
rect 3400 3040 3402 3057
rect 3442 3040 3464 3057
rect 3464 3040 3476 3057
rect 3476 3040 3498 3057
rect 3538 3040 3540 3057
rect 3540 3040 3592 3057
rect 3592 3040 3594 3057
rect 3154 3005 3156 3015
rect 3156 3005 3208 3015
rect 3208 3005 3210 3015
rect 3250 3005 3272 3015
rect 3272 3005 3284 3015
rect 3284 3005 3306 3015
rect 3346 3005 3348 3015
rect 3348 3005 3400 3015
rect 3400 3005 3402 3015
rect 3442 3005 3464 3015
rect 3464 3005 3476 3015
rect 3476 3005 3498 3015
rect 3538 3005 3540 3015
rect 3540 3005 3592 3015
rect 3592 3005 3594 3015
rect 3154 2981 3210 3005
rect 3250 2981 3306 3005
rect 3346 2981 3402 3005
rect 3442 2981 3498 3005
rect 3538 2981 3594 3005
rect 3154 2959 3156 2981
rect 3156 2959 3208 2981
rect 3208 2959 3210 2981
rect 3250 2959 3272 2981
rect 3272 2959 3284 2981
rect 3284 2959 3306 2981
rect 3346 2959 3348 2981
rect 3348 2959 3400 2981
rect 3400 2959 3402 2981
rect 3442 2959 3464 2981
rect 3464 2959 3476 2981
rect 3476 2959 3498 2981
rect 3538 2959 3540 2981
rect 3540 2959 3592 2981
rect 3592 2959 3594 2981
rect 3154 2929 3156 2934
rect 3156 2929 3208 2934
rect 3208 2929 3210 2934
rect 3250 2929 3272 2934
rect 3272 2929 3284 2934
rect 3284 2929 3306 2934
rect 3346 2929 3348 2934
rect 3348 2929 3400 2934
rect 3400 2929 3402 2934
rect 3442 2929 3464 2934
rect 3464 2929 3476 2934
rect 3476 2929 3498 2934
rect 3538 2929 3540 2934
rect 3540 2929 3592 2934
rect 3592 2929 3594 2934
rect 3154 2878 3210 2929
rect 3250 2878 3306 2929
rect 3346 2878 3402 2929
rect 3442 2878 3498 2929
rect 3538 2878 3594 2929
rect 3154 2797 3210 2853
rect 3250 2797 3306 2853
rect 3346 2797 3402 2853
rect 3442 2797 3498 2853
rect 3538 2797 3594 2853
rect 3154 2716 3210 2772
rect 3250 2716 3306 2772
rect 3346 2716 3402 2772
rect 3442 2716 3498 2772
rect 3538 2716 3594 2772
rect 3154 2635 3210 2691
rect 3250 2635 3306 2691
rect 3346 2635 3402 2691
rect 3442 2635 3498 2691
rect 3538 2635 3594 2691
rect 3154 2554 3210 2610
rect 3250 2554 3306 2610
rect 3346 2554 3402 2610
rect 3442 2554 3498 2610
rect 3538 2554 3594 2610
rect 3154 2473 3210 2529
rect 3250 2473 3306 2529
rect 3346 2473 3402 2529
rect 3442 2473 3498 2529
rect 3538 2473 3594 2529
rect 3154 2442 3210 2447
rect 3250 2442 3306 2447
rect 3346 2442 3402 2447
rect 3442 2442 3498 2447
rect 3538 2442 3594 2447
rect 3154 2391 3156 2442
rect 3156 2391 3208 2442
rect 3208 2391 3210 2442
rect 3250 2391 3272 2442
rect 3272 2391 3284 2442
rect 3284 2391 3306 2442
rect 3346 2391 3348 2442
rect 3348 2391 3400 2442
rect 3400 2391 3402 2442
rect 3442 2391 3464 2442
rect 3464 2391 3476 2442
rect 3476 2391 3498 2442
rect 3538 2391 3540 2442
rect 3540 2391 3592 2442
rect 3592 2391 3594 2442
rect 3154 2364 3210 2365
rect 3250 2364 3306 2365
rect 3346 2364 3402 2365
rect 3442 2364 3498 2365
rect 3538 2364 3594 2365
rect 3154 2312 3156 2364
rect 3156 2312 3208 2364
rect 3208 2312 3210 2364
rect 3250 2312 3272 2364
rect 3272 2312 3284 2364
rect 3284 2312 3306 2364
rect 3346 2312 3348 2364
rect 3348 2312 3400 2364
rect 3400 2312 3402 2364
rect 3442 2312 3464 2364
rect 3464 2312 3476 2364
rect 3476 2312 3498 2364
rect 3538 2312 3540 2364
rect 3540 2312 3592 2364
rect 3592 2312 3594 2364
rect 3154 2309 3210 2312
rect 3250 2309 3306 2312
rect 3346 2309 3402 2312
rect 3442 2309 3498 2312
rect 3538 2309 3594 2312
rect 3154 2227 3210 2283
rect 3250 2227 3306 2283
rect 3346 2227 3402 2283
rect 3442 2227 3498 2283
rect 3538 2227 3594 2283
rect 3154 2145 3210 2201
rect 3250 2145 3306 2201
rect 3346 2145 3402 2201
rect 3442 2145 3498 2201
rect 3538 2145 3594 2201
rect 3154 2063 3210 2119
rect 3250 2063 3306 2119
rect 3346 2063 3402 2119
rect 3442 2063 3498 2119
rect 3538 2063 3594 2119
rect 3154 2029 3210 2037
rect 3250 2029 3306 2037
rect 3346 2029 3402 2037
rect 3442 2029 3498 2037
rect 3538 2029 3594 2037
rect 3154 1981 3156 2029
rect 3156 1981 3208 2029
rect 3208 1981 3210 2029
rect 3250 1981 3272 2029
rect 3272 1981 3284 2029
rect 3284 1981 3306 2029
rect 3346 1981 3348 2029
rect 3348 1981 3400 2029
rect 3400 1981 3402 2029
rect 3442 1981 3464 2029
rect 3464 1981 3476 2029
rect 3476 1981 3498 2029
rect 3538 1981 3540 2029
rect 3540 1981 3592 2029
rect 3592 1981 3594 2029
rect 3154 1903 3156 1955
rect 3156 1903 3208 1955
rect 3208 1903 3210 1955
rect 3250 1903 3272 1955
rect 3272 1903 3284 1955
rect 3284 1903 3306 1955
rect 3346 1903 3348 1955
rect 3348 1903 3400 1955
rect 3400 1903 3402 1955
rect 3442 1903 3464 1955
rect 3464 1903 3476 1955
rect 3476 1903 3498 1955
rect 3538 1903 3540 1955
rect 3540 1903 3592 1955
rect 3592 1903 3594 1955
rect 3154 1899 3210 1903
rect 3250 1899 3306 1903
rect 3346 1899 3402 1903
rect 3442 1899 3498 1903
rect 3538 1899 3594 1903
rect 3154 1829 3156 1873
rect 3156 1829 3208 1873
rect 3208 1829 3210 1873
rect 3250 1829 3272 1873
rect 3272 1829 3284 1873
rect 3284 1829 3306 1873
rect 3346 1829 3348 1873
rect 3348 1829 3400 1873
rect 3400 1829 3402 1873
rect 3442 1829 3464 1873
rect 3464 1829 3476 1873
rect 3476 1829 3498 1873
rect 3538 1829 3540 1873
rect 3540 1829 3592 1873
rect 3592 1829 3594 1873
rect 3154 1817 3210 1829
rect 3250 1817 3306 1829
rect 3346 1817 3402 1829
rect 3442 1817 3498 1829
rect 3538 1817 3594 1829
rect 3154 1735 3210 1791
rect 3250 1735 3306 1791
rect 3346 1735 3402 1791
rect 3442 1735 3498 1791
rect 3538 1735 3594 1791
rect 3154 1653 3210 1709
rect 3250 1653 3306 1709
rect 3346 1653 3402 1709
rect 3442 1653 3498 1709
rect 3538 1653 3594 1709
rect 8981 3029 9037 3085
rect 9061 3029 9117 3085
rect 10425 1794 10481 1850
rect 10505 1794 10561 1850
rect 12264 591 12320 647
rect 12344 592 12400 647
rect 12344 591 12363 592
rect 12363 591 12400 592
rect -389 -6 -333 50
rect -389 -86 -333 -30
rect 12334 306 12390 362
rect 12334 226 12390 282
rect 11357 -371 11413 -315
rect 11437 -371 11493 -315
rect -191 -1588 -135 -1532
rect -111 -1588 -55 -1532
<< metal3 >>
rect -272 4709 -206 4714
rect -272 4653 -267 4709
rect -211 4653 -206 4709
rect -272 4629 -206 4653
rect -272 4573 -267 4629
rect -211 4573 -206 4629
rect -272 3128 -206 4573
rect 3146 3987 3602 3992
rect 3146 3931 3154 3987
rect 3210 3931 3250 3987
rect 3306 3931 3346 3987
rect 3402 3931 3442 3987
rect 3498 3931 3538 3987
rect 3594 3931 3602 3987
rect 3146 3906 3602 3931
rect 3146 3850 3154 3906
rect 3210 3850 3250 3906
rect 3306 3850 3346 3906
rect 3402 3850 3442 3906
rect 3498 3850 3538 3906
rect 3594 3850 3602 3906
rect 3146 3825 3602 3850
rect 3146 3769 3154 3825
rect 3210 3769 3250 3825
rect 3306 3769 3346 3825
rect 3402 3769 3442 3825
rect 3498 3769 3538 3825
rect 3594 3769 3602 3825
rect 3146 3744 3602 3769
rect 3146 3688 3154 3744
rect 3210 3688 3250 3744
rect 3306 3688 3346 3744
rect 3402 3688 3442 3744
rect 3498 3688 3538 3744
rect 3594 3688 3602 3744
rect 131 3666 197 3671
rect 131 3610 136 3666
rect 192 3610 197 3666
rect 131 3586 197 3610
rect 131 3530 136 3586
rect 192 3530 197 3586
tri -206 3128 -192 3142 sw
tri -279 3121 -272 3128 se
rect -272 3121 -192 3128
tri -192 3121 -185 3128 sw
tri -304 3096 -279 3121 se
rect -279 3096 -185 3121
tri -185 3096 -160 3121 sw
tri -310 3090 -304 3096 se
rect -304 3090 -160 3096
tri -160 3090 -154 3096 sw
rect -310 3026 -304 3090
rect -240 3026 -224 3090
rect -160 3026 -154 3090
tri 81 1899 131 1949 se
rect 131 1899 197 3530
tri 55 1873 81 1899 se
rect 81 1873 197 1899
tri 41 1859 55 1873 se
rect 55 1859 197 1873
rect 41 1795 47 1859
rect 111 1795 127 1859
rect 191 1795 197 1859
rect 3146 3663 3602 3688
rect 3146 3607 3154 3663
rect 3210 3607 3250 3663
rect 3306 3607 3346 3663
rect 3402 3607 3442 3663
rect 3498 3607 3538 3663
rect 3594 3607 3602 3663
rect 3146 3582 3602 3607
rect 3146 3526 3154 3582
rect 3210 3526 3250 3582
rect 3306 3526 3346 3582
rect 3402 3526 3442 3582
rect 3498 3526 3538 3582
rect 3594 3526 3602 3582
rect 3146 3501 3602 3526
rect 3146 3445 3154 3501
rect 3210 3445 3250 3501
rect 3306 3445 3346 3501
rect 3402 3445 3442 3501
rect 3498 3445 3538 3501
rect 3594 3445 3602 3501
rect 3146 3420 3602 3445
rect 3146 3364 3154 3420
rect 3210 3364 3250 3420
rect 3306 3364 3346 3420
rect 3402 3364 3442 3420
rect 3498 3364 3538 3420
rect 3594 3364 3602 3420
rect 3146 3339 3602 3364
rect 3146 3283 3154 3339
rect 3210 3283 3250 3339
rect 3306 3283 3346 3339
rect 3402 3283 3442 3339
rect 3498 3283 3538 3339
rect 3594 3283 3602 3339
rect 3146 3258 3602 3283
rect 3146 3202 3154 3258
rect 3210 3202 3250 3258
rect 3306 3202 3346 3258
rect 3402 3202 3442 3258
rect 3498 3202 3538 3258
rect 3594 3202 3602 3258
rect 3146 3177 3602 3202
rect 3146 3121 3154 3177
rect 3210 3121 3250 3177
rect 3306 3121 3346 3177
rect 3402 3121 3442 3177
rect 3498 3121 3538 3177
rect 3594 3121 3602 3177
rect 3146 3096 3602 3121
rect 3146 3040 3154 3096
rect 3210 3040 3250 3096
rect 3306 3040 3346 3096
rect 3402 3040 3442 3096
rect 3498 3040 3538 3096
rect 3594 3040 3602 3096
rect 3146 3015 3602 3040
rect 8960 3026 8971 3090
rect 9035 3085 9051 3090
rect 9115 3085 9122 3090
rect 9037 3029 9051 3085
rect 9117 3029 9122 3085
rect 9035 3026 9051 3029
rect 9115 3026 9122 3029
rect 8960 3024 9122 3026
rect 3146 2959 3154 3015
rect 3210 2959 3250 3015
rect 3306 2959 3346 3015
rect 3402 2959 3442 3015
rect 3498 2959 3538 3015
rect 3594 2959 3602 3015
rect 3146 2934 3602 2959
rect 3146 2554 3154 2934
rect 3210 2895 3250 2934
rect 3306 2895 3346 2934
rect 3402 2895 3442 2934
rect 3498 2895 3538 2934
rect 3218 2831 3248 2895
rect 3312 2831 3342 2895
rect 3406 2831 3436 2895
rect 3500 2831 3530 2895
rect 3210 2809 3250 2831
rect 3306 2809 3346 2831
rect 3402 2809 3442 2831
rect 3498 2809 3538 2831
rect 3218 2745 3248 2809
rect 3312 2745 3342 2809
rect 3406 2745 3436 2809
rect 3500 2745 3530 2809
rect 3210 2723 3250 2745
rect 3306 2723 3346 2745
rect 3402 2723 3442 2745
rect 3498 2723 3538 2745
rect 3218 2659 3248 2723
rect 3312 2659 3342 2723
rect 3406 2659 3436 2723
rect 3500 2659 3530 2723
rect 3210 2637 3250 2659
rect 3306 2637 3346 2659
rect 3402 2637 3442 2659
rect 3498 2637 3538 2659
rect 3218 2573 3248 2637
rect 3312 2573 3342 2637
rect 3406 2573 3436 2637
rect 3500 2573 3530 2637
rect 3210 2554 3250 2573
rect 3306 2554 3346 2573
rect 3402 2554 3442 2573
rect 3498 2554 3538 2573
rect 3594 2554 3602 2934
rect 3146 2551 3602 2554
rect 3146 2473 3154 2551
rect 3218 2487 3248 2551
rect 3312 2487 3342 2551
rect 3406 2487 3436 2551
rect 3500 2487 3530 2551
rect 3210 2473 3250 2487
rect 3306 2473 3346 2487
rect 3402 2473 3442 2487
rect 3498 2473 3538 2487
rect 3594 2473 3602 2551
rect 3146 2465 3602 2473
rect 3146 2391 3154 2465
rect 3218 2401 3248 2465
rect 3312 2401 3342 2465
rect 3406 2401 3436 2465
rect 3500 2401 3530 2465
rect 3210 2391 3250 2401
rect 3306 2391 3346 2401
rect 3402 2391 3442 2401
rect 3498 2391 3538 2401
rect 3594 2391 3602 2465
rect 3146 2379 3602 2391
rect 3146 2309 3154 2379
rect 3218 2315 3248 2379
rect 3312 2315 3342 2379
rect 3406 2315 3436 2379
rect 3500 2315 3530 2379
rect 3210 2309 3250 2315
rect 3306 2309 3346 2315
rect 3402 2309 3442 2315
rect 3498 2309 3538 2315
rect 3594 2309 3602 2379
rect 3146 2292 3602 2309
rect 3146 2227 3154 2292
rect 3218 2228 3248 2292
rect 3312 2228 3342 2292
rect 3406 2228 3436 2292
rect 3500 2228 3530 2292
rect 3210 2227 3250 2228
rect 3306 2227 3346 2228
rect 3402 2227 3442 2228
rect 3498 2227 3538 2228
rect 3594 2227 3602 2292
rect 3146 2205 3602 2227
rect 3146 2141 3154 2205
rect 3218 2141 3248 2205
rect 3312 2141 3342 2205
rect 3406 2141 3436 2205
rect 3500 2141 3530 2205
rect 3594 2141 3602 2205
rect 3146 2119 3602 2141
rect 3146 2054 3154 2119
rect 3210 2118 3250 2119
rect 3306 2118 3346 2119
rect 3402 2118 3442 2119
rect 3498 2118 3538 2119
rect 3218 2054 3248 2118
rect 3312 2054 3342 2118
rect 3406 2054 3436 2118
rect 3500 2054 3530 2118
rect 3594 2054 3602 2119
rect 3146 2037 3602 2054
rect 3146 1967 3154 2037
rect 3210 2031 3250 2037
rect 3306 2031 3346 2037
rect 3402 2031 3442 2037
rect 3498 2031 3538 2037
rect 3218 1967 3248 2031
rect 3312 1967 3342 2031
rect 3406 1967 3436 2031
rect 3500 1967 3530 2031
rect 3594 1967 3602 2037
rect 3146 1955 3602 1967
rect 3146 1899 3154 1955
rect 3210 1899 3250 1955
rect 3306 1899 3346 1955
rect 3402 1899 3442 1955
rect 3498 1899 3538 1955
rect 3594 1899 3602 1955
rect 3146 1873 3602 1899
rect 3146 1817 3154 1873
rect 3210 1817 3250 1873
rect 3306 1817 3346 1873
rect 3402 1817 3442 1873
rect 3498 1817 3538 1873
rect 3594 1817 3602 1873
rect 3146 1791 3602 1817
rect 10410 1795 10416 1859
rect 10480 1850 10496 1859
rect 10560 1850 10566 1859
rect 10481 1795 10496 1850
rect 3146 1735 3154 1791
rect 3210 1735 3250 1791
rect 3306 1735 3346 1791
rect 3402 1735 3442 1791
rect 3498 1735 3538 1791
rect 3594 1735 3602 1791
rect 10420 1794 10425 1795
rect 10481 1794 10505 1795
rect 10561 1794 10566 1850
rect 10420 1789 10566 1794
rect 3146 1709 3602 1735
rect 3146 1653 3154 1709
rect 3210 1653 3250 1709
rect 3306 1653 3346 1709
rect 3402 1653 3442 1709
rect 3498 1653 3538 1709
rect 3594 1653 3602 1709
rect 3146 1648 3602 1653
rect -413 687 -257 692
rect -413 650 -374 687
rect -318 650 -257 687
rect -413 586 -407 650
rect -343 607 -327 631
rect -263 586 -257 650
rect 12249 650 12405 652
rect 12249 586 12255 650
rect 12319 647 12335 650
rect 12399 647 12405 650
rect 12320 591 12335 647
rect 12400 591 12405 647
rect 12319 586 12335 591
rect 12399 586 12405 591
rect -413 551 -374 586
rect -318 551 -257 586
rect -413 545 -257 551
rect 12329 362 12395 367
rect 12329 306 12334 362
rect 12390 306 12395 362
rect 12329 282 12395 306
rect 12329 226 12334 282
rect 12390 226 12395 282
rect -394 50 -328 55
rect -394 -6 -389 50
rect -333 -6 -328 50
rect -394 -30 -328 -6
rect -394 -86 -389 -30
rect -333 -86 -328 -30
tri -412 -273 -394 -255 se
rect -394 -273 -328 -86
tri -448 -309 -412 -273 se
rect -412 -309 -328 -273
tri -328 -309 -292 -273 sw
rect -448 -373 -442 -309
rect -378 -373 -362 -309
rect -298 -373 -292 -309
rect 11348 -373 11357 -309
rect 11421 -373 11437 -309
rect 11501 -373 11516 -309
rect 11348 -376 11516 -373
tri 12240 -1527 12329 -1438 se
rect 12329 -1527 12395 226
rect -204 -1528 -47 -1527
rect -204 -1592 -198 -1528
rect -134 -1592 -118 -1528
rect -54 -1592 -47 -1528
tri 12239 -1528 12240 -1527 se
rect 12240 -1528 12395 -1527
rect 12239 -1592 12245 -1528
rect 12309 -1592 12325 -1528
rect 12389 -1592 12395 -1528
rect -204 -1593 -47 -1592
<< via3 >>
rect -304 3026 -240 3090
rect -224 3026 -160 3090
rect 47 1795 111 1859
rect 127 1795 191 1859
rect 8971 3085 9035 3090
rect 9051 3085 9115 3090
rect 8971 3029 8981 3085
rect 8981 3029 9035 3085
rect 9051 3029 9061 3085
rect 9061 3029 9115 3085
rect 8971 3026 9035 3029
rect 9051 3026 9115 3029
rect 3154 2878 3210 2895
rect 3210 2878 3218 2895
rect 3154 2853 3218 2878
rect 3154 2831 3210 2853
rect 3210 2831 3218 2853
rect 3248 2878 3250 2895
rect 3250 2878 3306 2895
rect 3306 2878 3312 2895
rect 3248 2853 3312 2878
rect 3248 2831 3250 2853
rect 3250 2831 3306 2853
rect 3306 2831 3312 2853
rect 3342 2878 3346 2895
rect 3346 2878 3402 2895
rect 3402 2878 3406 2895
rect 3342 2853 3406 2878
rect 3342 2831 3346 2853
rect 3346 2831 3402 2853
rect 3402 2831 3406 2853
rect 3436 2878 3442 2895
rect 3442 2878 3498 2895
rect 3498 2878 3500 2895
rect 3436 2853 3500 2878
rect 3436 2831 3442 2853
rect 3442 2831 3498 2853
rect 3498 2831 3500 2853
rect 3530 2878 3538 2895
rect 3538 2878 3594 2895
rect 3530 2853 3594 2878
rect 3530 2831 3538 2853
rect 3538 2831 3594 2853
rect 3154 2797 3210 2809
rect 3210 2797 3218 2809
rect 3154 2772 3218 2797
rect 3154 2745 3210 2772
rect 3210 2745 3218 2772
rect 3248 2797 3250 2809
rect 3250 2797 3306 2809
rect 3306 2797 3312 2809
rect 3248 2772 3312 2797
rect 3248 2745 3250 2772
rect 3250 2745 3306 2772
rect 3306 2745 3312 2772
rect 3342 2797 3346 2809
rect 3346 2797 3402 2809
rect 3402 2797 3406 2809
rect 3342 2772 3406 2797
rect 3342 2745 3346 2772
rect 3346 2745 3402 2772
rect 3402 2745 3406 2772
rect 3436 2797 3442 2809
rect 3442 2797 3498 2809
rect 3498 2797 3500 2809
rect 3436 2772 3500 2797
rect 3436 2745 3442 2772
rect 3442 2745 3498 2772
rect 3498 2745 3500 2772
rect 3530 2797 3538 2809
rect 3538 2797 3594 2809
rect 3530 2772 3594 2797
rect 3530 2745 3538 2772
rect 3538 2745 3594 2772
rect 3154 2716 3210 2723
rect 3210 2716 3218 2723
rect 3154 2691 3218 2716
rect 3154 2659 3210 2691
rect 3210 2659 3218 2691
rect 3248 2716 3250 2723
rect 3250 2716 3306 2723
rect 3306 2716 3312 2723
rect 3248 2691 3312 2716
rect 3248 2659 3250 2691
rect 3250 2659 3306 2691
rect 3306 2659 3312 2691
rect 3342 2716 3346 2723
rect 3346 2716 3402 2723
rect 3402 2716 3406 2723
rect 3342 2691 3406 2716
rect 3342 2659 3346 2691
rect 3346 2659 3402 2691
rect 3402 2659 3406 2691
rect 3436 2716 3442 2723
rect 3442 2716 3498 2723
rect 3498 2716 3500 2723
rect 3436 2691 3500 2716
rect 3436 2659 3442 2691
rect 3442 2659 3498 2691
rect 3498 2659 3500 2691
rect 3530 2716 3538 2723
rect 3538 2716 3594 2723
rect 3530 2691 3594 2716
rect 3530 2659 3538 2691
rect 3538 2659 3594 2691
rect 3154 2635 3210 2637
rect 3210 2635 3218 2637
rect 3154 2610 3218 2635
rect 3154 2573 3210 2610
rect 3210 2573 3218 2610
rect 3248 2635 3250 2637
rect 3250 2635 3306 2637
rect 3306 2635 3312 2637
rect 3248 2610 3312 2635
rect 3248 2573 3250 2610
rect 3250 2573 3306 2610
rect 3306 2573 3312 2610
rect 3342 2635 3346 2637
rect 3346 2635 3402 2637
rect 3402 2635 3406 2637
rect 3342 2610 3406 2635
rect 3342 2573 3346 2610
rect 3346 2573 3402 2610
rect 3402 2573 3406 2610
rect 3436 2635 3442 2637
rect 3442 2635 3498 2637
rect 3498 2635 3500 2637
rect 3436 2610 3500 2635
rect 3436 2573 3442 2610
rect 3442 2573 3498 2610
rect 3498 2573 3500 2610
rect 3530 2635 3538 2637
rect 3538 2635 3594 2637
rect 3530 2610 3594 2635
rect 3530 2573 3538 2610
rect 3538 2573 3594 2610
rect 3154 2529 3218 2551
rect 3154 2487 3210 2529
rect 3210 2487 3218 2529
rect 3248 2529 3312 2551
rect 3248 2487 3250 2529
rect 3250 2487 3306 2529
rect 3306 2487 3312 2529
rect 3342 2529 3406 2551
rect 3342 2487 3346 2529
rect 3346 2487 3402 2529
rect 3402 2487 3406 2529
rect 3436 2529 3500 2551
rect 3436 2487 3442 2529
rect 3442 2487 3498 2529
rect 3498 2487 3500 2529
rect 3530 2529 3594 2551
rect 3530 2487 3538 2529
rect 3538 2487 3594 2529
rect 3154 2447 3218 2465
rect 3154 2401 3210 2447
rect 3210 2401 3218 2447
rect 3248 2447 3312 2465
rect 3248 2401 3250 2447
rect 3250 2401 3306 2447
rect 3306 2401 3312 2447
rect 3342 2447 3406 2465
rect 3342 2401 3346 2447
rect 3346 2401 3402 2447
rect 3402 2401 3406 2447
rect 3436 2447 3500 2465
rect 3436 2401 3442 2447
rect 3442 2401 3498 2447
rect 3498 2401 3500 2447
rect 3530 2447 3594 2465
rect 3530 2401 3538 2447
rect 3538 2401 3594 2447
rect 3154 2365 3218 2379
rect 3154 2315 3210 2365
rect 3210 2315 3218 2365
rect 3248 2365 3312 2379
rect 3248 2315 3250 2365
rect 3250 2315 3306 2365
rect 3306 2315 3312 2365
rect 3342 2365 3406 2379
rect 3342 2315 3346 2365
rect 3346 2315 3402 2365
rect 3402 2315 3406 2365
rect 3436 2365 3500 2379
rect 3436 2315 3442 2365
rect 3442 2315 3498 2365
rect 3498 2315 3500 2365
rect 3530 2365 3594 2379
rect 3530 2315 3538 2365
rect 3538 2315 3594 2365
rect 3154 2283 3218 2292
rect 3154 2228 3210 2283
rect 3210 2228 3218 2283
rect 3248 2283 3312 2292
rect 3248 2228 3250 2283
rect 3250 2228 3306 2283
rect 3306 2228 3312 2283
rect 3342 2283 3406 2292
rect 3342 2228 3346 2283
rect 3346 2228 3402 2283
rect 3402 2228 3406 2283
rect 3436 2283 3500 2292
rect 3436 2228 3442 2283
rect 3442 2228 3498 2283
rect 3498 2228 3500 2283
rect 3530 2283 3594 2292
rect 3530 2228 3538 2283
rect 3538 2228 3594 2283
rect 3154 2201 3218 2205
rect 3154 2145 3210 2201
rect 3210 2145 3218 2201
rect 3154 2141 3218 2145
rect 3248 2201 3312 2205
rect 3248 2145 3250 2201
rect 3250 2145 3306 2201
rect 3306 2145 3312 2201
rect 3248 2141 3312 2145
rect 3342 2201 3406 2205
rect 3342 2145 3346 2201
rect 3346 2145 3402 2201
rect 3402 2145 3406 2201
rect 3342 2141 3406 2145
rect 3436 2201 3500 2205
rect 3436 2145 3442 2201
rect 3442 2145 3498 2201
rect 3498 2145 3500 2201
rect 3436 2141 3500 2145
rect 3530 2201 3594 2205
rect 3530 2145 3538 2201
rect 3538 2145 3594 2201
rect 3530 2141 3594 2145
rect 3154 2063 3210 2118
rect 3210 2063 3218 2118
rect 3154 2054 3218 2063
rect 3248 2063 3250 2118
rect 3250 2063 3306 2118
rect 3306 2063 3312 2118
rect 3248 2054 3312 2063
rect 3342 2063 3346 2118
rect 3346 2063 3402 2118
rect 3402 2063 3406 2118
rect 3342 2054 3406 2063
rect 3436 2063 3442 2118
rect 3442 2063 3498 2118
rect 3498 2063 3500 2118
rect 3436 2054 3500 2063
rect 3530 2063 3538 2118
rect 3538 2063 3594 2118
rect 3530 2054 3594 2063
rect 3154 1981 3210 2031
rect 3210 1981 3218 2031
rect 3154 1967 3218 1981
rect 3248 1981 3250 2031
rect 3250 1981 3306 2031
rect 3306 1981 3312 2031
rect 3248 1967 3312 1981
rect 3342 1981 3346 2031
rect 3346 1981 3402 2031
rect 3402 1981 3406 2031
rect 3342 1967 3406 1981
rect 3436 1981 3442 2031
rect 3442 1981 3498 2031
rect 3498 1981 3500 2031
rect 3436 1967 3500 1981
rect 3530 1981 3538 2031
rect 3538 1981 3594 2031
rect 3530 1967 3594 1981
rect 10416 1850 10480 1859
rect 10496 1850 10560 1859
rect 10416 1795 10425 1850
rect 10425 1795 10480 1850
rect 10496 1795 10505 1850
rect 10505 1795 10560 1850
rect -407 631 -374 650
rect -374 631 -343 650
rect -327 631 -318 650
rect -318 631 -263 650
rect -407 607 -343 631
rect -327 607 -263 631
rect -407 586 -374 607
rect -374 586 -343 607
rect -327 586 -318 607
rect -318 586 -263 607
rect 12255 647 12319 650
rect 12335 647 12399 650
rect 12255 591 12264 647
rect 12264 591 12319 647
rect 12335 591 12344 647
rect 12344 591 12399 647
rect 12255 586 12319 591
rect 12335 586 12399 591
rect -442 -373 -378 -309
rect -362 -373 -298 -309
rect 11357 -315 11421 -309
rect 11357 -371 11413 -315
rect 11413 -371 11421 -315
rect 11357 -373 11421 -371
rect 11437 -315 11501 -309
rect 11437 -371 11493 -315
rect 11493 -371 11501 -315
rect 11437 -373 11501 -371
rect -198 -1532 -134 -1528
rect -198 -1588 -191 -1532
rect -191 -1588 -135 -1532
rect -135 -1588 -134 -1532
rect -198 -1592 -134 -1588
rect -118 -1532 -54 -1528
rect -118 -1588 -111 -1532
rect -111 -1588 -55 -1532
rect -55 -1588 -54 -1532
rect -118 -1592 -54 -1588
rect 12245 -1592 12309 -1528
rect 12325 -1592 12389 -1528
<< metal4 >>
rect -357 3090 9116 3091
rect -357 3026 -304 3090
rect -240 3026 -224 3090
rect -160 3026 8971 3090
rect 9035 3026 9051 3090
rect 9115 3026 9116 3090
rect -357 3025 9116 3026
rect 3150 2895 3598 2896
rect 3150 2831 3154 2895
rect 3218 2831 3248 2895
rect 3312 2831 3342 2895
rect 3406 2831 3436 2895
rect 3500 2831 3530 2895
rect 3594 2831 3598 2895
rect 3150 2809 3598 2831
rect 3150 2745 3154 2809
rect 3218 2745 3248 2809
rect 3312 2745 3342 2809
rect 3406 2745 3436 2809
rect 3500 2745 3530 2809
rect 3594 2745 3598 2809
rect 3150 2723 3598 2745
rect 3150 2659 3154 2723
rect 3218 2659 3248 2723
rect 3312 2659 3342 2723
rect 3406 2659 3436 2723
rect 3500 2659 3530 2723
rect 3594 2659 3598 2723
rect 3150 2637 3598 2659
rect 3150 2573 3154 2637
rect 3218 2573 3248 2637
rect 3312 2573 3342 2637
rect 3406 2573 3436 2637
rect 3500 2573 3530 2637
rect 3594 2573 3598 2637
rect 3150 2551 3598 2573
rect 3150 2487 3154 2551
rect 3218 2487 3248 2551
rect 3312 2487 3342 2551
rect 3406 2487 3436 2551
rect 3500 2487 3530 2551
rect 3594 2487 3598 2551
rect 3150 2465 3598 2487
rect 3150 2401 3154 2465
rect 3218 2401 3248 2465
rect 3312 2401 3342 2465
rect 3406 2401 3436 2465
rect 3500 2401 3530 2465
rect 3594 2401 3598 2465
rect 3150 2379 3598 2401
rect 3150 2315 3154 2379
rect 3218 2315 3248 2379
rect 3312 2315 3342 2379
rect 3406 2315 3436 2379
rect 3500 2315 3530 2379
rect 3594 2315 3598 2379
rect 3150 2292 3598 2315
rect 3150 2228 3154 2292
rect 3218 2228 3248 2292
rect 3312 2228 3342 2292
rect 3406 2228 3436 2292
rect 3500 2228 3530 2292
rect 3594 2228 3598 2292
rect 3150 2205 3598 2228
rect 3150 2141 3154 2205
rect 3218 2141 3248 2205
rect 3312 2141 3342 2205
rect 3406 2141 3436 2205
rect 3500 2141 3530 2205
rect 3594 2141 3598 2205
rect 3150 2118 3598 2141
rect 3150 2054 3154 2118
rect 3218 2054 3248 2118
rect 3312 2054 3342 2118
rect 3406 2054 3436 2118
rect 3500 2054 3530 2118
rect 3594 2054 3598 2118
rect 3150 2031 3598 2054
rect 3150 1967 3154 2031
rect 3218 1967 3248 2031
rect 3312 1967 3342 2031
rect 3406 1967 3436 2031
rect 3500 1967 3530 2031
rect 3594 1967 3598 2031
rect 3150 1966 3598 1967
rect 46 1859 10561 1860
rect 46 1795 47 1859
rect 111 1795 127 1859
rect 191 1795 10416 1859
rect 10480 1795 10496 1859
rect 10560 1795 10561 1859
rect 46 1794 10561 1795
rect -408 650 12400 651
rect -408 586 -407 650
rect -343 586 -327 650
rect -263 586 12255 650
rect 12319 586 12335 650
rect 12399 586 12400 650
rect -408 585 12400 586
rect -443 -309 11502 -308
rect -443 -373 -442 -309
rect -378 -373 -362 -309
rect -298 -373 11357 -309
rect 11421 -373 11437 -309
rect 11501 -373 11502 -309
rect -443 -374 11502 -373
rect -199 -1528 12394 -1527
rect -199 -1592 -198 -1528
rect -134 -1592 -118 -1528
rect -54 -1592 12245 -1528
rect 12309 -1592 12325 -1528
rect 12389 -1592 12394 -1528
rect -199 -1593 12394 -1592
use sky130_fd_io__com_opath_datoev2  sky130_fd_io__com_opath_datoev2_0
timestamp 1694700623
transform 1 0 467 0 -1 6943
box -349 -1098 12658 2562
use sky130_fd_io__gpiov2_obpredrvr  sky130_fd_io__gpiov2_obpredrvr_0
timestamp 1694700623
transform 1 0 288 0 -1 5207
box -714 451 12112 4765
use sky130_fd_io__gpiov2_octl  sky130_fd_io__gpiov2_octl_0
timestamp 1694700623
transform 1 0 8821 0 -1 7867
box -9346 1177 6467 7642
<< labels >>
flabel metal1 s 14854 6410 14989 6527 3 FreeSans 520 180 0 0 VPWR
port 2 nsew
flabel metal1 s 12123 2928 12165 3058 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 9029 3979 9071 4181 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 470 3979 512 4181 3 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 1264 2928 1306 3058 3 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 1264 2312 1306 2442 3 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 12634 1302 12676 1504 7 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 12639 644 12676 790 7 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 12634 3453 12676 3655 7 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 1264 3453 1306 3655 3 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 288 644 325 790 3 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 288 1302 330 1504 3 FreeSans 300 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 12158 1828 12200 2030 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 12258 2312 12300 2442 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 12140 2928 12182 3058 7 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 491 4080 491 4080 3 FreeSans 300 0 0 0 VGND_IO
flabel metal1 s 1285 2993 1285 2993 3 FreeSans 300 0 0 0 VGND_IO
flabel metal1 s 1285 2377 1285 2377 3 FreeSans 300 0 0 0 VGND_IO
flabel metal1 s 951 1828 993 2030 3 FreeSans 300 0 0 0 VGND_IO
port 3 nsew
flabel metal1 s 12655 1403 12655 1403 7 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 12657 717 12657 717 7 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 12655 3554 12655 3554 7 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 1285 3554 1285 3554 3 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 306 717 306 717 3 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 309 1403 309 1403 3 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 5854 6502 5921 6850 3 FreeSans 520 0 0 0 VPWR_KA
port 5 nsew
flabel metal1 s 524 4938 564 5068 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 288 5857 328 6059 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 288 4708 328 4910 3 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 12991 4708 13031 4910 3 FreeSans 300 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 5900 6502 5967 6850 3 FreeSans 520 0 0 0 VPWR_KA
port 5 nsew
flabel metal1 s 544 5003 544 5003 3 FreeSans 300 180 0 0 VGND
flabel metal1 s 12900 4938 12940 5068 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 308 5958 308 5958 3 FreeSans 300 180 0 0 VGND
flabel metal1 s 13102 5787 13142 5989 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 308 4809 308 4809 3 FreeSans 300 180 0 0 VCC_IO
flabel metal1 s 13011 4809 13011 4809 3 FreeSans 300 180 0 0 VCC_IO
flabel metal1 s 13170 5809 13337 5965 3 FreeSans 520 180 0 0 VGND
port 6 nsew
flabel metal1 s 14840 4258 15007 4414 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 14840 2226 15007 2382 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 14840 260 15007 416 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 13251 4812 13562 4987 3 FreeSans 520 180 0 0 VCC_IO
port 4 nsew
flabel metal1 s 14697 3248 15008 3480 3 FreeSans 520 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 14697 1137 15008 1369 3 FreeSans 520 0 0 0 VCC_IO
port 4 nsew
flabel metal1 s 14923 4336 14923 4336 3 FreeSans 520 0 0 0 VGND
flabel metal1 s 14923 2304 14923 2304 3 FreeSans 520 0 0 0 VGND
flabel metal1 s 14923 338 14923 338 3 FreeSans 520 0 0 0 VGND
flabel metal1 s 13406 4899 13406 4899 3 FreeSans 520 180 0 0 VCC_IO
flabel metal1 s 14852 3364 14852 3364 3 FreeSans 520 0 0 0 VCC_IO
flabel metal1 s 14852 1253 14852 1253 3 FreeSans 520 0 0 0 VCC_IO
flabel metal1 s 15042 5345 15116 5380 3 FreeSans 520 180 0 0 SLOW
port 7 nsew
flabel metal1 s 14478 5304 14522 5348 3 FreeSans 520 180 0 0 HLD_I_H_N
port 8 nsew
flabel metal1 s 15079 5362 15079 5362 3 FreeSans 520 180 0 0 SLOW
flabel metal1 s 14501 5326 14501 5326 3 FreeSans 520 180 0 0 HLD_I_H_N
flabel metal1 s 5095 6957 5128 6995 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 9 nsew
flabel metal1 s 5111 6976 5111 6976 3 FreeSans 520 0 0 0 HLD_I_OVR_H
flabel metal1 s 15079 5362 15079 5362 3 FreeSans 520 180 0 0 SLOW
flabel metal1 s 14824 6126 14868 6164 3 FreeSans 520 180 0 0 OD_H
port 10 nsew
flabel metal1 s 14501 5326 14501 5326 3 FreeSans 520 180 0 0 HLD_I_H_N
flabel metal1 s 13425 5630 13492 5674 3 FreeSans 520 180 0 0 SLOW_H_N
port 11 nsew
flabel metal1 s 8283 5096 8333 5148 3 FreeSans 300 180 0 0 DRVHI_H
port 12 nsew
flabel metal1 s 8308 5122 8308 5122 3 FreeSans 300 180 0 0 DRVHI_H
flabel metal1 s 6190 1228 6231 1274 3 FreeSans 300 0 0 0 PU_H_N[3]
port 13 nsew
flabel metal1 s 6054 1228 6094 1274 7 FreeSans 300 0 0 0 PU_H_N[2]
port 14 nsew
flabel metal1 s 10362 1072 10402 1118 3 FreeSans 300 0 0 0 PU_H_N[1]
port 15 nsew
flabel metal1 s 7956 1148 7996 1194 3 FreeSans 300 0 0 0 PU_H_N[0]
port 16 nsew
flabel metal1 s 9390 1030 9436 1076 3 FreeSans 300 0 0 0 PD_H[1]
port 17 nsew
flabel metal1 s 8148 1030 8194 1076 3 FreeSans 300 0 0 0 PD_H[0]
port 18 nsew
flabel metal1 s 11863 2475 11928 2502 3 FreeSans 520 0 0 0 PD_H[4]
port 19 nsew
flabel metal1 s 8242 4238 8242 4238 0 FreeSans 440 0 0 0 DRVLO_H_N
flabel metal2 s 13617 397 13652 442 3 FreeSans 520 90 0 0 DM_H_N[2]
port 21 nsew
flabel metal2 s 14263 399 14307 448 3 FreeSans 520 90 0 0 DM_H_N[0]
port 22 nsew
flabel metal2 s 12786 514 12812 563 3 FreeSans 520 90 0 0 DM_H[2]
port 23 nsew
flabel metal2 s 13425 445 13474 498 3 FreeSans 520 90 0 0 DM_H[1]
port 24 nsew
flabel metal2 s 13257 437 13306 500 3 FreeSans 520 90 0 0 DM_H[0]
port 25 nsew
flabel metal2 s 13634 419 13634 419 3 FreeSans 520 90 0 0 DM_H_N[2]
flabel metal2 s 14285 423 14285 423 3 FreeSans 520 90 0 0 DM_H_N[0]
flabel metal2 s 13449 471 13449 471 3 FreeSans 520 90 0 0 DM_H[1]
flabel metal2 s 3827 6885 3879 6924 3 FreeSans 520 0 0 0 OUT
port 26 nsew
flabel metal2 s 3354 6878 3400 6924 7 FreeSans 300 0 0 0 OE_N
port 27 nsew
flabel metal2 s 3848 6898 3848 6898 3 FreeSans 520 0 0 0 OUT
flabel metal2 s 3377 6901 3377 6901 7 FreeSans 300 0 0 0 OE_N
flabel metal2 s -367 5535 -318 5598 3 FreeSans 520 90 0 0 DM_H[0]
port 25 nsew
flabel metal2 s 13634 419 13634 419 3 FreeSans 520 90 0 0 DM_H_N[2]
flabel metal2 s 13789 394 13823 443 3 FreeSans 520 90 0 0 DM_H_N[1]
port 28 nsew
flabel metal2 s 14285 423 14285 423 3 FreeSans 520 90 0 0 DM_H_N[0]
flabel metal2 s 13449 471 13449 471 3 FreeSans 520 90 0 0 DM_H[1]
flabel metal2 s 11401 2065 11449 2117 3 FreeSans 300 0 0 0 PD_H[3]
port 29 nsew
flabel metal2 s 1 5402 27 5451 3 FreeSans 520 90 0 0 DM_H[2]
port 23 nsew
flabel metal2 s -193 5390 -144 5443 3 FreeSans 520 90 0 0 DM_H[1]
port 24 nsew
flabel metal2 s 10919 2470 10967 2522 3 FreeSans 300 0 0 0 PD_H[2]
port 30 nsew
<< properties >>
string GDS_END 7685534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7611198
<< end >>
