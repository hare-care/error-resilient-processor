magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< obsli1 >>
rect 199 1140 207 1174
rect 241 1140 279 1174
rect 313 1140 351 1174
rect 385 1140 423 1174
rect 457 1140 495 1174
rect 529 1140 567 1174
rect 601 1140 639 1174
rect 673 1140 711 1174
rect 745 1140 783 1174
rect 817 1140 855 1174
rect 889 1140 927 1174
rect 961 1140 999 1174
rect 1033 1140 1071 1174
rect 1105 1140 1143 1174
rect 1177 1140 1215 1174
rect 1249 1140 1287 1174
rect 1321 1140 1359 1174
rect 1393 1140 1431 1174
rect 1465 1140 1503 1174
rect 1537 1140 1575 1174
rect 1609 1140 1647 1174
rect 1681 1140 1719 1174
rect 1753 1140 1761 1174
rect 48 1010 82 1048
rect 48 938 82 976
rect 48 866 82 904
rect 48 794 82 832
rect 48 722 82 760
rect 48 650 82 688
rect 48 578 82 616
rect 48 506 82 544
rect 48 434 82 472
rect 48 362 82 400
rect 48 290 82 328
rect 48 218 82 256
rect 48 112 82 184
rect 183 88 217 1106
rect 339 88 373 1106
rect 495 88 529 1106
rect 651 88 685 1106
rect 807 88 841 1106
rect 963 88 997 1106
rect 1119 88 1153 1106
rect 1275 88 1309 1106
rect 1431 88 1465 1106
rect 1587 88 1621 1106
rect 1743 88 1777 1106
rect 1878 1010 1912 1048
rect 1878 938 1912 976
rect 1878 866 1912 904
rect 1878 794 1912 832
rect 1878 722 1912 760
rect 1878 650 1912 688
rect 1878 578 1912 616
rect 1878 506 1912 544
rect 1878 434 1912 472
rect 1878 362 1912 400
rect 1878 290 1912 328
rect 1878 218 1912 256
rect 1878 112 1912 184
rect 199 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1761 54
<< obsli1c >>
rect 207 1140 241 1174
rect 279 1140 313 1174
rect 351 1140 385 1174
rect 423 1140 457 1174
rect 495 1140 529 1174
rect 567 1140 601 1174
rect 639 1140 673 1174
rect 711 1140 745 1174
rect 783 1140 817 1174
rect 855 1140 889 1174
rect 927 1140 961 1174
rect 999 1140 1033 1174
rect 1071 1140 1105 1174
rect 1143 1140 1177 1174
rect 1215 1140 1249 1174
rect 1287 1140 1321 1174
rect 1359 1140 1393 1174
rect 1431 1140 1465 1174
rect 1503 1140 1537 1174
rect 1575 1140 1609 1174
rect 1647 1140 1681 1174
rect 1719 1140 1753 1174
rect 48 1048 82 1082
rect 48 976 82 1010
rect 48 904 82 938
rect 48 832 82 866
rect 48 760 82 794
rect 48 688 82 722
rect 48 616 82 650
rect 48 544 82 578
rect 48 472 82 506
rect 48 400 82 434
rect 48 328 82 362
rect 48 256 82 290
rect 48 184 82 218
rect 1878 1048 1912 1082
rect 1878 976 1912 1010
rect 1878 904 1912 938
rect 1878 832 1912 866
rect 1878 760 1912 794
rect 1878 688 1912 722
rect 1878 616 1912 650
rect 1878 544 1912 578
rect 1878 472 1912 506
rect 1878 400 1912 434
rect 1878 328 1912 362
rect 1878 256 1912 290
rect 1878 184 1912 218
rect 207 20 241 54
rect 279 20 313 54
rect 351 20 385 54
rect 423 20 457 54
rect 495 20 529 54
rect 567 20 601 54
rect 639 20 673 54
rect 711 20 745 54
rect 783 20 817 54
rect 855 20 889 54
rect 927 20 961 54
rect 999 20 1033 54
rect 1071 20 1105 54
rect 1143 20 1177 54
rect 1215 20 1249 54
rect 1287 20 1321 54
rect 1359 20 1393 54
rect 1431 20 1465 54
rect 1503 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1681 54
rect 1719 20 1753 54
<< metal1 >>
rect 195 1174 1765 1194
rect 195 1140 207 1174
rect 241 1140 279 1174
rect 313 1140 351 1174
rect 385 1140 423 1174
rect 457 1140 495 1174
rect 529 1140 567 1174
rect 601 1140 639 1174
rect 673 1140 711 1174
rect 745 1140 783 1174
rect 817 1140 855 1174
rect 889 1140 927 1174
rect 961 1140 999 1174
rect 1033 1140 1071 1174
rect 1105 1140 1143 1174
rect 1177 1140 1215 1174
rect 1249 1140 1287 1174
rect 1321 1140 1359 1174
rect 1393 1140 1431 1174
rect 1465 1140 1503 1174
rect 1537 1140 1575 1174
rect 1609 1140 1647 1174
rect 1681 1140 1719 1174
rect 1753 1140 1765 1174
rect 195 1128 1765 1140
rect 36 1082 95 1094
rect 36 1048 48 1082
rect 82 1048 95 1082
rect 36 1010 95 1048
rect 36 976 48 1010
rect 82 976 95 1010
rect 36 938 95 976
rect 36 904 48 938
rect 82 904 95 938
rect 36 866 95 904
rect 36 832 48 866
rect 82 832 95 866
rect 36 794 95 832
rect 36 760 48 794
rect 82 760 95 794
rect 36 722 95 760
rect 36 688 48 722
rect 82 688 95 722
rect 36 650 95 688
rect 36 616 48 650
rect 82 616 95 650
rect 36 578 95 616
rect 36 544 48 578
rect 82 544 95 578
rect 36 506 95 544
rect 36 472 48 506
rect 82 472 95 506
rect 36 434 95 472
rect 36 400 48 434
rect 82 400 95 434
rect 36 362 95 400
rect 36 328 48 362
rect 82 328 95 362
rect 36 290 95 328
rect 36 256 48 290
rect 82 256 95 290
rect 36 218 95 256
rect 36 184 48 218
rect 82 184 95 218
rect 36 100 95 184
rect 1866 1082 1925 1094
rect 1866 1048 1878 1082
rect 1912 1048 1925 1082
rect 1866 1010 1925 1048
rect 1866 976 1878 1010
rect 1912 976 1925 1010
rect 1866 938 1925 976
rect 1866 904 1878 938
rect 1912 904 1925 938
rect 1866 866 1925 904
rect 1866 832 1878 866
rect 1912 832 1925 866
rect 1866 794 1925 832
rect 1866 760 1878 794
rect 1912 760 1925 794
rect 1866 722 1925 760
rect 1866 688 1878 722
rect 1912 688 1925 722
rect 1866 650 1925 688
rect 1866 616 1878 650
rect 1912 616 1925 650
rect 1866 578 1925 616
rect 1866 544 1878 578
rect 1912 544 1925 578
rect 1866 506 1925 544
rect 1866 472 1878 506
rect 1912 472 1925 506
rect 1866 434 1925 472
rect 1866 400 1878 434
rect 1912 400 1925 434
rect 1866 362 1925 400
rect 1866 328 1878 362
rect 1912 328 1925 362
rect 1866 290 1925 328
rect 1866 256 1878 290
rect 1912 256 1925 290
rect 1866 218 1925 256
rect 1866 184 1878 218
rect 1912 184 1925 218
rect 1866 100 1925 184
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< obsm1 >>
rect 174 100 226 1094
rect 330 100 382 1094
rect 486 100 538 1094
rect 642 100 694 1094
rect 798 100 850 1094
rect 954 100 1006 1094
rect 1110 100 1162 1094
rect 1266 100 1318 1094
rect 1422 100 1474 1094
rect 1578 100 1630 1094
rect 1734 100 1786 1094
<< metal2 >>
rect 14 622 1946 1094
rect 14 100 1946 572
<< labels >>
rlabel metal2 s 14 622 1946 1094 6 DRAIN
port 1 nsew
rlabel metal1 s 195 1128 1765 1194 6 GATE
port 2 nsew
rlabel metal1 s 195 0 1765 66 6 GATE
port 2 nsew
rlabel metal2 s 14 100 1946 572 6 SOURCE
port 3 nsew
rlabel metal1 s 36 100 95 1094 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1866 100 1925 1094 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1946 1194
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7173406
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7130710
<< end >>
