VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO dcache_data_ram
   CLASS BLOCK ;
   SIZE 372.1 BY 288.02 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  100.54 0.0 100.92 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.38 0.0 106.76 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.22 0.0 112.6 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.06 0.0 118.44 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.9 0.0 124.28 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.74 0.0 130.12 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  135.58 0.0 135.96 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.42 0.0 141.8 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.26 0.0 147.64 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.1 0.0 153.48 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  158.94 0.0 159.32 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  164.78 0.0 165.16 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.62 0.0 171.0 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.46 0.0 176.84 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.3 0.0 182.68 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.14 0.0 188.52 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.98 0.0 194.36 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.82 0.0 200.2 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  205.66 0.0 206.04 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  211.5 0.0 211.88 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.34 0.0 217.72 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.18 0.0 223.56 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.02 0.0 229.4 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  234.86 0.0 235.24 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  240.7 0.0 241.08 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.54 0.0 246.92 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  252.38 0.0 252.76 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  258.22 0.0 258.6 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.06 0.0 264.44 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.9 0.0 270.28 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  275.74 0.0 276.12 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  281.58 0.0 281.96 0.38 ;
      END
   END din0[31]
   PIN din1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.16 287.64 80.54 288.02 ;
      END
   END din1[0]
   PIN din1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.0 287.64 86.38 288.02 ;
      END
   END din1[1]
   PIN din1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.84 287.64 92.22 288.02 ;
      END
   END din1[2]
   PIN din1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.68 287.64 98.06 288.02 ;
      END
   END din1[3]
   PIN din1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.52 287.64 103.9 288.02 ;
      END
   END din1[4]
   PIN din1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  109.36 287.64 109.74 288.02 ;
      END
   END din1[5]
   PIN din1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.2 287.64 115.58 288.02 ;
      END
   END din1[6]
   PIN din1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.04 287.64 121.42 288.02 ;
      END
   END din1[7]
   PIN din1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  126.88 287.64 127.26 288.02 ;
      END
   END din1[8]
   PIN din1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.72 287.64 133.1 288.02 ;
      END
   END din1[9]
   PIN din1[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.56 287.64 138.94 288.02 ;
      END
   END din1[10]
   PIN din1[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.4 287.64 144.78 288.02 ;
      END
   END din1[11]
   PIN din1[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.24 287.64 150.62 288.02 ;
      END
   END din1[12]
   PIN din1[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.08 287.64 156.46 288.02 ;
      END
   END din1[13]
   PIN din1[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.92 287.64 162.3 288.02 ;
      END
   END din1[14]
   PIN din1[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.76 287.64 168.14 288.02 ;
      END
   END din1[15]
   PIN din1[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.6 287.64 173.98 288.02 ;
      END
   END din1[16]
   PIN din1[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.44 287.64 179.82 288.02 ;
      END
   END din1[17]
   PIN din1[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.28 287.64 185.66 288.02 ;
      END
   END din1[18]
   PIN din1[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.12 287.64 191.5 288.02 ;
      END
   END din1[19]
   PIN din1[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.96 287.64 197.34 288.02 ;
      END
   END din1[20]
   PIN din1[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.8 287.64 203.18 288.02 ;
      END
   END din1[21]
   PIN din1[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.64 287.64 209.02 288.02 ;
      END
   END din1[22]
   PIN din1[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.48 287.64 214.86 288.02 ;
      END
   END din1[23]
   PIN din1[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.32 287.64 220.7 288.02 ;
      END
   END din1[24]
   PIN din1[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.16 287.64 226.54 288.02 ;
      END
   END din1[25]
   PIN din1[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.0 287.64 232.38 288.02 ;
      END
   END din1[26]
   PIN din1[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.84 287.64 238.22 288.02 ;
      END
   END din1[27]
   PIN din1[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.68 287.64 244.06 288.02 ;
      END
   END din1[28]
   PIN din1[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  249.52 287.64 249.9 288.02 ;
      END
   END din1[29]
   PIN din1[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.36 287.64 255.74 288.02 ;
      END
   END din1[30]
   PIN din1[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.2 287.64 261.58 288.02 ;
      END
   END din1[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 109.585 0.38 109.965 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 117.985 0.38 118.365 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 123.85 0.38 124.23 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 132.35 0.38 132.73 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 137.99 0.38 138.37 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 146.49 0.38 146.87 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  371.72 72.47 372.1 72.85 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  304.095 0.0 304.475 0.38 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  307.76 0.0 308.14 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  304.785 0.0 305.165 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  305.475 0.0 305.855 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.22 0.0 306.6 0.38 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 16.73 0.38 17.11 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  371.72 260.0 372.1 260.38 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 25.23 0.38 25.61 ;
      END
   END web0
   PIN web1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  371.72 251.5 372.1 251.88 ;
      END
   END web1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  340.62 287.64 341.0 288.02 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  77.18 0.0 77.56 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.02 0.0 83.4 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.86 0.0 89.24 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  94.7 0.0 95.08 0.38 ;
      END
   END wmask0[3]
   PIN wmask1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.04 287.64 267.42 288.02 ;
      END
   END wmask1[0]
   PIN wmask1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.88 287.64 273.26 288.02 ;
      END
   END wmask1[1]
   PIN wmask1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.72 287.64 279.1 288.02 ;
      END
   END wmask1[2]
   PIN wmask1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.56 287.64 284.94 288.02 ;
      END
   END wmask1[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.685 0.0 138.065 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.11 0.0 142.49 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.925 0.0 144.305 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.95 0.0 148.33 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.785 0.0 149.165 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.815 0.0 154.195 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.025 0.0 155.405 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.0 0.0 160.38 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.645 0.0 163.025 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.295 0.0 166.675 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.505 0.0 167.885 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.535 0.0 172.915 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.745 0.0 174.125 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.775 0.0 179.155 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.985 0.0 180.365 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.285 0.0 186.665 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.255 0.0 191.635 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.175 0.0 192.555 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.495 0.0 197.875 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  200.51 0.0 200.89 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.735 0.0 204.115 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.35 0.0 206.73 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.695 0.0 210.075 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.565 0.0 212.945 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.535 0.0 215.915 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.03 0.0 218.41 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.515 0.0 220.895 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.87 0.0 224.25 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.71 0.0 230.09 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.285 0.0 231.665 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.68 0.0 236.06 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.56 287.64 136.94 288.02 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.335 287.64 141.715 288.02 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.545 287.64 142.925 288.02 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.575 287.64 147.955 288.02 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.435 287.64 148.815 288.02 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.815 287.64 154.195 288.02 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  156.77 287.64 157.15 288.02 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.0 287.64 160.38 288.02 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.645 287.64 163.025 288.02 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.955 287.64 166.335 288.02 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.885 287.64 169.265 288.02 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  171.795 287.64 172.175 288.02 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.29 287.64 174.67 288.02 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.835 287.64 177.215 288.02 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.13 287.64 180.51 288.02 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.075 287.64 183.455 288.02 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.605 287.64 187.985 288.02 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.81 287.64 192.19 288.02 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.525 287.64 192.905 288.02 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.65 287.64 198.03 288.02 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.705 287.64 199.085 288.02 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.735 287.64 204.115 288.02 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.945 287.64 205.325 288.02 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.92 287.64 210.3 288.02 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.565 287.64 212.945 288.02 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.215 287.64 216.595 288.02 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.425 287.64 217.805 288.02 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.455 287.64 222.835 288.02 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.665 287.64 224.045 288.02 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.695 287.64 229.075 288.02 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.905 287.64 230.285 288.02 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.935 287.64 235.315 288.02 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 286.28 372.1 288.02 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 288.02 ;
         LAYER met4 ;
         RECT  370.36 0.0 372.1 288.02 ;
         LAYER met3 ;
         RECT  0.0 0.0 372.1 1.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 3.48 368.62 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 284.54 ;
         LAYER met3 ;
         RECT  3.48 282.8 368.62 284.54 ;
         LAYER met4 ;
         RECT  366.88 3.48 368.62 284.54 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 371.48 287.4 ;
   LAYER  met2 ;
      RECT  0.62 0.62 371.48 287.4 ;
   LAYER  met3 ;
      RECT  0.98 108.985 371.48 110.565 ;
      RECT  0.62 110.565 0.98 117.385 ;
      RECT  0.62 118.965 0.98 123.25 ;
      RECT  0.62 124.83 0.98 131.75 ;
      RECT  0.62 133.33 0.98 137.39 ;
      RECT  0.62 138.97 0.98 145.89 ;
      RECT  0.98 71.87 371.12 73.45 ;
      RECT  0.98 73.45 371.12 108.985 ;
      RECT  371.12 73.45 371.48 108.985 ;
      RECT  0.98 110.565 371.12 259.4 ;
      RECT  0.98 259.4 371.12 260.98 ;
      RECT  0.62 17.71 0.98 24.63 ;
      RECT  0.62 26.21 0.98 108.985 ;
      RECT  371.12 110.565 371.48 250.9 ;
      RECT  371.12 252.48 371.48 259.4 ;
      RECT  0.62 147.47 0.98 285.68 ;
      RECT  371.12 260.98 371.48 285.68 ;
      RECT  371.12 2.34 371.48 71.87 ;
      RECT  0.62 2.34 0.98 16.13 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 71.87 ;
      RECT  2.88 2.34 369.22 2.88 ;
      RECT  2.88 5.82 369.22 71.87 ;
      RECT  369.22 2.34 371.12 2.88 ;
      RECT  369.22 2.88 371.12 5.82 ;
      RECT  369.22 5.82 371.12 71.87 ;
      RECT  0.98 260.98 2.88 282.2 ;
      RECT  0.98 282.2 2.88 285.14 ;
      RECT  0.98 285.14 2.88 285.68 ;
      RECT  2.88 260.98 369.22 282.2 ;
      RECT  2.88 285.14 369.22 285.68 ;
      RECT  369.22 260.98 371.12 282.2 ;
      RECT  369.22 282.2 371.12 285.14 ;
      RECT  369.22 285.14 371.12 285.68 ;
   LAYER  met4 ;
      RECT  99.94 0.98 101.52 287.4 ;
      RECT  101.52 0.62 105.78 0.98 ;
      RECT  107.36 0.62 111.62 0.98 ;
      RECT  113.2 0.62 117.46 0.98 ;
      RECT  119.04 0.62 123.3 0.98 ;
      RECT  124.88 0.62 129.14 0.98 ;
      RECT  130.72 0.62 134.98 0.98 ;
      RECT  241.68 0.62 245.94 0.98 ;
      RECT  247.52 0.62 251.78 0.98 ;
      RECT  253.36 0.62 257.62 0.98 ;
      RECT  259.2 0.62 263.46 0.98 ;
      RECT  265.04 0.62 269.3 0.98 ;
      RECT  270.88 0.62 275.14 0.98 ;
      RECT  276.72 0.62 280.98 0.98 ;
      RECT  79.56 0.98 81.14 287.04 ;
      RECT  81.14 0.98 99.94 287.04 ;
      RECT  81.14 287.04 85.4 287.4 ;
      RECT  86.98 287.04 91.24 287.4 ;
      RECT  92.82 287.04 97.08 287.4 ;
      RECT  98.66 287.04 99.94 287.4 ;
      RECT  101.52 0.98 102.92 287.04 ;
      RECT  101.52 287.04 102.92 287.4 ;
      RECT  102.92 0.98 104.5 287.04 ;
      RECT  104.5 287.04 108.76 287.4 ;
      RECT  110.34 287.04 114.6 287.4 ;
      RECT  116.18 287.04 120.44 287.4 ;
      RECT  122.02 287.04 126.28 287.4 ;
      RECT  127.86 287.04 132.12 287.4 ;
      RECT  238.82 287.04 243.08 287.4 ;
      RECT  244.66 287.04 248.92 287.4 ;
      RECT  250.5 287.04 254.76 287.4 ;
      RECT  256.34 287.04 260.6 287.4 ;
      RECT  282.56 0.62 303.495 0.98 ;
      RECT  32.08 0.62 76.58 0.98 ;
      RECT  78.16 0.62 82.42 0.98 ;
      RECT  84.0 0.62 88.26 0.98 ;
      RECT  89.84 0.62 94.1 0.98 ;
      RECT  95.68 0.62 99.94 0.98 ;
      RECT  262.18 287.04 266.44 287.4 ;
      RECT  268.02 287.04 272.28 287.4 ;
      RECT  273.86 287.04 278.12 287.4 ;
      RECT  279.7 287.04 283.96 287.4 ;
      RECT  285.54 287.04 340.02 287.4 ;
      RECT  136.56 0.62 137.085 0.98 ;
      RECT  138.665 0.62 140.82 0.98 ;
      RECT  143.09 0.62 143.325 0.98 ;
      RECT  144.905 0.62 146.66 0.98 ;
      RECT  149.765 0.62 152.5 0.98 ;
      RECT  156.005 0.62 158.34 0.98 ;
      RECT  160.98 0.62 162.045 0.98 ;
      RECT  163.625 0.62 164.18 0.98 ;
      RECT  168.485 0.62 170.02 0.98 ;
      RECT  171.6 0.62 171.935 0.98 ;
      RECT  174.725 0.62 175.86 0.98 ;
      RECT  177.44 0.62 178.175 0.98 ;
      RECT  180.965 0.62 181.7 0.98 ;
      RECT  183.28 0.62 184.36 0.98 ;
      RECT  187.265 0.62 187.54 0.98 ;
      RECT  189.12 0.62 190.655 0.98 ;
      RECT  193.155 0.62 193.38 0.98 ;
      RECT  194.96 0.62 196.895 0.98 ;
      RECT  198.475 0.62 199.22 0.98 ;
      RECT  201.49 0.62 203.135 0.98 ;
      RECT  204.715 0.62 205.06 0.98 ;
      RECT  207.33 0.62 209.095 0.98 ;
      RECT  210.675 0.62 210.9 0.98 ;
      RECT  213.545 0.62 214.935 0.98 ;
      RECT  216.515 0.62 216.74 0.98 ;
      RECT  219.01 0.62 219.915 0.98 ;
      RECT  221.495 0.62 222.58 0.98 ;
      RECT  224.85 0.62 228.42 0.98 ;
      RECT  232.265 0.62 234.26 0.98 ;
      RECT  236.66 0.62 240.1 0.98 ;
      RECT  133.7 287.04 135.96 287.4 ;
      RECT  137.54 287.04 137.96 287.4 ;
      RECT  139.54 287.04 140.735 287.4 ;
      RECT  143.525 287.04 143.8 287.4 ;
      RECT  145.38 287.04 146.975 287.4 ;
      RECT  149.415 287.04 149.64 287.4 ;
      RECT  151.22 287.04 153.215 287.4 ;
      RECT  154.795 287.04 155.48 287.4 ;
      RECT  157.75 287.04 159.4 287.4 ;
      RECT  160.98 287.04 161.32 287.4 ;
      RECT  163.625 287.04 165.355 287.4 ;
      RECT  166.935 287.04 167.16 287.4 ;
      RECT  169.865 287.04 171.195 287.4 ;
      RECT  172.775 287.04 173.0 287.4 ;
      RECT  175.27 287.04 176.235 287.4 ;
      RECT  177.815 287.04 178.84 287.4 ;
      RECT  181.11 287.04 182.475 287.4 ;
      RECT  184.055 287.04 184.68 287.4 ;
      RECT  186.26 287.04 187.005 287.4 ;
      RECT  188.585 287.04 190.52 287.4 ;
      RECT  193.505 287.04 196.36 287.4 ;
      RECT  199.685 287.04 202.2 287.4 ;
      RECT  205.925 287.04 208.04 287.4 ;
      RECT  210.9 287.04 211.965 287.4 ;
      RECT  213.545 287.04 213.88 287.4 ;
      RECT  215.46 287.04 215.615 287.4 ;
      RECT  218.405 287.04 219.72 287.4 ;
      RECT  221.3 287.04 221.855 287.4 ;
      RECT  224.645 287.04 225.56 287.4 ;
      RECT  227.14 287.04 228.095 287.4 ;
      RECT  230.885 287.04 231.4 287.4 ;
      RECT  232.98 287.04 234.335 287.4 ;
      RECT  235.915 287.04 237.24 287.4 ;
      RECT  2.34 287.04 79.56 287.4 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  308.74 0.62 369.76 0.98 ;
      RECT  341.6 287.04 369.76 287.4 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 285.14 ;
      RECT  2.34 285.14 2.88 287.04 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 285.14 5.82 287.04 ;
      RECT  5.82 0.98 79.56 2.88 ;
      RECT  5.82 2.88 79.56 285.14 ;
      RECT  5.82 285.14 79.56 287.04 ;
      RECT  104.5 0.98 366.28 2.88 ;
      RECT  104.5 2.88 366.28 285.14 ;
      RECT  104.5 285.14 366.28 287.04 ;
      RECT  366.28 0.98 369.22 2.88 ;
      RECT  366.28 285.14 369.22 287.04 ;
      RECT  369.22 0.98 369.76 2.88 ;
      RECT  369.22 2.88 369.76 285.14 ;
      RECT  369.22 285.14 369.76 287.04 ;
   END
END    dcache_data_ram
END    LIBRARY
