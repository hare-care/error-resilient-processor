VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO icache_tag_ram
   CLASS BLOCK ;
   SIZE 337.22 BY 188.98 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  69.86 0.0 70.24 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.7 0.0 76.08 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.54 0.0 81.92 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.38 0.0 87.76 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.22 0.0 93.6 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.06 0.0 99.44 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.9 0.0 105.28 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.74 0.0 111.12 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.58 0.0 116.96 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.42 0.0 122.8 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.26 0.0 128.64 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.1 0.0 134.48 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.94 0.0 140.32 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.78 0.0 146.16 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.62 0.0 152.0 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.46 0.0 157.84 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.3 0.0 163.68 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.14 0.0 169.52 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.98 0.0 175.36 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.82 0.0 181.2 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.66 0.0 187.04 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.5 0.0 192.88 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  198.34 0.0 198.72 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.18 0.0 204.56 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.02 0.0 210.4 0.38 ;
      END
   END din0[24]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 107.58 0.38 107.96 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 116.08 0.38 116.46 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 121.72 0.38 122.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 130.22 0.38 130.6 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  58.18 188.6 58.56 188.98 ;
      END
   END addr0[4]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  336.84 63.54 337.22 63.92 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.2 0.0 280.58 0.38 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  277.225 0.0 277.605 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  277.915 0.0 278.295 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.66 0.0 279.04 0.38 ;
      END
   END addr1[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  336.84 173.73 337.22 174.11 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.26 0.0 30.64 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.58 188.6 306.96 188.98 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  129.845 188.6 130.225 188.98 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  134.815 188.6 135.195 188.98 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.085 188.6 136.465 188.98 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.055 188.6 141.435 188.98 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.325 188.6 142.705 188.98 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.295 188.6 147.675 188.98 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.565 188.6 148.945 188.98 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.535 188.6 153.915 188.98 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  154.805 188.6 155.185 188.98 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.775 188.6 160.155 188.98 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.045 188.6 161.425 188.98 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.015 188.6 166.395 188.98 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.285 188.6 167.665 188.98 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.255 188.6 172.635 188.98 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.525 188.6 173.905 188.98 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.495 188.6 178.875 188.98 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.765 188.6 180.145 188.98 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.735 188.6 185.115 188.98 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.005 188.6 186.385 188.98 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.975 188.6 191.355 188.98 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.245 188.6 192.625 188.98 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.215 188.6 197.595 188.98 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.485 188.6 198.865 188.98 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.455 188.6 203.835 188.98 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.725 188.6 205.105 188.98 ;
      END
   END dout1[24]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 188.98 ;
         LAYER met3 ;
         RECT  0.0 187.24 337.22 188.98 ;
         LAYER met3 ;
         RECT  0.0 0.0 337.22 1.74 ;
         LAYER met4 ;
         RECT  335.48 0.0 337.22 188.98 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 185.5 ;
         LAYER met3 ;
         RECT  3.48 183.76 333.74 185.5 ;
         LAYER met4 ;
         RECT  332.0 3.48 333.74 185.5 ;
         LAYER met3 ;
         RECT  3.48 3.48 333.74 5.22 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 336.6 188.36 ;
   LAYER  met2 ;
      RECT  0.62 0.62 336.6 188.36 ;
   LAYER  met3 ;
      RECT  0.98 106.98 336.6 108.56 ;
      RECT  0.62 108.56 0.98 115.48 ;
      RECT  0.62 117.06 0.98 121.12 ;
      RECT  0.62 122.7 0.98 129.62 ;
      RECT  0.98 62.94 336.24 64.52 ;
      RECT  0.98 64.52 336.24 106.98 ;
      RECT  336.24 64.52 336.6 106.98 ;
      RECT  0.62 15.85 0.98 106.98 ;
      RECT  0.98 108.56 336.24 173.13 ;
      RECT  0.98 173.13 336.24 174.71 ;
      RECT  336.24 108.56 336.6 173.13 ;
      RECT  0.62 131.2 0.98 186.64 ;
      RECT  336.24 174.71 336.6 186.64 ;
      RECT  336.24 2.34 336.6 62.94 ;
      RECT  0.62 2.34 0.98 14.27 ;
      RECT  0.98 174.71 2.88 183.16 ;
      RECT  0.98 183.16 2.88 186.1 ;
      RECT  0.98 186.1 2.88 186.64 ;
      RECT  2.88 174.71 334.34 183.16 ;
      RECT  2.88 186.1 334.34 186.64 ;
      RECT  334.34 174.71 336.24 183.16 ;
      RECT  334.34 183.16 336.24 186.1 ;
      RECT  334.34 186.1 336.24 186.64 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 62.94 ;
      RECT  2.88 2.34 334.34 2.88 ;
      RECT  2.88 5.82 334.34 62.94 ;
      RECT  334.34 2.34 336.24 2.88 ;
      RECT  334.34 2.88 336.24 5.82 ;
      RECT  334.34 5.82 336.24 62.94 ;
   LAYER  met4 ;
      RECT  69.26 0.98 70.84 188.36 ;
      RECT  70.84 0.62 75.1 0.98 ;
      RECT  76.68 0.62 80.94 0.98 ;
      RECT  82.52 0.62 86.78 0.98 ;
      RECT  88.36 0.62 92.62 0.98 ;
      RECT  94.2 0.62 98.46 0.98 ;
      RECT  100.04 0.62 104.3 0.98 ;
      RECT  105.88 0.62 110.14 0.98 ;
      RECT  111.72 0.62 115.98 0.98 ;
      RECT  117.56 0.62 121.82 0.98 ;
      RECT  123.4 0.62 127.66 0.98 ;
      RECT  129.24 0.62 133.5 0.98 ;
      RECT  135.08 0.62 139.34 0.98 ;
      RECT  140.92 0.62 145.18 0.98 ;
      RECT  146.76 0.62 151.02 0.98 ;
      RECT  152.6 0.62 156.86 0.98 ;
      RECT  158.44 0.62 162.7 0.98 ;
      RECT  164.28 0.62 168.54 0.98 ;
      RECT  170.12 0.62 174.38 0.98 ;
      RECT  175.96 0.62 180.22 0.98 ;
      RECT  181.8 0.62 186.06 0.98 ;
      RECT  187.64 0.62 191.9 0.98 ;
      RECT  193.48 0.62 197.74 0.98 ;
      RECT  199.32 0.62 203.58 0.98 ;
      RECT  205.16 0.62 209.42 0.98 ;
      RECT  57.58 0.98 59.16 188.0 ;
      RECT  59.16 0.98 69.26 188.0 ;
      RECT  59.16 188.0 69.26 188.36 ;
      RECT  211.0 0.62 276.625 0.98 ;
      RECT  31.24 0.62 69.26 0.98 ;
      RECT  70.84 0.98 305.98 188.0 ;
      RECT  305.98 0.98 307.56 188.0 ;
      RECT  70.84 188.0 129.245 188.36 ;
      RECT  130.825 188.0 134.215 188.36 ;
      RECT  137.065 188.0 140.455 188.36 ;
      RECT  143.305 188.0 146.695 188.36 ;
      RECT  149.545 188.0 152.935 188.36 ;
      RECT  155.785 188.0 159.175 188.36 ;
      RECT  162.025 188.0 165.415 188.36 ;
      RECT  168.265 188.0 171.655 188.36 ;
      RECT  174.505 188.0 177.895 188.36 ;
      RECT  180.745 188.0 184.135 188.36 ;
      RECT  186.985 188.0 190.375 188.36 ;
      RECT  193.225 188.0 196.615 188.36 ;
      RECT  199.465 188.0 202.855 188.36 ;
      RECT  205.705 188.0 305.98 188.36 ;
      RECT  2.34 188.0 57.58 188.36 ;
      RECT  2.34 0.62 29.66 0.98 ;
      RECT  281.18 0.62 334.88 0.98 ;
      RECT  307.56 188.0 334.88 188.36 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 186.1 ;
      RECT  2.34 186.1 2.88 188.0 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 186.1 5.82 188.0 ;
      RECT  5.82 0.98 57.58 2.88 ;
      RECT  5.82 2.88 57.58 186.1 ;
      RECT  5.82 186.1 57.58 188.0 ;
      RECT  307.56 0.98 331.4 2.88 ;
      RECT  307.56 2.88 331.4 186.1 ;
      RECT  307.56 186.1 331.4 188.0 ;
      RECT  331.4 0.98 334.34 2.88 ;
      RECT  331.4 186.1 334.34 188.0 ;
      RECT  334.34 0.98 334.88 2.88 ;
      RECT  334.34 2.88 334.88 186.1 ;
      RECT  334.34 186.1 334.88 188.0 ;
   END
END    icache_tag_ram
END    LIBRARY
