magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 2850 897
<< pwell >>
rect 2073 287 2780 315
rect 4 221 422 222
rect 1159 221 1417 287
rect 1807 221 2780 287
rect 4 43 2780 221
rect -26 -43 2810 43
<< locali >>
rect 112 310 178 444
rect 505 309 670 425
rect 2091 439 2178 747
rect 2137 293 2178 439
rect 2692 435 2762 751
rect 2091 135 2178 293
rect 2696 135 2762 435
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2784 831
rect 114 735 232 741
rect 114 701 120 735
rect 154 701 192 735
rect 226 701 232 735
rect 494 735 600 741
rect 22 274 76 646
rect 114 480 232 701
rect 268 682 458 716
rect 268 374 302 682
rect 338 480 388 646
rect 243 274 309 374
rect 22 240 309 274
rect 350 273 388 480
rect 424 495 458 682
rect 528 701 566 735
rect 1053 735 1243 743
rect 1053 701 1059 735
rect 1093 701 1131 735
rect 1165 701 1203 735
rect 1237 701 1243 735
rect 494 531 600 701
rect 636 667 1017 701
rect 636 495 670 667
rect 424 461 670 495
rect 706 531 754 631
rect 22 108 88 240
rect 350 239 668 273
rect 124 113 314 204
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 350 104 384 239
rect 420 113 598 203
rect 124 73 314 79
rect 454 79 492 113
rect 526 79 564 113
rect 420 73 598 79
rect 634 87 668 239
rect 706 187 740 531
rect 790 357 824 667
rect 776 223 824 357
rect 860 415 910 631
rect 951 561 1017 667
rect 1053 597 1243 701
rect 1279 727 1649 761
rect 1279 561 1313 727
rect 951 527 1313 561
rect 951 451 1017 527
rect 1349 491 1383 691
rect 1087 457 1383 491
rect 1087 451 1153 457
rect 1242 415 1308 421
rect 860 381 1308 415
rect 860 203 894 381
rect 930 283 996 345
rect 1242 319 1308 381
rect 930 249 1297 283
rect 1349 265 1383 457
rect 1419 499 1453 727
rect 1489 535 1559 691
rect 1419 441 1485 499
rect 930 239 996 249
rect 704 123 770 187
rect 860 123 926 203
rect 962 87 996 239
rect 634 53 996 87
rect 1037 113 1227 213
rect 1037 79 1043 113
rect 1077 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1227 113
rect 1037 73 1227 79
rect 1263 87 1297 249
rect 1333 123 1399 265
rect 1435 239 1489 373
rect 1435 87 1469 239
rect 1525 203 1559 535
rect 1595 221 1649 727
rect 1701 737 1891 743
rect 1701 703 1707 737
rect 1741 703 1779 737
rect 1813 703 1851 737
rect 1885 703 1891 737
rect 1701 535 1891 703
rect 1685 465 1945 499
rect 1508 137 1559 203
rect 1685 137 1719 465
rect 1755 335 1821 429
rect 1879 371 1945 465
rect 1981 395 2047 743
rect 2214 735 2321 747
rect 2248 701 2286 735
rect 2320 701 2321 735
rect 2214 439 2321 701
rect 2459 735 2649 751
rect 2459 701 2465 735
rect 2499 701 2537 735
rect 2571 701 2609 735
rect 2643 701 2649 735
rect 2357 439 2423 597
rect 1981 335 2101 395
rect 1755 329 2101 335
rect 1755 301 2047 329
rect 1508 103 1719 137
rect 1755 113 1945 265
rect 1263 53 1469 87
rect 1755 79 1761 113
rect 1795 79 1833 113
rect 1867 79 1905 113
rect 1939 79 1945 113
rect 1981 107 2047 301
rect 2361 399 2423 439
rect 2459 435 2649 701
rect 2361 333 2660 399
rect 2214 113 2325 297
rect 2361 201 2427 333
rect 1755 73 1945 79
rect 2214 79 2216 113
rect 2250 79 2288 113
rect 2322 79 2325 113
rect 2214 73 2325 79
rect 2463 113 2653 297
rect 2463 79 2469 113
rect 2503 79 2541 113
rect 2575 79 2613 113
rect 2647 79 2653 113
rect 2463 73 2653 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 120 701 154 735
rect 192 701 226 735
rect 494 701 528 735
rect 566 701 600 735
rect 1059 701 1093 735
rect 1131 701 1165 735
rect 1203 701 1237 735
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 420 79 454 113
rect 492 79 526 113
rect 564 79 598 113
rect 1043 79 1077 113
rect 1115 79 1149 113
rect 1187 79 1221 113
rect 1707 703 1741 737
rect 1779 703 1813 737
rect 1851 703 1885 737
rect 2214 701 2248 735
rect 2286 701 2320 735
rect 2465 701 2499 735
rect 2537 701 2571 735
rect 2609 701 2643 735
rect 1761 79 1795 113
rect 1833 79 1867 113
rect 1905 79 1939 113
rect 2216 79 2250 113
rect 2288 79 2322 113
rect 2469 79 2503 113
rect 2541 79 2575 113
rect 2613 79 2647 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 831 2784 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2784 831
rect 0 791 2784 797
rect 0 737 2784 763
rect 0 735 1707 737
rect 0 701 120 735
rect 154 701 192 735
rect 226 701 494 735
rect 528 701 566 735
rect 600 701 1059 735
rect 1093 701 1131 735
rect 1165 701 1203 735
rect 1237 703 1707 735
rect 1741 703 1779 737
rect 1813 703 1851 737
rect 1885 735 2784 737
rect 1885 703 2214 735
rect 1237 701 2214 703
rect 2248 701 2286 735
rect 2320 701 2465 735
rect 2499 701 2537 735
rect 2571 701 2609 735
rect 2643 701 2784 735
rect 0 689 2784 701
rect 0 113 2784 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 420 113
rect 454 79 492 113
rect 526 79 564 113
rect 598 79 1043 113
rect 1077 79 1115 113
rect 1149 79 1187 113
rect 1221 79 1761 113
rect 1795 79 1833 113
rect 1867 79 1905 113
rect 1939 79 2216 113
rect 2250 79 2288 113
rect 2322 79 2469 113
rect 2503 79 2541 113
rect 2575 79 2613 113
rect 2647 79 2784 113
rect 0 51 2784 79
rect 0 17 2784 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -23 2784 -17
<< labels >>
rlabel locali s 112 310 178 444 6 CLK
port 1 nsew clock input
rlabel locali s 505 309 670 425 6 D
port 2 nsew signal input
rlabel metal1 s 0 51 2784 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 2784 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 2810 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 2780 221 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1807 221 2780 287 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1159 221 1417 287 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 221 422 222 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 2073 287 2780 315 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 2784 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 2850 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 2784 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 2091 135 2178 293 6 Q
port 7 nsew signal output
rlabel locali s 2137 293 2178 439 6 Q
port 7 nsew signal output
rlabel locali s 2091 439 2178 747 6 Q
port 7 nsew signal output
rlabel locali s 2696 135 2762 435 6 Q_N
port 8 nsew signal output
rlabel locali s 2692 435 2762 751 6 Q_N
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2784 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 889718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 861306
<< end >>
