magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal2 >>
rect 99 0 4879 148
rect 5179 0 5579 107
rect 10078 0 14858 148
<< metal3 >>
rect 632 37072 5002 40000
rect 640 37064 5002 37072
rect 670 37034 5002 37064
rect 700 37004 5002 37034
rect 730 36974 5002 37004
rect 760 36944 5002 36974
rect 790 36914 5002 36944
rect 820 36884 5002 36914
rect 850 36854 5002 36884
rect 880 36824 5002 36854
rect 910 36794 5002 36824
rect 940 36764 5002 36794
rect 970 36734 5002 36764
rect 1000 36704 5002 36734
rect 1030 36674 5002 36704
rect 1060 36644 5002 36674
rect 1090 36614 5002 36644
rect 1120 36584 5002 36614
rect 1150 36554 5002 36584
rect 1180 36524 5002 36554
rect 1210 36494 5002 36524
rect 1240 36464 5002 36494
rect 1270 36434 5002 36464
rect 1300 36404 5002 36434
rect 1330 36374 5002 36404
rect 1360 36344 5002 36374
rect 1390 36314 5002 36344
rect 1420 36284 5002 36314
rect 1450 36254 5002 36284
rect 1480 36224 5002 36254
rect 1510 36194 5002 36224
rect 1540 36164 5002 36194
rect 1570 36134 5002 36164
rect 1600 36104 5002 36134
rect 1630 36074 5002 36104
rect 1660 36044 5002 36074
rect 1690 36014 5002 36044
rect 1720 35984 5002 36014
rect 1750 35954 5002 35984
rect 1780 35924 5002 35954
rect 1810 35894 5002 35924
rect 1840 35864 5002 35894
rect 1870 35834 5002 35864
rect 1900 35804 5002 35834
rect 1930 35774 5002 35804
rect 1960 35744 5002 35774
rect 1990 35714 5002 35744
rect 2020 35684 5002 35714
rect 2050 35654 5002 35684
rect 2080 35624 5002 35654
rect 2110 35594 5002 35624
rect 2140 35564 5002 35594
rect 2170 35534 5002 35564
rect 2200 35504 5002 35534
rect 2230 35474 5002 35504
rect 2260 35444 5002 35474
rect 2290 35414 5002 35444
rect 2320 35384 5002 35414
rect 2350 35354 5002 35384
rect 2380 35324 5002 35354
rect 2410 35294 5002 35324
rect 2440 35264 5002 35294
rect 2470 35234 5002 35264
rect 2500 35204 5002 35234
rect 2530 35174 5002 35204
rect 2560 35144 5002 35174
rect 2590 35114 5002 35144
rect 2620 35084 5002 35114
rect 2650 35054 5002 35084
rect 2680 35024 5002 35054
rect 2710 34994 5002 35024
rect 2740 34964 5002 34994
rect 2770 34934 5002 34964
rect 2800 34904 5002 34934
rect 2830 34874 5002 34904
rect 2860 34844 5002 34874
rect 2890 34814 5002 34844
rect 2920 34784 5002 34814
rect 2950 34754 5002 34784
rect 2980 34724 5002 34754
rect 3010 34694 5002 34724
rect 3040 34664 5002 34694
rect 3070 34634 5002 34664
rect 3100 34528 5002 34634
rect 5186 35070 7364 40000
rect 7593 35070 9771 38004
rect 5186 35052 7346 35070
rect 7611 35052 9771 35070
rect 5186 35022 7316 35052
rect 7641 35022 9771 35052
rect 5186 34992 7286 35022
rect 7671 34992 9771 35022
rect 5186 34962 7256 34992
rect 7701 34962 9771 34992
rect 5186 34932 7226 34962
rect 7731 34932 9771 34962
rect 5186 34902 7196 34932
rect 7761 34902 9771 34932
rect 5186 34872 7166 34902
rect 7791 34872 9771 34902
rect 5186 34842 7136 34872
rect 7821 34842 9771 34872
rect 5186 34812 7106 34842
rect 7851 34812 9771 34842
rect 5186 34782 7076 34812
rect 7881 34782 9771 34812
rect 5186 34752 7046 34782
rect 7911 34752 9771 34782
rect 5186 34722 7016 34752
rect 7941 34722 9771 34752
rect 5186 34692 6986 34722
rect 7971 34692 9771 34722
rect 5186 34662 6956 34692
rect 8001 34662 9771 34692
rect 5186 34632 6926 34662
rect 8031 34632 9771 34662
rect 5186 34602 6896 34632
rect 8061 34602 9771 34632
rect 5186 34572 6866 34602
rect 8091 34572 9771 34602
rect 5186 34542 6836 34572
rect 8121 34542 9771 34572
rect 3100 34516 4990 34528
rect 3100 34486 4960 34516
rect 5186 34512 6806 34542
rect 8151 34512 9771 34542
rect 9955 37072 14325 38008
rect 9955 37064 14317 37072
rect 9955 37034 14287 37064
rect 9955 37004 14257 37034
rect 9955 36974 14227 37004
rect 9955 36944 14197 36974
rect 9955 36914 14167 36944
rect 9955 36884 14137 36914
rect 9955 36854 14107 36884
rect 9955 36824 14077 36854
rect 9955 36794 14047 36824
rect 9955 36764 14017 36794
rect 9955 36734 13987 36764
rect 9955 36704 13957 36734
rect 9955 36674 13927 36704
rect 9955 36644 13897 36674
rect 9955 36614 13867 36644
rect 9955 36584 13837 36614
rect 9955 36554 13807 36584
rect 9955 36524 13777 36554
rect 9955 36494 13747 36524
rect 9955 36464 13717 36494
rect 9955 36434 13687 36464
rect 9955 36404 13657 36434
rect 9955 36374 13627 36404
rect 9955 36344 13597 36374
rect 9955 36314 13567 36344
rect 9955 36284 13537 36314
rect 9955 36254 13507 36284
rect 9955 36224 13477 36254
rect 9955 36194 13447 36224
rect 9955 36164 13417 36194
rect 9955 36134 13387 36164
rect 9955 36104 13357 36134
rect 9955 36074 13327 36104
rect 9955 36044 13297 36074
rect 9955 36014 13267 36044
rect 9955 35984 13237 36014
rect 9955 35954 13207 35984
rect 9955 35924 13177 35954
rect 9955 35894 13147 35924
rect 9955 35864 13117 35894
rect 9955 35834 13087 35864
rect 9955 35804 13057 35834
rect 9955 35774 13027 35804
rect 9955 35744 12997 35774
rect 9955 35714 12967 35744
rect 9955 35684 12937 35714
rect 9955 35654 12907 35684
rect 9955 35624 12877 35654
rect 9955 35594 12847 35624
rect 9955 35564 12817 35594
rect 9955 35534 12787 35564
rect 9955 35504 12757 35534
rect 9955 35474 12727 35504
rect 9955 35444 12697 35474
rect 9955 35414 12667 35444
rect 9955 35384 12637 35414
rect 9955 35354 12607 35384
rect 9955 35324 12577 35354
rect 9955 35294 12547 35324
rect 9955 35264 12517 35294
rect 9955 35234 12487 35264
rect 9955 35204 12457 35234
rect 9955 35174 12427 35204
rect 9955 35144 12397 35174
rect 9955 35114 12367 35144
rect 9955 35084 12337 35114
rect 9955 35054 12307 35084
rect 9955 35024 12277 35054
rect 9955 34994 12247 35024
rect 9955 34964 12217 34994
rect 9955 34934 12187 34964
rect 9955 34904 12157 34934
rect 9955 34874 12127 34904
rect 9955 34844 12097 34874
rect 9955 34814 12067 34844
rect 9955 34784 12037 34814
rect 9955 34754 12007 34784
rect 9955 34724 11977 34754
rect 9955 34694 11947 34724
rect 9955 34664 11917 34694
rect 9955 34634 11887 34664
rect 9955 34529 11857 34634
rect 9967 34517 11857 34529
rect 3100 34456 4930 34486
rect 5186 34482 6776 34512
rect 8181 34482 9771 34512
rect 9997 34487 11857 34517
rect 3100 34426 4900 34456
rect 5186 34452 6746 34482
rect 8211 34452 9771 34482
rect 10027 34457 11857 34487
rect 3100 34396 4870 34426
rect 5186 34422 6716 34452
rect 8241 34422 9771 34452
rect 10057 34427 11857 34457
rect 3100 34366 4840 34396
rect 5186 34392 6686 34422
rect 8271 34392 9771 34422
rect 10087 34397 11857 34427
rect 3100 34336 4810 34366
rect 5186 34362 6656 34392
rect 8301 34362 9771 34392
rect 10117 34367 11857 34397
rect 3100 34306 4780 34336
rect 5186 34332 6626 34362
rect 8331 34332 9771 34362
rect 10147 34337 11857 34367
rect 3100 34276 4750 34306
rect 5186 34302 6596 34332
rect 8361 34302 9771 34332
rect 10177 34307 11857 34337
rect 3100 34246 4720 34276
rect 5186 34272 6566 34302
rect 8391 34272 9771 34302
rect 10207 34277 11857 34307
rect 3100 34216 4690 34246
rect 5186 34242 6536 34272
rect 8421 34242 9771 34272
rect 10237 34247 11857 34277
rect 3100 34186 4660 34216
rect 5186 34212 6506 34242
rect 8451 34212 9771 34242
rect 10267 34217 11857 34247
rect 3100 34156 4630 34186
rect 5186 34182 6476 34212
rect 8481 34182 9771 34212
rect 10297 34187 11857 34217
rect 3100 34126 4600 34156
rect 5186 34152 6446 34182
rect 8511 34152 9771 34182
rect 10327 34157 11857 34187
rect 3100 34096 4570 34126
rect 5186 34122 6416 34152
rect 8541 34122 9771 34152
rect 10357 34127 11857 34157
rect 3100 34066 4540 34096
rect 3100 34036 4510 34066
rect 3100 34006 4480 34036
rect 3100 33976 4450 34006
rect 3100 33946 4420 33976
rect 3100 33916 4390 33946
rect 3100 33886 4360 33916
rect 3100 33856 4330 33886
rect 3100 20920 4300 33856
rect 5186 20958 6386 34122
rect 8571 22110 9771 34122
rect 10387 34097 11857 34127
rect 10417 34067 11857 34097
rect 10447 34037 11857 34067
rect 10477 34007 11857 34037
rect 10507 33977 11857 34007
rect 10537 33947 11857 33977
rect 10567 33917 11857 33947
rect 10597 33887 11857 33917
rect 10627 33857 11857 33887
rect 8557 22080 9771 22110
rect 8527 22050 9771 22080
rect 10657 22072 11857 33857
rect 8497 22020 9771 22050
rect 10641 22042 11857 22072
rect 8467 21990 9771 22020
rect 10611 22012 11857 22042
rect 8437 21960 9771 21990
rect 10581 21982 11857 22012
rect 8407 21930 9771 21960
rect 10551 21952 11857 21982
rect 8377 21900 9771 21930
rect 10521 21922 11857 21952
rect 8347 21870 9771 21900
rect 10491 21892 11857 21922
rect 8317 21840 9771 21870
rect 10461 21862 11857 21892
rect 8287 21810 9771 21840
rect 10431 21832 11857 21862
rect 8257 21780 9771 21810
rect 10401 21802 11857 21832
rect 8227 21750 9771 21780
rect 10371 21772 11857 21802
rect 8197 21720 9771 21750
rect 10341 21742 11857 21772
rect 8167 21690 9771 21720
rect 10311 21712 11857 21742
rect 8137 21660 9771 21690
rect 10281 21682 11857 21712
rect 8107 21630 9771 21660
rect 10251 21652 11857 21682
rect 8077 21611 9752 21630
rect 10221 21622 11857 21652
rect 8058 21581 9722 21611
rect 10191 21592 11857 21622
rect 8028 21551 9692 21581
rect 10161 21563 11828 21592
rect 7998 21521 9662 21551
rect 10132 21533 11798 21563
rect 7968 21491 9632 21521
rect 10102 21503 11768 21533
rect 7938 21461 9602 21491
rect 10072 21473 11738 21503
rect 7908 21431 9572 21461
rect 10042 21443 11708 21473
rect 7878 21401 9542 21431
rect 10012 21413 11678 21443
rect 7848 21371 9512 21401
rect 9982 21383 11648 21413
rect 7818 21341 9482 21371
rect 9952 21353 11618 21383
rect 7788 21311 9452 21341
rect 9922 21323 11588 21353
rect 7758 21281 9422 21311
rect 9892 21293 11558 21323
rect 7728 21251 9392 21281
rect 9862 21263 11528 21293
rect 7698 21221 9362 21251
rect 9832 21233 11498 21263
rect 7668 21191 9332 21221
rect 9802 21203 11468 21233
rect 7638 21161 9302 21191
rect 9772 21173 11438 21203
rect 7608 21131 9272 21161
rect 9742 21143 11408 21173
rect 7578 21117 9258 21131
rect 7578 21087 9228 21117
rect 9712 21113 11378 21143
rect 7578 21057 9198 21087
rect 9682 21083 11348 21113
rect 7578 21027 9168 21057
rect 9652 21053 11318 21083
rect 7578 20997 9138 21027
rect 9622 21023 11288 21053
rect 7578 20967 9108 20997
rect 9592 20993 11258 21023
rect 5186 20928 6400 20958
rect 7578 20937 9078 20967
rect 9562 20963 11228 20993
rect 3100 20890 4316 20920
rect 5186 20898 6430 20928
rect 7578 20907 9048 20937
rect 9532 20933 11198 20963
rect 3100 20860 4346 20890
rect 5186 20868 6460 20898
rect 7578 20877 9018 20907
rect 9502 20903 11168 20933
rect 3100 20830 4376 20860
rect 5186 20838 6490 20868
rect 7578 20847 8988 20877
rect 9472 20873 11138 20903
rect 3100 20800 4406 20830
rect 5186 20808 6520 20838
rect 7578 20817 8958 20847
rect 9442 20843 11108 20873
rect 3100 20770 4436 20800
rect 5186 20778 6550 20808
rect 7578 20787 8928 20817
rect 9412 20813 11078 20843
rect 3100 20740 4466 20770
rect 5186 20748 6580 20778
rect 7578 20757 8898 20787
rect 9382 20783 11048 20813
rect 3100 20710 4496 20740
rect 5186 20718 6610 20748
rect 7578 20727 8868 20757
rect 9352 20753 11018 20783
rect 3100 20680 4526 20710
rect 5186 20688 6640 20718
rect 7578 20697 8838 20727
rect 9322 20723 10988 20753
rect 3100 20650 4556 20680
rect 5186 20658 6670 20688
rect 7578 20667 8808 20697
rect 9292 20693 10958 20723
rect 3100 20620 4586 20650
rect 5186 20628 6700 20658
rect 7578 20637 8778 20667
rect 9262 20663 10928 20693
rect 3100 20590 4616 20620
rect 5186 20598 6730 20628
rect 7578 20607 8748 20637
rect 9232 20633 10898 20663
rect 3100 20560 4646 20590
rect 5186 20568 6760 20598
rect 7578 20577 8718 20607
rect 9202 20603 10868 20633
rect 3100 20530 4676 20560
rect 5186 20538 6790 20568
rect 7578 20547 8688 20577
rect 9172 20573 10838 20603
rect 3100 20500 4706 20530
rect 5186 20508 6820 20538
rect 7578 20517 8658 20547
rect 9142 20543 10808 20573
rect 3100 20470 4736 20500
rect 5186 20478 6850 20508
rect 7578 20487 8628 20517
rect 9112 20513 10778 20543
rect 3100 20440 4766 20470
rect 5205 20459 6880 20478
rect 3129 20411 4796 20440
rect 5235 20429 6899 20459
rect 7578 20457 8598 20487
rect 9082 20483 10748 20513
rect 9052 20463 10728 20483
rect 3159 20381 4825 20411
rect 5265 20399 6929 20429
rect 3189 20351 4855 20381
rect 5295 20369 6959 20399
rect 3219 20321 4885 20351
rect 5325 20339 6989 20369
rect 3249 20291 4915 20321
rect 5355 20309 7019 20339
rect 3279 20261 4945 20291
rect 5385 20279 7049 20309
rect 3309 20231 4975 20261
rect 5415 20249 7079 20279
rect 3339 20201 5005 20231
rect 5445 20219 7109 20249
rect 3369 20171 5035 20201
rect 5475 20189 7139 20219
rect 3399 20141 5065 20171
rect 5505 20159 7169 20189
rect 3429 20111 5095 20141
rect 5535 20129 7199 20159
rect 3459 20081 5125 20111
rect 5565 20099 7229 20129
rect 3489 20051 5155 20081
rect 5595 20069 7259 20099
rect 3519 20021 5185 20051
rect 5625 20039 7289 20069
rect 3549 19991 5215 20021
rect 5655 20009 7319 20039
rect 7578 20021 8568 20457
rect 9052 20433 10698 20463
rect 9052 20403 10668 20433
rect 9052 20373 10638 20403
rect 9052 20343 10608 20373
rect 9052 20313 10578 20343
rect 9052 20283 10548 20313
rect 9052 20253 10518 20283
rect 12300 20257 14858 34664
rect 9052 20223 10488 20253
rect 12298 20227 14858 20257
rect 9052 20193 10458 20223
rect 12268 20197 14858 20227
rect 9052 20163 10428 20193
rect 12238 20167 14858 20197
rect 9052 20133 10398 20163
rect 12208 20137 14858 20167
rect 9052 20103 10368 20133
rect 12178 20107 14858 20137
rect 9052 20073 10338 20103
rect 12148 20077 14858 20107
rect 9052 20043 10308 20073
rect 12118 20047 14858 20077
rect 9052 20033 10298 20043
rect 3579 19961 5245 19991
rect 5685 19979 7349 20009
rect 7578 19991 8590 20021
rect 9042 20003 10268 20033
rect 12088 20017 14858 20047
rect 5699 19965 7379 19979
rect 3609 19931 5275 19961
rect 5729 19935 7379 19965
rect 3639 19901 5305 19931
rect 5759 19905 7379 19935
rect 3669 19871 5335 19901
rect 5789 19875 7379 19905
rect 3699 19841 5365 19871
rect 5819 19845 7379 19875
rect 3729 19811 5395 19841
rect 5849 19815 7379 19845
rect 3759 19781 5425 19811
rect 5879 19785 7379 19815
rect 3789 19751 5455 19781
rect 5909 19755 7379 19785
rect 3819 19721 5485 19751
rect 5939 19725 7379 19755
rect 3849 19691 5515 19721
rect 5969 19695 7379 19725
rect 3879 19661 5545 19691
rect 5999 19665 7379 19695
rect 3909 19631 5575 19661
rect 6029 19635 7379 19665
rect 3939 19601 5605 19631
rect 6059 19605 7379 19635
rect 3969 19571 5635 19601
rect 6089 19575 7379 19605
rect 3999 19541 5665 19571
rect 6119 19545 7379 19575
rect 4029 19511 5695 19541
rect 6149 19515 7379 19545
rect 4059 19481 5725 19511
rect 6179 19485 7379 19515
rect 4089 19451 5755 19481
rect 6209 19455 7379 19485
rect 4119 19421 5785 19451
rect 6239 19425 7379 19455
rect 4149 19391 5815 19421
rect 6269 19395 7379 19425
rect 4179 19361 5845 19391
rect 6299 19365 7379 19395
rect 4209 19331 5875 19361
rect 6329 19335 7379 19365
rect 4239 19301 5905 19331
rect 6359 19305 7379 19335
rect 4269 19271 5905 19301
rect 4299 19241 5905 19271
rect 4329 19211 5905 19241
rect 4359 19181 5905 19211
rect 4389 19151 5905 19181
rect 4419 19121 5905 19151
rect 4449 19091 5905 19121
rect 4479 19061 5905 19091
rect 4509 19031 5905 19061
rect 4539 19001 5905 19031
rect 4569 18971 5905 19001
rect 4599 18941 5905 18971
rect 4629 18911 5905 18941
rect 4659 18881 5905 18911
rect 4689 18851 5905 18881
rect 4719 18821 5905 18851
rect 4749 18598 5905 18821
rect 6389 18598 7379 19305
rect 4749 18568 5927 18598
rect 6367 18568 7379 18598
rect 4749 18538 5957 18568
rect 6337 18538 7379 18568
rect 4749 18508 5987 18538
rect 6307 18508 7379 18538
rect 4764 18493 6017 18508
rect 4779 18478 6032 18493
rect 6277 18478 7379 18508
rect 4789 18468 7379 18478
rect 4819 18438 7379 18468
rect 4849 18408 7379 18438
rect 4879 18378 7379 18408
rect 4909 18348 7379 18378
rect 4939 18318 7379 18348
rect 4969 18288 7379 18318
rect 4999 18258 7379 18288
rect 5029 18228 7379 18258
rect 5059 18198 7379 18228
rect 5089 18168 7379 18198
rect 5119 18138 7379 18168
rect 5149 18108 7379 18138
rect 99 0 4879 391
rect 5179 0 7379 18108
rect 7578 19961 8620 19991
rect 9012 19973 10238 20003
rect 12058 19987 14858 20017
rect 7578 19931 8650 19961
rect 8982 19943 10208 19973
rect 12028 19957 14858 19987
rect 7578 19901 8680 19931
rect 8952 19922 10208 19943
rect 11998 19927 14858 19957
rect 8931 19901 10208 19922
rect 7578 19660 10208 19901
rect 11968 19897 14858 19927
rect 11938 19867 14858 19897
rect 11908 19837 14858 19867
rect 11878 19807 14858 19837
rect 11848 19777 14858 19807
rect 11818 19747 14858 19777
rect 11788 19717 14858 19747
rect 11758 19687 14858 19717
rect 7578 19650 10198 19660
rect 11728 19657 14858 19687
rect 7578 19620 10168 19650
rect 11698 19627 14858 19657
rect 7578 19590 10138 19620
rect 11668 19597 14858 19627
rect 7578 19560 10108 19590
rect 11638 19567 14858 19597
rect 7578 19530 10078 19560
rect 11608 19537 14858 19567
rect 7578 19500 10048 19530
rect 11578 19507 14858 19537
rect 7578 19470 10018 19500
rect 11548 19477 14858 19507
rect 7578 19440 9988 19470
rect 11518 19447 14858 19477
rect 7578 19410 9958 19440
rect 11488 19417 14858 19447
rect 7578 19380 9928 19410
rect 11458 19387 14858 19417
rect 7578 19350 9898 19380
rect 11428 19357 14858 19387
rect 7578 19320 9868 19350
rect 11398 19327 14858 19357
rect 7578 19290 9838 19320
rect 11368 19297 14858 19327
rect 7578 19260 9808 19290
rect 11338 19267 14858 19297
rect 7578 0 9778 19260
rect 11308 19237 14858 19267
rect 11278 19207 14858 19237
rect 11248 19177 14858 19207
rect 11218 19147 14858 19177
rect 11188 19117 14858 19147
rect 11158 19087 14858 19117
rect 11128 19057 14858 19087
rect 11098 19027 14858 19057
rect 11068 18997 14858 19027
rect 11038 18967 14858 18997
rect 11008 18937 14858 18967
rect 10978 18907 14858 18937
rect 10948 18877 14858 18907
rect 10918 18847 14858 18877
rect 10888 18817 14858 18847
rect 10858 18787 14858 18817
rect 10828 18757 14858 18787
rect 10798 18727 14858 18757
rect 10768 18697 14858 18727
rect 10738 18667 14858 18697
rect 10708 18637 14858 18667
rect 10678 18607 14858 18637
rect 10648 18577 14858 18607
rect 10618 18547 14858 18577
rect 10588 18517 14858 18547
rect 10558 18487 14858 18517
rect 10528 18457 14858 18487
rect 10498 18427 14858 18457
rect 10468 18397 14858 18427
rect 10438 18367 14858 18397
rect 10408 18337 14858 18367
rect 10378 18307 14858 18337
rect 10348 18277 14858 18307
rect 10318 18247 14858 18277
rect 10288 18217 14858 18247
rect 10258 18187 14858 18217
rect 10228 18157 14858 18187
rect 10198 18127 14858 18157
rect 10168 18097 14858 18127
rect 10138 18067 14858 18097
rect 10108 18037 14858 18067
rect 10078 0 14858 391
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 7329 27865 7594 29187
rect 0 14007 15000 18997
rect 0 12837 15000 13687
rect 0 11667 15000 12517
rect 0 9547 15000 11347
rect 0 8337 15000 9227
rect 0 7367 15000 8017
rect 0 6397 15000 7047
rect 0 5187 15000 6077
rect 0 3977 15000 4867
rect 0 3007 15000 3657
rect 0 1797 15000 2687
rect 0 427 15000 1477
use sky130_fd_io__hvc_clampv2  sky130_fd_io__hvc_clampv2_0
timestamp 1694700623
transform 1 0 0 0 1 0
box 0 0 15000 40000
<< labels >>
flabel metal3 s 99 0 4879 391 0 FreeSans 96 0 0 0 P_CORE
port 3 nsew power bidirectional
flabel metal3 s 13490 13244 13490 13244 0 FreeSans 596 0 0 0 PADISOR
port 1 nsew
flabel metal3 s 1010 13244 1010 13244 0 FreeSans 596 0 0 0 PADISOL
port 2 nsew
flabel metal3 s 7578 0 9778 318 0 FreeSans 96 0 0 0 DRN_HVC
port 4 nsew power bidirectional
flabel metal3 s 10078 0 14858 391 0 FreeSans 96 0 0 0 P_CORE
port 3 nsew power bidirectional
flabel metal3 s 5179 0 7379 148 2 FreeSans 96 90 0 0 SRC_BDY_HVC
port 5 nsew ground bidirectional
flabel metal2 s 10078 0 14858 148 2 FreeSans 44 90 0 0 DRN_HVC
port 4 nsew power bidirectional
flabel metal2 s 99 0 4879 148 2 FreeSans 44 90 0 0 SRC_BDY_HVC
port 5 nsew ground bidirectional
flabel metal2 s 5179 0 5579 107 2 FreeSans 1000 90 0 0 OGC_HVC
port 6 nsew power bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 9 nsew ground bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 10 nsew signal bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 14 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 16 nsew power bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 17 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 18 nsew power bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 19 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 9 nsew ground bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 10 nsew signal bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 14 nsew power bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 16 nsew power bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 17 nsew power bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 18 nsew power bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 19 nsew ground bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal4 s 127 38321 127 38321 3 FreeSans 520 0 0 0 VSSIO
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal4 s 14873 38321 14873 38321 3 FreeSans 520 180 0 0 VSSIO
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 7329 27865 7594 29187 0 FreeSans 512 0 0 0 P_PAD
port 21 nsew signal bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 19 nsew ground bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 14 nsew power bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 17 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 18 nsew power bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 16 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 9 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 15 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 14 nsew power bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 19 nsew ground bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 17 nsew power bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 18 nsew power bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 16 nsew power bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 13 nsew power bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 9 nsew ground bidirectional
rlabel metal3 s 10657 33827 11857 33857 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 22088 11857 33827 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 22072 11857 22088 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10641 22042 11857 22072 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10627 33857 11857 33887 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10611 22012 11857 22042 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10597 33887 11857 33917 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10581 21982 11857 22012 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10567 33917 11857 33947 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10551 21952 11857 21982 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10537 33947 11857 33977 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10521 21922 11857 21952 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10507 33977 11857 34007 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10491 21892 11857 21922 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10477 34007 11857 34037 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10461 21862 11857 21892 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10447 34037 11857 34067 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10431 21832 11857 21862 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10417 34067 11857 34097 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10401 21802 11857 21832 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10387 34097 11857 34127 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10371 21772 11857 21802 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10357 34127 11857 34157 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10341 21742 11857 21772 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10327 34157 11857 34187 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10311 21712 11857 21742 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10297 34187 11857 34217 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10281 21682 11857 21712 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10267 34217 11857 34247 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10251 21652 11857 21682 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10237 34247 11857 34277 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10221 21622 11857 21652 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10207 34277 11857 34307 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10191 21592 11857 21622 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10177 34307 11857 34337 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10161 21563 11828 21592 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10147 34337 11857 34367 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10132 21533 11798 21563 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10117 34367 11857 34397 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10102 21503 11768 21533 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10087 34397 11857 34427 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10072 21473 11738 21503 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10057 34427 11857 34457 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10042 21443 11708 21473 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10027 34457 11857 34487 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10012 21413 11678 21443 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9997 34487 11857 34517 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9982 21383 11648 21413 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9967 34517 11857 34529 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37072 14325 38008 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37064 14317 37072 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37034 14287 37064 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 37004 14257 37034 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36974 14227 37004 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36944 14197 36974 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36914 14167 36944 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36884 14137 36914 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36854 14107 36884 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36824 14077 36854 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36794 14047 36824 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36764 14017 36794 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36734 13987 36764 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36704 13957 36734 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36674 13927 36704 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36644 13897 36674 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36614 13867 36644 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36584 13837 36614 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36554 13807 36584 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36524 13777 36554 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36494 13747 36524 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36464 13717 36494 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36434 13687 36464 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36404 13657 36434 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36374 13627 36404 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36344 13597 36374 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36314 13567 36344 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36284 13537 36314 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36254 13507 36284 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36224 13477 36254 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36194 13447 36224 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36164 13417 36194 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36134 13387 36164 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36104 13357 36134 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36074 13327 36104 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36044 13297 36074 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 36014 13267 36044 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35984 13237 36014 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35954 13207 35984 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35924 13177 35954 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35894 13147 35924 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35864 13117 35894 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35834 13087 35864 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35804 13057 35834 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35774 13027 35804 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35744 12997 35774 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35714 12967 35744 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35684 12937 35714 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35654 12907 35684 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35624 12877 35654 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35594 12847 35624 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35564 12817 35594 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35534 12787 35564 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35504 12757 35534 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35474 12727 35504 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35444 12697 35474 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35414 12667 35444 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35384 12637 35414 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35354 12607 35384 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35324 12577 35354 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35294 12547 35324 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35264 12517 35294 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35234 12487 35264 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35204 12457 35234 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35174 12427 35204 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35144 12397 35174 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35114 12367 35144 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35084 12337 35114 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35054 12307 35084 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 35024 12277 35054 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34994 12247 35024 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34964 12217 34994 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34934 12187 34964 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34904 12157 34934 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34874 12127 34904 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34844 12097 34874 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34814 12067 34844 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34784 12037 34814 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34754 12007 34784 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34724 11977 34754 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34694 11947 34724 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34664 11917 34694 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34634 11887 34664 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34604 11857 34634 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34529 11857 34604 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9952 21353 11618 21383 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9922 21323 11588 21353 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9892 21293 11558 21323 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9862 21263 11528 21293 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9832 21233 11498 21263 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9802 21203 11468 21233 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9772 21173 11438 21203 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9742 21143 11408 21173 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9712 21113 11378 21143 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9682 21083 11348 21113 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9652 21053 11318 21083 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9622 21023 11288 21053 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9592 20993 11258 21023 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9562 20963 11228 20993 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9532 20933 11198 20963 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9502 20903 11168 20933 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9472 20873 11138 20903 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9442 20843 11108 20873 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9412 20813 11078 20843 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9382 20783 11048 20813 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9352 20753 11018 20783 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9322 20723 10988 20753 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9292 20693 10958 20723 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9262 20663 10928 20693 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9232 20633 10898 20663 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9202 20603 10868 20633 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9172 20573 10838 20603 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9142 20543 10808 20573 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9112 20513 10778 20543 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9082 20483 10748 20513 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20463 10728 20483 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20433 10698 20463 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20403 10668 20433 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20373 10638 20403 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20343 10608 20373 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20313 10578 20343 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20283 10548 20313 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20253 10518 20283 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20223 10488 20253 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20193 10458 20223 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20163 10428 20193 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20133 10398 20163 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20103 10368 20133 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20073 10338 20103 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20043 10308 20073 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20033 10298 20043 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9042 20003 10268 20033 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9012 19973 10238 20003 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8982 19943 10208 19973 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8952 19922 10208 19943 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8931 19901 10208 19922 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 34092 9771 34122 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 22124 9771 34092 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 22110 9771 22124 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8557 22080 9771 22110 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8541 34122 9771 34152 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8527 22050 9771 22080 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8511 34152 9771 34182 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8497 22020 9771 22050 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8481 34182 9771 34212 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8467 21990 9771 22020 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8451 34212 9771 34242 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8437 21960 9771 21990 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8421 34242 9771 34272 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8407 21930 9771 21960 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8391 34272 9771 34302 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8377 21900 9771 21930 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8361 34302 9771 34332 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8347 21870 9771 21900 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8331 34332 9771 34362 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8317 21840 9771 21870 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8301 34362 9771 34392 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8287 21810 9771 21840 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8271 34392 9771 34422 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8257 21780 9771 21810 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8241 34422 9771 34452 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8227 21750 9771 21780 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8211 34452 9771 34482 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8197 21720 9771 21750 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8181 34482 9771 34512 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8167 21690 9771 21720 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8151 34512 9771 34542 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8137 21660 9771 21690 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8121 34542 9771 34572 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8107 21630 9771 21660 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8091 34572 9771 34602 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8077 21611 9752 21630 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8061 34602 9771 34632 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8058 21581 9722 21611 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8031 34632 9771 34662 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8028 21551 9692 21581 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8001 34662 9771 34692 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7998 21521 9662 21551 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7971 34692 9771 34722 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7968 21491 9632 21521 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7941 34722 9771 34752 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7938 21461 9602 21491 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7911 34752 9771 34782 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7908 21431 9572 21461 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7881 34782 9771 34812 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7878 21401 9542 21431 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7851 34812 9771 34842 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7848 21371 9512 21401 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7821 34842 9771 34872 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7818 21341 9482 21371 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7791 34872 9771 34902 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7788 21311 9452 21341 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7761 34902 9771 34932 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7758 21281 9422 21311 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7731 34932 9771 34962 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7728 21251 9392 21281 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7701 34962 9771 34992 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7698 21221 9362 21251 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7671 34992 9771 35022 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7668 21191 9332 21221 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7641 35022 9771 35052 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7638 21161 9302 21191 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7611 35052 9771 35070 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7608 21131 9272 21161 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7593 35070 9771 38004 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21117 9258 21131 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21087 9228 21117 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21057 9198 21087 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21027 9168 21057 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20997 9138 21027 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20967 9108 20997 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20937 9078 20967 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20907 9048 20937 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20877 9018 20907 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20847 8988 20877 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20817 8958 20847 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20787 8928 20817 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20757 8898 20787 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20727 8868 20757 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20697 8838 20727 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20667 8808 20697 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20637 8778 20667 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20607 8748 20637 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20577 8718 20607 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20547 8688 20577 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20517 8658 20547 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20487 8628 20517 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20457 8598 20487 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20427 8568 20457 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20043 8568 20427 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20021 8568 20043 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19991 8590 20021 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19961 8620 19991 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19931 8650 19961 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19901 8680 19931 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19660 10208 19901 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19650 10198 19660 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19620 10168 19650 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19590 10138 19620 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19560 10108 19590 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19530 10078 19560 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19500 10048 19530 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19470 10018 19500 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19440 9988 19470 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19410 9958 19440 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19380 9928 19410 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19350 9898 19380 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19320 9868 19350 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19290 9838 19320 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19260 9808 19290 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19230 9778 19260 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 0 9778 19230 1 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 12300 20259 14858 34664 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12300 20257 14858 20259 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12298 20227 14858 20257 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12268 20197 14858 20227 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12238 20167 14858 20197 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12208 20137 14858 20167 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12178 20107 14858 20137 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12148 20077 14858 20107 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12118 20047 14858 20077 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12088 20017 14858 20047 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12058 19987 14858 20017 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 12028 19957 14858 19987 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11998 19927 14858 19957 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11968 19897 14858 19927 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11938 19867 14858 19897 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11908 19837 14858 19867 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11878 19807 14858 19837 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11848 19777 14858 19807 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11818 19747 14858 19777 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11788 19717 14858 19747 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11758 19687 14858 19717 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11728 19657 14858 19687 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11698 19627 14858 19657 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11668 19597 14858 19627 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11638 19567 14858 19597 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11608 19537 14858 19567 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11578 19507 14858 19537 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11548 19477 14858 19507 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11518 19447 14858 19477 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11488 19417 14858 19447 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11458 19387 14858 19417 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11428 19357 14858 19387 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11398 19327 14858 19357 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11368 19297 14858 19327 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11338 19267 14858 19297 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11308 19237 14858 19267 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11278 19207 14858 19237 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11248 19177 14858 19207 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11218 19147 14858 19177 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11188 19117 14858 19147 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11158 19087 14858 19117 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11128 19057 14858 19087 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11098 19027 14858 19057 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11068 18997 14858 19027 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11038 18967 14858 18997 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 11008 18937 14858 18967 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10978 18907 14858 18937 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10948 18877 14858 18907 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10918 18847 14858 18877 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10888 18817 14858 18847 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10858 18787 14858 18817 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10828 18757 14858 18787 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10798 18727 14858 18757 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10768 18697 14858 18727 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10738 18667 14858 18697 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10708 18637 14858 18667 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10678 18607 14858 18637 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10648 18577 14858 18607 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10618 18547 14858 18577 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10588 18517 14858 18547 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10558 18487 14858 18517 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10528 18457 14858 18487 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10498 18427 14858 18457 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10468 18397 14858 18427 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10438 18367 14858 18397 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10408 18337 14858 18367 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10378 18307 14858 18337 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10348 18277 14858 18307 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10318 18247 14858 18277 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10288 18217 14858 18247 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10258 18187 14858 18217 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10228 18157 14858 18187 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10198 18127 14858 18157 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10168 18097 14858 18127 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10138 18067 14858 18097 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 10108 18037 14858 18067 1 P_CORE
port 3 nsew power bidirectional
rlabel metal3 s 6389 19275 7379 19305 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6389 18620 7379 19275 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6389 18598 7379 18620 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6367 18568 7379 18598 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6359 19305 7379 19335 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6337 18538 7379 18568 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6329 19335 7379 19365 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6307 18508 7379 18538 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6299 19365 7379 19395 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6277 18478 7379 18508 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6269 19395 7379 19425 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6239 19425 7379 19455 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6209 19455 7379 19485 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6179 19485 7379 19515 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6149 19515 7379 19545 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6119 19545 7379 19575 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6089 19575 7379 19605 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6059 19605 7379 19635 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 6029 19635 7379 19665 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5999 19665 7379 19695 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5969 19695 7379 19725 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5939 19725 7379 19755 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5909 19755 7379 19785 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5879 19785 7379 19815 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5849 19815 7379 19845 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5819 19845 7379 19875 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5789 19875 7379 19905 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5759 19905 7379 19935 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5729 19935 7379 19965 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5699 19965 7379 19979 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5685 19979 7349 20009 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5655 20009 7319 20039 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5625 20039 7289 20069 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5595 20069 7259 20099 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5565 20099 7229 20129 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5535 20129 7199 20159 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5505 20159 7169 20189 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5475 20189 7139 20219 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5445 20219 7109 20249 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5415 20249 7079 20279 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5385 20279 7049 20309 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5355 20309 7019 20339 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5325 20339 6989 20369 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5295 20369 6959 20399 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5265 20399 6929 20429 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5235 20429 6899 20459 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5205 20459 6880 20478 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 35070 7364 40000 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 35052 7346 35070 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 35022 7316 35052 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34992 7286 35022 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34962 7256 34992 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34932 7226 34962 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34902 7196 34932 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34872 7166 34902 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34842 7136 34872 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34812 7106 34842 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34782 7076 34812 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34752 7046 34782 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34722 7016 34752 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34692 6986 34722 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34662 6956 34692 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34632 6926 34662 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34602 6896 34632 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34572 6866 34602 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34542 6836 34572 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34512 6806 34542 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34482 6776 34512 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34452 6746 34482 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34422 6716 34452 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34392 6686 34422 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34362 6656 34392 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34332 6626 34362 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34302 6596 34332 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34272 6566 34302 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34242 6536 34272 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34212 6506 34242 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34182 6476 34212 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34152 6446 34182 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34122 6416 34152 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 34092 6386 34122 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20972 6386 34092 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20958 6386 20972 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20928 6400 20958 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20898 6430 20928 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20868 6460 20898 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20838 6490 20868 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20808 6520 20838 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20778 6550 20808 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20748 6580 20778 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20718 6610 20748 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20688 6640 20718 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20658 6670 20688 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20628 6700 20658 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20598 6730 20628 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20568 6760 20598 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20538 6790 20568 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20508 6820 20538 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5186 20478 6850 20508 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5179 18078 7379 18108 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5179 0 7379 18078 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5149 18108 7379 18138 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5119 18138 7379 18168 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5089 18168 7379 18198 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5059 18198 7379 18228 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 5029 18228 7379 18258 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4999 18258 7379 18288 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4969 18288 7379 18318 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4939 18318 7379 18348 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4909 18348 7379 18378 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4879 18378 7379 18408 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4849 18408 7379 18438 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4819 18438 7379 18468 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4789 18468 7379 18478 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4779 18478 6032 18493 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4764 18493 6017 18508 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18791 5905 18821 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18620 5905 18791 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18598 5905 18620 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18568 5927 18598 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18538 5957 18568 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4749 18508 5987 18538 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4719 18821 5905 18851 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4689 18851 5905 18881 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4659 18881 5905 18911 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4629 18911 5905 18941 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4599 18941 5905 18971 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4569 18971 5905 19001 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4539 19001 5905 19031 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4509 19031 5905 19061 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4479 19061 5905 19091 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4449 19091 5905 19121 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4419 19121 5905 19151 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4389 19151 5905 19181 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4359 19181 5905 19211 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4329 19211 5905 19241 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4299 19241 5905 19271 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4269 19271 5905 19301 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4239 19301 5905 19331 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4209 19331 5875 19361 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4179 19361 5845 19391 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4149 19391 5815 19421 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4119 19421 5785 19451 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4089 19451 5755 19481 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4059 19481 5725 19511 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 4029 19511 5695 19541 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3999 19541 5665 19571 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3969 19571 5635 19601 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3939 19601 5605 19631 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3909 19631 5575 19661 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3879 19661 5545 19691 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3849 19691 5515 19721 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3819 19721 5485 19751 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3789 19751 5455 19781 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3759 19781 5425 19811 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3729 19811 5395 19841 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3699 19841 5365 19871 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3669 19871 5335 19901 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3639 19901 5305 19931 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3609 19931 5275 19961 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3579 19961 5245 19991 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3549 19991 5215 20021 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3519 20021 5185 20051 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3489 20051 5155 20081 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3459 20081 5125 20111 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3429 20111 5095 20141 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3399 20141 5065 20171 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3369 20171 5035 20201 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3339 20201 5005 20231 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3309 20231 4975 20261 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3279 20261 4945 20291 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3249 20291 4915 20321 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3219 20321 4885 20351 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3189 20351 4855 20381 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3159 20381 4825 20411 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3129 20411 4796 20440 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34604 5002 34634 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34528 5002 34604 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34516 4990 34528 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34486 4960 34516 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34456 4930 34486 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34426 4900 34456 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34396 4870 34426 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34366 4840 34396 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34336 4810 34366 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34306 4780 34336 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34276 4750 34306 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34246 4720 34276 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34216 4690 34246 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34186 4660 34216 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34156 4630 34186 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34126 4600 34156 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34096 4570 34126 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34066 4540 34096 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34036 4510 34066 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 34006 4480 34036 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33976 4450 34006 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33946 4420 33976 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33916 4390 33946 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33886 4360 33916 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33856 4330 33886 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 33826 4300 33856 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20936 4300 33826 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20920 4300 20936 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20890 4316 20920 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20860 4346 20890 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20830 4376 20860 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20800 4406 20830 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20770 4436 20800 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20740 4466 20770 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20710 4496 20740 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20680 4526 20710 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20650 4556 20680 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20620 4586 20650 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20590 4616 20620 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20560 4646 20590 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20530 4676 20560 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20500 4706 20530 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20470 4736 20500 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3100 20440 4766 20470 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3070 34634 5002 34664 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3040 34664 5002 34694 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 3010 34694 5002 34724 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2980 34724 5002 34754 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2950 34754 5002 34784 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2920 34784 5002 34814 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2890 34814 5002 34844 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2860 34844 5002 34874 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2830 34874 5002 34904 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2800 34904 5002 34934 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2770 34934 5002 34964 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2740 34964 5002 34994 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2710 34994 5002 35024 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2680 35024 5002 35054 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2650 35054 5002 35084 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2620 35084 5002 35114 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2590 35114 5002 35144 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2560 35144 5002 35174 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2530 35174 5002 35204 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2500 35204 5002 35234 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2470 35234 5002 35264 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2440 35264 5002 35294 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2410 35294 5002 35324 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2380 35324 5002 35354 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2350 35354 5002 35384 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2320 35384 5002 35414 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2290 35414 5002 35444 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2260 35444 5002 35474 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2230 35474 5002 35504 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2200 35504 5002 35534 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2170 35534 5002 35564 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2140 35564 5002 35594 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2110 35594 5002 35624 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2080 35624 5002 35654 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2050 35654 5002 35684 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 2020 35684 5002 35714 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1990 35714 5002 35744 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1960 35744 5002 35774 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1930 35774 5002 35804 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1900 35804 5002 35834 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1870 35834 5002 35864 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1840 35864 5002 35894 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1810 35894 5002 35924 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1780 35924 5002 35954 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1750 35954 5002 35984 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1720 35984 5002 36014 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1690 36014 5002 36044 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1660 36044 5002 36074 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1630 36074 5002 36104 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1600 36104 5002 36134 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1570 36134 5002 36164 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1540 36164 5002 36194 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1510 36194 5002 36224 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1480 36224 5002 36254 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1450 36254 5002 36284 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1420 36284 5002 36314 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1390 36314 5002 36344 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1360 36344 5002 36374 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1330 36374 5002 36404 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1300 36404 5002 36434 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1270 36434 5002 36464 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1240 36464 5002 36494 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1210 36494 5002 36524 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1180 36524 5002 36554 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1150 36554 5002 36584 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1120 36584 5002 36614 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1090 36614 5002 36644 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1060 36644 5002 36674 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1030 36674 5002 36704 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 1000 36704 5002 36734 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 970 36734 5002 36764 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 940 36764 5002 36794 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 910 36794 5002 36824 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 880 36824 5002 36854 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 850 36854 5002 36884 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 820 36884 5002 36914 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 790 36914 5002 36944 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 760 36944 5002 36974 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 730 36974 5002 37004 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 700 37004 5002 37034 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 670 37034 5002 37064 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 640 37064 5002 37072 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal3 s 632 37072 5002 40000 1 SRC_BDY_HVC
port 5 nsew ground bidirectional
rlabel metal5 s 0 1797 15000 2687 1 VCCD
port 17 nsew power bidirectional
rlabel metal5 s 0 427 15000 1477 1 VCCHIB
port 18 nsew power bidirectional
rlabel metal5 s 0 3007 15000 3657 1 VDDA
port 16 nsew power bidirectional
rlabel metal4 s 0 14007 15000 19000 1 VDDIO
port 13 nsew power bidirectional
rlabel metal5 s 0 3977 15000 4867 1 VDDIO
port 13 nsew power bidirectional
rlabel metal5 s 0 14007 15000 18997 1 VDDIO
port 13 nsew power bidirectional
rlabel metal5 s 0 12837 15000 13687 1 VDDIO_Q
port 12 nsew power bidirectional
rlabel metal4 s 0 9547 15000 9613 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 10329 15000 10565 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 7367 15000 8017 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 9547 15000 11347 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 8337 15000 9227 1 VSSD
port 9 nsew ground bidirectional
rlabel metal5 s 0 5187 15000 6077 1 VSSIO
port 15 nsew ground bidirectional
rlabel metal5 s 0 11667 15000 12517 1 VSSIO_Q
port 19 nsew ground bidirectional
rlabel metal5 s 0 6397 15000 7047 1 VSWITCH
port 14 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string GDS_END 24125096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24115484
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
