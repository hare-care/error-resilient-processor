magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< locali >>
rect 400 1777 962 1796
rect 400 1671 412 1777
rect 950 1671 962 1777
rect 400 1659 962 1671
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< viali >>
rect 412 1671 950 1777
rect 412 19 950 125
<< obsli1 >>
rect 190 1633 256 1699
rect 1106 1633 1172 1699
rect 190 1611 230 1633
rect 1132 1611 1172 1633
rect 41 1563 230 1611
rect 41 1529 60 1563
rect 94 1529 230 1563
rect 41 1491 230 1529
rect 41 1457 60 1491
rect 94 1457 230 1491
rect 41 1419 230 1457
rect 41 1385 60 1419
rect 94 1385 230 1419
rect 41 1347 230 1385
rect 41 1313 60 1347
rect 94 1313 230 1347
rect 41 1275 230 1313
rect 41 1241 60 1275
rect 94 1241 230 1275
rect 41 1203 230 1241
rect 41 1169 60 1203
rect 94 1169 230 1203
rect 41 1131 230 1169
rect 41 1097 60 1131
rect 94 1097 230 1131
rect 41 1059 230 1097
rect 41 1025 60 1059
rect 94 1025 230 1059
rect 41 987 230 1025
rect 41 953 60 987
rect 94 953 230 987
rect 41 915 230 953
rect 41 881 60 915
rect 94 881 230 915
rect 41 843 230 881
rect 41 809 60 843
rect 94 809 230 843
rect 41 771 230 809
rect 41 737 60 771
rect 94 737 230 771
rect 41 699 230 737
rect 41 665 60 699
rect 94 665 230 699
rect 41 627 230 665
rect 41 593 60 627
rect 94 593 230 627
rect 41 555 230 593
rect 41 521 60 555
rect 94 521 230 555
rect 41 483 230 521
rect 41 449 60 483
rect 94 449 230 483
rect 41 411 230 449
rect 41 377 60 411
rect 94 377 230 411
rect 41 339 230 377
rect 41 305 60 339
rect 94 305 230 339
rect 41 267 230 305
rect 41 233 60 267
rect 94 233 230 267
rect 41 185 230 233
rect 352 185 386 1611
rect 508 185 542 1611
rect 664 185 698 1611
rect 820 185 854 1611
rect 976 185 1010 1611
rect 1132 1563 1321 1611
rect 1132 1529 1268 1563
rect 1302 1529 1321 1563
rect 1132 1491 1321 1529
rect 1132 1457 1268 1491
rect 1302 1457 1321 1491
rect 1132 1419 1321 1457
rect 1132 1385 1268 1419
rect 1302 1385 1321 1419
rect 1132 1347 1321 1385
rect 1132 1313 1268 1347
rect 1302 1313 1321 1347
rect 1132 1275 1321 1313
rect 1132 1241 1268 1275
rect 1302 1241 1321 1275
rect 1132 1203 1321 1241
rect 1132 1169 1268 1203
rect 1302 1169 1321 1203
rect 1132 1131 1321 1169
rect 1132 1097 1268 1131
rect 1302 1097 1321 1131
rect 1132 1059 1321 1097
rect 1132 1025 1268 1059
rect 1302 1025 1321 1059
rect 1132 987 1321 1025
rect 1132 953 1268 987
rect 1302 953 1321 987
rect 1132 915 1321 953
rect 1132 881 1268 915
rect 1302 881 1321 915
rect 1132 843 1321 881
rect 1132 809 1268 843
rect 1302 809 1321 843
rect 1132 771 1321 809
rect 1132 737 1268 771
rect 1302 737 1321 771
rect 1132 699 1321 737
rect 1132 665 1268 699
rect 1302 665 1321 699
rect 1132 627 1321 665
rect 1132 593 1268 627
rect 1302 593 1321 627
rect 1132 555 1321 593
rect 1132 521 1268 555
rect 1302 521 1321 555
rect 1132 483 1321 521
rect 1132 449 1268 483
rect 1302 449 1321 483
rect 1132 411 1321 449
rect 1132 377 1268 411
rect 1302 377 1321 411
rect 1132 339 1321 377
rect 1132 305 1268 339
rect 1302 305 1321 339
rect 1132 267 1321 305
rect 1132 233 1268 267
rect 1302 233 1321 267
rect 1132 185 1321 233
rect 190 163 230 185
rect 1132 163 1172 185
rect 190 97 256 163
rect 1106 97 1172 163
<< obsli1c >>
rect 60 1529 94 1563
rect 60 1457 94 1491
rect 60 1385 94 1419
rect 60 1313 94 1347
rect 60 1241 94 1275
rect 60 1169 94 1203
rect 60 1097 94 1131
rect 60 1025 94 1059
rect 60 953 94 987
rect 60 881 94 915
rect 60 809 94 843
rect 60 737 94 771
rect 60 665 94 699
rect 60 593 94 627
rect 60 521 94 555
rect 60 449 94 483
rect 60 377 94 411
rect 60 305 94 339
rect 60 233 94 267
rect 1268 1529 1302 1563
rect 1268 1457 1302 1491
rect 1268 1385 1302 1419
rect 1268 1313 1302 1347
rect 1268 1241 1302 1275
rect 1268 1169 1302 1203
rect 1268 1097 1302 1131
rect 1268 1025 1302 1059
rect 1268 953 1302 987
rect 1268 881 1302 915
rect 1268 809 1302 843
rect 1268 737 1302 771
rect 1268 665 1302 699
rect 1268 593 1302 627
rect 1268 521 1302 555
rect 1268 449 1302 483
rect 1268 377 1302 411
rect 1268 305 1302 339
rect 1268 233 1302 267
<< metal1 >>
rect 400 1777 962 1796
rect 400 1671 412 1777
rect 950 1671 962 1777
rect 400 1659 962 1671
rect 41 1563 100 1594
rect 41 1529 60 1563
rect 94 1529 100 1563
rect 41 1491 100 1529
rect 41 1457 60 1491
rect 94 1457 100 1491
rect 41 1419 100 1457
rect 41 1385 60 1419
rect 94 1385 100 1419
rect 41 1347 100 1385
rect 41 1313 60 1347
rect 94 1313 100 1347
rect 41 1275 100 1313
rect 41 1241 60 1275
rect 94 1241 100 1275
rect 41 1203 100 1241
rect 41 1169 60 1203
rect 94 1169 100 1203
rect 41 1131 100 1169
rect 41 1097 60 1131
rect 94 1097 100 1131
rect 41 1059 100 1097
rect 41 1025 60 1059
rect 94 1025 100 1059
rect 41 987 100 1025
rect 41 953 60 987
rect 94 953 100 987
rect 41 915 100 953
rect 41 881 60 915
rect 94 881 100 915
rect 41 843 100 881
rect 41 809 60 843
rect 94 809 100 843
rect 41 771 100 809
rect 41 737 60 771
rect 94 737 100 771
rect 41 699 100 737
rect 41 665 60 699
rect 94 665 100 699
rect 41 627 100 665
rect 41 593 60 627
rect 94 593 100 627
rect 41 555 100 593
rect 41 521 60 555
rect 94 521 100 555
rect 41 483 100 521
rect 41 449 60 483
rect 94 449 100 483
rect 41 411 100 449
rect 41 377 60 411
rect 94 377 100 411
rect 41 339 100 377
rect 41 305 60 339
rect 94 305 100 339
rect 41 267 100 305
rect 41 233 60 267
rect 94 233 100 267
rect 41 202 100 233
rect 1262 1563 1321 1594
rect 1262 1529 1268 1563
rect 1302 1529 1321 1563
rect 1262 1491 1321 1529
rect 1262 1457 1268 1491
rect 1302 1457 1321 1491
rect 1262 1419 1321 1457
rect 1262 1385 1268 1419
rect 1302 1385 1321 1419
rect 1262 1347 1321 1385
rect 1262 1313 1268 1347
rect 1302 1313 1321 1347
rect 1262 1275 1321 1313
rect 1262 1241 1268 1275
rect 1302 1241 1321 1275
rect 1262 1203 1321 1241
rect 1262 1169 1268 1203
rect 1302 1169 1321 1203
rect 1262 1131 1321 1169
rect 1262 1097 1268 1131
rect 1302 1097 1321 1131
rect 1262 1059 1321 1097
rect 1262 1025 1268 1059
rect 1302 1025 1321 1059
rect 1262 987 1321 1025
rect 1262 953 1268 987
rect 1302 953 1321 987
rect 1262 915 1321 953
rect 1262 881 1268 915
rect 1302 881 1321 915
rect 1262 843 1321 881
rect 1262 809 1268 843
rect 1302 809 1321 843
rect 1262 771 1321 809
rect 1262 737 1268 771
rect 1302 737 1321 771
rect 1262 699 1321 737
rect 1262 665 1268 699
rect 1302 665 1321 699
rect 1262 627 1321 665
rect 1262 593 1268 627
rect 1302 593 1321 627
rect 1262 555 1321 593
rect 1262 521 1268 555
rect 1302 521 1321 555
rect 1262 483 1321 521
rect 1262 449 1268 483
rect 1302 449 1321 483
rect 1262 411 1321 449
rect 1262 377 1268 411
rect 1302 377 1321 411
rect 1262 339 1321 377
rect 1262 305 1268 339
rect 1302 305 1321 339
rect 1262 267 1321 305
rect 1262 233 1268 267
rect 1302 233 1321 267
rect 1262 202 1321 233
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< obsm1 >>
rect 343 202 395 1594
rect 499 202 551 1594
rect 655 202 707 1594
rect 811 202 863 1594
rect 967 202 1019 1594
<< metal2 >>
rect 14 1274 1348 1594
rect 14 578 1348 1218
rect 14 202 1348 522
<< labels >>
rlabel metal2 s 14 578 1348 1218 6 DRAIN
port 1 nsew
rlabel viali s 412 1671 950 1777 6 GATE
port 2 nsew
rlabel viali s 412 19 950 125 6 GATE
port 2 nsew
rlabel locali s 400 1659 962 1796 6 GATE
port 2 nsew
rlabel locali s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal1 s 400 1659 962 1796 6 GATE
port 2 nsew
rlabel metal1 s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal2 s 14 1274 1348 1594 6 SOURCE
port 3 nsew
rlabel metal2 s 14 202 1348 522 6 SOURCE
port 3 nsew
rlabel metal1 s 41 202 100 1594 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1262 202 1321 1594 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1348 1796
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8523062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8484878
string device primitive
<< end >>
