magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 78 2718 2336 3529
rect 78 2318 412 2718
rect 715 1816 1956 2310
<< pwell >>
rect 137 -43 2179 309
rect 475 -457 2179 -43
<< nmos >>
rect 554 -317 604 283
rect 660 -317 710 283
rect 876 -317 926 283
rect 982 -317 1032 283
rect 1088 -317 1138 283
rect 1194 -317 1244 283
rect 1410 -317 1460 283
rect 1516 -317 1566 283
rect 1732 -317 1782 283
rect 1838 -317 1888 283
rect 1944 -317 1994 283
rect 2050 -317 2100 283
<< pmos >>
rect 167 2354 217 3354
rect 273 2354 323 3354
rect 489 2754 539 3354
rect 595 2754 645 3354
rect 701 2754 751 3354
rect 807 2754 857 3354
rect 1023 2754 1073 3354
rect 1129 2754 1179 3354
rect 1235 2754 1285 3354
rect 1341 2754 1391 3354
rect 1557 2754 1607 3354
rect 1663 2754 1713 3354
rect 1769 2754 1819 3354
rect 1875 2754 1925 3354
rect 2091 2754 2141 3354
rect 2197 2754 2247 3354
<< mvnmos >>
rect 216 -17 316 283
<< mvpmos >>
rect 781 2091 1781 2191
rect 781 1935 1781 2035
<< ndiff >>
rect 501 205 554 283
rect 501 171 509 205
rect 543 171 554 205
rect 501 137 554 171
rect 501 103 509 137
rect 543 103 554 137
rect 501 69 554 103
rect 501 35 509 69
rect 543 35 554 69
rect 501 1 554 35
rect 501 -33 509 1
rect 543 -33 554 1
rect 501 -67 554 -33
rect 501 -101 509 -67
rect 543 -101 554 -67
rect 501 -135 554 -101
rect 501 -169 509 -135
rect 543 -169 554 -135
rect 501 -203 554 -169
rect 501 -237 509 -203
rect 543 -237 554 -203
rect 501 -271 554 -237
rect 501 -305 509 -271
rect 543 -305 554 -271
rect 501 -317 554 -305
rect 604 205 660 283
rect 604 171 615 205
rect 649 171 660 205
rect 604 137 660 171
rect 604 103 615 137
rect 649 103 660 137
rect 604 69 660 103
rect 604 35 615 69
rect 649 35 660 69
rect 604 1 660 35
rect 604 -33 615 1
rect 649 -33 660 1
rect 604 -67 660 -33
rect 604 -101 615 -67
rect 649 -101 660 -67
rect 604 -135 660 -101
rect 604 -169 615 -135
rect 649 -169 660 -135
rect 604 -203 660 -169
rect 604 -237 615 -203
rect 649 -237 660 -203
rect 604 -271 660 -237
rect 604 -305 615 -271
rect 649 -305 660 -271
rect 604 -317 660 -305
rect 710 205 763 283
rect 710 171 721 205
rect 755 171 763 205
rect 710 137 763 171
rect 710 103 721 137
rect 755 103 763 137
rect 710 69 763 103
rect 710 35 721 69
rect 755 35 763 69
rect 710 1 763 35
rect 710 -33 721 1
rect 755 -33 763 1
rect 710 -67 763 -33
rect 710 -101 721 -67
rect 755 -101 763 -67
rect 710 -135 763 -101
rect 710 -169 721 -135
rect 755 -169 763 -135
rect 710 -203 763 -169
rect 710 -237 721 -203
rect 755 -237 763 -203
rect 710 -271 763 -237
rect 710 -305 721 -271
rect 755 -305 763 -271
rect 710 -317 763 -305
rect 823 205 876 283
rect 823 171 831 205
rect 865 171 876 205
rect 823 137 876 171
rect 823 103 831 137
rect 865 103 876 137
rect 823 69 876 103
rect 823 35 831 69
rect 865 35 876 69
rect 823 1 876 35
rect 823 -33 831 1
rect 865 -33 876 1
rect 823 -67 876 -33
rect 823 -101 831 -67
rect 865 -101 876 -67
rect 823 -135 876 -101
rect 823 -169 831 -135
rect 865 -169 876 -135
rect 823 -203 876 -169
rect 823 -237 831 -203
rect 865 -237 876 -203
rect 823 -271 876 -237
rect 823 -305 831 -271
rect 865 -305 876 -271
rect 823 -317 876 -305
rect 926 205 982 283
rect 926 171 937 205
rect 971 171 982 205
rect 926 137 982 171
rect 926 103 937 137
rect 971 103 982 137
rect 926 69 982 103
rect 926 35 937 69
rect 971 35 982 69
rect 926 1 982 35
rect 926 -33 937 1
rect 971 -33 982 1
rect 926 -67 982 -33
rect 926 -101 937 -67
rect 971 -101 982 -67
rect 926 -135 982 -101
rect 926 -169 937 -135
rect 971 -169 982 -135
rect 926 -203 982 -169
rect 926 -237 937 -203
rect 971 -237 982 -203
rect 926 -271 982 -237
rect 926 -305 937 -271
rect 971 -305 982 -271
rect 926 -317 982 -305
rect 1032 205 1088 283
rect 1032 171 1043 205
rect 1077 171 1088 205
rect 1032 137 1088 171
rect 1032 103 1043 137
rect 1077 103 1088 137
rect 1032 69 1088 103
rect 1032 35 1043 69
rect 1077 35 1088 69
rect 1032 1 1088 35
rect 1032 -33 1043 1
rect 1077 -33 1088 1
rect 1032 -67 1088 -33
rect 1032 -101 1043 -67
rect 1077 -101 1088 -67
rect 1032 -135 1088 -101
rect 1032 -169 1043 -135
rect 1077 -169 1088 -135
rect 1032 -203 1088 -169
rect 1032 -237 1043 -203
rect 1077 -237 1088 -203
rect 1032 -271 1088 -237
rect 1032 -305 1043 -271
rect 1077 -305 1088 -271
rect 1032 -317 1088 -305
rect 1138 205 1194 283
rect 1138 171 1149 205
rect 1183 171 1194 205
rect 1138 137 1194 171
rect 1138 103 1149 137
rect 1183 103 1194 137
rect 1138 69 1194 103
rect 1138 35 1149 69
rect 1183 35 1194 69
rect 1138 1 1194 35
rect 1138 -33 1149 1
rect 1183 -33 1194 1
rect 1138 -67 1194 -33
rect 1138 -101 1149 -67
rect 1183 -101 1194 -67
rect 1138 -135 1194 -101
rect 1138 -169 1149 -135
rect 1183 -169 1194 -135
rect 1138 -203 1194 -169
rect 1138 -237 1149 -203
rect 1183 -237 1194 -203
rect 1138 -271 1194 -237
rect 1138 -305 1149 -271
rect 1183 -305 1194 -271
rect 1138 -317 1194 -305
rect 1244 205 1297 283
rect 1244 171 1255 205
rect 1289 171 1297 205
rect 1244 137 1297 171
rect 1244 103 1255 137
rect 1289 103 1297 137
rect 1244 69 1297 103
rect 1244 35 1255 69
rect 1289 35 1297 69
rect 1244 1 1297 35
rect 1244 -33 1255 1
rect 1289 -33 1297 1
rect 1244 -67 1297 -33
rect 1244 -101 1255 -67
rect 1289 -101 1297 -67
rect 1244 -135 1297 -101
rect 1244 -169 1255 -135
rect 1289 -169 1297 -135
rect 1244 -203 1297 -169
rect 1244 -237 1255 -203
rect 1289 -237 1297 -203
rect 1244 -271 1297 -237
rect 1244 -305 1255 -271
rect 1289 -305 1297 -271
rect 1244 -317 1297 -305
rect 1357 205 1410 283
rect 1357 171 1365 205
rect 1399 171 1410 205
rect 1357 137 1410 171
rect 1357 103 1365 137
rect 1399 103 1410 137
rect 1357 69 1410 103
rect 1357 35 1365 69
rect 1399 35 1410 69
rect 1357 1 1410 35
rect 1357 -33 1365 1
rect 1399 -33 1410 1
rect 1357 -67 1410 -33
rect 1357 -101 1365 -67
rect 1399 -101 1410 -67
rect 1357 -135 1410 -101
rect 1357 -169 1365 -135
rect 1399 -169 1410 -135
rect 1357 -203 1410 -169
rect 1357 -237 1365 -203
rect 1399 -237 1410 -203
rect 1357 -271 1410 -237
rect 1357 -305 1365 -271
rect 1399 -305 1410 -271
rect 1357 -317 1410 -305
rect 1460 205 1516 283
rect 1460 171 1471 205
rect 1505 171 1516 205
rect 1460 137 1516 171
rect 1460 103 1471 137
rect 1505 103 1516 137
rect 1460 69 1516 103
rect 1460 35 1471 69
rect 1505 35 1516 69
rect 1460 1 1516 35
rect 1460 -33 1471 1
rect 1505 -33 1516 1
rect 1460 -67 1516 -33
rect 1460 -101 1471 -67
rect 1505 -101 1516 -67
rect 1460 -135 1516 -101
rect 1460 -169 1471 -135
rect 1505 -169 1516 -135
rect 1460 -203 1516 -169
rect 1460 -237 1471 -203
rect 1505 -237 1516 -203
rect 1460 -271 1516 -237
rect 1460 -305 1471 -271
rect 1505 -305 1516 -271
rect 1460 -317 1516 -305
rect 1566 205 1619 283
rect 1566 171 1577 205
rect 1611 171 1619 205
rect 1566 137 1619 171
rect 1566 103 1577 137
rect 1611 103 1619 137
rect 1566 69 1619 103
rect 1566 35 1577 69
rect 1611 35 1619 69
rect 1566 1 1619 35
rect 1566 -33 1577 1
rect 1611 -33 1619 1
rect 1566 -67 1619 -33
rect 1566 -101 1577 -67
rect 1611 -101 1619 -67
rect 1566 -135 1619 -101
rect 1566 -169 1577 -135
rect 1611 -169 1619 -135
rect 1566 -203 1619 -169
rect 1566 -237 1577 -203
rect 1611 -237 1619 -203
rect 1566 -271 1619 -237
rect 1566 -305 1577 -271
rect 1611 -305 1619 -271
rect 1566 -317 1619 -305
rect 1679 205 1732 283
rect 1679 171 1687 205
rect 1721 171 1732 205
rect 1679 137 1732 171
rect 1679 103 1687 137
rect 1721 103 1732 137
rect 1679 69 1732 103
rect 1679 35 1687 69
rect 1721 35 1732 69
rect 1679 1 1732 35
rect 1679 -33 1687 1
rect 1721 -33 1732 1
rect 1679 -67 1732 -33
rect 1679 -101 1687 -67
rect 1721 -101 1732 -67
rect 1679 -135 1732 -101
rect 1679 -169 1687 -135
rect 1721 -169 1732 -135
rect 1679 -203 1732 -169
rect 1679 -237 1687 -203
rect 1721 -237 1732 -203
rect 1679 -271 1732 -237
rect 1679 -305 1687 -271
rect 1721 -305 1732 -271
rect 1679 -317 1732 -305
rect 1782 205 1838 283
rect 1782 171 1793 205
rect 1827 171 1838 205
rect 1782 137 1838 171
rect 1782 103 1793 137
rect 1827 103 1838 137
rect 1782 69 1838 103
rect 1782 35 1793 69
rect 1827 35 1838 69
rect 1782 1 1838 35
rect 1782 -33 1793 1
rect 1827 -33 1838 1
rect 1782 -67 1838 -33
rect 1782 -101 1793 -67
rect 1827 -101 1838 -67
rect 1782 -135 1838 -101
rect 1782 -169 1793 -135
rect 1827 -169 1838 -135
rect 1782 -203 1838 -169
rect 1782 -237 1793 -203
rect 1827 -237 1838 -203
rect 1782 -271 1838 -237
rect 1782 -305 1793 -271
rect 1827 -305 1838 -271
rect 1782 -317 1838 -305
rect 1888 205 1944 283
rect 1888 171 1899 205
rect 1933 171 1944 205
rect 1888 137 1944 171
rect 1888 103 1899 137
rect 1933 103 1944 137
rect 1888 69 1944 103
rect 1888 35 1899 69
rect 1933 35 1944 69
rect 1888 1 1944 35
rect 1888 -33 1899 1
rect 1933 -33 1944 1
rect 1888 -67 1944 -33
rect 1888 -101 1899 -67
rect 1933 -101 1944 -67
rect 1888 -135 1944 -101
rect 1888 -169 1899 -135
rect 1933 -169 1944 -135
rect 1888 -203 1944 -169
rect 1888 -237 1899 -203
rect 1933 -237 1944 -203
rect 1888 -271 1944 -237
rect 1888 -305 1899 -271
rect 1933 -305 1944 -271
rect 1888 -317 1944 -305
rect 1994 205 2050 283
rect 1994 171 2005 205
rect 2039 171 2050 205
rect 1994 137 2050 171
rect 1994 103 2005 137
rect 2039 103 2050 137
rect 1994 69 2050 103
rect 1994 35 2005 69
rect 2039 35 2050 69
rect 1994 1 2050 35
rect 1994 -33 2005 1
rect 2039 -33 2050 1
rect 1994 -67 2050 -33
rect 1994 -101 2005 -67
rect 2039 -101 2050 -67
rect 1994 -135 2050 -101
rect 1994 -169 2005 -135
rect 2039 -169 2050 -135
rect 1994 -203 2050 -169
rect 1994 -237 2005 -203
rect 2039 -237 2050 -203
rect 1994 -271 2050 -237
rect 1994 -305 2005 -271
rect 2039 -305 2050 -271
rect 1994 -317 2050 -305
rect 2100 205 2153 283
rect 2100 171 2111 205
rect 2145 171 2153 205
rect 2100 137 2153 171
rect 2100 103 2111 137
rect 2145 103 2153 137
rect 2100 69 2153 103
rect 2100 35 2111 69
rect 2145 35 2153 69
rect 2100 1 2153 35
rect 2100 -33 2111 1
rect 2145 -33 2153 1
rect 2100 -67 2153 -33
rect 2100 -101 2111 -67
rect 2145 -101 2153 -67
rect 2100 -135 2153 -101
rect 2100 -169 2111 -135
rect 2145 -169 2153 -135
rect 2100 -203 2153 -169
rect 2100 -237 2111 -203
rect 2145 -237 2153 -203
rect 2100 -271 2153 -237
rect 2100 -305 2111 -271
rect 2145 -305 2153 -271
rect 2100 -317 2153 -305
<< pdiff >>
rect 114 3342 167 3354
rect 114 3308 122 3342
rect 156 3308 167 3342
rect 114 3274 167 3308
rect 114 3240 122 3274
rect 156 3240 167 3274
rect 114 3206 167 3240
rect 114 3172 122 3206
rect 156 3172 167 3206
rect 114 3138 167 3172
rect 114 3104 122 3138
rect 156 3104 167 3138
rect 114 3070 167 3104
rect 114 3036 122 3070
rect 156 3036 167 3070
rect 114 3002 167 3036
rect 114 2968 122 3002
rect 156 2968 167 3002
rect 114 2934 167 2968
rect 114 2900 122 2934
rect 156 2900 167 2934
rect 114 2866 167 2900
rect 114 2832 122 2866
rect 156 2832 167 2866
rect 114 2798 167 2832
rect 114 2764 122 2798
rect 156 2764 167 2798
rect 114 2730 167 2764
rect 114 2696 122 2730
rect 156 2696 167 2730
rect 114 2662 167 2696
rect 114 2628 122 2662
rect 156 2628 167 2662
rect 114 2594 167 2628
rect 114 2560 122 2594
rect 156 2560 167 2594
rect 114 2526 167 2560
rect 114 2492 122 2526
rect 156 2492 167 2526
rect 114 2458 167 2492
rect 114 2424 122 2458
rect 156 2424 167 2458
rect 114 2354 167 2424
rect 217 3342 273 3354
rect 217 3308 228 3342
rect 262 3308 273 3342
rect 217 3274 273 3308
rect 217 3240 228 3274
rect 262 3240 273 3274
rect 217 3206 273 3240
rect 217 3172 228 3206
rect 262 3172 273 3206
rect 217 3138 273 3172
rect 217 3104 228 3138
rect 262 3104 273 3138
rect 217 3070 273 3104
rect 217 3036 228 3070
rect 262 3036 273 3070
rect 217 3002 273 3036
rect 217 2968 228 3002
rect 262 2968 273 3002
rect 217 2934 273 2968
rect 217 2900 228 2934
rect 262 2900 273 2934
rect 217 2866 273 2900
rect 217 2832 228 2866
rect 262 2832 273 2866
rect 217 2798 273 2832
rect 217 2764 228 2798
rect 262 2764 273 2798
rect 217 2730 273 2764
rect 217 2696 228 2730
rect 262 2696 273 2730
rect 217 2662 273 2696
rect 217 2628 228 2662
rect 262 2628 273 2662
rect 217 2594 273 2628
rect 217 2560 228 2594
rect 262 2560 273 2594
rect 217 2526 273 2560
rect 217 2492 228 2526
rect 262 2492 273 2526
rect 217 2458 273 2492
rect 217 2424 228 2458
rect 262 2424 273 2458
rect 217 2354 273 2424
rect 323 3342 376 3354
rect 323 3308 334 3342
rect 368 3308 376 3342
rect 323 3274 376 3308
rect 323 3240 334 3274
rect 368 3240 376 3274
rect 323 3206 376 3240
rect 323 3172 334 3206
rect 368 3172 376 3206
rect 323 3138 376 3172
rect 323 3104 334 3138
rect 368 3104 376 3138
rect 323 3070 376 3104
rect 323 3036 334 3070
rect 368 3036 376 3070
rect 323 3002 376 3036
rect 323 2968 334 3002
rect 368 2968 376 3002
rect 323 2934 376 2968
rect 323 2900 334 2934
rect 368 2900 376 2934
rect 323 2866 376 2900
rect 323 2832 334 2866
rect 368 2832 376 2866
rect 323 2798 376 2832
rect 323 2764 334 2798
rect 368 2764 376 2798
rect 323 2730 376 2764
rect 436 3276 489 3354
rect 436 3242 444 3276
rect 478 3242 489 3276
rect 436 3208 489 3242
rect 436 3174 444 3208
rect 478 3174 489 3208
rect 436 3140 489 3174
rect 436 3106 444 3140
rect 478 3106 489 3140
rect 436 3072 489 3106
rect 436 3038 444 3072
rect 478 3038 489 3072
rect 436 3004 489 3038
rect 436 2970 444 3004
rect 478 2970 489 3004
rect 436 2936 489 2970
rect 436 2902 444 2936
rect 478 2902 489 2936
rect 436 2868 489 2902
rect 436 2834 444 2868
rect 478 2834 489 2868
rect 436 2800 489 2834
rect 436 2766 444 2800
rect 478 2766 489 2800
rect 436 2754 489 2766
rect 539 3276 595 3354
rect 539 3242 550 3276
rect 584 3242 595 3276
rect 539 3208 595 3242
rect 539 3174 550 3208
rect 584 3174 595 3208
rect 539 3140 595 3174
rect 539 3106 550 3140
rect 584 3106 595 3140
rect 539 3072 595 3106
rect 539 3038 550 3072
rect 584 3038 595 3072
rect 539 3004 595 3038
rect 539 2970 550 3004
rect 584 2970 595 3004
rect 539 2936 595 2970
rect 539 2902 550 2936
rect 584 2902 595 2936
rect 539 2868 595 2902
rect 539 2834 550 2868
rect 584 2834 595 2868
rect 539 2800 595 2834
rect 539 2766 550 2800
rect 584 2766 595 2800
rect 539 2754 595 2766
rect 645 3276 701 3354
rect 645 3242 656 3276
rect 690 3242 701 3276
rect 645 3208 701 3242
rect 645 3174 656 3208
rect 690 3174 701 3208
rect 645 3140 701 3174
rect 645 3106 656 3140
rect 690 3106 701 3140
rect 645 3072 701 3106
rect 645 3038 656 3072
rect 690 3038 701 3072
rect 645 3004 701 3038
rect 645 2970 656 3004
rect 690 2970 701 3004
rect 645 2936 701 2970
rect 645 2902 656 2936
rect 690 2902 701 2936
rect 645 2868 701 2902
rect 645 2834 656 2868
rect 690 2834 701 2868
rect 645 2800 701 2834
rect 645 2766 656 2800
rect 690 2766 701 2800
rect 645 2754 701 2766
rect 751 3276 807 3354
rect 751 3242 762 3276
rect 796 3242 807 3276
rect 751 3208 807 3242
rect 751 3174 762 3208
rect 796 3174 807 3208
rect 751 3140 807 3174
rect 751 3106 762 3140
rect 796 3106 807 3140
rect 751 3072 807 3106
rect 751 3038 762 3072
rect 796 3038 807 3072
rect 751 3004 807 3038
rect 751 2970 762 3004
rect 796 2970 807 3004
rect 751 2936 807 2970
rect 751 2902 762 2936
rect 796 2902 807 2936
rect 751 2868 807 2902
rect 751 2834 762 2868
rect 796 2834 807 2868
rect 751 2800 807 2834
rect 751 2766 762 2800
rect 796 2766 807 2800
rect 751 2754 807 2766
rect 857 3276 910 3354
rect 857 3242 868 3276
rect 902 3242 910 3276
rect 857 3208 910 3242
rect 857 3174 868 3208
rect 902 3174 910 3208
rect 857 3140 910 3174
rect 857 3106 868 3140
rect 902 3106 910 3140
rect 857 3072 910 3106
rect 857 3038 868 3072
rect 902 3038 910 3072
rect 857 3004 910 3038
rect 857 2970 868 3004
rect 902 2970 910 3004
rect 857 2936 910 2970
rect 857 2902 868 2936
rect 902 2902 910 2936
rect 857 2868 910 2902
rect 857 2834 868 2868
rect 902 2834 910 2868
rect 857 2800 910 2834
rect 857 2766 868 2800
rect 902 2766 910 2800
rect 857 2754 910 2766
rect 970 3276 1023 3354
rect 970 3242 978 3276
rect 1012 3242 1023 3276
rect 970 3208 1023 3242
rect 970 3174 978 3208
rect 1012 3174 1023 3208
rect 970 3140 1023 3174
rect 970 3106 978 3140
rect 1012 3106 1023 3140
rect 970 3072 1023 3106
rect 970 3038 978 3072
rect 1012 3038 1023 3072
rect 970 3004 1023 3038
rect 970 2970 978 3004
rect 1012 2970 1023 3004
rect 970 2936 1023 2970
rect 970 2902 978 2936
rect 1012 2902 1023 2936
rect 970 2868 1023 2902
rect 970 2834 978 2868
rect 1012 2834 1023 2868
rect 970 2800 1023 2834
rect 970 2766 978 2800
rect 1012 2766 1023 2800
rect 970 2754 1023 2766
rect 1073 3276 1129 3354
rect 1073 3242 1084 3276
rect 1118 3242 1129 3276
rect 1073 3208 1129 3242
rect 1073 3174 1084 3208
rect 1118 3174 1129 3208
rect 1073 3140 1129 3174
rect 1073 3106 1084 3140
rect 1118 3106 1129 3140
rect 1073 3072 1129 3106
rect 1073 3038 1084 3072
rect 1118 3038 1129 3072
rect 1073 3004 1129 3038
rect 1073 2970 1084 3004
rect 1118 2970 1129 3004
rect 1073 2936 1129 2970
rect 1073 2902 1084 2936
rect 1118 2902 1129 2936
rect 1073 2868 1129 2902
rect 1073 2834 1084 2868
rect 1118 2834 1129 2868
rect 1073 2800 1129 2834
rect 1073 2766 1084 2800
rect 1118 2766 1129 2800
rect 1073 2754 1129 2766
rect 1179 3276 1235 3354
rect 1179 3242 1190 3276
rect 1224 3242 1235 3276
rect 1179 3208 1235 3242
rect 1179 3174 1190 3208
rect 1224 3174 1235 3208
rect 1179 3140 1235 3174
rect 1179 3106 1190 3140
rect 1224 3106 1235 3140
rect 1179 3072 1235 3106
rect 1179 3038 1190 3072
rect 1224 3038 1235 3072
rect 1179 3004 1235 3038
rect 1179 2970 1190 3004
rect 1224 2970 1235 3004
rect 1179 2936 1235 2970
rect 1179 2902 1190 2936
rect 1224 2902 1235 2936
rect 1179 2868 1235 2902
rect 1179 2834 1190 2868
rect 1224 2834 1235 2868
rect 1179 2800 1235 2834
rect 1179 2766 1190 2800
rect 1224 2766 1235 2800
rect 1179 2754 1235 2766
rect 1285 3276 1341 3354
rect 1285 3242 1296 3276
rect 1330 3242 1341 3276
rect 1285 3208 1341 3242
rect 1285 3174 1296 3208
rect 1330 3174 1341 3208
rect 1285 3140 1341 3174
rect 1285 3106 1296 3140
rect 1330 3106 1341 3140
rect 1285 3072 1341 3106
rect 1285 3038 1296 3072
rect 1330 3038 1341 3072
rect 1285 3004 1341 3038
rect 1285 2970 1296 3004
rect 1330 2970 1341 3004
rect 1285 2936 1341 2970
rect 1285 2902 1296 2936
rect 1330 2902 1341 2936
rect 1285 2868 1341 2902
rect 1285 2834 1296 2868
rect 1330 2834 1341 2868
rect 1285 2800 1341 2834
rect 1285 2766 1296 2800
rect 1330 2766 1341 2800
rect 1285 2754 1341 2766
rect 1391 3276 1444 3354
rect 1391 3242 1402 3276
rect 1436 3242 1444 3276
rect 1391 3208 1444 3242
rect 1391 3174 1402 3208
rect 1436 3174 1444 3208
rect 1391 3140 1444 3174
rect 1391 3106 1402 3140
rect 1436 3106 1444 3140
rect 1391 3072 1444 3106
rect 1391 3038 1402 3072
rect 1436 3038 1444 3072
rect 1391 3004 1444 3038
rect 1391 2970 1402 3004
rect 1436 2970 1444 3004
rect 1391 2936 1444 2970
rect 1391 2902 1402 2936
rect 1436 2902 1444 2936
rect 1391 2868 1444 2902
rect 1391 2834 1402 2868
rect 1436 2834 1444 2868
rect 1391 2800 1444 2834
rect 1391 2766 1402 2800
rect 1436 2766 1444 2800
rect 1391 2754 1444 2766
rect 1504 3276 1557 3354
rect 1504 3242 1512 3276
rect 1546 3242 1557 3276
rect 1504 3208 1557 3242
rect 1504 3174 1512 3208
rect 1546 3174 1557 3208
rect 1504 3140 1557 3174
rect 1504 3106 1512 3140
rect 1546 3106 1557 3140
rect 1504 3072 1557 3106
rect 1504 3038 1512 3072
rect 1546 3038 1557 3072
rect 1504 3004 1557 3038
rect 1504 2970 1512 3004
rect 1546 2970 1557 3004
rect 1504 2936 1557 2970
rect 1504 2902 1512 2936
rect 1546 2902 1557 2936
rect 1504 2868 1557 2902
rect 1504 2834 1512 2868
rect 1546 2834 1557 2868
rect 1504 2800 1557 2834
rect 1504 2766 1512 2800
rect 1546 2766 1557 2800
rect 1504 2754 1557 2766
rect 1607 3276 1663 3354
rect 1607 3242 1618 3276
rect 1652 3242 1663 3276
rect 1607 3208 1663 3242
rect 1607 3174 1618 3208
rect 1652 3174 1663 3208
rect 1607 3140 1663 3174
rect 1607 3106 1618 3140
rect 1652 3106 1663 3140
rect 1607 3072 1663 3106
rect 1607 3038 1618 3072
rect 1652 3038 1663 3072
rect 1607 3004 1663 3038
rect 1607 2970 1618 3004
rect 1652 2970 1663 3004
rect 1607 2936 1663 2970
rect 1607 2902 1618 2936
rect 1652 2902 1663 2936
rect 1607 2868 1663 2902
rect 1607 2834 1618 2868
rect 1652 2834 1663 2868
rect 1607 2800 1663 2834
rect 1607 2766 1618 2800
rect 1652 2766 1663 2800
rect 1607 2754 1663 2766
rect 1713 3276 1769 3354
rect 1713 3242 1724 3276
rect 1758 3242 1769 3276
rect 1713 3208 1769 3242
rect 1713 3174 1724 3208
rect 1758 3174 1769 3208
rect 1713 3140 1769 3174
rect 1713 3106 1724 3140
rect 1758 3106 1769 3140
rect 1713 3072 1769 3106
rect 1713 3038 1724 3072
rect 1758 3038 1769 3072
rect 1713 3004 1769 3038
rect 1713 2970 1724 3004
rect 1758 2970 1769 3004
rect 1713 2936 1769 2970
rect 1713 2902 1724 2936
rect 1758 2902 1769 2936
rect 1713 2868 1769 2902
rect 1713 2834 1724 2868
rect 1758 2834 1769 2868
rect 1713 2800 1769 2834
rect 1713 2766 1724 2800
rect 1758 2766 1769 2800
rect 1713 2754 1769 2766
rect 1819 3276 1875 3354
rect 1819 3242 1830 3276
rect 1864 3242 1875 3276
rect 1819 3208 1875 3242
rect 1819 3174 1830 3208
rect 1864 3174 1875 3208
rect 1819 3140 1875 3174
rect 1819 3106 1830 3140
rect 1864 3106 1875 3140
rect 1819 3072 1875 3106
rect 1819 3038 1830 3072
rect 1864 3038 1875 3072
rect 1819 3004 1875 3038
rect 1819 2970 1830 3004
rect 1864 2970 1875 3004
rect 1819 2936 1875 2970
rect 1819 2902 1830 2936
rect 1864 2902 1875 2936
rect 1819 2868 1875 2902
rect 1819 2834 1830 2868
rect 1864 2834 1875 2868
rect 1819 2800 1875 2834
rect 1819 2766 1830 2800
rect 1864 2766 1875 2800
rect 1819 2754 1875 2766
rect 1925 3276 1978 3354
rect 1925 3242 1936 3276
rect 1970 3242 1978 3276
rect 1925 3208 1978 3242
rect 1925 3174 1936 3208
rect 1970 3174 1978 3208
rect 1925 3140 1978 3174
rect 1925 3106 1936 3140
rect 1970 3106 1978 3140
rect 1925 3072 1978 3106
rect 1925 3038 1936 3072
rect 1970 3038 1978 3072
rect 1925 3004 1978 3038
rect 1925 2970 1936 3004
rect 1970 2970 1978 3004
rect 1925 2936 1978 2970
rect 1925 2902 1936 2936
rect 1970 2902 1978 2936
rect 1925 2868 1978 2902
rect 1925 2834 1936 2868
rect 1970 2834 1978 2868
rect 1925 2800 1978 2834
rect 1925 2766 1936 2800
rect 1970 2766 1978 2800
rect 1925 2754 1978 2766
rect 2038 3342 2091 3354
rect 2038 3308 2046 3342
rect 2080 3308 2091 3342
rect 2038 3274 2091 3308
rect 2038 3240 2046 3274
rect 2080 3240 2091 3274
rect 2038 3206 2091 3240
rect 2038 3172 2046 3206
rect 2080 3172 2091 3206
rect 2038 3138 2091 3172
rect 2038 3104 2046 3138
rect 2080 3104 2091 3138
rect 2038 3070 2091 3104
rect 2038 3036 2046 3070
rect 2080 3036 2091 3070
rect 2038 3002 2091 3036
rect 2038 2968 2046 3002
rect 2080 2968 2091 3002
rect 2038 2934 2091 2968
rect 2038 2900 2046 2934
rect 2080 2900 2091 2934
rect 2038 2866 2091 2900
rect 2038 2832 2046 2866
rect 2080 2832 2091 2866
rect 2038 2754 2091 2832
rect 2141 3342 2197 3354
rect 2141 3308 2152 3342
rect 2186 3308 2197 3342
rect 2141 3274 2197 3308
rect 2141 3240 2152 3274
rect 2186 3240 2197 3274
rect 2141 3206 2197 3240
rect 2141 3172 2152 3206
rect 2186 3172 2197 3206
rect 2141 3138 2197 3172
rect 2141 3104 2152 3138
rect 2186 3104 2197 3138
rect 2141 3070 2197 3104
rect 2141 3036 2152 3070
rect 2186 3036 2197 3070
rect 2141 3002 2197 3036
rect 2141 2968 2152 3002
rect 2186 2968 2197 3002
rect 2141 2934 2197 2968
rect 2141 2900 2152 2934
rect 2186 2900 2197 2934
rect 2141 2866 2197 2900
rect 2141 2832 2152 2866
rect 2186 2832 2197 2866
rect 2141 2754 2197 2832
rect 2247 3342 2300 3354
rect 2247 3308 2258 3342
rect 2292 3308 2300 3342
rect 2247 3274 2300 3308
rect 2247 3240 2258 3274
rect 2292 3240 2300 3274
rect 2247 3206 2300 3240
rect 2247 3172 2258 3206
rect 2292 3172 2300 3206
rect 2247 3138 2300 3172
rect 2247 3104 2258 3138
rect 2292 3104 2300 3138
rect 2247 3070 2300 3104
rect 2247 3036 2258 3070
rect 2292 3036 2300 3070
rect 2247 3002 2300 3036
rect 2247 2968 2258 3002
rect 2292 2968 2300 3002
rect 2247 2934 2300 2968
rect 2247 2900 2258 2934
rect 2292 2900 2300 2934
rect 2247 2866 2300 2900
rect 2247 2832 2258 2866
rect 2292 2832 2300 2866
rect 2247 2754 2300 2832
rect 323 2696 334 2730
rect 368 2696 376 2730
rect 323 2662 376 2696
rect 323 2628 334 2662
rect 368 2628 376 2662
rect 323 2594 376 2628
rect 323 2560 334 2594
rect 368 2560 376 2594
rect 323 2526 376 2560
rect 323 2492 334 2526
rect 368 2492 376 2526
rect 323 2458 376 2492
rect 323 2424 334 2458
rect 368 2424 376 2458
rect 323 2354 376 2424
<< mvndiff >>
rect 163 233 216 283
rect 163 199 171 233
rect 205 199 216 233
rect 163 165 216 199
rect 163 131 171 165
rect 205 131 216 165
rect 163 97 216 131
rect 163 63 171 97
rect 205 63 216 97
rect 163 29 216 63
rect 163 -5 171 29
rect 205 -5 216 29
rect 163 -17 216 -5
rect 316 233 369 283
rect 316 199 327 233
rect 361 199 369 233
rect 316 165 369 199
rect 316 131 327 165
rect 361 131 369 165
rect 316 97 369 131
rect 316 63 327 97
rect 361 63 369 97
rect 316 29 369 63
rect 316 -5 327 29
rect 361 -5 369 29
rect 316 -17 369 -5
<< mvpdiff >>
rect 781 2236 1781 2244
rect 781 2202 851 2236
rect 885 2202 919 2236
rect 953 2202 987 2236
rect 1021 2202 1055 2236
rect 1089 2202 1123 2236
rect 1157 2202 1191 2236
rect 1225 2202 1259 2236
rect 1293 2202 1327 2236
rect 1361 2202 1395 2236
rect 1429 2202 1463 2236
rect 1497 2202 1531 2236
rect 1565 2202 1599 2236
rect 1633 2202 1667 2236
rect 1701 2202 1735 2236
rect 1769 2202 1781 2236
rect 781 2191 1781 2202
rect 781 2080 1781 2091
rect 781 2046 851 2080
rect 885 2046 919 2080
rect 953 2046 987 2080
rect 1021 2046 1055 2080
rect 1089 2046 1123 2080
rect 1157 2046 1191 2080
rect 1225 2046 1259 2080
rect 1293 2046 1327 2080
rect 1361 2046 1395 2080
rect 1429 2046 1463 2080
rect 1497 2046 1531 2080
rect 1565 2046 1599 2080
rect 1633 2046 1667 2080
rect 1701 2046 1735 2080
rect 1769 2046 1781 2080
rect 781 2035 1781 2046
rect 781 1924 1781 1935
rect 781 1890 851 1924
rect 885 1890 919 1924
rect 953 1890 987 1924
rect 1021 1890 1055 1924
rect 1089 1890 1123 1924
rect 1157 1890 1191 1924
rect 1225 1890 1259 1924
rect 1293 1890 1327 1924
rect 1361 1890 1395 1924
rect 1429 1890 1463 1924
rect 1497 1890 1531 1924
rect 1565 1890 1599 1924
rect 1633 1890 1667 1924
rect 1701 1890 1735 1924
rect 1769 1890 1781 1924
rect 781 1882 1781 1890
<< ndiffc >>
rect 509 171 543 205
rect 509 103 543 137
rect 509 35 543 69
rect 509 -33 543 1
rect 509 -101 543 -67
rect 509 -169 543 -135
rect 509 -237 543 -203
rect 509 -305 543 -271
rect 615 171 649 205
rect 615 103 649 137
rect 615 35 649 69
rect 615 -33 649 1
rect 615 -101 649 -67
rect 615 -169 649 -135
rect 615 -237 649 -203
rect 615 -305 649 -271
rect 721 171 755 205
rect 721 103 755 137
rect 721 35 755 69
rect 721 -33 755 1
rect 721 -101 755 -67
rect 721 -169 755 -135
rect 721 -237 755 -203
rect 721 -305 755 -271
rect 831 171 865 205
rect 831 103 865 137
rect 831 35 865 69
rect 831 -33 865 1
rect 831 -101 865 -67
rect 831 -169 865 -135
rect 831 -237 865 -203
rect 831 -305 865 -271
rect 937 171 971 205
rect 937 103 971 137
rect 937 35 971 69
rect 937 -33 971 1
rect 937 -101 971 -67
rect 937 -169 971 -135
rect 937 -237 971 -203
rect 937 -305 971 -271
rect 1043 171 1077 205
rect 1043 103 1077 137
rect 1043 35 1077 69
rect 1043 -33 1077 1
rect 1043 -101 1077 -67
rect 1043 -169 1077 -135
rect 1043 -237 1077 -203
rect 1043 -305 1077 -271
rect 1149 171 1183 205
rect 1149 103 1183 137
rect 1149 35 1183 69
rect 1149 -33 1183 1
rect 1149 -101 1183 -67
rect 1149 -169 1183 -135
rect 1149 -237 1183 -203
rect 1149 -305 1183 -271
rect 1255 171 1289 205
rect 1255 103 1289 137
rect 1255 35 1289 69
rect 1255 -33 1289 1
rect 1255 -101 1289 -67
rect 1255 -169 1289 -135
rect 1255 -237 1289 -203
rect 1255 -305 1289 -271
rect 1365 171 1399 205
rect 1365 103 1399 137
rect 1365 35 1399 69
rect 1365 -33 1399 1
rect 1365 -101 1399 -67
rect 1365 -169 1399 -135
rect 1365 -237 1399 -203
rect 1365 -305 1399 -271
rect 1471 171 1505 205
rect 1471 103 1505 137
rect 1471 35 1505 69
rect 1471 -33 1505 1
rect 1471 -101 1505 -67
rect 1471 -169 1505 -135
rect 1471 -237 1505 -203
rect 1471 -305 1505 -271
rect 1577 171 1611 205
rect 1577 103 1611 137
rect 1577 35 1611 69
rect 1577 -33 1611 1
rect 1577 -101 1611 -67
rect 1577 -169 1611 -135
rect 1577 -237 1611 -203
rect 1577 -305 1611 -271
rect 1687 171 1721 205
rect 1687 103 1721 137
rect 1687 35 1721 69
rect 1687 -33 1721 1
rect 1687 -101 1721 -67
rect 1687 -169 1721 -135
rect 1687 -237 1721 -203
rect 1687 -305 1721 -271
rect 1793 171 1827 205
rect 1793 103 1827 137
rect 1793 35 1827 69
rect 1793 -33 1827 1
rect 1793 -101 1827 -67
rect 1793 -169 1827 -135
rect 1793 -237 1827 -203
rect 1793 -305 1827 -271
rect 1899 171 1933 205
rect 1899 103 1933 137
rect 1899 35 1933 69
rect 1899 -33 1933 1
rect 1899 -101 1933 -67
rect 1899 -169 1933 -135
rect 1899 -237 1933 -203
rect 1899 -305 1933 -271
rect 2005 171 2039 205
rect 2005 103 2039 137
rect 2005 35 2039 69
rect 2005 -33 2039 1
rect 2005 -101 2039 -67
rect 2005 -169 2039 -135
rect 2005 -237 2039 -203
rect 2005 -305 2039 -271
rect 2111 171 2145 205
rect 2111 103 2145 137
rect 2111 35 2145 69
rect 2111 -33 2145 1
rect 2111 -101 2145 -67
rect 2111 -169 2145 -135
rect 2111 -237 2145 -203
rect 2111 -305 2145 -271
<< pdiffc >>
rect 122 3308 156 3342
rect 122 3240 156 3274
rect 122 3172 156 3206
rect 122 3104 156 3138
rect 122 3036 156 3070
rect 122 2968 156 3002
rect 122 2900 156 2934
rect 122 2832 156 2866
rect 122 2764 156 2798
rect 122 2696 156 2730
rect 122 2628 156 2662
rect 122 2560 156 2594
rect 122 2492 156 2526
rect 122 2424 156 2458
rect 228 3308 262 3342
rect 228 3240 262 3274
rect 228 3172 262 3206
rect 228 3104 262 3138
rect 228 3036 262 3070
rect 228 2968 262 3002
rect 228 2900 262 2934
rect 228 2832 262 2866
rect 228 2764 262 2798
rect 228 2696 262 2730
rect 228 2628 262 2662
rect 228 2560 262 2594
rect 228 2492 262 2526
rect 228 2424 262 2458
rect 334 3308 368 3342
rect 334 3240 368 3274
rect 334 3172 368 3206
rect 334 3104 368 3138
rect 334 3036 368 3070
rect 334 2968 368 3002
rect 334 2900 368 2934
rect 334 2832 368 2866
rect 334 2764 368 2798
rect 444 3242 478 3276
rect 444 3174 478 3208
rect 444 3106 478 3140
rect 444 3038 478 3072
rect 444 2970 478 3004
rect 444 2902 478 2936
rect 444 2834 478 2868
rect 444 2766 478 2800
rect 550 3242 584 3276
rect 550 3174 584 3208
rect 550 3106 584 3140
rect 550 3038 584 3072
rect 550 2970 584 3004
rect 550 2902 584 2936
rect 550 2834 584 2868
rect 550 2766 584 2800
rect 656 3242 690 3276
rect 656 3174 690 3208
rect 656 3106 690 3140
rect 656 3038 690 3072
rect 656 2970 690 3004
rect 656 2902 690 2936
rect 656 2834 690 2868
rect 656 2766 690 2800
rect 762 3242 796 3276
rect 762 3174 796 3208
rect 762 3106 796 3140
rect 762 3038 796 3072
rect 762 2970 796 3004
rect 762 2902 796 2936
rect 762 2834 796 2868
rect 762 2766 796 2800
rect 868 3242 902 3276
rect 868 3174 902 3208
rect 868 3106 902 3140
rect 868 3038 902 3072
rect 868 2970 902 3004
rect 868 2902 902 2936
rect 868 2834 902 2868
rect 868 2766 902 2800
rect 978 3242 1012 3276
rect 978 3174 1012 3208
rect 978 3106 1012 3140
rect 978 3038 1012 3072
rect 978 2970 1012 3004
rect 978 2902 1012 2936
rect 978 2834 1012 2868
rect 978 2766 1012 2800
rect 1084 3242 1118 3276
rect 1084 3174 1118 3208
rect 1084 3106 1118 3140
rect 1084 3038 1118 3072
rect 1084 2970 1118 3004
rect 1084 2902 1118 2936
rect 1084 2834 1118 2868
rect 1084 2766 1118 2800
rect 1190 3242 1224 3276
rect 1190 3174 1224 3208
rect 1190 3106 1224 3140
rect 1190 3038 1224 3072
rect 1190 2970 1224 3004
rect 1190 2902 1224 2936
rect 1190 2834 1224 2868
rect 1190 2766 1224 2800
rect 1296 3242 1330 3276
rect 1296 3174 1330 3208
rect 1296 3106 1330 3140
rect 1296 3038 1330 3072
rect 1296 2970 1330 3004
rect 1296 2902 1330 2936
rect 1296 2834 1330 2868
rect 1296 2766 1330 2800
rect 1402 3242 1436 3276
rect 1402 3174 1436 3208
rect 1402 3106 1436 3140
rect 1402 3038 1436 3072
rect 1402 2970 1436 3004
rect 1402 2902 1436 2936
rect 1402 2834 1436 2868
rect 1402 2766 1436 2800
rect 1512 3242 1546 3276
rect 1512 3174 1546 3208
rect 1512 3106 1546 3140
rect 1512 3038 1546 3072
rect 1512 2970 1546 3004
rect 1512 2902 1546 2936
rect 1512 2834 1546 2868
rect 1512 2766 1546 2800
rect 1618 3242 1652 3276
rect 1618 3174 1652 3208
rect 1618 3106 1652 3140
rect 1618 3038 1652 3072
rect 1618 2970 1652 3004
rect 1618 2902 1652 2936
rect 1618 2834 1652 2868
rect 1618 2766 1652 2800
rect 1724 3242 1758 3276
rect 1724 3174 1758 3208
rect 1724 3106 1758 3140
rect 1724 3038 1758 3072
rect 1724 2970 1758 3004
rect 1724 2902 1758 2936
rect 1724 2834 1758 2868
rect 1724 2766 1758 2800
rect 1830 3242 1864 3276
rect 1830 3174 1864 3208
rect 1830 3106 1864 3140
rect 1830 3038 1864 3072
rect 1830 2970 1864 3004
rect 1830 2902 1864 2936
rect 1830 2834 1864 2868
rect 1830 2766 1864 2800
rect 1936 3242 1970 3276
rect 1936 3174 1970 3208
rect 1936 3106 1970 3140
rect 1936 3038 1970 3072
rect 1936 2970 1970 3004
rect 1936 2902 1970 2936
rect 1936 2834 1970 2868
rect 1936 2766 1970 2800
rect 2046 3308 2080 3342
rect 2046 3240 2080 3274
rect 2046 3172 2080 3206
rect 2046 3104 2080 3138
rect 2046 3036 2080 3070
rect 2046 2968 2080 3002
rect 2046 2900 2080 2934
rect 2046 2832 2080 2866
rect 2152 3308 2186 3342
rect 2152 3240 2186 3274
rect 2152 3172 2186 3206
rect 2152 3104 2186 3138
rect 2152 3036 2186 3070
rect 2152 2968 2186 3002
rect 2152 2900 2186 2934
rect 2152 2832 2186 2866
rect 2258 3308 2292 3342
rect 2258 3240 2292 3274
rect 2258 3172 2292 3206
rect 2258 3104 2292 3138
rect 2258 3036 2292 3070
rect 2258 2968 2292 3002
rect 2258 2900 2292 2934
rect 2258 2832 2292 2866
rect 334 2696 368 2730
rect 334 2628 368 2662
rect 334 2560 368 2594
rect 334 2492 368 2526
rect 334 2424 368 2458
<< mvndiffc >>
rect 171 199 205 233
rect 171 131 205 165
rect 171 63 205 97
rect 171 -5 205 29
rect 327 199 361 233
rect 327 131 361 165
rect 327 63 361 97
rect 327 -5 361 29
<< mvpdiffc >>
rect 851 2202 885 2236
rect 919 2202 953 2236
rect 987 2202 1021 2236
rect 1055 2202 1089 2236
rect 1123 2202 1157 2236
rect 1191 2202 1225 2236
rect 1259 2202 1293 2236
rect 1327 2202 1361 2236
rect 1395 2202 1429 2236
rect 1463 2202 1497 2236
rect 1531 2202 1565 2236
rect 1599 2202 1633 2236
rect 1667 2202 1701 2236
rect 1735 2202 1769 2236
rect 851 2046 885 2080
rect 919 2046 953 2080
rect 987 2046 1021 2080
rect 1055 2046 1089 2080
rect 1123 2046 1157 2080
rect 1191 2046 1225 2080
rect 1259 2046 1293 2080
rect 1327 2046 1361 2080
rect 1395 2046 1429 2080
rect 1463 2046 1497 2080
rect 1531 2046 1565 2080
rect 1599 2046 1633 2080
rect 1667 2046 1701 2080
rect 1735 2046 1769 2080
rect 851 1890 885 1924
rect 919 1890 953 1924
rect 987 1890 1021 1924
rect 1055 1890 1089 1924
rect 1123 1890 1157 1924
rect 1191 1890 1225 1924
rect 1259 1890 1293 1924
rect 1327 1890 1361 1924
rect 1395 1890 1429 1924
rect 1463 1890 1497 1924
rect 1531 1890 1565 1924
rect 1599 1890 1633 1924
rect 1667 1890 1701 1924
rect 1735 1890 1769 1924
<< psubdiff >>
rect 501 -431 525 -397
rect 559 -431 594 -397
rect 628 -431 663 -397
rect 697 -431 732 -397
rect 766 -431 801 -397
rect 835 -431 870 -397
rect 904 -431 939 -397
rect 973 -431 1007 -397
rect 1041 -431 1075 -397
rect 1109 -431 1143 -397
rect 1177 -431 1211 -397
rect 1245 -431 1279 -397
rect 1313 -431 1347 -397
rect 1381 -431 1415 -397
rect 1449 -431 1483 -397
rect 1517 -431 1551 -397
rect 1585 -431 1619 -397
rect 1653 -431 1687 -397
rect 1721 -431 1755 -397
rect 1789 -431 1823 -397
rect 1857 -431 1891 -397
rect 1925 -431 1959 -397
rect 1993 -431 2027 -397
rect 2061 -431 2095 -397
rect 2129 -431 2153 -397
<< nsubdiff >>
rect 145 3428 179 3462
rect 213 3428 247 3462
rect 281 3428 315 3462
rect 349 3428 383 3462
rect 417 3428 451 3462
rect 485 3428 519 3462
rect 553 3428 587 3462
rect 621 3428 655 3462
rect 689 3428 723 3462
rect 757 3428 791 3462
rect 825 3428 859 3462
rect 893 3428 927 3462
rect 961 3428 995 3462
rect 1029 3428 1063 3462
rect 1097 3428 1131 3462
rect 1165 3428 1199 3462
rect 1233 3428 1267 3462
rect 1301 3428 1335 3462
rect 1369 3428 1403 3462
rect 1437 3428 1471 3462
rect 1505 3428 1539 3462
rect 1573 3428 1607 3462
rect 1641 3428 1675 3462
rect 1709 3428 1743 3462
rect 1777 3428 1811 3462
rect 1845 3428 1879 3462
rect 1913 3428 1947 3462
rect 1981 3428 2015 3462
rect 2049 3428 2083 3462
rect 2117 3428 2151 3462
rect 2185 3428 2269 3462
<< mvnsubdiff >>
rect 1855 2155 1889 2243
rect 1855 2087 1889 2121
rect 1855 2019 1889 2053
rect 1855 1951 1889 1985
rect 1855 1883 1889 1917
<< psubdiffcont >>
rect 525 -431 559 -397
rect 594 -431 628 -397
rect 663 -431 697 -397
rect 732 -431 766 -397
rect 801 -431 835 -397
rect 870 -431 904 -397
rect 939 -431 973 -397
rect 1007 -431 1041 -397
rect 1075 -431 1109 -397
rect 1143 -431 1177 -397
rect 1211 -431 1245 -397
rect 1279 -431 1313 -397
rect 1347 -431 1381 -397
rect 1415 -431 1449 -397
rect 1483 -431 1517 -397
rect 1551 -431 1585 -397
rect 1619 -431 1653 -397
rect 1687 -431 1721 -397
rect 1755 -431 1789 -397
rect 1823 -431 1857 -397
rect 1891 -431 1925 -397
rect 1959 -431 1993 -397
rect 2027 -431 2061 -397
rect 2095 -431 2129 -397
<< nsubdiffcont >>
rect 179 3428 213 3462
rect 247 3428 281 3462
rect 315 3428 349 3462
rect 383 3428 417 3462
rect 451 3428 485 3462
rect 519 3428 553 3462
rect 587 3428 621 3462
rect 655 3428 689 3462
rect 723 3428 757 3462
rect 791 3428 825 3462
rect 859 3428 893 3462
rect 927 3428 961 3462
rect 995 3428 1029 3462
rect 1063 3428 1097 3462
rect 1131 3428 1165 3462
rect 1199 3428 1233 3462
rect 1267 3428 1301 3462
rect 1335 3428 1369 3462
rect 1403 3428 1437 3462
rect 1471 3428 1505 3462
rect 1539 3428 1573 3462
rect 1607 3428 1641 3462
rect 1675 3428 1709 3462
rect 1743 3428 1777 3462
rect 1811 3428 1845 3462
rect 1879 3428 1913 3462
rect 1947 3428 1981 3462
rect 2015 3428 2049 3462
rect 2083 3428 2117 3462
rect 2151 3428 2185 3462
<< mvnsubdiffcont >>
rect 1855 2121 1889 2155
rect 1855 2053 1889 2087
rect 1855 1985 1889 2019
rect 1855 1917 1889 1951
<< poly >>
rect 167 3354 217 3386
rect 273 3354 323 3386
rect 489 3354 539 3386
rect 595 3354 645 3386
rect 701 3354 751 3386
rect 807 3354 857 3386
rect 1023 3354 1073 3386
rect 1129 3354 1179 3386
rect 1235 3354 1285 3386
rect 1341 3354 1391 3386
rect 1557 3354 1607 3386
rect 1663 3354 1713 3386
rect 1769 3354 1819 3386
rect 1875 3354 1925 3386
rect 2091 3354 2141 3386
rect 2197 3354 2247 3386
rect 489 2722 539 2754
rect 595 2722 645 2754
rect 489 2706 645 2722
rect 489 2672 505 2706
rect 539 2672 595 2706
rect 629 2672 645 2706
rect 489 2656 645 2672
rect 701 2722 751 2754
rect 807 2722 857 2754
rect 701 2706 857 2722
rect 701 2672 717 2706
rect 751 2672 807 2706
rect 841 2672 857 2706
rect 701 2656 857 2672
rect 1023 2722 1073 2754
rect 1129 2722 1179 2754
rect 1235 2722 1285 2754
rect 1341 2722 1391 2754
rect 1023 2706 1391 2722
rect 1023 2672 1039 2706
rect 1073 2672 1115 2706
rect 1149 2672 1191 2706
rect 1225 2672 1266 2706
rect 1300 2672 1341 2706
rect 1375 2672 1391 2706
rect 1023 2656 1391 2672
rect 1557 2722 1607 2754
rect 1663 2722 1713 2754
rect 1557 2706 1713 2722
rect 1557 2672 1573 2706
rect 1607 2672 1663 2706
rect 1697 2672 1713 2706
rect 1557 2656 1713 2672
rect 1769 2722 1819 2754
rect 1875 2722 1925 2754
rect 2091 2722 2141 2754
rect 1769 2706 1925 2722
rect 1769 2672 1785 2706
rect 1819 2672 1875 2706
rect 1909 2672 1925 2706
rect 1769 2656 1925 2672
rect 2075 2706 2141 2722
rect 2075 2672 2091 2706
rect 2125 2672 2141 2706
rect 2075 2616 2141 2672
rect 2075 2582 2091 2616
rect 2125 2582 2141 2616
rect 2075 2566 2141 2582
rect 2197 2722 2247 2754
rect 2197 2706 2263 2722
rect 2197 2672 2213 2706
rect 2247 2672 2263 2706
rect 2197 2616 2263 2672
rect 2197 2582 2213 2616
rect 2247 2582 2263 2616
rect 2197 2566 2263 2582
rect 167 2322 217 2354
rect 151 2306 217 2322
rect 151 2272 167 2306
rect 201 2272 217 2306
rect 151 2238 217 2272
rect 151 2204 167 2238
rect 201 2204 217 2238
rect 151 2188 217 2204
rect 273 2322 323 2354
rect 273 2306 339 2322
rect 273 2272 289 2306
rect 323 2272 339 2306
rect 273 2238 339 2272
rect 273 2204 289 2238
rect 323 2204 339 2238
rect 273 2188 339 2204
rect 683 2175 781 2191
rect 683 2141 699 2175
rect 733 2141 781 2175
rect 683 2091 781 2141
rect 1781 2091 1813 2191
rect 683 2080 749 2091
rect 683 2046 699 2080
rect 733 2046 749 2080
rect 683 2035 749 2046
rect 683 1985 781 2035
rect 683 1951 699 1985
rect 733 1951 781 1985
rect 683 1935 781 1951
rect 1781 1935 1813 2035
rect 216 365 350 381
rect 216 331 232 365
rect 266 331 300 365
rect 334 331 350 365
rect 216 315 350 331
rect 470 365 604 381
rect 470 331 486 365
rect 520 331 554 365
rect 588 331 604 365
rect 470 315 604 331
rect 216 283 316 315
rect 554 283 604 315
rect 660 365 794 381
rect 660 331 676 365
rect 710 331 744 365
rect 778 331 794 365
rect 660 315 794 331
rect 876 365 1032 381
rect 876 331 892 365
rect 926 331 982 365
rect 1016 331 1032 365
rect 876 315 1032 331
rect 660 283 710 315
rect 876 283 926 315
rect 982 283 1032 315
rect 1088 365 1244 381
rect 1088 331 1104 365
rect 1138 331 1194 365
rect 1228 331 1244 365
rect 1088 315 1244 331
rect 1088 283 1138 315
rect 1194 283 1244 315
rect 1410 365 1566 381
rect 1410 331 1426 365
rect 1460 331 1516 365
rect 1550 331 1566 365
rect 1410 315 1566 331
rect 1410 283 1460 315
rect 1516 283 1566 315
rect 1732 365 1888 381
rect 1732 331 1748 365
rect 1782 331 1838 365
rect 1872 331 1888 365
rect 1732 315 1888 331
rect 1732 283 1782 315
rect 1838 283 1888 315
rect 1944 365 2100 381
rect 1944 331 1960 365
rect 1994 331 2050 365
rect 2084 331 2100 365
rect 1944 315 2100 331
rect 1944 283 1994 315
rect 2050 283 2100 315
rect 216 -49 316 -17
rect 554 -349 604 -317
rect 660 -349 710 -317
rect 876 -349 926 -317
rect 982 -349 1032 -317
rect 1088 -349 1138 -317
rect 1194 -349 1244 -317
rect 1410 -349 1460 -317
rect 1516 -349 1566 -317
rect 1732 -349 1782 -317
rect 1838 -349 1888 -317
rect 1944 -349 1994 -317
rect 2050 -349 2100 -317
<< polycont >>
rect 505 2672 539 2706
rect 595 2672 629 2706
rect 717 2672 751 2706
rect 807 2672 841 2706
rect 1039 2672 1073 2706
rect 1115 2672 1149 2706
rect 1191 2672 1225 2706
rect 1266 2672 1300 2706
rect 1341 2672 1375 2706
rect 1573 2672 1607 2706
rect 1663 2672 1697 2706
rect 1785 2672 1819 2706
rect 1875 2672 1909 2706
rect 2091 2672 2125 2706
rect 2091 2582 2125 2616
rect 2213 2672 2247 2706
rect 2213 2582 2247 2616
rect 167 2272 201 2306
rect 167 2204 201 2238
rect 289 2272 323 2306
rect 289 2204 323 2238
rect 699 2141 733 2175
rect 699 2046 733 2080
rect 699 1951 733 1985
rect 232 331 266 365
rect 300 331 334 365
rect 486 331 520 365
rect 554 331 588 365
rect 676 331 710 365
rect 744 331 778 365
rect 892 331 926 365
rect 982 331 1016 365
rect 1104 331 1138 365
rect 1194 331 1228 365
rect 1426 331 1460 365
rect 1516 331 1550 365
rect 1748 331 1782 365
rect 1838 331 1872 365
rect 1960 331 1994 365
rect 2050 331 2084 365
<< locali >>
rect 145 3428 157 3462
rect 213 3428 231 3462
rect 281 3428 305 3462
rect 349 3428 379 3462
rect 417 3428 451 3462
rect 487 3428 519 3462
rect 561 3428 587 3462
rect 635 3428 655 3462
rect 709 3428 723 3462
rect 783 3428 791 3462
rect 857 3428 859 3462
rect 893 3428 897 3462
rect 961 3428 971 3462
rect 1029 3428 1045 3462
rect 1097 3428 1119 3462
rect 1165 3428 1193 3462
rect 1233 3428 1267 3462
rect 1301 3428 1335 3462
rect 1375 3428 1403 3462
rect 1449 3428 1471 3462
rect 1523 3428 1539 3462
rect 1597 3428 1607 3462
rect 1671 3428 1675 3462
rect 1709 3428 1711 3462
rect 1777 3428 1785 3462
rect 1845 3428 1858 3462
rect 1913 3428 1931 3462
rect 1981 3428 2004 3462
rect 2049 3428 2077 3462
rect 2117 3428 2150 3462
rect 2185 3428 2223 3462
rect 2257 3428 2269 3462
rect 122 3342 156 3358
rect 122 3274 156 3308
rect 122 3206 156 3240
rect 122 3138 156 3154
rect 122 3070 156 3081
rect 122 3002 156 3008
rect 122 2934 156 2935
rect 122 2896 156 2900
rect 122 2823 156 2832
rect 122 2749 156 2764
rect 122 2675 156 2696
rect 122 2601 156 2628
rect 122 2527 156 2560
rect 122 2458 156 2492
rect 122 2408 156 2424
rect 228 3342 262 3358
rect 228 3274 262 3308
rect 228 3206 262 3232
rect 228 3138 262 3156
rect 228 3070 262 3080
rect 228 3002 262 3004
rect 228 2961 262 2968
rect 228 2884 262 2900
rect 228 2807 262 2832
rect 228 2730 262 2764
rect 228 2662 262 2696
rect 228 2594 262 2619
rect 228 2526 262 2542
rect 228 2458 262 2465
rect 228 2408 262 2424
rect 334 3342 368 3358
rect 2046 3342 2080 3358
rect 334 3274 368 3308
rect 334 3206 368 3240
rect 334 3138 368 3154
rect 334 3070 368 3078
rect 334 2960 368 2968
rect 334 2884 368 2900
rect 334 2807 368 2832
rect 334 2730 368 2764
rect 444 3276 478 3292
rect 444 3208 478 3242
rect 444 3140 478 3156
rect 444 3072 478 3078
rect 444 3034 478 3038
rect 444 2956 478 2970
rect 444 2878 478 2902
rect 444 2800 478 2834
rect 444 2750 478 2766
rect 550 3276 584 3292
rect 550 3224 584 3242
rect 550 3146 584 3174
rect 550 3072 584 3106
rect 550 3004 584 3034
rect 550 2936 584 2956
rect 550 2868 584 2878
rect 550 2800 584 2834
rect 550 2750 584 2766
rect 656 3276 690 3292
rect 656 3208 690 3242
rect 656 3140 690 3156
rect 656 3072 690 3078
rect 656 3034 690 3038
rect 656 2956 690 2970
rect 656 2878 690 2902
rect 656 2800 690 2834
rect 656 2750 690 2766
rect 762 3276 796 3308
rect 762 3208 796 3222
rect 762 3170 796 3174
rect 762 3084 796 3106
rect 762 3004 796 3038
rect 762 2936 796 2964
rect 762 2868 796 2878
rect 762 2800 796 2834
rect 762 2750 796 2766
rect 868 3276 902 3292
rect 868 3208 902 3242
rect 868 3140 902 3156
rect 868 3072 902 3078
rect 868 3034 902 3038
rect 868 2956 902 2970
rect 868 2878 902 2902
rect 868 2800 902 2834
rect 868 2750 902 2766
rect 978 3276 1012 3308
rect 978 3208 1012 3235
rect 978 3140 1012 3162
rect 978 3072 1012 3089
rect 978 3004 1012 3015
rect 978 2936 1012 2941
rect 978 2901 1012 2902
rect 978 2800 1012 2834
rect 978 2750 1012 2766
rect 1084 3276 1118 3292
rect 1084 3208 1118 3242
rect 1084 3140 1118 3156
rect 1084 3072 1118 3078
rect 1084 3034 1118 3038
rect 1084 2956 1118 2970
rect 1084 2878 1118 2902
rect 1084 2800 1118 2834
rect 1084 2750 1118 2766
rect 1190 3276 1224 3308
rect 1190 3208 1224 3235
rect 1190 3140 1224 3162
rect 1190 3072 1224 3089
rect 1190 3004 1224 3015
rect 1190 2936 1224 2941
rect 1190 2901 1224 2902
rect 1190 2800 1224 2834
rect 1190 2750 1224 2766
rect 1296 3276 1330 3292
rect 1296 3208 1330 3242
rect 1296 3140 1330 3156
rect 1296 3072 1330 3078
rect 1296 3034 1330 3038
rect 1296 2956 1330 2970
rect 1296 2878 1330 2902
rect 1296 2800 1330 2834
rect 1296 2750 1330 2766
rect 1402 3276 1436 3308
rect 1402 3208 1436 3235
rect 1402 3140 1436 3162
rect 1402 3072 1436 3089
rect 1402 3004 1436 3015
rect 1402 2936 1436 2941
rect 1402 2901 1436 2902
rect 1402 2800 1436 2834
rect 1402 2750 1436 2766
rect 1512 3276 1546 3292
rect 1512 3208 1546 3242
rect 1512 3140 1546 3156
rect 1512 3072 1546 3078
rect 1512 3034 1546 3038
rect 1512 2956 1546 2970
rect 1512 2878 1546 2902
rect 1512 2800 1546 2834
rect 1512 2750 1546 2766
rect 1618 3276 1652 3308
rect 1618 3208 1652 3222
rect 1618 3170 1652 3174
rect 1618 3084 1652 3106
rect 1618 3004 1652 3038
rect 1618 2936 1652 2964
rect 1618 2868 1652 2878
rect 1618 2800 1652 2834
rect 1618 2750 1652 2766
rect 1724 3276 1758 3292
rect 1724 3208 1758 3242
rect 1724 3140 1758 3156
rect 1724 3072 1758 3078
rect 1724 3034 1758 3038
rect 1724 2956 1758 2970
rect 1724 2878 1758 2902
rect 1724 2800 1758 2834
rect 1724 2750 1758 2766
rect 1830 3276 1864 3292
rect 1830 3224 1864 3242
rect 1830 3146 1864 3174
rect 1830 3072 1864 3106
rect 1830 3004 1864 3034
rect 1830 2936 1864 2956
rect 1830 2868 1864 2878
rect 1830 2800 1864 2834
rect 1830 2750 1864 2766
rect 1936 3276 1970 3292
rect 1936 3208 1970 3242
rect 1936 3140 1970 3156
rect 1936 3072 1970 3078
rect 1936 3034 1970 3038
rect 1936 2956 1970 2970
rect 1936 2878 1970 2902
rect 1936 2800 1970 2834
rect 2046 3274 2080 3308
rect 2046 3206 2080 3240
rect 2046 3138 2080 3156
rect 2046 3070 2080 3078
rect 2046 3034 2080 3036
rect 2046 2956 2080 2968
rect 2046 2878 2080 2900
rect 2046 2800 2080 2832
rect 2152 3342 2186 3358
rect 2152 3274 2186 3308
rect 2152 3206 2186 3240
rect 2152 3138 2186 3156
rect 2152 3070 2186 3078
rect 2152 3034 2186 3036
rect 2152 2956 2186 2968
rect 2152 2878 2186 2900
rect 2152 2800 2186 2832
rect 2258 3342 2292 3358
rect 2258 3274 2292 3308
rect 2258 3206 2292 3235
rect 2258 3138 2292 3162
rect 2258 3070 2292 3089
rect 2258 3002 2292 3015
rect 2258 2934 2292 2941
rect 2258 2866 2292 2867
rect 2258 2816 2292 2832
rect 1936 2750 1970 2766
rect 2091 2706 2125 2722
rect 334 2662 368 2696
rect 489 2672 500 2706
rect 539 2672 572 2706
rect 629 2672 645 2706
rect 701 2672 717 2706
rect 773 2672 807 2706
rect 845 2672 857 2706
rect 1023 2672 1039 2706
rect 1079 2672 1115 2706
rect 1175 2672 1191 2706
rect 1225 2672 1236 2706
rect 1300 2672 1331 2706
rect 1375 2672 1391 2706
rect 1557 2672 1573 2706
rect 1611 2672 1649 2706
rect 1697 2672 1713 2706
rect 1769 2672 1782 2706
rect 1819 2672 1854 2706
rect 1909 2672 1925 2706
rect 2213 2706 2247 2722
rect 334 2594 368 2619
rect 2091 2650 2092 2672
rect 2091 2616 2126 2650
rect 2125 2612 2126 2616
rect 2091 2578 2092 2582
rect 2213 2616 2247 2650
rect 2091 2566 2125 2578
rect 2213 2566 2247 2578
rect 334 2526 368 2542
rect 334 2458 368 2465
rect 334 2408 368 2424
rect 167 2310 201 2322
rect 198 2306 201 2310
rect 164 2272 167 2276
rect 164 2238 201 2272
rect 167 2188 201 2204
rect 289 2310 323 2322
rect 289 2238 323 2272
rect 289 2188 323 2204
rect 835 2202 846 2236
rect 885 2202 919 2236
rect 955 2202 987 2236
rect 1030 2202 1055 2236
rect 1105 2202 1123 2236
rect 1180 2202 1191 2236
rect 1255 2202 1259 2236
rect 1293 2202 1295 2236
rect 1361 2202 1369 2236
rect 1429 2202 1443 2236
rect 1497 2202 1517 2236
rect 1565 2202 1591 2236
rect 1633 2202 1665 2236
rect 1701 2202 1735 2236
rect 1773 2202 1785 2236
rect 1855 2230 1889 2243
rect 699 2179 733 2191
rect 732 2175 733 2179
rect 698 2141 699 2145
rect 698 2080 733 2141
rect 1855 2155 1889 2196
rect 1855 2087 1889 2121
rect 835 2046 846 2080
rect 885 2046 919 2080
rect 959 2046 987 2080
rect 1038 2046 1055 2080
rect 1117 2046 1123 2080
rect 1157 2046 1162 2080
rect 1225 2046 1240 2080
rect 1293 2046 1318 2080
rect 1361 2046 1395 2080
rect 1430 2046 1463 2080
rect 1508 2046 1531 2080
rect 1586 2046 1599 2080
rect 1664 2046 1667 2080
rect 1701 2046 1735 2080
rect 1769 2046 1785 2080
rect 698 1985 733 2046
rect 698 1981 699 1985
rect 732 1947 733 1951
rect 699 1935 733 1947
rect 1855 2019 1889 2046
rect 1855 1951 1889 1971
rect 880 1924 921 1926
rect 955 1924 996 1926
rect 1030 1924 1071 1926
rect 1105 1924 1146 1926
rect 1180 1924 1221 1926
rect 1255 1924 1295 1926
rect 1329 1924 1369 1926
rect 1403 1924 1443 1926
rect 1477 1924 1517 1926
rect 1551 1924 1591 1926
rect 1625 1924 1665 1926
rect 1699 1924 1739 1926
rect 835 1892 846 1924
rect 835 1890 851 1892
rect 885 1890 919 1924
rect 955 1892 987 1924
rect 1030 1892 1055 1924
rect 1105 1892 1123 1924
rect 1180 1892 1191 1924
rect 1255 1892 1259 1924
rect 953 1890 987 1892
rect 1021 1890 1055 1892
rect 1089 1890 1123 1892
rect 1157 1890 1191 1892
rect 1225 1890 1259 1892
rect 1293 1892 1295 1924
rect 1361 1892 1369 1924
rect 1429 1892 1443 1924
rect 1497 1892 1517 1924
rect 1565 1892 1591 1924
rect 1633 1892 1665 1924
rect 1293 1890 1327 1892
rect 1361 1890 1395 1892
rect 1429 1890 1463 1892
rect 1497 1890 1531 1892
rect 1565 1890 1599 1892
rect 1633 1890 1667 1892
rect 1701 1890 1735 1924
rect 1773 1892 1785 1924
rect 1769 1890 1785 1892
rect 1855 1883 1889 1896
rect 216 331 228 365
rect 266 331 300 365
rect 334 331 350 365
rect 470 331 477 365
rect 520 331 549 365
rect 588 331 604 365
rect 660 331 672 365
rect 710 331 744 365
rect 778 331 794 365
rect 876 331 892 365
rect 931 331 969 365
rect 1016 331 1032 365
rect 1088 331 1104 365
rect 1152 331 1190 365
rect 1228 331 1244 365
rect 1410 331 1426 365
rect 1472 331 1510 365
rect 1550 331 1566 365
rect 1732 331 1748 365
rect 1797 331 1835 365
rect 1872 331 1888 365
rect 1944 331 1960 365
rect 2016 331 2050 365
rect 2088 331 2100 365
rect 171 237 205 249
rect 171 165 205 199
rect 171 97 205 99
rect 171 29 205 63
rect 171 -21 205 -5
rect 327 233 361 249
rect 327 191 361 199
rect 327 110 361 131
rect 327 29 361 63
rect 327 -21 361 -5
rect 509 205 543 221
rect 509 137 543 157
rect 509 69 543 81
rect 509 1 543 5
rect 509 -37 543 -33
rect 509 -113 543 -101
rect 509 -189 543 -169
rect 509 -271 543 -237
rect 509 -321 543 -305
rect 615 205 649 221
rect 615 145 649 171
rect 615 73 649 103
rect 615 1 649 35
rect 615 -67 649 -33
rect 615 -135 649 -105
rect 615 -203 649 -177
rect 615 -271 649 -249
rect 721 209 755 221
rect 721 137 755 171
rect 721 69 755 96
rect 721 1 755 17
rect 721 -67 755 -63
rect 721 -109 755 -101
rect 721 -189 755 -169
rect 721 -271 755 -237
rect 721 -321 755 -305
rect 831 209 865 221
rect 831 137 865 171
rect 831 69 865 96
rect 831 1 865 17
rect 831 -67 865 -63
rect 831 -109 865 -101
rect 831 -189 865 -169
rect 831 -271 865 -237
rect 831 -321 865 -305
rect 937 205 971 221
rect 937 161 971 171
rect 937 74 971 103
rect 937 1 971 35
rect 937 -67 971 -47
rect 937 -189 971 -169
rect 937 -271 971 -237
rect 937 -321 971 -305
rect 1043 209 1077 221
rect 1043 137 1077 171
rect 1043 69 1077 96
rect 1043 1 1077 17
rect 1043 -67 1077 -63
rect 1043 -109 1077 -101
rect 1043 -189 1077 -169
rect 1043 -271 1077 -237
rect 1043 -321 1077 -305
rect 1149 205 1183 221
rect 1149 137 1183 171
rect 1149 69 1183 101
rect 1149 1 1183 17
rect 1149 -117 1183 -101
rect 1149 -202 1183 -169
rect 1149 -271 1183 -237
rect 1255 209 1289 221
rect 1255 137 1289 171
rect 1255 69 1289 96
rect 1255 1 1289 17
rect 1255 -67 1289 -63
rect 1255 -109 1289 -101
rect 1255 -189 1289 -169
rect 1255 -271 1289 -237
rect 1255 -321 1289 -305
rect 1365 205 1399 221
rect 1365 137 1399 171
rect 1365 69 1399 101
rect 1365 1 1399 17
rect 1365 -117 1399 -101
rect 1365 -202 1399 -169
rect 1365 -271 1399 -237
rect 1471 209 1505 221
rect 1471 137 1505 171
rect 1471 69 1505 96
rect 1471 1 1505 17
rect 1471 -67 1505 -63
rect 1471 -109 1505 -101
rect 1471 -189 1505 -169
rect 1471 -271 1505 -237
rect 1471 -321 1505 -305
rect 1577 205 1611 221
rect 1577 137 1611 171
rect 1577 69 1611 101
rect 1577 1 1611 17
rect 1577 -117 1611 -101
rect 1577 -202 1611 -169
rect 1577 -271 1611 -237
rect 1687 209 1721 221
rect 1687 137 1721 171
rect 1687 69 1721 96
rect 1687 1 1721 17
rect 1687 -67 1721 -63
rect 1687 -109 1721 -101
rect 1687 -189 1721 -169
rect 1687 -271 1721 -237
rect 1687 -321 1721 -305
rect 1793 205 1827 221
rect 1793 161 1827 171
rect 1793 74 1827 103
rect 1793 1 1827 35
rect 1793 -67 1827 -47
rect 1793 -189 1827 -169
rect 1793 -271 1827 -237
rect 1793 -321 1827 -305
rect 1899 209 1933 221
rect 1899 137 1933 171
rect 1899 69 1933 96
rect 1899 1 1933 17
rect 1899 -67 1933 -63
rect 1899 -109 1933 -101
rect 1899 -189 1933 -169
rect 1899 -271 1933 -237
rect 1899 -321 1933 -305
rect 2005 205 2039 221
rect 2005 137 2039 171
rect 2005 69 2039 101
rect 2005 1 2039 17
rect 2005 -117 2039 -101
rect 2005 -202 2039 -169
rect 2005 -271 2039 -237
rect 2111 209 2145 221
rect 2111 137 2145 171
rect 2111 69 2145 96
rect 2111 1 2145 17
rect 2111 -67 2145 -63
rect 2111 -109 2145 -101
rect 2111 -189 2145 -169
rect 2111 -271 2145 -237
rect 2111 -321 2145 -305
rect 559 -431 575 -397
rect 628 -431 649 -397
rect 697 -431 723 -397
rect 766 -431 797 -397
rect 835 -431 870 -397
rect 905 -431 939 -397
rect 979 -431 1007 -397
rect 1053 -431 1075 -397
rect 1127 -431 1143 -397
rect 1201 -431 1211 -397
rect 1275 -431 1279 -397
rect 1313 -431 1315 -397
rect 1381 -431 1388 -397
rect 1449 -431 1461 -397
rect 1517 -431 1534 -397
rect 1585 -431 1607 -397
rect 1653 -431 1680 -397
rect 1721 -431 1753 -397
rect 1789 -431 1823 -397
rect 1860 -431 1891 -397
rect 1933 -431 1959 -397
rect 2006 -431 2027 -397
rect 2079 -431 2095 -397
rect 2152 -431 2153 -397
<< viali >>
rect 157 3428 179 3462
rect 179 3428 191 3462
rect 231 3428 247 3462
rect 247 3428 265 3462
rect 305 3428 315 3462
rect 315 3428 339 3462
rect 379 3428 383 3462
rect 383 3428 413 3462
rect 453 3428 485 3462
rect 485 3428 487 3462
rect 527 3428 553 3462
rect 553 3428 561 3462
rect 601 3428 621 3462
rect 621 3428 635 3462
rect 675 3428 689 3462
rect 689 3428 709 3462
rect 749 3428 757 3462
rect 757 3428 783 3462
rect 823 3428 825 3462
rect 825 3428 857 3462
rect 897 3428 927 3462
rect 927 3428 931 3462
rect 971 3428 995 3462
rect 995 3428 1005 3462
rect 1045 3428 1063 3462
rect 1063 3428 1079 3462
rect 1119 3428 1131 3462
rect 1131 3428 1153 3462
rect 1193 3428 1199 3462
rect 1199 3428 1227 3462
rect 1267 3428 1301 3462
rect 1341 3428 1369 3462
rect 1369 3428 1375 3462
rect 1415 3428 1437 3462
rect 1437 3428 1449 3462
rect 1489 3428 1505 3462
rect 1505 3428 1523 3462
rect 1563 3428 1573 3462
rect 1573 3428 1597 3462
rect 1637 3428 1641 3462
rect 1641 3428 1671 3462
rect 1711 3428 1743 3462
rect 1743 3428 1745 3462
rect 1785 3428 1811 3462
rect 1811 3428 1819 3462
rect 1858 3428 1879 3462
rect 1879 3428 1892 3462
rect 1931 3428 1947 3462
rect 1947 3428 1965 3462
rect 2004 3428 2015 3462
rect 2015 3428 2038 3462
rect 2077 3428 2083 3462
rect 2083 3428 2111 3462
rect 2150 3428 2151 3462
rect 2151 3428 2184 3462
rect 2223 3428 2257 3462
rect 122 3172 156 3188
rect 122 3154 156 3172
rect 122 3104 156 3115
rect 122 3081 156 3104
rect 122 3036 156 3042
rect 122 3008 156 3036
rect 122 2968 156 2969
rect 122 2935 156 2968
rect 122 2866 156 2896
rect 122 2862 156 2866
rect 122 2798 156 2823
rect 122 2789 156 2798
rect 122 2730 156 2749
rect 122 2715 156 2730
rect 122 2662 156 2675
rect 122 2641 156 2662
rect 122 2594 156 2601
rect 122 2567 156 2594
rect 122 2526 156 2527
rect 122 2493 156 2526
rect 228 3308 262 3342
rect 228 3240 262 3266
rect 228 3232 262 3240
rect 228 3172 262 3190
rect 228 3156 262 3172
rect 228 3104 262 3114
rect 228 3080 262 3104
rect 228 3036 262 3038
rect 228 3004 262 3036
rect 228 2934 262 2961
rect 228 2927 262 2934
rect 228 2866 262 2884
rect 228 2850 262 2866
rect 228 2798 262 2807
rect 228 2773 262 2798
rect 228 2696 262 2730
rect 228 2628 262 2653
rect 228 2619 262 2628
rect 228 2560 262 2576
rect 228 2542 262 2560
rect 228 2492 262 2499
rect 228 2465 262 2492
rect 762 3308 796 3342
rect 334 3172 368 3188
rect 334 3154 368 3172
rect 334 3104 368 3112
rect 334 3078 368 3104
rect 334 3002 368 3036
rect 334 2934 368 2960
rect 334 2926 368 2934
rect 334 2866 368 2884
rect 334 2850 368 2866
rect 334 2798 368 2807
rect 334 2773 368 2798
rect 444 3174 478 3190
rect 444 3156 478 3174
rect 444 3106 478 3112
rect 444 3078 478 3106
rect 444 3004 478 3034
rect 444 3000 478 3004
rect 444 2936 478 2956
rect 444 2922 478 2936
rect 444 2868 478 2878
rect 444 2844 478 2868
rect 444 2766 478 2800
rect 550 3208 584 3224
rect 550 3190 584 3208
rect 550 3140 584 3146
rect 550 3112 584 3140
rect 550 3038 584 3068
rect 550 3034 584 3038
rect 550 2970 584 2990
rect 550 2956 584 2970
rect 550 2902 584 2912
rect 550 2878 584 2902
rect 656 3174 690 3190
rect 656 3156 690 3174
rect 656 3106 690 3112
rect 656 3078 690 3106
rect 656 3004 690 3034
rect 656 3000 690 3004
rect 656 2936 690 2956
rect 656 2922 690 2936
rect 656 2868 690 2878
rect 656 2844 690 2868
rect 656 2766 690 2800
rect 978 3308 1012 3342
rect 762 3242 796 3256
rect 762 3222 796 3242
rect 762 3140 796 3170
rect 762 3136 796 3140
rect 762 3072 796 3084
rect 762 3050 796 3072
rect 762 2970 796 2998
rect 762 2964 796 2970
rect 762 2902 796 2912
rect 762 2878 796 2902
rect 868 3174 902 3190
rect 868 3156 902 3174
rect 868 3106 902 3112
rect 868 3078 902 3106
rect 868 3004 902 3034
rect 868 3000 902 3004
rect 868 2936 902 2956
rect 868 2922 902 2936
rect 868 2868 902 2878
rect 868 2844 902 2868
rect 868 2766 902 2800
rect 1190 3308 1224 3342
rect 978 3242 1012 3269
rect 978 3235 1012 3242
rect 978 3174 1012 3196
rect 978 3162 1012 3174
rect 978 3106 1012 3123
rect 978 3089 1012 3106
rect 978 3038 1012 3049
rect 978 3015 1012 3038
rect 978 2970 1012 2975
rect 978 2941 1012 2970
rect 978 2868 1012 2901
rect 978 2867 1012 2868
rect 1084 3174 1118 3190
rect 1084 3156 1118 3174
rect 1084 3106 1118 3112
rect 1084 3078 1118 3106
rect 1084 3004 1118 3034
rect 1084 3000 1118 3004
rect 1084 2936 1118 2956
rect 1084 2922 1118 2936
rect 1084 2868 1118 2878
rect 1084 2844 1118 2868
rect 1084 2766 1118 2800
rect 1402 3308 1436 3342
rect 1190 3242 1224 3269
rect 1190 3235 1224 3242
rect 1190 3174 1224 3196
rect 1190 3162 1224 3174
rect 1190 3106 1224 3123
rect 1190 3089 1224 3106
rect 1190 3038 1224 3049
rect 1190 3015 1224 3038
rect 1190 2970 1224 2975
rect 1190 2941 1224 2970
rect 1190 2868 1224 2901
rect 1190 2867 1224 2868
rect 1296 3174 1330 3190
rect 1296 3156 1330 3174
rect 1296 3106 1330 3112
rect 1296 3078 1330 3106
rect 1296 3004 1330 3034
rect 1296 3000 1330 3004
rect 1296 2936 1330 2956
rect 1296 2922 1330 2936
rect 1296 2868 1330 2878
rect 1296 2844 1330 2868
rect 1296 2766 1330 2800
rect 1618 3308 1652 3342
rect 1402 3242 1436 3269
rect 1402 3235 1436 3242
rect 1402 3174 1436 3196
rect 1402 3162 1436 3174
rect 1402 3106 1436 3123
rect 1402 3089 1436 3106
rect 1402 3038 1436 3049
rect 1402 3015 1436 3038
rect 1402 2970 1436 2975
rect 1402 2941 1436 2970
rect 1402 2868 1436 2901
rect 1402 2867 1436 2868
rect 1512 3174 1546 3190
rect 1512 3156 1546 3174
rect 1512 3106 1546 3112
rect 1512 3078 1546 3106
rect 1512 3004 1546 3034
rect 1512 3000 1546 3004
rect 1512 2936 1546 2956
rect 1512 2922 1546 2936
rect 1512 2868 1546 2878
rect 1512 2844 1546 2868
rect 1512 2766 1546 2800
rect 1618 3242 1652 3256
rect 1618 3222 1652 3242
rect 1618 3140 1652 3170
rect 1618 3136 1652 3140
rect 1618 3072 1652 3084
rect 1618 3050 1652 3072
rect 1618 2970 1652 2998
rect 1618 2964 1652 2970
rect 1618 2902 1652 2912
rect 1618 2878 1652 2902
rect 1724 3174 1758 3190
rect 1724 3156 1758 3174
rect 1724 3106 1758 3112
rect 1724 3078 1758 3106
rect 1724 3004 1758 3034
rect 1724 3000 1758 3004
rect 1724 2936 1758 2956
rect 1724 2922 1758 2936
rect 1724 2868 1758 2878
rect 1724 2844 1758 2868
rect 1724 2766 1758 2800
rect 1830 3208 1864 3224
rect 1830 3190 1864 3208
rect 1830 3140 1864 3146
rect 1830 3112 1864 3140
rect 1830 3038 1864 3068
rect 1830 3034 1864 3038
rect 1830 2970 1864 2990
rect 1830 2956 1864 2970
rect 1830 2902 1864 2912
rect 1830 2878 1864 2902
rect 1936 3174 1970 3190
rect 1936 3156 1970 3174
rect 1936 3106 1970 3112
rect 1936 3078 1970 3106
rect 1936 3004 1970 3034
rect 1936 3000 1970 3004
rect 1936 2936 1970 2956
rect 1936 2922 1970 2936
rect 1936 2868 1970 2878
rect 1936 2844 1970 2868
rect 1936 2766 1970 2800
rect 2046 3172 2080 3190
rect 2046 3156 2080 3172
rect 2046 3104 2080 3112
rect 2046 3078 2080 3104
rect 2046 3002 2080 3034
rect 2046 3000 2080 3002
rect 2046 2934 2080 2956
rect 2046 2922 2080 2934
rect 2046 2866 2080 2878
rect 2046 2844 2080 2866
rect 2046 2766 2080 2800
rect 2152 3172 2186 3190
rect 2152 3156 2186 3172
rect 2152 3104 2186 3112
rect 2152 3078 2186 3104
rect 2152 3002 2186 3034
rect 2152 3000 2186 3002
rect 2152 2934 2186 2956
rect 2152 2922 2186 2934
rect 2152 2866 2186 2878
rect 2152 2844 2186 2866
rect 2258 3308 2292 3342
rect 2258 3240 2292 3269
rect 2258 3235 2292 3240
rect 2258 3172 2292 3196
rect 2258 3162 2292 3172
rect 2258 3104 2292 3123
rect 2258 3089 2292 3104
rect 2258 3036 2292 3049
rect 2258 3015 2292 3036
rect 2258 2968 2292 2975
rect 2258 2941 2292 2968
rect 2258 2900 2292 2901
rect 2258 2867 2292 2900
rect 2152 2766 2186 2800
rect 334 2696 368 2730
rect 500 2672 505 2706
rect 505 2672 534 2706
rect 572 2672 595 2706
rect 595 2672 606 2706
rect 739 2672 751 2706
rect 751 2672 773 2706
rect 811 2672 841 2706
rect 841 2672 845 2706
rect 1045 2672 1073 2706
rect 1073 2672 1079 2706
rect 1141 2672 1149 2706
rect 1149 2672 1175 2706
rect 1236 2672 1266 2706
rect 1266 2672 1270 2706
rect 1331 2672 1341 2706
rect 1341 2672 1365 2706
rect 1577 2672 1607 2706
rect 1607 2672 1611 2706
rect 1649 2672 1663 2706
rect 1663 2672 1683 2706
rect 1782 2672 1785 2706
rect 1785 2672 1816 2706
rect 1854 2672 1875 2706
rect 1875 2672 1888 2706
rect 2092 2672 2125 2684
rect 2125 2672 2126 2684
rect 334 2628 368 2653
rect 334 2619 368 2628
rect 334 2560 368 2576
rect 2092 2650 2126 2672
rect 2092 2582 2125 2612
rect 2125 2582 2126 2612
rect 2092 2578 2126 2582
rect 2213 2672 2247 2684
rect 2213 2650 2247 2672
rect 2213 2582 2247 2612
rect 2213 2578 2247 2582
rect 334 2542 368 2560
rect 334 2492 368 2499
rect 334 2465 368 2492
rect 164 2306 198 2310
rect 164 2276 167 2306
rect 167 2276 198 2306
rect 164 2204 167 2238
rect 167 2204 198 2238
rect 289 2306 323 2310
rect 289 2276 323 2306
rect 289 2204 323 2238
rect 846 2202 851 2236
rect 851 2202 880 2236
rect 921 2202 953 2236
rect 953 2202 955 2236
rect 996 2202 1021 2236
rect 1021 2202 1030 2236
rect 1071 2202 1089 2236
rect 1089 2202 1105 2236
rect 1146 2202 1157 2236
rect 1157 2202 1180 2236
rect 1221 2202 1225 2236
rect 1225 2202 1255 2236
rect 1295 2202 1327 2236
rect 1327 2202 1329 2236
rect 1369 2202 1395 2236
rect 1395 2202 1403 2236
rect 1443 2202 1463 2236
rect 1463 2202 1477 2236
rect 1517 2202 1531 2236
rect 1531 2202 1551 2236
rect 1591 2202 1599 2236
rect 1599 2202 1625 2236
rect 1665 2202 1667 2236
rect 1667 2202 1699 2236
rect 1739 2202 1769 2236
rect 1769 2202 1773 2236
rect 1855 2196 1889 2230
rect 698 2175 732 2179
rect 698 2145 699 2175
rect 699 2145 732 2175
rect 1855 2121 1889 2155
rect 698 2046 699 2080
rect 699 2046 732 2080
rect 846 2046 851 2080
rect 851 2046 880 2080
rect 925 2046 953 2080
rect 953 2046 959 2080
rect 1004 2046 1021 2080
rect 1021 2046 1038 2080
rect 1083 2046 1089 2080
rect 1089 2046 1117 2080
rect 1162 2046 1191 2080
rect 1191 2046 1196 2080
rect 1240 2046 1259 2080
rect 1259 2046 1274 2080
rect 1318 2046 1327 2080
rect 1327 2046 1352 2080
rect 1396 2046 1429 2080
rect 1429 2046 1430 2080
rect 1474 2046 1497 2080
rect 1497 2046 1508 2080
rect 1552 2046 1565 2080
rect 1565 2046 1586 2080
rect 1630 2046 1633 2080
rect 1633 2046 1664 2080
rect 1855 2053 1889 2080
rect 1855 2046 1889 2053
rect 698 1951 699 1981
rect 699 1951 732 1981
rect 698 1947 732 1951
rect 1855 1985 1889 2005
rect 1855 1971 1889 1985
rect 846 1924 880 1926
rect 921 1924 955 1926
rect 996 1924 1030 1926
rect 1071 1924 1105 1926
rect 1146 1924 1180 1926
rect 1221 1924 1255 1926
rect 1295 1924 1329 1926
rect 1369 1924 1403 1926
rect 1443 1924 1477 1926
rect 1517 1924 1551 1926
rect 1591 1924 1625 1926
rect 1665 1924 1699 1926
rect 1739 1924 1773 1926
rect 846 1892 851 1924
rect 851 1892 880 1924
rect 921 1892 953 1924
rect 953 1892 955 1924
rect 996 1892 1021 1924
rect 1021 1892 1030 1924
rect 1071 1892 1089 1924
rect 1089 1892 1105 1924
rect 1146 1892 1157 1924
rect 1157 1892 1180 1924
rect 1221 1892 1225 1924
rect 1225 1892 1255 1924
rect 1295 1892 1327 1924
rect 1327 1892 1329 1924
rect 1369 1892 1395 1924
rect 1395 1892 1403 1924
rect 1443 1892 1463 1924
rect 1463 1892 1477 1924
rect 1517 1892 1531 1924
rect 1531 1892 1551 1924
rect 1591 1892 1599 1924
rect 1599 1892 1625 1924
rect 1665 1892 1667 1924
rect 1667 1892 1699 1924
rect 1739 1892 1769 1924
rect 1769 1892 1773 1924
rect 1855 1917 1889 1930
rect 1855 1896 1889 1917
rect 228 331 232 365
rect 232 331 262 365
rect 300 331 334 365
rect 477 331 486 365
rect 486 331 511 365
rect 549 331 554 365
rect 554 331 583 365
rect 672 331 676 365
rect 676 331 706 365
rect 744 331 778 365
rect 897 331 926 365
rect 926 331 931 365
rect 969 331 982 365
rect 982 331 1003 365
rect 1118 331 1138 365
rect 1138 331 1152 365
rect 1190 331 1194 365
rect 1194 331 1224 365
rect 1438 331 1460 365
rect 1460 331 1472 365
rect 1510 331 1516 365
rect 1516 331 1544 365
rect 1763 331 1782 365
rect 1782 331 1797 365
rect 1835 331 1838 365
rect 1838 331 1869 365
rect 1982 331 1994 365
rect 1994 331 2016 365
rect 2054 331 2084 365
rect 2084 331 2088 365
rect 171 233 205 237
rect 171 203 205 233
rect 171 131 205 133
rect 171 99 205 131
rect 171 -5 205 29
rect 327 165 361 191
rect 327 157 361 165
rect 327 97 361 110
rect 327 76 361 97
rect 327 -5 361 29
rect 509 171 543 191
rect 509 157 543 171
rect 509 103 543 115
rect 509 81 543 103
rect 509 35 543 39
rect 509 5 543 35
rect 509 -67 543 -37
rect 509 -71 543 -67
rect 509 -135 543 -113
rect 509 -147 543 -135
rect 509 -203 543 -189
rect 509 -223 543 -203
rect 615 137 649 145
rect 615 111 649 137
rect 615 69 649 73
rect 615 39 649 69
rect 615 -33 649 1
rect 615 -101 649 -71
rect 615 -105 649 -101
rect 615 -169 649 -143
rect 615 -177 649 -169
rect 615 -237 649 -215
rect 615 -249 649 -237
rect 615 -305 649 -287
rect 615 -321 649 -305
rect 721 205 755 209
rect 721 175 755 205
rect 721 103 755 130
rect 721 96 755 103
rect 721 35 755 51
rect 721 17 755 35
rect 721 -33 755 -29
rect 721 -63 755 -33
rect 721 -135 755 -109
rect 721 -143 755 -135
rect 721 -203 755 -189
rect 721 -223 755 -203
rect 831 205 865 209
rect 831 175 865 205
rect 831 103 865 130
rect 831 96 865 103
rect 831 35 865 51
rect 831 17 865 35
rect 831 -33 865 -29
rect 831 -63 865 -33
rect 831 -135 865 -109
rect 831 -143 865 -135
rect 831 -203 865 -189
rect 831 -223 865 -203
rect 937 137 971 161
rect 937 127 971 137
rect 937 69 971 74
rect 937 40 971 69
rect 937 -33 971 -13
rect 937 -47 971 -33
rect 937 -135 971 -101
rect 937 -203 971 -189
rect 937 -223 971 -203
rect 1043 205 1077 209
rect 1043 175 1077 205
rect 1043 103 1077 130
rect 1043 96 1077 103
rect 1043 35 1077 51
rect 1043 17 1077 35
rect 1043 -33 1077 -29
rect 1043 -63 1077 -33
rect 1043 -135 1077 -109
rect 1043 -143 1077 -135
rect 1043 -203 1077 -189
rect 1043 -223 1077 -203
rect 1149 103 1183 135
rect 1149 101 1183 103
rect 1149 35 1183 51
rect 1149 17 1183 35
rect 1149 -67 1183 -33
rect 1149 -135 1183 -117
rect 1149 -151 1183 -135
rect 1149 -203 1183 -202
rect 1149 -236 1183 -203
rect 1149 -305 1183 -287
rect 1149 -321 1183 -305
rect 1255 205 1289 209
rect 1255 175 1289 205
rect 1255 103 1289 130
rect 1255 96 1289 103
rect 1255 35 1289 51
rect 1255 17 1289 35
rect 1255 -33 1289 -29
rect 1255 -63 1289 -33
rect 1255 -135 1289 -109
rect 1255 -143 1289 -135
rect 1255 -203 1289 -189
rect 1255 -223 1289 -203
rect 1365 103 1399 135
rect 1365 101 1399 103
rect 1365 35 1399 51
rect 1365 17 1399 35
rect 1365 -67 1399 -33
rect 1365 -135 1399 -117
rect 1365 -151 1399 -135
rect 1365 -203 1399 -202
rect 1365 -236 1399 -203
rect 1365 -305 1399 -287
rect 1365 -321 1399 -305
rect 1471 205 1505 209
rect 1471 175 1505 205
rect 1471 103 1505 130
rect 1471 96 1505 103
rect 1471 35 1505 51
rect 1471 17 1505 35
rect 1471 -33 1505 -29
rect 1471 -63 1505 -33
rect 1471 -135 1505 -109
rect 1471 -143 1505 -135
rect 1471 -203 1505 -189
rect 1471 -223 1505 -203
rect 1577 103 1611 135
rect 1577 101 1611 103
rect 1577 35 1611 51
rect 1577 17 1611 35
rect 1577 -67 1611 -33
rect 1577 -135 1611 -117
rect 1577 -151 1611 -135
rect 1577 -203 1611 -202
rect 1577 -236 1611 -203
rect 1577 -305 1611 -287
rect 1577 -321 1611 -305
rect 1687 205 1721 209
rect 1687 175 1721 205
rect 1687 103 1721 130
rect 1687 96 1721 103
rect 1687 35 1721 51
rect 1687 17 1721 35
rect 1687 -33 1721 -29
rect 1687 -63 1721 -33
rect 1687 -135 1721 -109
rect 1687 -143 1721 -135
rect 1687 -203 1721 -189
rect 1687 -223 1721 -203
rect 1793 137 1827 161
rect 1793 127 1827 137
rect 1793 69 1827 74
rect 1793 40 1827 69
rect 1793 -33 1827 -13
rect 1793 -47 1827 -33
rect 1793 -135 1827 -101
rect 1793 -203 1827 -189
rect 1793 -223 1827 -203
rect 1899 205 1933 209
rect 1899 175 1933 205
rect 1899 103 1933 130
rect 1899 96 1933 103
rect 1899 35 1933 51
rect 1899 17 1933 35
rect 1899 -33 1933 -29
rect 1899 -63 1933 -33
rect 1899 -135 1933 -109
rect 1899 -143 1933 -135
rect 1899 -203 1933 -189
rect 1899 -223 1933 -203
rect 2005 103 2039 135
rect 2005 101 2039 103
rect 2005 35 2039 51
rect 2005 17 2039 35
rect 2005 -67 2039 -33
rect 2005 -135 2039 -117
rect 2005 -151 2039 -135
rect 2005 -203 2039 -202
rect 2005 -236 2039 -203
rect 2005 -305 2039 -287
rect 2005 -321 2039 -305
rect 2111 205 2145 209
rect 2111 175 2145 205
rect 2111 103 2145 130
rect 2111 96 2145 103
rect 2111 35 2145 51
rect 2111 17 2145 35
rect 2111 -33 2145 -29
rect 2111 -63 2145 -33
rect 2111 -135 2145 -109
rect 2111 -143 2145 -135
rect 2111 -203 2145 -189
rect 2111 -223 2145 -203
rect 501 -431 525 -397
rect 525 -431 535 -397
rect 575 -431 594 -397
rect 594 -431 609 -397
rect 649 -431 663 -397
rect 663 -431 683 -397
rect 723 -431 732 -397
rect 732 -431 757 -397
rect 797 -431 801 -397
rect 801 -431 831 -397
rect 871 -431 904 -397
rect 904 -431 905 -397
rect 945 -431 973 -397
rect 973 -431 979 -397
rect 1019 -431 1041 -397
rect 1041 -431 1053 -397
rect 1093 -431 1109 -397
rect 1109 -431 1127 -397
rect 1167 -431 1177 -397
rect 1177 -431 1201 -397
rect 1241 -431 1245 -397
rect 1245 -431 1275 -397
rect 1315 -431 1347 -397
rect 1347 -431 1349 -397
rect 1388 -431 1415 -397
rect 1415 -431 1422 -397
rect 1461 -431 1483 -397
rect 1483 -431 1495 -397
rect 1534 -431 1551 -397
rect 1551 -431 1568 -397
rect 1607 -431 1619 -397
rect 1619 -431 1641 -397
rect 1680 -431 1687 -397
rect 1687 -431 1714 -397
rect 1753 -431 1755 -397
rect 1755 -431 1787 -397
rect 1826 -431 1857 -397
rect 1857 -431 1860 -397
rect 1899 -431 1925 -397
rect 1925 -431 1933 -397
rect 1972 -431 1993 -397
rect 1993 -431 2006 -397
rect 2045 -431 2061 -397
rect 2061 -431 2079 -397
rect 2118 -431 2129 -397
rect 2129 -431 2152 -397
<< metal1 >>
rect 145 3462 2336 3529
rect 145 3428 157 3462
rect 191 3428 231 3462
rect 265 3428 305 3462
rect 339 3428 379 3462
rect 413 3428 453 3462
rect 487 3428 527 3462
rect 561 3428 601 3462
rect 635 3428 675 3462
rect 709 3428 749 3462
rect 783 3428 823 3462
rect 857 3428 897 3462
rect 931 3428 971 3462
rect 1005 3428 1045 3462
rect 1079 3428 1119 3462
rect 1153 3428 1193 3462
rect 1227 3428 1267 3462
rect 1301 3428 1341 3462
rect 1375 3428 1415 3462
rect 1449 3428 1489 3462
rect 1523 3428 1563 3462
rect 1597 3428 1637 3462
rect 1671 3428 1711 3462
rect 1745 3428 1785 3462
rect 1819 3428 1858 3462
rect 1892 3428 1914 3462
rect 1966 3428 2004 3462
rect 2038 3428 2077 3462
rect 2111 3428 2150 3462
rect 2184 3428 2223 3462
rect 2257 3428 2336 3462
rect 145 3410 1914 3428
rect 1966 3410 2336 3428
rect 145 3394 2336 3410
rect 145 3342 1914 3394
rect 1966 3342 2336 3394
rect 145 3308 228 3342
rect 262 3308 762 3342
rect 796 3308 978 3342
rect 1012 3308 1190 3342
rect 1224 3308 1402 3342
rect 1436 3308 1618 3342
rect 1652 3326 2258 3342
rect 1652 3308 1914 3326
rect 145 3274 1914 3308
rect 1966 3308 2258 3326
rect 2292 3308 2336 3342
rect 1966 3274 2336 3308
rect 145 3269 2336 3274
rect 145 3268 978 3269
tri 188 3266 190 3268 ne
rect 190 3266 290 3268
tri 190 3234 222 3266 ne
rect 222 3232 228 3266
rect 262 3256 290 3266
tri 290 3256 302 3268 nw
tri 722 3256 734 3268 ne
rect 734 3256 803 3268
rect 262 3236 270 3256
tri 270 3236 290 3256 nw
tri 734 3236 754 3256 ne
rect 754 3236 762 3256
rect 262 3232 268 3236
tri 268 3234 270 3236 nw
rect 116 3188 162 3200
rect 116 3154 122 3188
rect 156 3154 162 3188
rect 116 3115 162 3154
rect 116 3081 122 3115
rect 156 3081 162 3115
rect 116 3042 162 3081
rect 116 3008 122 3042
rect 156 3008 162 3042
rect 116 2969 162 3008
rect 116 2935 122 2969
rect 156 2935 162 2969
rect 116 2896 162 2935
rect 116 2862 122 2896
rect 156 2862 162 2896
rect 116 2823 162 2862
rect 116 2789 122 2823
rect 156 2789 162 2823
rect 116 2749 162 2789
rect 116 2715 122 2749
rect 156 2715 162 2749
rect 116 2675 162 2715
rect 116 2641 122 2675
rect 156 2641 162 2675
rect 116 2601 162 2641
rect 116 2567 122 2601
rect 156 2567 162 2601
rect 116 2527 162 2567
rect 116 2493 122 2527
rect 156 2493 162 2527
rect 116 2453 162 2493
rect 222 3190 268 3232
rect 541 3224 593 3236
tri 754 3234 756 3236 ne
rect 222 3156 228 3190
rect 262 3156 268 3190
rect 222 3114 268 3156
rect 222 3080 228 3114
rect 262 3080 268 3114
rect 222 3038 268 3080
rect 222 3004 228 3038
rect 262 3004 268 3038
rect 222 2961 268 3004
rect 222 2927 228 2961
rect 262 2927 268 2961
rect 222 2884 268 2927
rect 222 2850 228 2884
rect 262 2850 268 2884
rect 222 2807 268 2850
rect 222 2773 228 2807
rect 262 2773 268 2807
rect 222 2730 268 2773
rect 222 2696 228 2730
rect 262 2696 268 2730
rect 222 2653 268 2696
rect 222 2619 228 2653
rect 262 2619 268 2653
rect 222 2576 268 2619
rect 222 2542 228 2576
rect 262 2542 268 2576
rect 222 2499 268 2542
rect 222 2465 228 2499
rect 262 2465 268 2499
tri 162 2453 163 2454 sw
rect 222 2453 268 2465
rect 325 3188 377 3200
rect 325 3154 334 3188
rect 368 3154 377 3188
rect 325 3112 377 3154
rect 325 3078 334 3112
rect 368 3078 377 3112
rect 325 3036 377 3078
rect 325 3002 334 3036
rect 368 3002 377 3036
rect 325 2960 377 3002
rect 325 2926 334 2960
rect 368 2926 377 2960
rect 325 2884 377 2926
rect 325 2850 334 2884
rect 368 2850 377 2884
rect 325 2807 377 2850
rect 325 2773 334 2807
rect 368 2773 377 2807
rect 325 2730 377 2773
rect 438 3190 484 3202
rect 438 3156 444 3190
rect 478 3156 484 3190
rect 438 3112 484 3156
rect 438 3078 444 3112
rect 478 3078 484 3112
rect 438 3034 484 3078
rect 438 3000 444 3034
rect 478 3000 484 3034
rect 438 2956 484 3000
rect 438 2922 444 2956
rect 478 2922 484 2956
rect 438 2878 484 2922
rect 438 2844 444 2878
rect 478 2865 484 2878
rect 541 3190 550 3224
rect 584 3190 593 3224
rect 756 3222 762 3236
rect 796 3235 803 3256
tri 803 3235 836 3268 nw
tri 938 3235 971 3268 ne
rect 971 3235 978 3268
rect 1012 3268 1190 3269
rect 1012 3235 1019 3268
tri 1019 3235 1052 3268 nw
tri 1150 3235 1183 3268 ne
rect 1183 3235 1190 3268
rect 1224 3268 1402 3269
rect 1224 3235 1231 3268
tri 1231 3235 1264 3268 nw
tri 1362 3235 1395 3268 ne
rect 1395 3235 1402 3268
rect 1436 3268 2258 3269
rect 1436 3256 1464 3268
tri 1464 3256 1476 3268 nw
tri 1578 3256 1590 3268 ne
rect 1590 3256 1660 3268
rect 1436 3235 1442 3256
rect 796 3222 802 3235
tri 802 3234 803 3235 nw
tri 971 3234 972 3235 ne
rect 541 3146 593 3190
rect 541 3112 550 3146
rect 584 3112 593 3146
rect 541 3068 593 3112
rect 541 3034 550 3068
rect 584 3034 593 3068
rect 541 2990 593 3034
rect 541 2987 550 2990
rect 584 2987 593 2990
rect 541 2923 593 2935
tri 484 2865 487 2868 sw
rect 541 2865 593 2871
rect 650 3190 696 3202
rect 650 3156 656 3190
rect 690 3156 696 3190
rect 650 3112 696 3156
rect 650 3078 656 3112
rect 690 3078 696 3112
rect 650 3034 696 3078
rect 650 3000 656 3034
rect 690 3000 696 3034
rect 650 2956 696 3000
rect 650 2922 656 2956
rect 690 2922 696 2956
rect 650 2878 696 2922
tri 647 2865 650 2868 se
rect 650 2865 656 2878
rect 478 2844 487 2865
tri 487 2844 508 2865 sw
tri 626 2844 647 2865 se
rect 647 2844 656 2865
rect 690 2866 696 2878
rect 756 3170 802 3222
rect 756 3136 762 3170
rect 796 3136 802 3170
rect 756 3084 802 3136
rect 756 3050 762 3084
rect 796 3050 802 3084
rect 756 2998 802 3050
rect 756 2964 762 2998
rect 796 2964 802 2998
rect 756 2912 802 2964
rect 756 2878 762 2912
rect 796 2878 802 2912
tri 696 2866 698 2868 sw
rect 756 2866 802 2878
rect 862 3190 908 3202
rect 862 3156 868 3190
rect 902 3156 908 3190
rect 862 3112 908 3156
rect 862 3078 868 3112
rect 902 3078 908 3112
rect 862 3034 908 3078
rect 862 3000 868 3034
rect 902 3000 908 3034
rect 862 2956 908 3000
rect 862 2922 868 2956
rect 902 2922 908 2956
rect 862 2878 908 2922
tri 860 2866 862 2868 se
rect 862 2866 868 2878
rect 690 2844 698 2866
tri 698 2844 720 2866 sw
tri 838 2844 860 2866 se
rect 860 2844 868 2866
rect 902 2844 908 2878
rect 972 3196 1018 3235
tri 1018 3234 1019 3235 nw
tri 1183 3234 1184 3235 ne
rect 972 3162 978 3196
rect 1012 3162 1018 3196
rect 972 3123 1018 3162
rect 972 3089 978 3123
rect 1012 3089 1018 3123
rect 972 3049 1018 3089
rect 972 3015 978 3049
rect 1012 3015 1018 3049
rect 972 2975 1018 3015
rect 972 2941 978 2975
rect 1012 2941 1018 2975
rect 972 2901 1018 2941
rect 972 2867 978 2901
rect 1012 2867 1018 2901
rect 972 2855 1018 2867
rect 1078 3190 1124 3202
rect 1078 3156 1084 3190
rect 1118 3156 1124 3190
rect 1078 3112 1124 3156
rect 1078 3078 1084 3112
rect 1118 3078 1124 3112
rect 1078 3034 1124 3078
rect 1078 3000 1084 3034
rect 1118 3000 1124 3034
rect 1078 2956 1124 3000
rect 1078 2922 1084 2956
rect 1118 2922 1124 2956
rect 1078 2878 1124 2922
rect 438 2834 508 2844
tri 508 2834 518 2844 sw
tri 616 2834 626 2844 se
rect 626 2834 720 2844
tri 720 2834 730 2844 sw
tri 828 2834 838 2844 se
rect 838 2834 908 2844
rect 438 2800 908 2834
rect 438 2766 444 2800
rect 478 2766 656 2800
rect 690 2766 868 2800
rect 902 2766 908 2800
rect 438 2754 908 2766
rect 1078 2844 1084 2878
rect 1118 2855 1124 2878
rect 1184 3196 1230 3235
tri 1230 3234 1231 3235 nw
tri 1395 3234 1396 3235 ne
rect 1184 3162 1190 3196
rect 1224 3162 1230 3196
rect 1184 3123 1230 3162
rect 1184 3089 1190 3123
rect 1224 3089 1230 3123
rect 1184 3049 1230 3089
rect 1184 3015 1190 3049
rect 1224 3015 1230 3049
rect 1184 2975 1230 3015
rect 1184 2941 1190 2975
rect 1224 2941 1230 2975
rect 1184 2901 1230 2941
rect 1184 2867 1190 2901
rect 1224 2867 1230 2901
tri 1124 2855 1126 2857 sw
rect 1184 2855 1230 2867
rect 1290 3190 1336 3202
rect 1290 3156 1296 3190
rect 1330 3156 1336 3190
rect 1290 3112 1336 3156
rect 1290 3078 1296 3112
rect 1330 3078 1336 3112
rect 1290 3034 1336 3078
rect 1290 3000 1296 3034
rect 1330 3000 1336 3034
rect 1290 2956 1336 3000
rect 1290 2922 1296 2956
rect 1330 2922 1336 2956
rect 1290 2878 1336 2922
tri 1288 2855 1290 2857 se
rect 1290 2855 1296 2878
rect 1118 2844 1126 2855
tri 1126 2844 1137 2855 sw
tri 1277 2844 1288 2855 se
rect 1288 2844 1296 2855
rect 1330 2844 1336 2878
rect 1396 3196 1442 3235
tri 1442 3234 1464 3256 nw
tri 1590 3234 1612 3256 ne
rect 1612 3222 1618 3256
rect 1652 3236 1660 3256
tri 1660 3236 1692 3268 nw
tri 2218 3236 2250 3268 ne
rect 2250 3236 2258 3268
rect 1652 3235 1659 3236
tri 1659 3235 1660 3236 nw
rect 1652 3222 1658 3235
tri 1658 3234 1659 3235 nw
rect 1396 3162 1402 3196
rect 1436 3162 1442 3196
rect 1396 3123 1442 3162
rect 1396 3089 1402 3123
rect 1436 3089 1442 3123
rect 1396 3049 1442 3089
rect 1396 3015 1402 3049
rect 1436 3015 1442 3049
rect 1396 2975 1442 3015
rect 1396 2941 1402 2975
rect 1436 2941 1442 2975
rect 1396 2901 1442 2941
rect 1396 2867 1402 2901
rect 1436 2867 1442 2901
rect 1396 2855 1442 2867
rect 1506 3190 1552 3202
rect 1506 3156 1512 3190
rect 1546 3156 1552 3190
rect 1506 3112 1552 3156
rect 1506 3078 1512 3112
rect 1546 3078 1552 3112
rect 1506 3034 1552 3078
rect 1506 3000 1512 3034
rect 1546 3000 1552 3034
rect 1506 2956 1552 3000
rect 1506 2922 1512 2956
rect 1546 2922 1552 2956
rect 1506 2878 1552 2922
rect 1078 2823 1137 2844
tri 1137 2823 1158 2844 sw
tri 1256 2823 1277 2844 se
rect 1277 2823 1336 2844
rect 1078 2806 1336 2823
rect 1078 2754 1084 2806
rect 1136 2754 1149 2806
rect 1201 2754 1214 2806
rect 1266 2754 1278 2806
rect 1330 2754 1336 2806
rect 1506 2844 1512 2878
rect 1546 2866 1552 2878
rect 1612 3170 1658 3222
rect 1821 3224 1873 3236
tri 2250 3235 2251 3236 ne
rect 2251 3235 2258 3236
rect 2292 3268 2336 3269
rect 2292 3235 2298 3268
tri 2251 3234 2252 3235 ne
rect 1612 3136 1618 3170
rect 1652 3136 1658 3170
rect 1612 3084 1658 3136
rect 1612 3050 1618 3084
rect 1652 3050 1658 3084
rect 1612 2998 1658 3050
rect 1612 2964 1618 2998
rect 1652 2964 1658 2998
rect 1612 2912 1658 2964
rect 1612 2878 1618 2912
rect 1652 2878 1658 2912
tri 1552 2866 1554 2868 sw
rect 1612 2866 1658 2878
rect 1718 3190 1764 3202
rect 1718 3156 1724 3190
rect 1758 3156 1764 3190
rect 1718 3112 1764 3156
rect 1718 3078 1724 3112
rect 1758 3078 1764 3112
rect 1718 3034 1764 3078
rect 1718 3000 1724 3034
rect 1758 3000 1764 3034
rect 1718 2956 1764 3000
rect 1718 2922 1724 2956
rect 1758 2922 1764 2956
rect 1718 2878 1764 2922
tri 1716 2866 1718 2868 se
rect 1718 2866 1724 2878
rect 1546 2844 1554 2866
tri 1554 2844 1576 2866 sw
tri 1694 2844 1716 2866 se
rect 1716 2844 1724 2866
rect 1758 2866 1764 2878
rect 1821 3190 1830 3224
rect 1864 3190 1873 3224
rect 1821 3146 1873 3190
rect 1821 3112 1830 3146
rect 1864 3112 1873 3146
rect 1821 3068 1873 3112
rect 1821 3034 1830 3068
rect 1864 3034 1873 3068
rect 1821 2990 1873 3034
rect 1821 2988 1830 2990
rect 1864 2988 1873 2990
rect 1821 2924 1873 2936
tri 1764 2866 1766 2868 sw
rect 1821 2866 1873 2872
rect 1930 3190 1976 3202
rect 1930 3156 1936 3190
rect 1970 3156 1976 3190
rect 1930 3112 1976 3156
rect 1930 3078 1936 3112
rect 1970 3078 1976 3112
rect 1930 3034 1976 3078
rect 1930 3000 1936 3034
rect 1970 3000 1976 3034
rect 1930 2956 1976 3000
rect 1930 2922 1936 2956
rect 1970 2922 1976 2956
rect 1930 2878 1976 2922
tri 1928 2866 1930 2868 se
rect 1930 2866 1936 2878
rect 1758 2844 1766 2866
tri 1766 2844 1788 2866 sw
tri 1906 2844 1928 2866 se
rect 1928 2844 1936 2866
rect 1970 2844 1976 2878
rect 1506 2834 1576 2844
tri 1576 2834 1586 2844 sw
tri 1684 2834 1694 2844 se
rect 1694 2834 1788 2844
tri 1788 2834 1798 2844 sw
tri 1896 2834 1906 2844 se
rect 1906 2834 1976 2844
rect 1506 2800 1976 2834
rect 1506 2766 1512 2800
rect 1546 2766 1724 2800
rect 1758 2766 1936 2800
rect 1970 2766 1976 2800
rect 1506 2754 1976 2766
rect 2037 3190 2089 3202
rect 2037 3156 2046 3190
rect 2080 3156 2089 3190
rect 2037 3112 2089 3156
rect 2037 3078 2046 3112
rect 2080 3078 2089 3112
rect 2037 3034 2089 3078
rect 2037 3000 2046 3034
rect 2080 3000 2089 3034
rect 2037 2982 2089 3000
rect 2037 2922 2046 2930
rect 2080 2922 2089 2930
rect 2037 2918 2089 2922
rect 2037 2844 2046 2866
rect 2080 2844 2089 2866
rect 2037 2800 2089 2844
rect 2037 2766 2046 2800
rect 2080 2766 2089 2800
rect 2037 2754 2089 2766
rect 2146 3190 2192 3202
rect 2146 3156 2152 3190
rect 2186 3156 2192 3190
rect 2146 3112 2192 3156
rect 2146 3078 2152 3112
rect 2186 3078 2192 3112
rect 2146 3034 2192 3078
rect 2146 3000 2152 3034
rect 2186 3000 2192 3034
rect 2146 2956 2192 3000
rect 2146 2922 2152 2956
rect 2186 2922 2192 2956
rect 2146 2878 2192 2922
rect 2146 2844 2152 2878
rect 2186 2844 2192 2878
rect 2252 3196 2298 3235
tri 2298 3234 2332 3268 nw
rect 2252 3162 2258 3196
rect 2292 3162 2298 3196
rect 2252 3123 2298 3162
rect 2252 3089 2258 3123
rect 2292 3089 2298 3123
rect 2252 3049 2298 3089
rect 2252 3015 2258 3049
rect 2292 3015 2298 3049
rect 2252 2975 2298 3015
rect 2252 2941 2258 2975
rect 2292 2941 2298 2975
rect 2252 2901 2298 2941
rect 2252 2867 2258 2901
rect 2292 2867 2298 2901
rect 2252 2855 2298 2867
rect 2146 2800 2192 2844
rect 2146 2766 2152 2800
rect 2186 2766 2192 2800
rect 2146 2754 2192 2766
rect 325 2706 334 2730
rect 368 2715 377 2730
tri 377 2715 408 2746 sw
rect 368 2712 408 2715
tri 408 2712 411 2715 sw
rect 368 2706 618 2712
rect 377 2672 500 2706
rect 534 2672 572 2706
rect 606 2672 618 2706
rect 377 2666 618 2672
rect 377 2663 408 2666
tri 408 2663 411 2666 nw
rect 727 2663 735 2715
rect 787 2663 799 2715
rect 851 2663 857 2715
rect 1033 2706 1173 2715
rect 1225 2706 1237 2715
rect 1289 2706 1377 2715
rect 1033 2672 1045 2706
rect 1079 2672 1141 2706
rect 1225 2672 1236 2706
rect 1289 2672 1331 2706
rect 1365 2672 1377 2706
rect 1033 2663 1173 2672
rect 1225 2663 1237 2672
rect 1289 2663 1377 2672
rect 1565 2663 1571 2715
rect 1623 2663 1635 2715
rect 1687 2663 1695 2715
rect 1735 2706 1900 2712
rect 1816 2672 1854 2706
rect 1888 2672 1900 2706
rect 377 2654 395 2663
rect 325 2653 395 2654
rect 325 2642 334 2653
rect 368 2650 395 2653
tri 395 2650 408 2663 nw
rect 1787 2666 1900 2672
rect 2083 2688 2135 2696
rect 1787 2654 1805 2666
rect 1735 2650 1805 2654
tri 1805 2650 1821 2666 nw
rect 368 2642 377 2650
tri 377 2632 395 2650 nw
rect 1735 2642 1787 2650
rect 325 2576 377 2590
tri 1787 2632 1805 2650 nw
rect 1735 2584 1787 2590
rect 2083 2624 2135 2636
rect 325 2542 334 2576
rect 368 2542 377 2576
rect 2083 2566 2135 2572
rect 2204 2688 2256 2696
rect 2204 2624 2256 2636
rect 2204 2566 2256 2572
rect 325 2499 377 2542
rect 325 2465 334 2499
rect 368 2465 377 2499
rect 325 2453 377 2465
rect 541 2529 2278 2530
rect 541 2477 547 2529
rect 599 2477 611 2529
rect 663 2524 2278 2529
rect 663 2505 1642 2524
rect 663 2477 1054 2505
rect 541 2453 1054 2477
rect 1106 2453 1118 2505
rect 1170 2472 1642 2505
rect 1694 2472 1821 2524
rect 1873 2472 2003 2524
rect 2055 2472 2278 2524
rect 1170 2460 2278 2472
rect 1170 2453 1642 2460
rect 116 2420 163 2453
tri 163 2420 196 2453 sw
rect 116 2417 266 2420
tri 266 2417 269 2420 sw
rect 116 2374 269 2417
tri 269 2374 312 2417 sw
rect 541 2408 1642 2453
rect 1694 2408 1821 2460
rect 1873 2408 2003 2460
rect 2055 2408 2278 2460
rect 541 2402 2278 2408
tri 246 2351 269 2374 ne
rect 269 2351 312 2374
tri 312 2351 335 2374 sw
tri 269 2337 283 2351 ne
rect 158 2310 210 2322
rect 158 2246 210 2258
rect 158 2188 210 2194
rect 283 2310 335 2351
rect 283 2246 335 2258
rect 834 2236 1975 2242
rect 834 2202 846 2236
rect 880 2202 921 2236
rect 955 2202 996 2236
rect 1030 2202 1071 2236
rect 1105 2202 1146 2236
rect 1180 2202 1221 2236
rect 1255 2202 1295 2236
rect 1329 2202 1369 2236
rect 1403 2202 1443 2236
rect 1477 2202 1517 2236
rect 1551 2202 1591 2236
rect 1625 2202 1665 2236
rect 1699 2202 1739 2236
rect 1773 2230 1914 2236
rect 1773 2202 1855 2230
rect 834 2196 1855 2202
rect 1889 2196 1914 2230
rect 283 2188 335 2194
tri 1680 2191 1685 2196 ne
rect 1685 2191 1914 2196
rect 692 2179 738 2191
rect 692 2145 698 2179
rect 732 2145 738 2179
tri 1685 2162 1714 2191 ne
rect 1714 2184 1914 2191
rect 1966 2184 1975 2236
tri 675 2080 692 2097 se
rect 692 2080 738 2145
rect 1714 2155 1975 2184
rect 1714 2121 1855 2155
rect 1889 2138 1975 2155
rect 1889 2121 1914 2138
tri 658 2063 675 2080 se
rect 675 2063 698 2080
rect 482 2057 698 2063
rect 534 2046 698 2057
rect 732 2046 738 2080
rect 534 2005 738 2046
rect 834 2080 1207 2089
rect 1259 2080 1271 2089
rect 1323 2080 1676 2089
rect 834 2046 846 2080
rect 880 2046 925 2080
rect 959 2046 1004 2080
rect 1038 2046 1083 2080
rect 1117 2046 1162 2080
rect 1196 2046 1207 2080
rect 1352 2046 1396 2080
rect 1430 2046 1474 2080
rect 1508 2046 1552 2080
rect 1586 2046 1630 2080
rect 1664 2046 1676 2080
rect 834 2037 1207 2046
rect 1259 2037 1271 2046
rect 1323 2037 1676 2046
rect 1714 2086 1914 2121
rect 1966 2086 1975 2138
rect 1714 2080 1975 2086
rect 1714 2046 1855 2080
rect 1889 2046 1975 2080
rect 1714 2040 1975 2046
rect 482 1993 738 2005
rect 534 1981 738 1993
rect 534 1947 698 1981
rect 732 1947 738 1981
rect 1714 2005 1914 2040
rect 1714 1971 1855 2005
rect 1889 1988 1914 2005
rect 1966 1988 1975 2040
rect 1889 1971 1975 1988
rect 534 1941 738 1947
rect 482 1935 738 1941
tri 1683 1935 1714 1966 se
rect 1714 1942 1975 1971
rect 1714 1935 1914 1942
tri 1680 1932 1683 1935 se
rect 1683 1932 1914 1935
rect 834 1930 1914 1932
rect 834 1926 1855 1930
rect 834 1892 846 1926
rect 880 1892 921 1926
rect 955 1892 996 1926
rect 1030 1892 1071 1926
rect 1105 1892 1146 1926
rect 1180 1892 1221 1926
rect 1255 1892 1295 1926
rect 1329 1892 1369 1926
rect 1403 1892 1443 1926
rect 1477 1892 1517 1926
rect 1551 1892 1591 1926
rect 1625 1892 1665 1926
rect 1699 1892 1739 1926
rect 1773 1896 1855 1926
rect 1889 1896 1914 1930
rect 1773 1892 1914 1896
rect 834 1890 1914 1892
rect 1966 1890 1975 1942
rect 834 1886 1975 1890
rect 1714 1884 1975 1886
rect 283 1726 289 1778
rect 341 1726 353 1778
rect 405 1726 1207 1778
rect 1259 1726 1271 1778
rect 1323 1726 1329 1778
rect 124 1646 130 1698
rect 182 1646 194 1698
rect 246 1646 694 1698
rect 746 1646 758 1698
rect 810 1646 1259 1698
rect 1311 1646 1323 1698
rect 1375 1646 2013 1698
rect 2065 1646 2077 1698
rect 2129 1646 2135 1698
rect 844 1566 850 1618
rect 902 1566 914 1618
rect 966 1566 972 1618
rect 260 1486 1395 1538
rect 1447 1486 1459 1538
rect 1511 1486 1703 1538
rect 260 1458 1703 1486
rect 260 1424 1597 1430
rect 260 1378 1545 1424
tri 1511 1344 1545 1378 ne
rect 1545 1360 1597 1372
rect 1545 1302 1597 1308
rect 260 1122 1741 1174
rect 1793 1122 1805 1174
rect 1857 1122 1903 1174
rect 260 1042 2134 1094
rect 2186 1042 2198 1094
rect 2250 1042 2256 1094
rect 406 894 412 946
rect 464 894 476 946
rect 528 894 2146 946
rect 566 819 824 825
rect 618 773 824 819
rect 876 773 888 825
rect 940 773 946 825
rect 566 755 618 767
rect 566 697 618 703
rect 551 447 603 453
tri 520 374 551 405 se
rect 551 383 603 395
rect 216 365 248 374
rect 300 365 312 374
rect 216 331 228 365
rect 216 323 248 331
rect 242 322 248 323
rect 300 322 312 331
rect 364 322 370 374
tri 517 371 520 374 se
rect 520 371 551 374
rect 465 365 551 371
rect 465 331 477 365
rect 511 331 549 365
rect 465 325 603 331
rect 660 365 790 371
rect 660 331 672 365
rect 706 331 744 365
rect 778 331 790 365
rect 660 325 790 331
rect 660 322 743 325
tri 743 322 746 325 nw
rect 818 322 824 374
rect 876 322 888 374
rect 940 365 1015 374
rect 940 331 969 365
rect 1003 331 1015 365
rect 940 322 1015 331
rect 1106 365 1122 374
rect 1106 331 1118 365
rect 1106 322 1122 331
rect 1174 322 1186 374
rect 1238 322 1244 374
rect 1426 322 1435 374
rect 1487 322 1499 374
rect 1551 322 1557 374
rect 1751 365 1781 374
rect 1833 365 1845 374
rect 1751 331 1763 365
rect 1833 331 1835 365
rect 1751 322 1781 331
rect 1833 322 1845 331
rect 1897 322 1903 374
rect 1970 322 1978 374
rect 2030 322 2042 374
rect 2094 322 2100 374
tri 626 283 660 317 se
rect 660 283 712 322
tri 712 291 743 322 nw
rect 162 279 712 283
rect 162 249 682 279
tri 682 249 712 279 nw
rect 162 238 671 249
tri 671 238 682 249 nw
rect 162 237 664 238
rect 162 232 171 237
rect 205 232 664 237
rect 214 231 664 232
tri 664 231 671 238 nw
rect 214 221 238 231
tri 238 221 248 231 nw
rect 214 209 226 221
tri 226 209 238 221 nw
rect 712 215 764 221
rect 214 203 220 209
tri 220 203 226 209 nw
tri 214 197 220 203 nw
rect 162 168 214 180
rect 162 99 171 116
rect 205 99 214 116
rect 162 29 214 99
rect 162 -5 171 29
rect 205 -5 214 29
rect 162 -17 214 -5
rect 321 191 549 203
rect 321 157 327 191
rect 361 157 509 191
rect 543 157 549 191
rect 321 115 549 157
rect 321 110 509 115
rect 321 76 327 110
rect 361 81 509 110
rect 543 81 549 115
rect 361 76 549 81
rect 321 39 549 76
rect 321 29 509 39
rect 321 -5 327 29
rect 361 5 509 29
rect 543 5 549 39
rect 361 -5 549 5
rect 321 -17 549 -5
tri 469 -33 485 -17 ne
rect 485 -33 549 -17
tri 485 -37 489 -33 ne
rect 489 -37 549 -33
tri 489 -51 503 -37 ne
rect 503 -71 509 -37
rect 543 -71 549 -37
rect 503 -113 549 -71
rect 503 -147 509 -113
rect 543 -147 549 -113
rect 503 -189 549 -147
rect 503 -223 509 -189
rect 543 -223 549 -189
rect 503 -235 549 -223
rect 609 145 655 157
rect 609 111 615 145
rect 649 111 655 145
rect 609 73 655 111
rect 609 39 615 73
rect 649 39 655 73
rect 609 1 655 39
rect 609 -33 615 1
rect 649 -33 655 1
rect 609 -71 655 -33
rect 609 -105 615 -71
rect 649 -105 655 -71
rect 609 -143 655 -105
rect 609 -177 615 -143
rect 649 -177 655 -143
rect 609 -215 655 -177
tri 602 -249 609 -242 se
rect 609 -249 615 -215
rect 649 -249 655 -215
rect 712 151 764 163
rect 712 96 721 99
rect 755 96 764 99
rect 712 51 764 96
rect 712 17 721 51
rect 755 17 764 51
rect 712 -29 764 17
rect 712 -63 721 -29
rect 755 -63 764 -29
rect 712 -109 764 -63
rect 712 -143 721 -109
rect 755 -143 764 -109
rect 712 -189 764 -143
rect 712 -223 721 -189
rect 755 -223 764 -189
rect 712 -235 764 -223
rect 825 209 1295 283
rect 825 175 831 209
rect 865 203 1043 209
rect 865 175 877 203
tri 877 175 905 203 nw
tri 1003 175 1031 203 ne
rect 1031 175 1043 203
rect 1077 203 1255 209
rect 1077 175 1089 203
tri 1089 175 1117 203 nw
tri 1215 175 1243 203 ne
rect 1243 175 1255 203
rect 1289 175 1295 209
rect 825 173 875 175
tri 875 173 877 175 nw
tri 1031 173 1033 175 ne
rect 1033 173 1083 175
rect 825 130 871 173
tri 871 169 875 173 nw
rect 825 96 831 130
rect 865 96 871 130
rect 825 51 871 96
rect 825 17 831 51
rect 865 17 871 51
rect 825 -29 871 17
rect 825 -63 831 -29
rect 865 -63 871 -29
rect 825 -109 871 -63
rect 825 -143 831 -109
rect 865 -143 871 -109
rect 825 -189 871 -143
rect 825 -223 831 -189
rect 865 -223 871 -189
rect 825 -235 871 -223
rect 928 163 980 173
tri 1033 169 1037 173 ne
rect 928 99 980 111
rect 928 40 937 47
rect 971 40 980 47
rect 928 -13 980 40
rect 928 -47 937 -13
rect 971 -47 980 -13
rect 928 -101 980 -47
rect 928 -135 937 -101
rect 971 -135 980 -101
rect 928 -189 980 -135
rect 928 -223 937 -189
rect 971 -223 980 -189
rect 928 -235 980 -223
rect 1037 130 1083 173
tri 1083 169 1089 175 nw
tri 1243 169 1249 175 ne
rect 1037 96 1043 130
rect 1077 96 1083 130
rect 1037 51 1083 96
rect 1037 17 1043 51
rect 1077 17 1083 51
rect 1037 -29 1083 17
rect 1037 -63 1043 -29
rect 1077 -63 1083 -29
rect 1037 -109 1083 -63
rect 1037 -143 1043 -109
rect 1077 -143 1083 -109
rect 1037 -189 1083 -143
rect 1037 -223 1043 -189
rect 1077 -223 1083 -189
rect 1037 -235 1083 -223
rect 1143 135 1189 147
rect 1143 101 1149 135
rect 1183 101 1189 135
rect 1143 51 1189 101
rect 1143 17 1149 51
rect 1183 17 1189 51
rect 1143 -33 1189 17
rect 1143 -67 1149 -33
rect 1183 -67 1189 -33
rect 1143 -117 1189 -67
rect 1143 -151 1149 -117
rect 1183 -151 1189 -117
rect 1143 -202 1189 -151
rect 1143 -236 1149 -202
rect 1183 -236 1189 -202
rect 1249 130 1295 175
rect 1462 209 1514 221
rect 1462 175 1471 209
rect 1505 175 1514 209
rect 1249 96 1255 130
rect 1289 96 1295 130
rect 1249 51 1295 96
rect 1249 17 1255 51
rect 1289 17 1295 51
rect 1249 -29 1295 17
rect 1249 -63 1255 -29
rect 1289 -63 1295 -29
rect 1249 -109 1295 -63
rect 1249 -143 1255 -109
rect 1289 -143 1295 -109
rect 1249 -189 1295 -143
rect 1249 -223 1255 -189
rect 1289 -223 1295 -189
rect 1249 -235 1295 -223
rect 1359 135 1405 147
rect 1359 101 1365 135
rect 1399 101 1405 135
rect 1359 51 1405 101
rect 1359 17 1365 51
rect 1399 17 1405 51
rect 1359 -33 1405 17
rect 1359 -67 1365 -33
rect 1399 -67 1405 -33
rect 1359 -117 1405 -67
rect 1359 -151 1365 -117
rect 1399 -151 1405 -117
rect 1359 -202 1405 -151
tri 575 -276 602 -249 se
rect 602 -276 655 -249
tri 655 -276 689 -242 sw
tri 1109 -276 1143 -242 se
rect 1143 -276 1189 -236
rect 1359 -236 1365 -202
rect 1399 -236 1405 -202
rect 1462 130 1514 175
rect 1681 209 2151 283
rect 1681 175 1687 209
rect 1721 203 1899 209
rect 1721 175 1733 203
tri 1733 175 1761 203 nw
tri 1859 175 1887 203 ne
rect 1887 175 1899 203
rect 1933 203 2111 209
rect 1933 175 1945 203
tri 1945 175 1973 203 nw
tri 2071 175 2099 203 ne
rect 2099 175 2111 203
rect 2145 175 2151 209
rect 1681 173 1731 175
tri 1731 173 1733 175 nw
tri 1887 173 1889 175 ne
rect 1889 173 1939 175
rect 1462 129 1471 130
rect 1505 129 1514 130
rect 1462 65 1514 77
rect 1462 -29 1514 13
rect 1462 -63 1471 -29
rect 1505 -63 1514 -29
rect 1462 -109 1514 -63
rect 1462 -143 1471 -109
rect 1505 -143 1514 -109
rect 1462 -189 1514 -143
rect 1462 -223 1471 -189
rect 1505 -223 1514 -189
rect 1462 -235 1514 -223
rect 1571 135 1617 147
rect 1571 101 1577 135
rect 1611 101 1617 135
rect 1571 51 1617 101
rect 1571 17 1577 51
rect 1611 17 1617 51
rect 1571 -33 1617 17
rect 1571 -67 1577 -33
rect 1611 -67 1617 -33
rect 1571 -117 1617 -67
rect 1571 -151 1577 -117
rect 1611 -151 1617 -117
rect 1571 -202 1617 -151
tri 1189 -276 1223 -242 sw
tri 1325 -276 1359 -242 se
rect 1359 -276 1405 -236
rect 1571 -236 1577 -202
rect 1611 -236 1617 -202
rect 1681 130 1727 173
tri 1727 169 1731 173 nw
rect 1681 96 1687 130
rect 1721 96 1727 130
rect 1681 51 1727 96
rect 1681 17 1687 51
rect 1721 17 1727 51
rect 1681 -29 1727 17
rect 1681 -63 1687 -29
rect 1721 -63 1727 -29
rect 1681 -109 1727 -63
rect 1681 -143 1687 -109
rect 1721 -143 1727 -109
rect 1681 -189 1727 -143
rect 1681 -223 1687 -189
rect 1721 -223 1727 -189
rect 1681 -235 1727 -223
rect 1784 167 1836 173
tri 1889 169 1893 173 ne
rect 1784 103 1836 115
rect 1784 40 1793 51
rect 1827 40 1836 51
rect 1784 -13 1836 40
rect 1784 -47 1793 -13
rect 1827 -47 1836 -13
rect 1784 -101 1836 -47
rect 1784 -135 1793 -101
rect 1827 -135 1836 -101
rect 1784 -189 1836 -135
rect 1784 -223 1793 -189
rect 1827 -223 1836 -189
rect 1784 -235 1836 -223
rect 1893 130 1939 173
tri 1939 169 1945 175 nw
tri 2099 169 2105 175 ne
rect 1893 96 1899 130
rect 1933 96 1939 130
rect 1893 51 1939 96
rect 1893 17 1899 51
rect 1933 17 1939 51
rect 1893 -29 1939 17
rect 1893 -63 1899 -29
rect 1933 -63 1939 -29
rect 1893 -109 1939 -63
rect 1893 -143 1899 -109
rect 1933 -143 1939 -109
rect 1893 -189 1939 -143
rect 1893 -223 1899 -189
rect 1933 -223 1939 -189
rect 1893 -235 1939 -223
rect 1999 135 2045 147
rect 1999 101 2005 135
rect 2039 101 2045 135
rect 1999 51 2045 101
rect 1999 17 2005 51
rect 2039 17 2045 51
rect 1999 -33 2045 17
rect 1999 -67 2005 -33
rect 2039 -67 2045 -33
rect 1999 -117 2045 -67
rect 1999 -151 2005 -117
rect 2039 -151 2045 -117
rect 1999 -202 2045 -151
tri 1405 -276 1439 -242 sw
tri 1537 -276 1571 -242 se
rect 1571 -276 1617 -236
rect 1999 -236 2005 -202
rect 2039 -236 2045 -202
rect 2105 130 2151 175
rect 2105 96 2111 130
rect 2145 96 2151 130
rect 2105 51 2151 96
rect 2105 17 2111 51
rect 2145 17 2151 51
rect 2105 -29 2151 17
rect 2105 -63 2111 -29
rect 2145 -63 2151 -29
rect 2105 -109 2151 -63
rect 2105 -143 2111 -109
rect 2145 -143 2151 -109
rect 2105 -189 2151 -143
rect 2105 -223 2111 -189
rect 2145 -223 2151 -189
rect 2105 -235 2151 -223
tri 1617 -276 1651 -242 sw
tri 1965 -276 1999 -242 se
rect 1999 -276 2045 -236
tri 2045 -276 2079 -242 sw
rect 74 -287 2179 -276
rect 74 -321 615 -287
rect 649 -321 1149 -287
rect 1183 -321 1365 -287
rect 1399 -321 1577 -287
rect 1611 -321 2005 -287
rect 2039 -321 2179 -287
rect 74 -397 2179 -321
rect 74 -431 501 -397
rect 535 -431 575 -397
rect 609 -431 649 -397
rect 683 -431 723 -397
rect 757 -431 797 -397
rect 831 -431 871 -397
rect 905 -431 945 -397
rect 979 -431 1019 -397
rect 1053 -431 1093 -397
rect 1127 -431 1167 -397
rect 1201 -431 1241 -397
rect 1275 -431 1315 -397
rect 1349 -431 1388 -397
rect 1422 -431 1461 -397
rect 1495 -431 1534 -397
rect 1568 -431 1607 -397
rect 1641 -431 1680 -397
rect 1714 -431 1753 -397
rect 1787 -431 1826 -397
rect 1860 -431 1899 -397
rect 1933 -431 1972 -397
rect 2006 -431 2045 -397
rect 2079 -431 2118 -397
rect 2152 -431 2179 -397
rect 74 -691 2179 -431
<< via1 >>
rect 1914 3428 1931 3462
rect 1931 3428 1965 3462
rect 1965 3428 1966 3462
rect 1914 3410 1966 3428
rect 1914 3342 1966 3394
rect 1914 3274 1966 3326
rect 541 2956 550 2987
rect 550 2956 584 2987
rect 584 2956 593 2987
rect 541 2935 593 2956
rect 541 2912 593 2923
rect 541 2878 550 2912
rect 550 2878 584 2912
rect 584 2878 593 2912
rect 541 2871 593 2878
rect 1084 2800 1136 2806
rect 1084 2766 1118 2800
rect 1118 2766 1136 2800
rect 1084 2754 1136 2766
rect 1149 2754 1201 2806
rect 1214 2754 1266 2806
rect 1278 2800 1330 2806
rect 1278 2766 1296 2800
rect 1296 2766 1330 2800
rect 1278 2754 1330 2766
rect 1821 2956 1830 2988
rect 1830 2956 1864 2988
rect 1864 2956 1873 2988
rect 1821 2936 1873 2956
rect 1821 2912 1873 2924
rect 1821 2878 1830 2912
rect 1830 2878 1864 2912
rect 1864 2878 1873 2912
rect 1821 2872 1873 2878
rect 2037 2956 2089 2982
rect 2037 2930 2046 2956
rect 2046 2930 2080 2956
rect 2080 2930 2089 2956
rect 2037 2878 2089 2918
rect 2037 2866 2046 2878
rect 2046 2866 2080 2878
rect 2080 2866 2089 2878
rect 325 2696 334 2706
rect 334 2696 368 2706
rect 368 2696 377 2706
rect 325 2654 377 2696
rect 735 2706 787 2715
rect 735 2672 739 2706
rect 739 2672 773 2706
rect 773 2672 787 2706
rect 735 2663 787 2672
rect 799 2706 851 2715
rect 799 2672 811 2706
rect 811 2672 845 2706
rect 845 2672 851 2706
rect 799 2663 851 2672
rect 1173 2706 1225 2715
rect 1237 2706 1289 2715
rect 1173 2672 1175 2706
rect 1175 2672 1225 2706
rect 1237 2672 1270 2706
rect 1270 2672 1289 2706
rect 1173 2663 1225 2672
rect 1237 2663 1289 2672
rect 1571 2706 1623 2715
rect 1571 2672 1577 2706
rect 1577 2672 1611 2706
rect 1611 2672 1623 2706
rect 1571 2663 1623 2672
rect 1635 2706 1687 2715
rect 1635 2672 1649 2706
rect 1649 2672 1683 2706
rect 1683 2672 1687 2706
rect 1635 2663 1687 2672
rect 1735 2672 1782 2706
rect 1782 2672 1787 2706
rect 1735 2654 1787 2672
rect 2083 2684 2135 2688
rect 2083 2650 2092 2684
rect 2092 2650 2126 2684
rect 2126 2650 2135 2684
rect 325 2619 334 2642
rect 334 2619 368 2642
rect 368 2619 377 2642
rect 325 2590 377 2619
rect 1735 2590 1787 2642
rect 2083 2636 2135 2650
rect 2083 2612 2135 2624
rect 2083 2578 2092 2612
rect 2092 2578 2126 2612
rect 2126 2578 2135 2612
rect 2083 2572 2135 2578
rect 2204 2684 2256 2688
rect 2204 2650 2213 2684
rect 2213 2650 2247 2684
rect 2247 2650 2256 2684
rect 2204 2636 2256 2650
rect 2204 2612 2256 2624
rect 2204 2578 2213 2612
rect 2213 2578 2247 2612
rect 2247 2578 2256 2612
rect 2204 2572 2256 2578
rect 547 2477 599 2529
rect 611 2477 663 2529
rect 1054 2453 1106 2505
rect 1118 2453 1170 2505
rect 1642 2472 1694 2524
rect 1821 2472 1873 2524
rect 2003 2472 2055 2524
rect 1642 2408 1694 2460
rect 1821 2408 1873 2460
rect 2003 2408 2055 2460
rect 158 2276 164 2310
rect 164 2276 198 2310
rect 198 2276 210 2310
rect 158 2258 210 2276
rect 158 2238 210 2246
rect 158 2204 164 2238
rect 164 2204 198 2238
rect 198 2204 210 2238
rect 158 2194 210 2204
rect 283 2276 289 2310
rect 289 2276 323 2310
rect 323 2276 335 2310
rect 283 2258 335 2276
rect 283 2238 335 2246
rect 283 2204 289 2238
rect 289 2204 323 2238
rect 323 2204 335 2238
rect 283 2194 335 2204
rect 1914 2184 1966 2236
rect 482 2005 534 2057
rect 1207 2080 1259 2089
rect 1271 2080 1323 2089
rect 1207 2046 1240 2080
rect 1240 2046 1259 2080
rect 1271 2046 1274 2080
rect 1274 2046 1318 2080
rect 1318 2046 1323 2080
rect 1207 2037 1259 2046
rect 1271 2037 1323 2046
rect 1914 2086 1966 2138
rect 482 1941 534 1993
rect 1914 1988 1966 2040
rect 1914 1890 1966 1942
rect 289 1726 341 1778
rect 353 1726 405 1778
rect 1207 1726 1259 1778
rect 1271 1726 1323 1778
rect 130 1646 182 1698
rect 194 1646 246 1698
rect 694 1646 746 1698
rect 758 1646 810 1698
rect 1259 1646 1311 1698
rect 1323 1646 1375 1698
rect 2013 1646 2065 1698
rect 2077 1646 2129 1698
rect 850 1566 902 1618
rect 914 1566 966 1618
rect 1395 1486 1447 1538
rect 1459 1486 1511 1538
rect 1545 1372 1597 1424
rect 1545 1308 1597 1360
rect 1741 1122 1793 1174
rect 1805 1122 1857 1174
rect 2134 1042 2186 1094
rect 2198 1042 2250 1094
rect 412 894 464 946
rect 476 894 528 946
rect 566 767 618 819
rect 824 773 876 825
rect 888 773 940 825
rect 566 703 618 755
rect 551 395 603 447
rect 248 365 300 374
rect 312 365 364 374
rect 248 331 262 365
rect 262 331 300 365
rect 312 331 334 365
rect 334 331 364 365
rect 248 322 300 331
rect 312 322 364 331
rect 551 365 603 383
rect 551 331 583 365
rect 583 331 603 365
rect 824 322 876 374
rect 888 365 940 374
rect 888 331 897 365
rect 897 331 931 365
rect 931 331 940 365
rect 888 322 940 331
rect 1122 365 1174 374
rect 1122 331 1152 365
rect 1152 331 1174 365
rect 1122 322 1174 331
rect 1186 365 1238 374
rect 1186 331 1190 365
rect 1190 331 1224 365
rect 1224 331 1238 365
rect 1186 322 1238 331
rect 1435 365 1487 374
rect 1435 331 1438 365
rect 1438 331 1472 365
rect 1472 331 1487 365
rect 1435 322 1487 331
rect 1499 365 1551 374
rect 1499 331 1510 365
rect 1510 331 1544 365
rect 1544 331 1551 365
rect 1499 322 1551 331
rect 1781 365 1833 374
rect 1845 365 1897 374
rect 1781 331 1797 365
rect 1797 331 1833 365
rect 1845 331 1869 365
rect 1869 331 1897 365
rect 1781 322 1833 331
rect 1845 322 1897 331
rect 1978 365 2030 374
rect 1978 331 1982 365
rect 1982 331 2016 365
rect 2016 331 2030 365
rect 1978 322 2030 331
rect 2042 365 2094 374
rect 2042 331 2054 365
rect 2054 331 2088 365
rect 2088 331 2094 365
rect 2042 322 2094 331
rect 162 203 171 232
rect 171 203 205 232
rect 205 203 214 232
rect 712 209 764 215
rect 162 180 214 203
rect 162 133 214 168
rect 162 116 171 133
rect 171 116 205 133
rect 205 116 214 133
rect 712 175 721 209
rect 721 175 755 209
rect 755 175 764 209
rect 712 163 764 175
rect 712 130 764 151
rect 712 99 721 130
rect 721 99 755 130
rect 755 99 764 130
rect 928 161 980 163
rect 928 127 937 161
rect 937 127 971 161
rect 971 127 980 161
rect 928 111 980 127
rect 928 74 980 99
rect 928 47 937 74
rect 937 47 971 74
rect 971 47 980 74
rect 1462 96 1471 129
rect 1471 96 1505 129
rect 1505 96 1514 129
rect 1462 77 1514 96
rect 1462 51 1514 65
rect 1462 17 1471 51
rect 1471 17 1505 51
rect 1505 17 1514 51
rect 1462 13 1514 17
rect 1784 161 1836 167
rect 1784 127 1793 161
rect 1793 127 1827 161
rect 1827 127 1836 161
rect 1784 115 1836 127
rect 1784 74 1836 103
rect 1784 51 1793 74
rect 1793 51 1827 74
rect 1827 51 1836 74
<< metal2 >>
rect 1905 3462 1975 3468
rect 1905 3410 1914 3462
rect 1966 3410 1975 3462
rect 1905 3394 1975 3410
rect 1905 3342 1914 3394
rect 1966 3342 1975 3394
rect 1905 3326 1975 3342
rect 1905 3274 1914 3326
rect 1966 3274 1975 3326
rect 541 2987 593 2993
rect 541 2923 593 2935
rect 325 2706 377 2712
rect 325 2642 377 2654
rect 325 2529 377 2590
tri 377 2529 385 2537 sw
rect 541 2529 593 2871
rect 1821 2988 1873 2994
rect 1821 2924 1873 2936
rect 1078 2754 1084 2806
rect 1136 2754 1149 2806
rect 1201 2754 1214 2806
rect 1266 2754 1278 2806
rect 1330 2764 1336 2806
tri 1336 2764 1369 2797 sw
rect 1330 2754 1369 2764
tri 1305 2715 1344 2754 ne
rect 1344 2715 1369 2754
tri 1369 2715 1418 2764 sw
rect 729 2663 735 2715
rect 787 2663 799 2715
rect 851 2663 896 2715
tri 810 2654 819 2663 ne
rect 819 2654 896 2663
tri 819 2642 831 2654 ne
rect 831 2642 896 2654
tri 831 2629 844 2642 ne
tri 593 2529 627 2563 sw
rect 325 2518 385 2529
tri 385 2518 396 2529 sw
rect 325 2515 396 2518
tri 325 2477 363 2515 ne
rect 363 2477 396 2515
tri 396 2477 437 2518 sw
rect 541 2477 547 2529
rect 599 2477 611 2529
rect 663 2477 669 2529
tri 363 2453 387 2477 ne
rect 387 2453 437 2477
tri 437 2453 461 2477 sw
tri 387 2444 396 2453 ne
rect 396 2444 461 2453
tri 461 2444 470 2453 sw
tri 396 2408 432 2444 ne
rect 432 2408 470 2444
tri 470 2408 506 2444 sw
tri 432 2370 470 2408 ne
rect 470 2370 506 2408
tri 506 2370 544 2408 sw
tri 470 2316 524 2370 ne
rect 524 2316 544 2370
tri 544 2316 598 2370 sw
rect 158 2310 210 2316
rect 158 2246 210 2258
tri 152 1726 158 1732 se
rect 158 1726 210 2194
rect 283 2310 335 2316
tri 524 2296 544 2316 ne
rect 544 2296 598 2316
tri 598 2296 618 2316 sw
tri 544 2274 566 2296 ne
rect 283 2246 335 2258
rect 283 1778 335 2194
rect 482 2057 534 2063
rect 482 1993 534 2005
tri 335 1778 369 1812 sw
tri 210 1726 216 1732 sw
rect 283 1726 289 1778
rect 341 1726 353 1778
rect 405 1726 411 1778
tri 124 1698 152 1726 se
rect 152 1710 216 1726
tri 216 1710 232 1726 sw
tri 283 1710 299 1726 ne
rect 152 1698 232 1710
tri 232 1698 244 1710 sw
rect 299 1698 357 1726
tri 357 1698 385 1726 nw
rect 124 1646 130 1698
rect 182 1646 194 1698
rect 246 1646 252 1698
tri 256 1122 299 1165 se
rect 299 1143 351 1698
tri 351 1692 357 1698 nw
rect 299 1122 330 1143
tri 330 1122 351 1143 nw
tri 228 1094 256 1122 se
rect 256 1094 302 1122
tri 302 1094 330 1122 nw
tri 225 1091 228 1094 se
rect 228 1091 299 1094
tri 299 1091 302 1094 nw
tri 176 1042 225 1091 se
rect 225 1042 250 1091
tri 250 1042 299 1091 nw
tri 162 1028 176 1042 se
rect 176 1028 236 1042
tri 236 1028 250 1042 nw
rect 162 232 214 1028
tri 214 1006 236 1028 nw
tri 448 946 482 980 se
rect 482 946 534 1941
rect 406 894 412 946
rect 464 894 476 946
rect 528 894 534 946
tri 431 860 465 894 ne
tri 452 395 465 408 se
rect 465 395 517 894
tri 517 877 534 894 nw
rect 566 819 618 2296
rect 566 755 618 767
rect 688 1646 694 1698
rect 746 1646 758 1698
rect 810 1646 816 1698
rect 844 1646 896 2642
rect 1167 2663 1173 2715
rect 1225 2663 1237 2715
rect 1289 2663 1295 2715
tri 1344 2690 1369 2715 ne
rect 1369 2690 1418 2715
tri 1418 2690 1443 2715 sw
tri 1369 2663 1396 2690 ne
rect 1396 2663 1443 2690
tri 1443 2663 1470 2690 sw
rect 1545 2663 1571 2715
rect 1623 2663 1635 2715
rect 1687 2663 1693 2715
rect 1735 2706 1787 2712
tri 1133 2529 1167 2563 se
rect 1167 2529 1295 2663
tri 1396 2654 1405 2663 ne
rect 1405 2654 1470 2663
tri 1470 2654 1479 2663 sw
rect 1545 2654 1622 2663
tri 1622 2654 1631 2663 nw
tri 1405 2642 1417 2654 ne
rect 1417 2642 1479 2654
tri 1479 2642 1491 2654 sw
rect 1545 2642 1610 2654
tri 1610 2642 1622 2654 nw
rect 1735 2642 1787 2654
tri 1417 2616 1443 2642 ne
rect 1443 2616 1491 2642
tri 1491 2616 1517 2642 sw
tri 1443 2594 1465 2616 ne
rect 1048 2505 1295 2529
rect 1048 2453 1054 2505
rect 1106 2453 1118 2505
rect 1170 2453 1295 2505
rect 1048 2429 1295 2453
rect 1048 2408 1113 2429
tri 1113 2408 1134 2429 nw
tri 896 1646 902 1652 sw
rect 688 1618 746 1646
tri 746 1618 774 1646 nw
rect 844 1618 902 1646
tri 902 1618 930 1646 sw
rect 566 697 618 703
tri 673 697 688 712 se
rect 688 697 740 1618
tri 740 1612 746 1618 nw
rect 844 1566 850 1618
rect 902 1566 914 1618
rect 966 1566 972 1618
rect 1048 1365 1100 2408
tri 1100 2395 1113 2408 nw
rect 1201 2037 1207 2089
rect 1259 2037 1271 2089
rect 1323 2037 1329 2089
rect 1201 1778 1329 2037
rect 1201 1726 1207 1778
rect 1259 1726 1271 1778
rect 1323 1726 1329 1778
rect 996 1268 1100 1365
rect 1253 1646 1259 1698
rect 1311 1646 1323 1698
rect 1375 1646 1381 1698
rect 818 773 824 825
rect 876 773 888 825
rect 940 773 946 825
tri 666 690 673 697 se
rect 673 690 740 697
tri 603 627 666 690 se
rect 666 627 677 690
tri 677 627 740 690 nw
tri 440 383 452 395 se
rect 452 383 517 395
tri 431 374 440 383 se
rect 440 374 517 383
rect 242 322 248 374
rect 300 322 312 374
rect 364 322 517 374
tri 551 575 603 627 se
rect 551 447 603 575
tri 603 553 677 627 nw
rect 551 383 603 395
rect 894 374 946 773
rect 551 325 603 331
rect 764 322 824 374
rect 876 322 888 374
rect 940 322 946 374
rect 764 296 878 322
tri 878 296 904 322 nw
tri 747 238 764 255 se
rect 764 238 870 296
tri 870 288 878 296 nw
tri 988 288 996 296 se
rect 996 288 1048 1268
tri 1231 1131 1253 1153 se
rect 1253 1131 1305 1646
tri 1305 1612 1339 1646 nw
tri 1431 1538 1465 1572 se
rect 1465 1538 1517 2616
rect 1389 1486 1395 1538
rect 1447 1486 1459 1538
rect 1511 1486 1517 1538
tri 1409 1452 1443 1486 ne
tri 1222 1122 1231 1131 se
rect 1231 1122 1296 1131
tri 1296 1122 1305 1131 nw
tri 1194 1094 1222 1122 se
rect 1222 1098 1272 1122
tri 1272 1098 1296 1122 nw
rect 1222 1094 1268 1098
tri 1268 1094 1272 1098 nw
tri 1439 1094 1443 1098 se
rect 1443 1094 1495 1486
tri 1495 1464 1517 1486 nw
rect 1545 1424 1597 2642
tri 1597 2629 1610 2642 nw
rect 1545 1360 1597 1372
rect 1545 1302 1597 1308
rect 1642 2524 1694 2530
rect 1642 2460 1694 2472
tri 1168 1068 1194 1094 se
rect 1194 1068 1242 1094
tri 1242 1068 1268 1094 nw
tri 1413 1068 1439 1094 se
rect 1439 1076 1495 1094
rect 1439 1068 1461 1076
tri 1142 1042 1168 1068 se
rect 1168 1042 1216 1068
tri 1216 1042 1242 1068 nw
tri 1387 1042 1413 1068 se
rect 1413 1042 1461 1068
tri 1461 1042 1495 1076 nw
tri 1116 1016 1142 1042 se
rect 1142 1024 1198 1042
tri 1198 1024 1216 1042 nw
tri 1369 1024 1387 1042 se
rect 1387 1024 1443 1042
tri 1443 1024 1461 1042 nw
tri 1630 1024 1642 1036 se
rect 1642 1024 1694 2408
rect 1735 1174 1787 2590
rect 1821 2524 1873 2872
rect 1821 2460 1873 2472
rect 1821 2402 1873 2408
rect 1905 2236 1975 3274
rect 2003 2982 2089 2988
rect 2003 2930 2037 2982
rect 2003 2918 2089 2930
rect 2003 2866 2037 2918
rect 2003 2860 2089 2866
rect 2003 2524 2055 2860
tri 2055 2826 2089 2860 nw
rect 2003 2460 2055 2472
rect 2003 2402 2055 2408
rect 2083 2688 2135 2694
rect 2083 2624 2135 2636
rect 1905 2184 1914 2236
rect 1966 2184 1975 2236
rect 1905 2138 1975 2184
rect 1905 2086 1914 2138
rect 1966 2086 1975 2138
rect 1905 2040 1975 2086
rect 1905 1988 1914 2040
rect 1966 1988 1975 2040
rect 1905 1942 1975 1988
rect 1905 1890 1914 1942
rect 1966 1890 1975 1942
rect 1905 1884 1975 1890
tri 2049 1698 2083 1732 se
rect 2083 1698 2135 2572
rect 2007 1646 2013 1698
rect 2065 1646 2077 1698
rect 2129 1646 2135 1698
rect 2204 2688 2256 2694
rect 2204 2624 2256 2636
tri 1787 1174 1821 1208 sw
rect 1735 1122 1741 1174
rect 1793 1122 1805 1174
rect 1857 1122 1903 1174
tri 2198 1122 2204 1128 se
rect 2204 1122 2256 2572
tri 1817 1094 1845 1122 ne
rect 1845 1094 1903 1122
tri 2170 1094 2198 1122 se
rect 2198 1094 2256 1122
tri 1845 1088 1851 1094 ne
rect 1142 1016 1168 1024
rect 1116 374 1168 1016
tri 1168 994 1198 1024 nw
tri 1339 994 1369 1024 se
rect 1369 994 1380 1024
tri 1306 961 1339 994 se
rect 1339 961 1380 994
tri 1380 961 1443 1024 nw
tri 1568 962 1630 1024 se
rect 1630 1014 1694 1024
rect 1630 962 1642 1014
tri 1642 962 1694 1014 nw
tri 1567 961 1568 962 se
rect 1568 961 1579 962
tri 1168 374 1202 408 sw
rect 1116 322 1122 374
rect 1174 322 1186 374
rect 1238 322 1244 374
tri 939 239 988 288 se
rect 988 274 1048 288
rect 988 239 1013 274
tri 1013 239 1048 274 nw
rect 1306 313 1358 961
tri 1358 939 1380 961 nw
tri 1545 939 1567 961 se
rect 1567 939 1579 961
tri 1505 899 1545 939 se
rect 1545 899 1579 939
tri 1579 899 1642 962 nw
tri 1471 374 1505 408 se
rect 1505 374 1557 899
tri 1557 877 1579 899 nw
tri 1557 374 1591 408 sw
tri 1817 374 1851 408 se
rect 1851 374 1903 1094
rect 2128 1042 2134 1094
rect 2186 1042 2198 1094
rect 2250 1042 2256 1094
tri 2170 1008 2204 1042 ne
tri 2197 899 2204 906 se
rect 2204 899 2256 1042
tri 2175 877 2197 899 se
rect 2197 884 2256 899
rect 2197 877 2204 884
tri 2130 832 2175 877 se
rect 2175 832 2204 877
tri 2204 832 2256 884 nw
tri 2067 769 2130 832 se
rect 2130 769 2141 832
tri 2141 769 2204 832 nw
tri 2033 374 2067 408 se
rect 2067 374 2119 769
tri 2119 747 2141 769 nw
rect 1429 322 1435 374
rect 1487 322 1499 374
rect 1551 322 1660 374
tri 1660 322 1712 374 sw
rect 1775 322 1781 374
rect 1833 322 1845 374
rect 1897 322 1903 374
rect 1972 322 1978 374
rect 2030 322 2042 374
rect 2094 322 2119 374
tri 1638 321 1639 322 ne
rect 1639 321 1712 322
tri 1358 313 1366 321 sw
tri 1639 313 1647 321 ne
rect 1647 313 1712 321
rect 1306 299 1366 313
tri 1306 239 1366 299 ne
tri 1366 239 1440 313 sw
tri 1647 248 1712 313 ne
tri 1712 250 1784 322 sw
rect 1712 248 1784 250
tri 1784 248 1786 250 sw
tri 1712 239 1721 248 ne
rect 1721 239 1786 248
tri 730 221 747 238 se
rect 747 221 870 238
rect 162 168 214 180
rect 162 110 214 116
rect 712 215 870 221
rect 764 163 870 215
rect 712 151 870 163
rect 764 99 870 151
rect 712 73 870 99
tri 928 228 939 239 se
rect 939 228 1002 239
tri 1002 228 1013 239 nw
tri 1366 228 1377 239 ne
rect 1377 228 1440 239
rect 928 163 980 228
tri 980 206 1002 228 nw
tri 1377 206 1399 228 ne
rect 1399 206 1440 228
tri 1399 169 1436 206 ne
rect 1436 169 1440 206
tri 1440 169 1510 239 sw
tri 1721 176 1784 239 ne
rect 1784 198 1786 239
tri 1786 198 1836 248 sw
tri 1436 167 1438 169 ne
rect 1438 167 1510 169
tri 1510 167 1512 169 sw
rect 1784 167 1836 198
tri 1438 165 1440 167 ne
rect 1440 165 1512 167
tri 1512 165 1514 167 sw
tri 1440 143 1462 165 ne
rect 928 99 980 111
rect 928 41 980 47
rect 1462 129 1514 165
rect 1462 65 1514 77
rect 1784 103 1836 115
rect 1784 45 1836 51
rect 1462 7 1514 13
use sky130_fd_pr__nfet_01v8__example_55959141808546  sky130_fd_pr__nfet_01v8__example_55959141808546_0
timestamp 1694700623
transform 1 0 660 0 1 -317
box -1 0 51 1
use sky130_fd_pr__nfet_01v8__example_55959141808546  sky130_fd_pr__nfet_01v8__example_55959141808546_1
timestamp 1694700623
transform 1 0 554 0 1 -317
box -1 0 51 1
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_0
timestamp 1694700623
transform 1 0 1732 0 1 -317
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_1
timestamp 1694700623
transform 1 0 1944 0 1 -317
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_2
timestamp 1694700623
transform 1 0 1410 0 1 -317
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_3
timestamp 1694700623
transform 1 0 876 0 1 -317
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808547  sky130_fd_pr__nfet_01v8__example_55959141808547_4
timestamp 1694700623
transform 1 0 1088 0 1 -317
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808600  sky130_fd_pr__nfet_01v8__example_55959141808600_0
timestamp 1694700623
transform 1 0 216 0 1 -17
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_0
timestamp 1694700623
transform 0 -1 1781 1 0 1935
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808596  sky130_fd_pr__pfet_01v8__example_55959141808596_0
timestamp 1694700623
transform -1 0 217 0 -1 3354
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808596  sky130_fd_pr__pfet_01v8__example_55959141808596_1
timestamp 1694700623
transform 1 0 273 0 -1 3354
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808597  sky130_fd_pr__pfet_01v8__example_55959141808597_0
timestamp 1694700623
transform 1 0 1023 0 1 2754
box -1 0 369 1
use sky130_fd_pr__pfet_01v8__example_55959141808598  sky130_fd_pr__pfet_01v8__example_55959141808598_0
timestamp 1694700623
transform 1 0 2197 0 -1 3354
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808598  sky130_fd_pr__pfet_01v8__example_55959141808598_1
timestamp 1694700623
transform 1 0 2091 0 -1 3354
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808599  sky130_fd_pr__pfet_01v8__example_55959141808599_0
timestamp 1694700623
transform 1 0 489 0 1 2754
box -1 0 157 1
use sky130_fd_pr__pfet_01v8__example_55959141808599  sky130_fd_pr__pfet_01v8__example_55959141808599_1
timestamp 1694700623
transform 1 0 1557 0 1 2754
box -1 0 157 1
use sky130_fd_pr__pfet_01v8__example_55959141808599  sky130_fd_pr__pfet_01v8__example_55959141808599_2
timestamp 1694700623
transform 1 0 701 0 1 2754
box -1 0 157 1
use sky130_fd_pr__pfet_01v8__example_55959141808599  sky130_fd_pr__pfet_01v8__example_55959141808599_3
timestamp 1694700623
transform 1 0 1769 0 1 2754
box -1 0 157 1
<< labels >>
flabel metal1 s 367 1129 452 1167 3 FreeSans 200 0 0 0 IN_VCCHIB
port 1 nsew
flabel metal1 s 548 911 656 940 3 FreeSans 200 0 0 0 IN_VDDIO
port 2 nsew
flabel metal1 s 225 1653 324 1691 3 FreeSans 200 0 0 0 MODE_NORMAL_LV
port 3 nsew
flabel metal1 s 844 1572 953 1613 3 FreeSans 200 0 0 0 MODE_NORMAL_LV_N
port 4 nsew
flabel metal1 s 367 1052 463 1086 3 FreeSans 200 0 0 0 MODE_VCCHIB_LV
port 5 nsew
flabel metal1 s 811 1389 932 1425 3 FreeSans 200 0 0 0 MODE_VCCHIB_LV_N
port 6 nsew
flabel metal1 s 244 3325 586 3440 3 FreeSans 200 0 0 0 VCCHIB
port 7 nsew
flabel metal1 s 553 -425 906 -307 3 FreeSans 200 0 0 0 VSSD
port 8 nsew
flabel metal1 s 860 1470 967 1525 3 FreeSans 200 0 0 0 OUT
port 9 nsew
flabel metal1 s 690 2436 845 2511 3 FreeSans 200 0 0 0 OUT_B
port 10 nsew
<< properties >>
string GDS_END 3669914
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3600366
<< end >>
