magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 79 21 1287 203
rect 29 -17 63 17
<< locali >>
rect 119 341 156 493
rect 290 341 328 493
rect 17 299 328 341
rect 17 175 68 299
rect 525 289 835 340
rect 525 265 561 289
rect 17 127 405 175
rect 197 123 405 127
rect 508 197 561 265
rect 595 197 729 255
rect 769 197 835 289
rect 899 302 1169 340
rect 899 204 965 302
rect 1007 204 1076 266
rect 1127 264 1169 302
rect 1127 204 1245 264
rect 197 51 235 123
rect 369 51 405 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 375 85 527
rect 190 375 256 527
rect 362 367 412 527
rect 464 442 890 493
rect 924 455 990 527
rect 824 421 890 442
rect 1032 421 1084 493
rect 1118 455 1184 527
rect 1218 421 1269 493
rect 456 374 702 408
rect 824 376 1269 421
rect 456 335 491 374
rect 437 301 491 335
rect 437 265 474 301
rect 105 209 474 265
rect 439 161 474 209
rect 1203 307 1269 376
rect 439 123 1098 161
rect 97 17 163 93
rect 269 17 335 89
rect 444 17 511 89
rect 545 51 594 123
rect 628 17 694 89
rect 728 51 804 123
rect 838 17 912 89
rect 1032 55 1098 123
rect 1203 17 1269 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1007 204 1076 266 6 A1
port 1 nsew signal input
rlabel locali s 1127 204 1245 264 6 A2
port 2 nsew signal input
rlabel locali s 1127 264 1169 302 6 A2
port 2 nsew signal input
rlabel locali s 899 204 965 302 6 A2
port 2 nsew signal input
rlabel locali s 899 302 1169 340 6 A2
port 2 nsew signal input
rlabel locali s 769 197 835 289 6 B1
port 3 nsew signal input
rlabel locali s 508 197 561 265 6 B1
port 3 nsew signal input
rlabel locali s 525 265 561 289 6 B1
port 3 nsew signal input
rlabel locali s 525 289 835 340 6 B1
port 3 nsew signal input
rlabel locali s 595 197 729 255 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 369 51 405 123 6 X
port 9 nsew signal output
rlabel locali s 197 51 235 123 6 X
port 9 nsew signal output
rlabel locali s 197 123 405 127 6 X
port 9 nsew signal output
rlabel locali s 17 127 405 175 6 X
port 9 nsew signal output
rlabel locali s 17 175 68 299 6 X
port 9 nsew signal output
rlabel locali s 17 299 328 341 6 X
port 9 nsew signal output
rlabel locali s 290 341 328 493 6 X
port 9 nsew signal output
rlabel locali s 119 341 156 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3628952
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3619892
<< end >>
