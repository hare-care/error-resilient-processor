magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 28 21 1078 203
rect 29 -17 63 21
<< scnmos >>
rect 106 47 136 177
rect 190 47 220 177
rect 274 47 304 177
rect 358 47 388 177
rect 442 47 472 177
rect 526 47 556 177
rect 714 47 744 177
rect 798 47 828 177
rect 882 47 912 177
rect 966 47 996 177
<< scpmoshvt >>
rect 106 297 136 497
rect 190 297 220 497
rect 274 297 304 497
rect 358 297 388 497
rect 442 297 472 497
rect 526 297 556 497
rect 714 297 744 497
rect 798 297 828 497
rect 882 297 912 497
rect 966 297 996 497
<< ndiff >>
rect 54 163 106 177
rect 54 129 62 163
rect 96 129 106 163
rect 54 95 106 129
rect 54 61 62 95
rect 96 61 106 95
rect 54 47 106 61
rect 136 163 190 177
rect 136 129 146 163
rect 180 129 190 163
rect 136 95 190 129
rect 136 61 146 95
rect 180 61 190 95
rect 136 47 190 61
rect 220 163 274 177
rect 220 129 230 163
rect 264 129 274 163
rect 220 47 274 129
rect 304 95 358 177
rect 304 61 314 95
rect 348 61 358 95
rect 304 47 358 61
rect 388 95 442 177
rect 388 61 398 95
rect 432 61 442 95
rect 388 47 442 61
rect 472 163 526 177
rect 472 129 482 163
rect 516 129 526 163
rect 472 95 526 129
rect 472 61 482 95
rect 516 61 526 95
rect 472 47 526 61
rect 556 95 714 177
rect 556 61 566 95
rect 600 61 670 95
rect 704 61 714 95
rect 556 47 714 61
rect 744 163 798 177
rect 744 129 754 163
rect 788 129 798 163
rect 744 95 798 129
rect 744 61 754 95
rect 788 61 798 95
rect 744 47 798 61
rect 828 95 882 177
rect 828 61 838 95
rect 872 61 882 95
rect 828 47 882 61
rect 912 163 966 177
rect 912 129 922 163
rect 956 129 966 163
rect 912 95 966 129
rect 912 61 922 95
rect 956 61 966 95
rect 912 47 966 61
rect 996 163 1052 177
rect 996 129 1006 163
rect 1040 129 1052 163
rect 996 95 1052 129
rect 996 61 1006 95
rect 1040 61 1052 95
rect 996 47 1052 61
<< pdiff >>
rect 54 477 106 497
rect 54 443 62 477
rect 96 443 106 477
rect 54 409 106 443
rect 54 375 62 409
rect 96 375 106 409
rect 54 297 106 375
rect 136 477 190 497
rect 136 443 146 477
rect 180 443 190 477
rect 136 297 190 443
rect 220 477 274 497
rect 220 443 230 477
rect 264 443 274 477
rect 220 409 274 443
rect 220 375 230 409
rect 264 375 274 409
rect 220 297 274 375
rect 304 477 358 497
rect 304 443 314 477
rect 348 443 358 477
rect 304 297 358 443
rect 388 477 442 497
rect 388 443 398 477
rect 432 443 442 477
rect 388 409 442 443
rect 388 375 398 409
rect 432 375 442 409
rect 388 297 442 375
rect 472 409 526 497
rect 472 375 482 409
rect 516 375 526 409
rect 472 341 526 375
rect 472 307 482 341
rect 516 307 526 341
rect 472 297 526 307
rect 556 477 608 497
rect 556 443 566 477
rect 600 443 608 477
rect 556 409 608 443
rect 556 375 566 409
rect 600 375 608 409
rect 556 297 608 375
rect 662 477 714 497
rect 662 443 670 477
rect 704 443 714 477
rect 662 409 714 443
rect 662 375 670 409
rect 704 375 714 409
rect 662 297 714 375
rect 744 477 798 497
rect 744 443 754 477
rect 788 443 798 477
rect 744 297 798 443
rect 828 477 882 497
rect 828 443 838 477
rect 872 443 882 477
rect 828 409 882 443
rect 828 375 838 409
rect 872 375 882 409
rect 828 297 882 375
rect 912 409 966 497
rect 912 375 922 409
rect 956 375 966 409
rect 912 341 966 375
rect 912 307 922 341
rect 956 307 966 341
rect 912 297 966 307
rect 996 477 1052 497
rect 996 443 1006 477
rect 1040 443 1052 477
rect 996 409 1052 443
rect 996 375 1006 409
rect 1040 375 1052 409
rect 996 341 1052 375
rect 996 307 1006 341
rect 1040 307 1052 341
rect 996 297 1052 307
<< ndiffc >>
rect 62 129 96 163
rect 62 61 96 95
rect 146 129 180 163
rect 146 61 180 95
rect 230 129 264 163
rect 314 61 348 95
rect 398 61 432 95
rect 482 129 516 163
rect 482 61 516 95
rect 566 61 600 95
rect 670 61 704 95
rect 754 129 788 163
rect 754 61 788 95
rect 838 61 872 95
rect 922 129 956 163
rect 922 61 956 95
rect 1006 129 1040 163
rect 1006 61 1040 95
<< pdiffc >>
rect 62 443 96 477
rect 62 375 96 409
rect 146 443 180 477
rect 230 443 264 477
rect 230 375 264 409
rect 314 443 348 477
rect 398 443 432 477
rect 398 375 432 409
rect 482 375 516 409
rect 482 307 516 341
rect 566 443 600 477
rect 566 375 600 409
rect 670 443 704 477
rect 670 375 704 409
rect 754 443 788 477
rect 838 443 872 477
rect 838 375 872 409
rect 922 375 956 409
rect 922 307 956 341
rect 1006 443 1040 477
rect 1006 375 1040 409
rect 1006 307 1040 341
<< poly >>
rect 106 497 136 523
rect 190 497 220 523
rect 274 497 304 523
rect 358 497 388 523
rect 442 497 472 523
rect 526 497 556 523
rect 714 497 744 523
rect 798 497 828 523
rect 882 497 912 523
rect 966 497 996 523
rect 106 265 136 297
rect 82 249 136 265
rect 82 215 92 249
rect 126 215 136 249
rect 82 199 136 215
rect 106 177 136 199
rect 190 265 220 297
rect 274 265 304 297
rect 358 265 388 297
rect 442 265 472 297
rect 526 265 556 297
rect 714 265 744 297
rect 798 265 828 297
rect 190 249 304 265
rect 190 215 230 249
rect 264 215 304 249
rect 190 199 304 215
rect 346 249 400 265
rect 346 215 356 249
rect 390 215 400 249
rect 346 199 400 215
rect 442 249 616 265
rect 442 215 566 249
rect 600 215 616 249
rect 442 199 616 215
rect 714 249 828 265
rect 714 215 752 249
rect 786 215 828 249
rect 714 199 828 215
rect 190 177 220 199
rect 274 177 304 199
rect 358 177 388 199
rect 442 177 472 199
rect 526 177 556 199
rect 714 177 744 199
rect 798 177 828 199
rect 882 265 912 297
rect 966 265 996 297
rect 882 249 996 265
rect 882 215 924 249
rect 958 215 996 249
rect 882 199 996 215
rect 882 177 912 199
rect 966 177 996 199
rect 106 21 136 47
rect 190 21 220 47
rect 274 21 304 47
rect 358 21 388 47
rect 442 21 472 47
rect 526 21 556 47
rect 714 21 744 47
rect 798 21 828 47
rect 882 21 912 47
rect 966 21 996 47
<< polycont >>
rect 92 215 126 249
rect 230 215 264 249
rect 356 215 390 249
rect 566 215 600 249
rect 752 215 786 249
rect 924 215 958 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 54 477 104 493
rect 54 443 62 477
rect 96 443 104 477
rect 54 409 104 443
rect 138 477 188 527
rect 138 443 146 477
rect 180 443 188 477
rect 138 427 188 443
rect 222 477 272 493
rect 222 443 230 477
rect 264 443 272 477
rect 54 375 62 409
rect 96 391 104 409
rect 222 409 272 443
rect 306 477 356 527
rect 306 443 314 477
rect 348 443 356 477
rect 306 427 356 443
rect 390 477 608 493
rect 390 443 398 477
rect 432 459 566 477
rect 432 443 440 459
rect 222 391 230 409
rect 96 375 230 391
rect 264 391 272 409
rect 390 409 440 443
rect 558 443 566 459
rect 600 443 608 477
rect 390 391 398 409
rect 264 375 398 391
rect 432 375 440 409
rect 54 357 440 375
rect 474 409 524 425
rect 474 375 482 409
rect 516 375 524 409
rect 474 341 524 375
rect 558 409 608 443
rect 558 375 566 409
rect 600 375 608 409
rect 558 359 608 375
rect 662 477 712 493
rect 662 443 670 477
rect 704 443 712 477
rect 662 409 712 443
rect 746 477 796 527
rect 746 443 754 477
rect 788 443 796 477
rect 746 427 796 443
rect 830 477 1048 493
rect 830 443 838 477
rect 872 459 1006 477
rect 872 443 880 459
rect 662 375 670 409
rect 704 393 712 409
rect 830 409 880 443
rect 998 443 1006 459
rect 1040 443 1048 477
rect 830 393 838 409
rect 704 375 838 393
rect 872 375 880 409
rect 662 357 880 375
rect 914 409 964 425
rect 914 375 922 409
rect 956 375 964 409
rect 17 289 406 323
rect 17 249 142 289
rect 17 215 92 249
rect 126 215 142 249
rect 188 249 296 255
rect 188 215 230 249
rect 264 215 296 249
rect 340 249 406 289
rect 340 215 356 249
rect 390 215 406 249
rect 474 307 482 341
rect 516 332 524 341
rect 914 341 964 375
rect 516 307 532 332
rect 914 323 922 341
rect 474 181 532 307
rect 590 307 922 323
rect 956 307 964 341
rect 590 289 964 307
rect 998 409 1048 443
rect 998 375 1006 409
rect 1040 375 1048 409
rect 998 341 1048 375
rect 998 307 1006 341
rect 1040 307 1048 341
rect 998 291 1048 307
rect 590 265 624 289
rect 566 249 624 265
rect 600 215 624 249
rect 662 249 841 255
rect 662 215 752 249
rect 786 215 841 249
rect 891 249 1087 255
rect 891 215 924 249
rect 958 215 1087 249
rect 566 199 624 215
rect 62 163 96 179
rect 62 95 96 129
rect 62 17 96 61
rect 130 163 180 179
rect 130 129 146 163
rect 214 163 532 181
rect 214 129 230 163
rect 264 145 482 163
rect 264 129 280 145
rect 466 129 482 145
rect 516 129 532 163
rect 590 181 624 199
rect 590 163 972 181
rect 590 145 754 163
rect 130 95 180 129
rect 398 95 432 111
rect 130 61 146 95
rect 180 61 314 95
rect 348 61 364 95
rect 130 51 364 61
rect 398 17 432 61
rect 466 95 532 129
rect 738 129 754 145
rect 788 145 922 163
rect 788 129 804 145
rect 466 61 482 95
rect 516 61 532 95
rect 466 51 532 61
rect 566 95 704 111
rect 600 61 670 95
rect 566 17 704 61
rect 738 95 804 129
rect 906 129 922 145
rect 956 129 972 163
rect 738 61 754 95
rect 788 61 804 95
rect 738 51 804 61
rect 838 95 872 111
rect 838 17 872 61
rect 906 95 972 129
rect 906 61 922 95
rect 956 61 972 95
rect 906 51 972 61
rect 1006 163 1040 181
rect 1006 95 1040 129
rect 1006 17 1040 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 953 221 987 255 0 FreeSans 400 180 0 0 A2_N
port 2 nsew signal input
flabel locali s 769 221 803 255 0 FreeSans 400 180 0 0 A1_N
port 1 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2bb2oi_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 3950548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3941750
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
