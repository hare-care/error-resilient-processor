magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 23790 36886 28084 37121
rect 26179 36716 28084 36886
rect 26788 36021 28084 36716
rect 26780 34970 28084 36021
rect 26635 32388 28084 34970
rect 26748 25618 28084 32388
rect 26500 24436 28084 25618
rect 23790 23485 28084 24436
rect 1231 21526 28211 21948
rect 27789 13586 28211 21526
rect 1231 13284 28211 13586
rect 26545 12731 28136 13003
rect 27864 10851 28136 12731
rect 26545 10579 28136 10851
rect -80 2099 2376 2385
rect -80 286 206 2099
rect -80 0 2376 286
<< pwell >>
rect 22823 22873 28026 23379
rect 26249 22054 28026 22873
rect 2294 3728 28026 4086
rect 6423 3404 28026 3728
<< obsli1 >>
rect 46 36935 28000 39956
rect 46 23538 28017 36935
rect 46 23353 28000 23538
rect 46 22080 28029 23353
rect 46 21822 28000 22080
rect 46 13434 28095 21822
rect 46 13350 28085 13434
rect 46 12937 28000 13350
rect 46 10645 28070 12937
rect 46 40 28000 10645
<< obsm1 >>
rect 16 36944 28000 39962
rect 16 36641 28029 36944
rect 16 23526 28023 36641
tri 28023 36635 28029 36641 nw
rect 16 21774 28000 23526
rect 16 13434 28095 21774
rect 16 12937 28000 13434
rect 16 10645 28070 12937
rect 16 0 28000 10645
<< obsm2 >>
rect 16 36944 28000 39991
rect 16 36578 28026 36944
rect 16 13628 28000 36578
rect 16 12743 28065 13628
rect 16 0 28000 12743
<< metal3 >>
rect 66 14276 144 14354
rect 248 14165 332 14249
rect 25995 12331 26058 12394
rect 25655 4036 25659 4040
rect 3927 3597 3990 3660
rect 15556 2973 15635 3052
rect 1586 2777 1623 2814
rect 5380 2720 5471 2811
rect 24916 2364 24982 2430
rect 8981 1522 9071 1612
rect 21456 1559 21509 1612
rect 24841 1564 24889 1612
rect 430 1153 529 1252
rect 1153 0 1273 129
rect 1422 0 1488 134
rect 1754 0 1820 134
rect 4076 0 4142 134
rect 4427 0 4493 134
rect 4876 0 4942 134
rect 8807 0 8873 134
rect 9241 0 9307 134
rect 10331 0 10397 156
rect 12997 183 13047 233
rect 13217 0 13283 134
rect 13387 0 13453 134
rect 17363 0 17429 134
rect 17533 0 17599 134
rect 19169 0 19243 74
rect 21679 0 21745 134
rect 23058 0 23178 166
rect 25825 0 25891 134
<< obsm3 >>
rect 66 14434 28000 39943
rect 224 14329 28000 14434
rect 66 14085 168 14196
rect 412 14085 28000 14329
rect 66 12474 28000 14085
rect 66 12251 25915 12474
rect 26138 12251 28000 12474
rect 66 4120 28000 12251
rect 66 3956 25575 4120
rect 25739 3956 28000 4120
rect 66 3740 28000 3956
rect 66 3517 3847 3740
rect 4070 3517 28000 3740
rect 66 3132 28000 3517
rect 66 2894 15476 3132
rect 66 2697 1506 2894
rect 1703 2893 15476 2894
rect 15715 2893 28000 3132
rect 1703 2891 28000 2893
rect 1703 2697 5300 2891
rect 66 2640 5300 2697
rect 5551 2640 28000 2891
rect 66 2510 28000 2640
rect 66 2284 24836 2510
rect 25062 2284 28000 2510
rect 66 1692 28000 2284
rect 66 1442 8901 1692
rect 9151 1479 21376 1692
rect 21589 1484 24761 1692
rect 24969 1484 28000 1692
rect 21589 1479 28000 1484
rect 9151 1442 28000 1479
rect 66 1332 28000 1442
rect 66 1073 350 1332
rect 609 1073 28000 1332
rect 66 313 28000 1073
rect 66 236 12917 313
rect 66 214 10251 236
rect 66 209 1342 214
rect 66 0 1073 209
rect 1568 0 1674 214
rect 1900 0 3996 214
rect 4222 0 4347 214
rect 4573 0 4796 214
rect 5022 0 8727 214
rect 8953 0 9161 214
rect 9387 0 10251 214
rect 10477 103 12917 236
rect 13127 246 28000 313
rect 13127 214 22978 246
rect 13127 103 13137 214
rect 10477 0 13137 103
rect 13533 0 17283 214
rect 17679 154 21599 214
rect 17679 0 19089 154
rect 19323 0 21599 154
rect 21825 0 22978 214
rect 23258 214 28000 246
rect 23258 0 25745 214
rect 25971 0 28000 214
<< metal4 >>
rect 0 35157 273 40000
rect 27746 35157 28000 40000
rect 0 14007 254 19000
rect 27746 14007 28000 19000
rect 0 12817 254 13707
rect 27746 12817 28000 13707
rect 0 11647 254 12537
rect 27746 11647 28000 12537
rect 0 11281 28000 11347
rect 0 10625 254 11221
rect 0 10329 408 10565
rect 0 9673 254 10269
rect 27746 10625 28000 11221
rect 27746 10329 28000 10565
rect 27746 9673 28000 10269
rect 0 9547 28000 9613
rect 0 8317 254 9247
rect 27746 8317 28000 9247
rect 0 7347 254 8037
rect 27746 7347 28000 8037
rect 0 6377 254 7067
rect 27746 6377 28000 7067
rect 0 5167 254 6097
rect 27746 5167 28000 6097
rect 0 3957 254 4887
rect 27746 3957 28000 4887
rect 0 2987 193 3677
rect 27807 2987 28000 3677
rect 0 1777 254 2707
rect 27746 1777 28000 2707
rect 0 407 254 1497
rect 27746 407 28000 1497
<< obsm4 >>
rect 353 35077 27666 40000
rect 193 19080 27807 35077
rect 334 13927 27666 19080
rect 193 13787 27807 13927
rect 334 12737 27666 13787
rect 193 12617 27807 12737
rect 334 11567 27666 12617
rect 193 11427 27807 11567
rect 334 10645 27666 11201
rect 488 10249 27666 10645
rect 334 9693 27666 10249
rect 193 9327 27807 9467
rect 334 8237 27666 9327
rect 193 8117 27807 8237
rect 334 7267 27666 8117
rect 193 7147 27807 7267
rect 334 6297 27666 7147
rect 193 6177 27807 6297
rect 334 5087 27666 6177
rect 193 4967 27807 5087
rect 334 3877 27666 4967
rect 193 3757 27807 3877
rect 273 2907 27727 3757
rect 193 2787 27807 2907
rect 334 1697 27666 2787
rect 193 1577 27807 1697
rect 334 327 27666 1577
rect 193 232 27807 327
<< metal5 >>
rect 0 35157 273 40000
rect 27746 35157 28000 40000
rect 8019 26541 12627 29546
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 27746 14007 28000 18997
rect 27746 12837 28000 13687
rect 27746 11667 28000 12517
rect 0 9547 408 11347
rect 27746 9547 28000 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 27746 8337 28000 9227
rect 27746 7368 28000 8017
rect 27746 6397 28000 7047
rect 27746 5187 28000 6077
rect 27746 3977 28000 4867
rect 0 3007 193 3657
rect 27807 3007 28000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 27746 1797 28000 2687
rect 27746 427 28000 1477
<< obsm5 >>
rect 593 34837 27426 40000
rect 0 29866 28000 34837
rect 0 26221 7699 29866
rect 12947 26221 28000 29866
rect 0 19317 28000 26221
rect 574 11667 27426 19317
rect 728 9227 27426 11667
rect 574 3657 27426 9227
rect 513 3007 27487 3657
rect 574 427 27426 3007
<< labels >>
rlabel metal5 s 27746 11667 28000 12517 6 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal4 s 27746 11647 28000 12537 6 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 1 nsew ground bidirectional
rlabel metal5 s 27746 6397 28000 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 27746 6377 28000 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 27746 5187 28000 6077 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 27746 35157 28000 40000 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 0 35157 273 40000 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 27746 35157 28000 40000 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 27746 5167 28000 6097 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 0 35157 273 40000 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 3 nsew ground bidirectional
rlabel metal5 s 27746 8337 28000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 27746 8317 28000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 27746 7368 28000 8017 6 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 27746 9547 28000 11347 6 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 0 9547 408 11347 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 10329 28000 10565 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 9547 28000 9613 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 11281 28000 11347 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 27746 7347 28000 8037 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 10329 408 10565 6 VSSA
port 5 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 5 nsew ground bidirectional
rlabel metal5 s 27746 12837 28000 13687 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 27746 12817 28000 13707 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 27746 14007 28000 18997 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 27746 3977 28000 4867 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 27746 3957 28000 4887 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 27746 14007 28000 19000 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 27807 3007 28000 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 27807 2987 28000 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 27746 427 28000 1477 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal4 s 27746 407 28000 1497 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 27746 1797 28000 2687 6 VCCD
port 10 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 27746 1777 28000 2707 6 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 10 nsew power bidirectional
rlabel metal5 s 8019 26541 12627 29546 6 PAD
port 11 nsew signal bidirectional
rlabel metal4 s 27746 10625 28000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 0 10625 254 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 27746 9673 28000 10269 6 AMUXBUS_B
port 13 nsew signal bidirectional
rlabel metal4 s 0 9673 254 10269 6 AMUXBUS_B
port 13 nsew signal bidirectional
rlabel metal3 s 25825 0 25891 134 6 DM[0]
port 14 nsew signal input
rlabel metal3 s 25655 4036 25659 4040 6 DM[1]
port 15 nsew signal input
rlabel metal3 s 21679 0 21745 134 6 DM[2]
port 16 nsew signal input
rlabel metal3 s 21456 1559 21509 1612 6 INP_DIS
port 17 nsew signal input
rlabel metal3 s 17533 0 17599 134 6 VTRIP_SEL
port 18 nsew signal input
rlabel metal3 s 17363 0 17429 134 6 IB_MODE_SEL[0]
port 19 nsew signal input
rlabel metal3 s 13387 0 13453 134 6 IB_MODE_SEL[1]
port 20 nsew signal input
rlabel metal3 s 13217 0 13283 134 6 SLEW_CTL[0]
port 21 nsew signal input
rlabel metal3 s 9241 0 9307 134 6 SLEW_CTL[1]
port 22 nsew signal input
rlabel metal3 s 8981 1522 9071 1612 6 HYS_TRIM
port 23 nsew signal input
rlabel metal3 s 5380 2720 5471 2811 6 HLD_OVR
port 24 nsew signal input
rlabel metal3 s 4427 0 4493 134 6 ENABLE_H
port 25 nsew signal input
rlabel metal3 s 3927 3597 3990 3660 6 HLD_H_N
port 26 nsew signal input
rlabel metal3 s 1754 0 1820 134 6 ENABLE_VDDA_H
port 27 nsew signal input
rlabel metal3 s 1586 2777 1623 2814 6 ANALOG_EN
port 28 nsew signal input
rlabel metal3 s 1422 0 1488 134 6 ENABLE_INP_H
port 29 nsew signal input
rlabel metal3 s 4076 0 4142 134 6 IN
port 30 nsew signal output
rlabel metal3 s 4876 0 4942 134 6 IN_H
port 31 nsew signal output
rlabel metal3 s 8807 0 8873 134 6 VINREF
port 32 nsew signal input
rlabel metal3 s 15556 2973 15635 3052 6 OUT
port 33 nsew signal input
rlabel metal3 s 12997 183 13047 233 6 ANALOG_POL
port 34 nsew signal input
rlabel metal3 s 10331 0 10397 156 6 ANALOG_SEL
port 35 nsew signal input
rlabel metal3 s 24916 2364 24982 2430 6 SLOW
port 36 nsew signal input
rlabel metal3 s 24841 1564 24889 1612 6 OE_N
port 37 nsew signal input
rlabel metal3 s 25995 12331 26058 12394 6 TIE_HI_ESD
port 38 nsew signal output
rlabel metal3 s 23058 0 23178 166 6 TIE_LO_ESD
port 39 nsew signal output
rlabel metal3 s 248 14165 332 14249 6 PAD_A_ESD_0_H
port 40 nsew signal bidirectional
rlabel metal3 s 66 14276 144 14354 6 PAD_A_ESD_1_H
port 41 nsew signal bidirectional
rlabel metal3 s 430 1153 529 1252 6 PAD_A_NOESD_H
port 42 nsew signal bidirectional
rlabel metal3 s 1153 0 1273 129 6 ENABLE_VSWITCH_H
port 43 nsew signal input
rlabel metal3 s 19169 0 19243 74 6 ENABLE_VDDIO
port 44 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 28000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 51049346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 50423142
<< end >>
