magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 39 79 513 203
rect 39 17 63 79
rect 29 -17 63 17
<< scnmos >>
rect 117 105 147 177
rect 189 105 219 177
rect 261 105 291 177
rect 333 105 363 177
rect 405 105 435 177
<< ndiff >>
rect 65 158 117 177
rect 65 124 73 158
rect 107 124 117 158
rect 65 105 117 124
rect 147 105 189 177
rect 219 105 261 177
rect 291 105 333 177
rect 363 105 405 177
rect 435 158 487 177
rect 435 124 445 158
rect 479 124 487 158
rect 435 105 487 124
<< ndiffc >>
rect 73 124 107 158
rect 445 124 479 158
<< poly >>
rect 117 249 435 265
rect 117 215 127 249
rect 161 215 195 249
rect 229 215 263 249
rect 297 215 331 249
rect 365 215 435 249
rect 117 199 435 215
rect 117 177 147 199
rect 189 177 219 199
rect 261 177 291 199
rect 333 177 363 199
rect 405 177 435 199
rect 117 79 147 105
rect 189 79 219 105
rect 261 79 291 105
rect 333 79 363 105
rect 405 79 435 105
<< polycont >>
rect 127 215 161 249
rect 195 215 229 249
rect 263 215 297 249
rect 331 215 365 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 55 249 395 346
rect 55 215 127 249
rect 161 215 195 249
rect 229 215 263 249
rect 297 215 331 249
rect 365 215 395 249
rect 55 208 395 215
rect 57 158 123 174
rect 57 124 73 158
rect 107 124 123 158
rect 57 17 123 124
rect 429 158 495 527
rect 429 124 445 158
rect 479 124 495 158
rect 429 108 495 124
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lpflow_bleeder_1
flabel nwell s 29 527 63 561 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel locali s 87 292 121 326 0 FreeSans 200 0 0 0 SHORT
port 1 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 2235430
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2232438
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
