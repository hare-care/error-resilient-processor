magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 145 457 157
rect 741 145 1011 203
rect 1 21 1011 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 446 47 476 119
rect 545 47 575 119
rect 629 47 659 119
rect 819 47 849 177
rect 903 47 933 177
<< scpmoshvt >>
rect 79 381 109 491
rect 163 381 193 491
rect 351 369 381 497
rect 446 413 476 497
rect 530 413 560 497
rect 629 413 659 497
rect 819 297 849 497
rect 903 297 933 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 767 133 819 177
rect 381 47 446 119
rect 476 107 545 119
rect 476 73 500 107
rect 534 73 545 107
rect 476 47 545 73
rect 575 47 629 119
rect 659 106 711 119
rect 659 72 669 106
rect 703 72 711 106
rect 659 47 711 72
rect 767 99 775 133
rect 809 99 819 133
rect 767 47 819 99
rect 849 127 903 177
rect 849 93 859 127
rect 893 93 903 127
rect 849 47 903 93
rect 933 133 985 177
rect 933 99 943 133
rect 977 99 985 133
rect 933 47 985 99
<< pdiff >>
rect 27 452 79 491
rect 27 418 35 452
rect 69 418 79 452
rect 27 381 79 418
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 381 163 427
rect 193 452 245 491
rect 193 418 203 452
rect 237 418 245 452
rect 193 381 245 418
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 369 351 451
rect 381 413 446 497
rect 476 485 530 497
rect 476 451 486 485
rect 520 451 530 485
rect 476 413 530 451
rect 560 413 629 497
rect 659 477 713 497
rect 659 443 671 477
rect 705 443 713 477
rect 659 413 713 443
rect 767 471 819 497
rect 767 437 775 471
rect 809 437 819 471
rect 381 369 431 413
rect 767 368 819 437
rect 767 334 775 368
rect 809 334 819 368
rect 767 297 819 334
rect 849 484 903 497
rect 849 450 859 484
rect 893 450 903 484
rect 849 364 903 450
rect 849 330 859 364
rect 893 330 903 364
rect 849 297 903 330
rect 933 475 985 497
rect 933 441 943 475
rect 977 441 985 475
rect 933 384 985 441
rect 933 350 943 384
rect 977 350 985 384
rect 933 297 985 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 500 73 534 107
rect 669 72 703 106
rect 775 99 809 133
rect 859 93 893 127
rect 943 99 977 133
<< pdiffc >>
rect 35 418 69 452
rect 119 427 153 461
rect 203 418 237 452
rect 307 451 341 485
rect 486 451 520 485
rect 671 443 705 477
rect 775 437 809 471
rect 775 334 809 368
rect 859 450 893 484
rect 859 330 893 364
rect 943 441 977 475
rect 943 350 977 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 446 497 476 523
rect 530 497 560 523
rect 629 497 659 523
rect 819 497 849 523
rect 903 497 933 523
rect 79 365 109 381
rect 46 335 109 365
rect 46 280 76 335
rect 163 316 193 381
rect 163 300 308 316
rect 163 292 264 300
rect 22 264 76 280
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 276 264 292
rect 118 242 128 276
rect 162 266 264 276
rect 298 266 308 300
rect 162 250 308 266
rect 162 242 193 250
rect 118 226 193 242
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 226
rect 351 219 381 369
rect 446 337 476 413
rect 530 375 560 413
rect 519 365 585 375
rect 423 321 477 337
rect 519 331 535 365
rect 569 331 585 365
rect 519 321 585 331
rect 629 373 659 413
rect 629 357 728 373
rect 629 323 684 357
rect 718 323 728 357
rect 423 287 433 321
rect 467 287 477 321
rect 423 279 477 287
rect 629 307 728 323
rect 423 271 575 279
rect 447 249 575 271
rect 340 203 394 219
rect 340 169 350 203
rect 384 169 394 203
rect 340 146 394 169
rect 446 191 503 207
rect 446 157 459 191
rect 493 157 503 191
rect 351 131 381 146
rect 446 141 503 157
rect 446 119 476 141
rect 545 119 575 249
rect 629 119 659 307
rect 819 265 849 297
rect 903 265 933 297
rect 704 249 933 265
rect 704 215 722 249
rect 756 215 933 249
rect 704 199 933 215
rect 819 177 849 199
rect 903 177 933 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 545 21 575 47
rect 629 21 659 47
rect 819 21 849 47
rect 903 21 933 47
<< polycont >>
rect 32 230 66 264
rect 128 242 162 276
rect 264 266 298 300
rect 535 331 569 365
rect 684 323 718 357
rect 433 287 467 321
rect 350 169 384 203
rect 459 157 493 191
rect 722 215 756 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 35 452 69 493
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 452 237 493
rect 35 393 69 418
rect 291 485 370 527
rect 291 451 307 485
rect 341 451 370 485
rect 462 451 486 485
rect 520 451 637 485
rect 203 417 237 418
rect 203 393 569 417
rect 35 359 156 393
rect 18 264 66 325
rect 18 230 32 264
rect 18 197 66 230
rect 122 292 156 359
rect 196 383 569 393
rect 196 365 237 383
rect 501 365 569 383
rect 122 276 162 292
rect 122 242 128 276
rect 122 226 162 242
rect 122 161 156 226
rect 35 127 156 161
rect 196 182 230 365
rect 264 321 467 339
rect 264 305 433 321
rect 264 300 298 305
rect 410 287 433 305
rect 410 271 467 287
rect 501 331 535 365
rect 501 315 569 331
rect 264 248 298 266
rect 350 203 425 219
rect 501 207 535 315
rect 603 265 637 451
rect 671 477 705 527
rect 671 427 705 443
rect 767 471 825 487
rect 767 437 775 471
rect 809 437 825 471
rect 767 373 825 437
rect 684 368 825 373
rect 684 357 775 368
rect 718 334 775 357
rect 809 334 825 368
rect 718 323 825 334
rect 684 307 825 323
rect 859 484 893 527
rect 859 364 893 450
rect 938 475 995 491
rect 938 441 943 475
rect 977 441 995 475
rect 938 384 995 441
rect 938 350 943 384
rect 977 350 995 384
rect 938 334 995 350
rect 859 314 893 330
rect 603 249 756 265
rect 603 233 722 249
rect 196 148 237 182
rect 384 169 425 203
rect 350 153 425 169
rect 459 191 535 207
rect 493 157 535 191
rect 35 119 69 127
rect 203 119 237 148
rect 459 141 535 157
rect 574 215 722 233
rect 574 199 756 215
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 574 107 608 199
rect 790 149 825 307
rect 961 149 995 334
rect 203 69 237 85
rect 103 17 169 59
rect 291 59 307 93
rect 341 59 357 93
rect 476 73 500 107
rect 534 73 608 107
rect 767 133 825 149
rect 291 17 357 59
rect 653 72 669 106
rect 703 72 719 106
rect 767 99 775 133
rect 809 99 825 133
rect 767 83 825 99
rect 859 127 893 143
rect 653 17 719 72
rect 859 17 893 93
rect 938 133 995 149
rect 938 99 943 133
rect 977 99 995 133
rect 938 83 995 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 28 244 55 267 0 FreeSans 200 0 0 0 SLEEP_B
port 2 nsew clock input
flabel locali s 366 167 401 203 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 954 357 988 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 954 425 988 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 954 85 988 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 lpflow_inputisolatch_1
flabel comment s 185 283 185 283 0 FreeSans 200 0 0 0 no_jumper_check
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 2376910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2367978
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
