magic
tech sky130A
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_1
timestamp 1694700623
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 6902134
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6901084
<< end >>
