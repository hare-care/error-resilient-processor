VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Top_multiplier
  CLASS BLOCK ;
  FOREIGN Top_multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 90.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.540 10.640 45.140 79.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.040 10.640 67.640 79.120 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END clk
  PIN data_sample
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END data_sample
  PIN error
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 86.000 47.640 90.000 48.240 ;
    END
  END error
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 86.000 44.240 90.000 44.840 ;
    END
  END nrst
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 84.180 78.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 85.030 79.120 ;
      LAYER met2 ;
        RECT 6.990 10.695 85.010 79.065 ;
      LAYER met3 ;
        RECT 4.000 48.640 86.000 79.045 ;
        RECT 4.400 47.240 85.600 48.640 ;
        RECT 4.000 45.240 86.000 47.240 ;
        RECT 4.400 43.840 85.600 45.240 ;
        RECT 4.000 10.715 86.000 43.840 ;
  END
END Top_multiplier
END LIBRARY

