magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 0 0 638 472
<< pmos >>
rect 89 36 119 436
rect 175 36 205 436
rect 261 36 291 436
rect 347 36 377 436
rect 433 36 463 436
rect 519 36 549 436
<< pdiff >>
rect 36 397 89 436
rect 36 363 44 397
rect 78 363 89 397
rect 36 325 89 363
rect 36 291 44 325
rect 78 291 89 325
rect 36 253 89 291
rect 36 219 44 253
rect 78 219 89 253
rect 36 181 89 219
rect 36 147 44 181
rect 78 147 89 181
rect 36 109 89 147
rect 36 75 44 109
rect 78 75 89 109
rect 36 36 89 75
rect 119 397 175 436
rect 119 363 130 397
rect 164 363 175 397
rect 119 325 175 363
rect 119 291 130 325
rect 164 291 175 325
rect 119 253 175 291
rect 119 219 130 253
rect 164 219 175 253
rect 119 181 175 219
rect 119 147 130 181
rect 164 147 175 181
rect 119 109 175 147
rect 119 75 130 109
rect 164 75 175 109
rect 119 36 175 75
rect 205 397 261 436
rect 205 363 216 397
rect 250 363 261 397
rect 205 325 261 363
rect 205 291 216 325
rect 250 291 261 325
rect 205 253 261 291
rect 205 219 216 253
rect 250 219 261 253
rect 205 181 261 219
rect 205 147 216 181
rect 250 147 261 181
rect 205 109 261 147
rect 205 75 216 109
rect 250 75 261 109
rect 205 36 261 75
rect 291 397 347 436
rect 291 363 302 397
rect 336 363 347 397
rect 291 325 347 363
rect 291 291 302 325
rect 336 291 347 325
rect 291 253 347 291
rect 291 219 302 253
rect 336 219 347 253
rect 291 181 347 219
rect 291 147 302 181
rect 336 147 347 181
rect 291 109 347 147
rect 291 75 302 109
rect 336 75 347 109
rect 291 36 347 75
rect 377 397 433 436
rect 377 363 388 397
rect 422 363 433 397
rect 377 325 433 363
rect 377 291 388 325
rect 422 291 433 325
rect 377 253 433 291
rect 377 219 388 253
rect 422 219 433 253
rect 377 181 433 219
rect 377 147 388 181
rect 422 147 433 181
rect 377 109 433 147
rect 377 75 388 109
rect 422 75 433 109
rect 377 36 433 75
rect 463 397 519 436
rect 463 363 474 397
rect 508 363 519 397
rect 463 325 519 363
rect 463 291 474 325
rect 508 291 519 325
rect 463 253 519 291
rect 463 219 474 253
rect 508 219 519 253
rect 463 181 519 219
rect 463 147 474 181
rect 508 147 519 181
rect 463 109 519 147
rect 463 75 474 109
rect 508 75 519 109
rect 463 36 519 75
rect 549 397 602 436
rect 549 363 560 397
rect 594 363 602 397
rect 549 325 602 363
rect 549 291 560 325
rect 594 291 602 325
rect 549 253 602 291
rect 549 219 560 253
rect 594 219 602 253
rect 549 181 602 219
rect 549 147 560 181
rect 594 147 602 181
rect 549 109 602 147
rect 549 75 560 109
rect 594 75 602 109
rect 549 36 602 75
<< pdiffc >>
rect 44 363 78 397
rect 44 291 78 325
rect 44 219 78 253
rect 44 147 78 181
rect 44 75 78 109
rect 130 363 164 397
rect 130 291 164 325
rect 130 219 164 253
rect 130 147 164 181
rect 130 75 164 109
rect 216 363 250 397
rect 216 291 250 325
rect 216 219 250 253
rect 216 147 250 181
rect 216 75 250 109
rect 302 363 336 397
rect 302 291 336 325
rect 302 219 336 253
rect 302 147 336 181
rect 302 75 336 109
rect 388 363 422 397
rect 388 291 422 325
rect 388 219 422 253
rect 388 147 422 181
rect 388 75 422 109
rect 474 363 508 397
rect 474 291 508 325
rect 474 219 508 253
rect 474 147 508 181
rect 474 75 508 109
rect 560 363 594 397
rect 560 291 594 325
rect 560 219 594 253
rect 560 147 594 181
rect 560 75 594 109
<< poly >>
rect 89 519 549 535
rect 89 485 132 519
rect 166 485 200 519
rect 234 485 268 519
rect 302 485 336 519
rect 370 485 404 519
rect 438 485 472 519
rect 506 485 549 519
rect 89 462 549 485
rect 89 436 119 462
rect 175 436 205 462
rect 261 436 291 462
rect 347 436 377 462
rect 433 436 463 462
rect 519 436 549 462
rect 89 10 119 36
rect 175 10 205 36
rect 261 10 291 36
rect 347 10 377 36
rect 433 10 463 36
rect 519 10 549 36
<< polycont >>
rect 132 485 166 519
rect 200 485 234 519
rect 268 485 302 519
rect 336 485 370 519
rect 404 485 438 519
rect 472 485 506 519
<< locali >>
rect 116 519 522 535
rect 116 485 122 519
rect 166 485 194 519
rect 234 485 266 519
rect 302 485 336 519
rect 372 485 404 519
rect 444 485 472 519
rect 516 485 522 519
rect 116 467 522 485
rect 44 397 78 421
rect 44 325 78 363
rect 44 253 78 291
rect 44 181 78 219
rect 44 109 78 147
rect 44 51 78 75
rect 130 397 164 421
rect 130 325 164 363
rect 130 253 164 291
rect 130 181 164 219
rect 130 109 164 147
rect 130 51 164 75
rect 216 397 250 421
rect 216 325 250 363
rect 216 253 250 291
rect 216 181 250 219
rect 216 109 250 147
rect 216 51 250 75
rect 302 397 336 421
rect 302 325 336 363
rect 302 253 336 291
rect 302 181 336 219
rect 302 109 336 147
rect 302 51 336 75
rect 388 397 422 421
rect 388 325 422 363
rect 388 253 422 291
rect 388 181 422 219
rect 388 109 422 147
rect 388 51 422 75
rect 474 397 508 421
rect 474 325 508 363
rect 474 253 508 291
rect 474 181 508 219
rect 474 109 508 147
rect 474 51 508 75
rect 560 397 594 421
rect 560 325 594 363
rect 560 253 594 291
rect 560 181 594 219
rect 560 109 594 147
rect 560 51 594 75
<< viali >>
rect 122 485 132 519
rect 132 485 156 519
rect 194 485 200 519
rect 200 485 228 519
rect 266 485 268 519
rect 268 485 300 519
rect 338 485 370 519
rect 370 485 372 519
rect 410 485 438 519
rect 438 485 444 519
rect 482 485 506 519
rect 506 485 516 519
rect 44 363 78 397
rect 44 291 78 325
rect 44 219 78 253
rect 44 147 78 181
rect 44 75 78 109
rect 130 363 164 397
rect 130 291 164 325
rect 130 219 164 253
rect 130 147 164 181
rect 130 75 164 109
rect 216 363 250 397
rect 216 291 250 325
rect 216 219 250 253
rect 216 147 250 181
rect 216 75 250 109
rect 302 363 336 397
rect 302 291 336 325
rect 302 219 336 253
rect 302 147 336 181
rect 302 75 336 109
rect 388 363 422 397
rect 388 291 422 325
rect 388 219 422 253
rect 388 147 422 181
rect 388 75 422 109
rect 474 363 508 397
rect 474 291 508 325
rect 474 219 508 253
rect 474 147 508 181
rect 474 75 508 109
rect 560 363 594 397
rect 560 291 594 325
rect 560 219 594 253
rect 560 147 594 181
rect 560 75 594 109
<< metal1 >>
rect 110 519 528 531
rect 110 485 122 519
rect 156 485 194 519
rect 228 485 266 519
rect 300 485 338 519
rect 372 485 410 519
rect 444 485 482 519
rect 516 485 528 519
rect 110 473 528 485
rect 38 397 84 421
rect 38 363 44 397
rect 78 363 84 397
rect 38 325 84 363
rect 38 291 44 325
rect 78 291 84 325
rect 38 253 84 291
rect 38 219 44 253
rect 78 219 84 253
rect 38 181 84 219
rect 38 147 44 181
rect 78 147 84 181
rect 38 109 84 147
rect 38 75 44 109
rect 78 75 84 109
rect 38 -29 84 75
rect 121 410 173 421
rect 121 346 173 358
rect 121 291 130 294
rect 164 291 173 294
rect 121 253 173 291
rect 121 219 130 253
rect 164 219 173 253
rect 121 181 173 219
rect 121 147 130 181
rect 164 147 173 181
rect 121 109 173 147
rect 121 75 130 109
rect 164 75 173 109
rect 121 51 173 75
rect 210 397 256 421
rect 210 363 216 397
rect 250 363 256 397
rect 210 325 256 363
rect 210 291 216 325
rect 250 291 256 325
rect 210 253 256 291
rect 210 219 216 253
rect 250 219 256 253
rect 210 181 256 219
rect 210 147 216 181
rect 250 147 256 181
rect 210 109 256 147
rect 210 75 216 109
rect 250 75 256 109
rect 210 -29 256 75
rect 293 410 345 421
rect 293 346 345 358
rect 293 291 302 294
rect 336 291 345 294
rect 293 253 345 291
rect 293 219 302 253
rect 336 219 345 253
rect 293 181 345 219
rect 293 147 302 181
rect 336 147 345 181
rect 293 109 345 147
rect 293 75 302 109
rect 336 75 345 109
rect 293 51 345 75
rect 382 397 428 421
rect 382 363 388 397
rect 422 363 428 397
rect 382 325 428 363
rect 382 291 388 325
rect 422 291 428 325
rect 382 253 428 291
rect 382 219 388 253
rect 422 219 428 253
rect 382 181 428 219
rect 382 147 388 181
rect 422 147 428 181
rect 382 109 428 147
rect 382 75 388 109
rect 422 75 428 109
rect 382 -29 428 75
rect 465 410 517 421
rect 465 346 517 358
rect 465 291 474 294
rect 508 291 517 294
rect 465 253 517 291
rect 465 219 474 253
rect 508 219 517 253
rect 465 181 517 219
rect 465 147 474 181
rect 508 147 517 181
rect 465 109 517 147
rect 465 75 474 109
rect 508 75 517 109
rect 465 51 517 75
rect 554 397 600 421
rect 554 363 560 397
rect 594 363 600 397
rect 554 325 600 363
rect 554 291 560 325
rect 594 291 600 325
rect 554 253 600 291
rect 554 219 560 253
rect 594 219 600 253
rect 554 181 600 219
rect 554 147 560 181
rect 594 147 600 181
rect 554 109 600 147
rect 554 75 560 109
rect 594 75 600 109
rect 554 -29 600 75
rect 38 -89 600 -29
<< via1 >>
rect 121 397 173 410
rect 121 363 130 397
rect 130 363 164 397
rect 164 363 173 397
rect 121 358 173 363
rect 121 325 173 346
rect 121 294 130 325
rect 130 294 164 325
rect 164 294 173 325
rect 293 397 345 410
rect 293 363 302 397
rect 302 363 336 397
rect 336 363 345 397
rect 293 358 345 363
rect 293 325 345 346
rect 293 294 302 325
rect 302 294 336 325
rect 336 294 345 325
rect 465 397 517 410
rect 465 363 474 397
rect 474 363 508 397
rect 508 363 517 397
rect 465 358 517 363
rect 465 325 517 346
rect 465 294 474 325
rect 474 294 508 325
rect 508 294 517 325
<< metal2 >>
rect 114 420 180 429
rect 114 364 119 420
rect 175 364 180 420
rect 114 358 121 364
rect 173 358 180 364
rect 114 346 180 358
rect 114 340 121 346
rect 173 340 180 346
rect 114 284 119 340
rect 175 284 180 340
rect 114 275 180 284
rect 286 420 352 429
rect 286 364 291 420
rect 347 364 352 420
rect 286 358 293 364
rect 345 358 352 364
rect 286 346 352 358
rect 286 340 293 346
rect 345 340 352 346
rect 286 284 291 340
rect 347 284 352 340
rect 286 275 352 284
rect 458 420 524 429
rect 458 364 463 420
rect 519 364 524 420
rect 458 358 465 364
rect 517 358 524 364
rect 458 346 524 358
rect 458 340 465 346
rect 517 340 524 346
rect 458 284 463 340
rect 519 284 524 340
rect 458 275 524 284
<< via2 >>
rect 119 410 175 420
rect 119 364 121 410
rect 121 364 173 410
rect 173 364 175 410
rect 119 294 121 340
rect 121 294 173 340
rect 173 294 175 340
rect 119 284 175 294
rect 291 410 347 420
rect 291 364 293 410
rect 293 364 345 410
rect 345 364 347 410
rect 291 294 293 340
rect 293 294 345 340
rect 345 294 347 340
rect 291 284 347 294
rect 463 410 519 420
rect 463 364 465 410
rect 465 364 517 410
rect 517 364 519 410
rect 463 294 465 340
rect 465 294 517 340
rect 517 294 519 340
rect 463 284 519 294
<< metal3 >>
rect 114 420 524 429
rect 114 364 119 420
rect 175 364 291 420
rect 347 364 463 420
rect 519 364 524 420
rect 114 363 524 364
rect 114 340 180 363
rect 114 284 119 340
rect 175 284 180 340
rect 114 275 180 284
rect 286 340 352 363
rect 286 284 291 340
rect 347 284 352 340
rect 286 275 352 284
rect 458 340 524 363
rect 458 284 463 340
rect 519 284 524 340
rect 458 275 524 284
<< labels >>
flabel metal3 s 114 363 524 429 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 110 473 528 531 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel metal1 s 38 -89 600 -29 0 FreeSans 400 0 0 0 SOURCE
port 4 nsew
flabel nwell s 85 463 88 471 0 FreeSans 400 0 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 9187710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9175750
string path 1.525 10.525 1.525 -2.225 
<< end >>
