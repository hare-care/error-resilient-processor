magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal1 >>
rect 1500 1959 1530 2011
rect 1702 1959 1732 2011
rect 2748 1959 2778 2011
rect 2950 1959 2980 2011
rect 3996 1959 4026 2011
rect 4198 1959 4228 2011
rect 5244 1959 5274 2011
rect 5446 1959 5476 2011
rect 6492 1959 6522 2011
rect 6694 1959 6724 2011
rect 7740 1959 7770 2011
rect 7942 1959 7972 2011
rect 8988 1959 9018 2011
rect 9190 1959 9220 2011
rect 10236 1959 10266 2011
rect 10438 1959 10468 2011
rect 11484 1959 11514 2011
rect 11686 1959 11716 2011
rect 12732 1959 12762 2011
rect 12934 1959 12964 2011
rect 13980 1959 14010 2011
rect 14182 1959 14212 2011
rect 15228 1959 15258 2011
rect 15430 1959 15460 2011
rect 16476 1959 16506 2011
rect 16678 1959 16708 2011
rect 17724 1959 17754 2011
rect 17926 1959 17956 2011
rect 18972 1959 19002 2011
rect 19174 1959 19204 2011
rect 20220 1959 20250 2011
rect 20422 1959 20452 2011
rect 21468 1959 21498 2011
rect 21670 1959 21700 2011
rect 22716 1959 22746 2011
rect 22918 1959 22948 2011
rect 23964 1959 23994 2011
rect 24166 1959 24196 2011
rect 25212 1959 25242 2011
rect 25414 1959 25444 2011
rect 26460 1959 26490 2011
rect 26662 1959 26692 2011
rect 27708 1959 27738 2011
rect 27910 1959 27940 2011
rect 28956 1959 28986 2011
rect 29158 1959 29188 2011
rect 30204 1959 30234 2011
rect 30406 1959 30436 2011
rect 31452 1959 31482 2011
rect 31654 1959 31684 2011
rect 32700 1959 32730 2011
rect 32902 1959 32932 2011
rect 33948 1959 33978 2011
rect 34150 1959 34180 2011
rect 35196 1959 35226 2011
rect 35398 1959 35428 2011
rect 36444 1959 36474 2011
rect 36646 1959 36676 2011
rect 37692 1959 37722 2011
rect 37894 1959 37924 2011
rect 38940 1959 38970 2011
rect 39142 1959 39172 2011
rect 40188 1959 40218 2011
rect 40390 1959 40420 2011
rect 1615 1604 1667 1610
rect 1615 1546 1667 1552
rect 2863 1604 2915 1610
rect 2863 1546 2915 1552
rect 4111 1604 4163 1610
rect 4111 1546 4163 1552
rect 5359 1604 5411 1610
rect 5359 1546 5411 1552
rect 6607 1604 6659 1610
rect 6607 1546 6659 1552
rect 7855 1604 7907 1610
rect 7855 1546 7907 1552
rect 9103 1604 9155 1610
rect 9103 1546 9155 1552
rect 10351 1604 10403 1610
rect 10351 1546 10403 1552
rect 11599 1604 11651 1610
rect 11599 1546 11651 1552
rect 12847 1604 12899 1610
rect 12847 1546 12899 1552
rect 14095 1604 14147 1610
rect 14095 1546 14147 1552
rect 15343 1604 15395 1610
rect 15343 1546 15395 1552
rect 16591 1604 16643 1610
rect 16591 1546 16643 1552
rect 17839 1604 17891 1610
rect 17839 1546 17891 1552
rect 19087 1604 19139 1610
rect 19087 1546 19139 1552
rect 20335 1604 20387 1610
rect 20335 1546 20387 1552
rect 21583 1604 21635 1610
rect 21583 1546 21635 1552
rect 22831 1604 22883 1610
rect 22831 1546 22883 1552
rect 24079 1604 24131 1610
rect 24079 1546 24131 1552
rect 25327 1604 25379 1610
rect 25327 1546 25379 1552
rect 26575 1604 26627 1610
rect 26575 1546 26627 1552
rect 27823 1604 27875 1610
rect 27823 1546 27875 1552
rect 29071 1604 29123 1610
rect 29071 1546 29123 1552
rect 30319 1604 30371 1610
rect 30319 1546 30371 1552
rect 31567 1604 31619 1610
rect 31567 1546 31619 1552
rect 32815 1604 32867 1610
rect 32815 1546 32867 1552
rect 34063 1604 34115 1610
rect 34063 1546 34115 1552
rect 35311 1604 35363 1610
rect 35311 1546 35363 1552
rect 36559 1604 36611 1610
rect 36559 1546 36611 1552
rect 37807 1604 37859 1610
rect 37807 1546 37859 1552
rect 39055 1604 39107 1610
rect 39055 1546 39107 1552
rect 40303 1604 40355 1610
rect 40303 1546 40355 1552
rect 1604 1167 1656 1173
rect 1604 1109 1656 1115
rect 2852 1167 2904 1173
rect 2852 1109 2904 1115
rect 4100 1167 4152 1173
rect 4100 1109 4152 1115
rect 5348 1167 5400 1173
rect 5348 1109 5400 1115
rect 6596 1167 6648 1173
rect 6596 1109 6648 1115
rect 7844 1167 7896 1173
rect 7844 1109 7896 1115
rect 9092 1167 9144 1173
rect 9092 1109 9144 1115
rect 10340 1167 10392 1173
rect 10340 1109 10392 1115
rect 11588 1167 11640 1173
rect 11588 1109 11640 1115
rect 12836 1167 12888 1173
rect 12836 1109 12888 1115
rect 14084 1167 14136 1173
rect 14084 1109 14136 1115
rect 15332 1167 15384 1173
rect 15332 1109 15384 1115
rect 16580 1167 16632 1173
rect 16580 1109 16632 1115
rect 17828 1167 17880 1173
rect 17828 1109 17880 1115
rect 19076 1167 19128 1173
rect 19076 1109 19128 1115
rect 20324 1167 20376 1173
rect 20324 1109 20376 1115
rect 21572 1167 21624 1173
rect 21572 1109 21624 1115
rect 22820 1167 22872 1173
rect 22820 1109 22872 1115
rect 24068 1167 24120 1173
rect 24068 1109 24120 1115
rect 25316 1167 25368 1173
rect 25316 1109 25368 1115
rect 26564 1167 26616 1173
rect 26564 1109 26616 1115
rect 27812 1167 27864 1173
rect 27812 1109 27864 1115
rect 29060 1167 29112 1173
rect 29060 1109 29112 1115
rect 30308 1167 30360 1173
rect 30308 1109 30360 1115
rect 31556 1167 31608 1173
rect 31556 1109 31608 1115
rect 32804 1167 32856 1173
rect 32804 1109 32856 1115
rect 34052 1167 34104 1173
rect 34052 1109 34104 1115
rect 35300 1167 35352 1173
rect 35300 1109 35352 1115
rect 36548 1167 36600 1173
rect 36548 1109 36600 1115
rect 37796 1167 37848 1173
rect 37796 1109 37848 1115
rect 39044 1167 39096 1173
rect 39044 1109 39096 1115
rect 40292 1167 40344 1173
rect 40292 1109 40344 1115
rect 1725 836 1777 842
rect 1725 778 1777 784
rect 2973 836 3025 842
rect 2973 778 3025 784
rect 4221 836 4273 842
rect 4221 778 4273 784
rect 5469 836 5521 842
rect 5469 778 5521 784
rect 6717 836 6769 842
rect 6717 778 6769 784
rect 7965 836 8017 842
rect 7965 778 8017 784
rect 9213 836 9265 842
rect 9213 778 9265 784
rect 10461 836 10513 842
rect 10461 778 10513 784
rect 11709 836 11761 842
rect 11709 778 11761 784
rect 12957 836 13009 842
rect 12957 778 13009 784
rect 14205 836 14257 842
rect 14205 778 14257 784
rect 15453 836 15505 842
rect 15453 778 15505 784
rect 16701 836 16753 842
rect 16701 778 16753 784
rect 17949 836 18001 842
rect 17949 778 18001 784
rect 19197 836 19249 842
rect 19197 778 19249 784
rect 20445 836 20497 842
rect 20445 778 20497 784
rect 21693 836 21745 842
rect 21693 778 21745 784
rect 22941 836 22993 842
rect 22941 778 22993 784
rect 24189 836 24241 842
rect 24189 778 24241 784
rect 25437 836 25489 842
rect 25437 778 25489 784
rect 26685 836 26737 842
rect 26685 778 26737 784
rect 27933 836 27985 842
rect 27933 778 27985 784
rect 29181 836 29233 842
rect 29181 778 29233 784
rect 30429 836 30481 842
rect 30429 778 30481 784
rect 31677 836 31729 842
rect 31677 778 31729 784
rect 32925 836 32977 842
rect 32925 778 32977 784
rect 34173 836 34225 842
rect 34173 778 34225 784
rect 35421 836 35473 842
rect 35421 778 35473 784
rect 36669 836 36721 842
rect 36669 778 36721 784
rect 37917 836 37969 842
rect 37917 778 37969 784
rect 39165 836 39217 842
rect 39165 778 39217 784
rect 40413 836 40465 842
rect 40413 778 40465 784
rect 1610 633 1662 639
rect 1610 575 1662 581
rect 2858 633 2910 639
rect 2858 575 2910 581
rect 4106 633 4158 639
rect 4106 575 4158 581
rect 5354 633 5406 639
rect 5354 575 5406 581
rect 6602 633 6654 639
rect 6602 575 6654 581
rect 7850 633 7902 639
rect 7850 575 7902 581
rect 9098 633 9150 639
rect 9098 575 9150 581
rect 10346 633 10398 639
rect 10346 575 10398 581
rect 11594 633 11646 639
rect 11594 575 11646 581
rect 12842 633 12894 639
rect 12842 575 12894 581
rect 14090 633 14142 639
rect 14090 575 14142 581
rect 15338 633 15390 639
rect 15338 575 15390 581
rect 16586 633 16638 639
rect 16586 575 16638 581
rect 17834 633 17886 639
rect 17834 575 17886 581
rect 19082 633 19134 639
rect 19082 575 19134 581
rect 20330 633 20382 639
rect 20330 575 20382 581
rect 21578 633 21630 639
rect 21578 575 21630 581
rect 22826 633 22878 639
rect 22826 575 22878 581
rect 24074 633 24126 639
rect 24074 575 24126 581
rect 25322 633 25374 639
rect 25322 575 25374 581
rect 26570 633 26622 639
rect 26570 575 26622 581
rect 27818 633 27870 639
rect 27818 575 27870 581
rect 29066 633 29118 639
rect 29066 575 29118 581
rect 30314 633 30366 639
rect 30314 575 30366 581
rect 31562 633 31614 639
rect 31562 575 31614 581
rect 32810 633 32862 639
rect 32810 575 32862 581
rect 34058 633 34110 639
rect 34058 575 34110 581
rect 35306 633 35358 639
rect 35306 575 35358 581
rect 36554 633 36606 639
rect 36554 575 36606 581
rect 37802 633 37854 639
rect 37802 575 37854 581
rect 39050 633 39102 639
rect 39050 575 39102 581
rect 40298 633 40350 639
rect 40298 575 40350 581
rect 1624 217 1676 223
rect 1624 159 1676 165
rect 2872 217 2924 223
rect 2872 159 2924 165
rect 4120 217 4172 223
rect 4120 159 4172 165
rect 5368 217 5420 223
rect 5368 159 5420 165
rect 6616 217 6668 223
rect 6616 159 6668 165
rect 7864 217 7916 223
rect 7864 159 7916 165
rect 9112 217 9164 223
rect 9112 159 9164 165
rect 10360 217 10412 223
rect 10360 159 10412 165
rect 11608 217 11660 223
rect 11608 159 11660 165
rect 12856 217 12908 223
rect 12856 159 12908 165
rect 14104 217 14156 223
rect 14104 159 14156 165
rect 15352 217 15404 223
rect 15352 159 15404 165
rect 16600 217 16652 223
rect 16600 159 16652 165
rect 17848 217 17900 223
rect 17848 159 17900 165
rect 19096 217 19148 223
rect 19096 159 19148 165
rect 20344 217 20396 223
rect 20344 159 20396 165
rect 21592 217 21644 223
rect 21592 159 21644 165
rect 22840 217 22892 223
rect 22840 159 22892 165
rect 24088 217 24140 223
rect 24088 159 24140 165
rect 25336 217 25388 223
rect 25336 159 25388 165
rect 26584 217 26636 223
rect 26584 159 26636 165
rect 27832 217 27884 223
rect 27832 159 27884 165
rect 29080 217 29132 223
rect 29080 159 29132 165
rect 30328 217 30380 223
rect 30328 159 30380 165
rect 31576 217 31628 223
rect 31576 159 31628 165
rect 32824 217 32876 223
rect 32824 159 32876 165
rect 34072 217 34124 223
rect 34072 159 34124 165
rect 35320 217 35372 223
rect 35320 159 35372 165
rect 36568 217 36620 223
rect 36568 159 36620 165
rect 37816 217 37868 223
rect 37816 159 37868 165
rect 39064 217 39116 223
rect 39064 159 39116 165
rect 40312 217 40364 223
rect 40312 159 40364 165
rect 1473 94 10833 128
rect 11457 94 20817 128
rect 21441 94 30801 128
rect 31425 94 40785 128
rect 1629 4 1689 60
rect 2877 4 2937 60
rect 4125 4 4185 60
rect 5373 4 5433 60
rect 6621 4 6681 60
rect 7869 4 7929 60
rect 9117 4 9177 60
rect 10365 4 10425 60
rect 11613 4 11673 60
rect 12861 4 12921 60
rect 14109 4 14169 60
rect 15357 4 15417 60
rect 16605 4 16665 60
rect 17853 4 17913 60
rect 19101 4 19161 60
rect 20349 4 20409 60
rect 21597 4 21657 60
rect 22845 4 22905 60
rect 24093 4 24153 60
rect 25341 4 25401 60
rect 26589 4 26649 60
rect 27837 4 27897 60
rect 29085 4 29145 60
rect 30333 4 30393 60
rect 31581 4 31641 60
rect 32829 4 32889 60
rect 34077 4 34137 60
rect 35325 4 35385 60
rect 36573 4 36633 60
rect 37821 4 37881 60
rect 39069 4 39129 60
rect 40317 4 40377 60
<< via1 >>
rect 1615 1552 1667 1604
rect 2863 1552 2915 1604
rect 4111 1552 4163 1604
rect 5359 1552 5411 1604
rect 6607 1552 6659 1604
rect 7855 1552 7907 1604
rect 9103 1552 9155 1604
rect 10351 1552 10403 1604
rect 11599 1552 11651 1604
rect 12847 1552 12899 1604
rect 14095 1552 14147 1604
rect 15343 1552 15395 1604
rect 16591 1552 16643 1604
rect 17839 1552 17891 1604
rect 19087 1552 19139 1604
rect 20335 1552 20387 1604
rect 21583 1552 21635 1604
rect 22831 1552 22883 1604
rect 24079 1552 24131 1604
rect 25327 1552 25379 1604
rect 26575 1552 26627 1604
rect 27823 1552 27875 1604
rect 29071 1552 29123 1604
rect 30319 1552 30371 1604
rect 31567 1552 31619 1604
rect 32815 1552 32867 1604
rect 34063 1552 34115 1604
rect 35311 1552 35363 1604
rect 36559 1552 36611 1604
rect 37807 1552 37859 1604
rect 39055 1552 39107 1604
rect 40303 1552 40355 1604
rect 1604 1115 1656 1167
rect 2852 1115 2904 1167
rect 4100 1115 4152 1167
rect 5348 1115 5400 1167
rect 6596 1115 6648 1167
rect 7844 1115 7896 1167
rect 9092 1115 9144 1167
rect 10340 1115 10392 1167
rect 11588 1115 11640 1167
rect 12836 1115 12888 1167
rect 14084 1115 14136 1167
rect 15332 1115 15384 1167
rect 16580 1115 16632 1167
rect 17828 1115 17880 1167
rect 19076 1115 19128 1167
rect 20324 1115 20376 1167
rect 21572 1115 21624 1167
rect 22820 1115 22872 1167
rect 24068 1115 24120 1167
rect 25316 1115 25368 1167
rect 26564 1115 26616 1167
rect 27812 1115 27864 1167
rect 29060 1115 29112 1167
rect 30308 1115 30360 1167
rect 31556 1115 31608 1167
rect 32804 1115 32856 1167
rect 34052 1115 34104 1167
rect 35300 1115 35352 1167
rect 36548 1115 36600 1167
rect 37796 1115 37848 1167
rect 39044 1115 39096 1167
rect 40292 1115 40344 1167
rect 1725 784 1777 836
rect 2973 784 3025 836
rect 4221 784 4273 836
rect 5469 784 5521 836
rect 6717 784 6769 836
rect 7965 784 8017 836
rect 9213 784 9265 836
rect 10461 784 10513 836
rect 11709 784 11761 836
rect 12957 784 13009 836
rect 14205 784 14257 836
rect 15453 784 15505 836
rect 16701 784 16753 836
rect 17949 784 18001 836
rect 19197 784 19249 836
rect 20445 784 20497 836
rect 21693 784 21745 836
rect 22941 784 22993 836
rect 24189 784 24241 836
rect 25437 784 25489 836
rect 26685 784 26737 836
rect 27933 784 27985 836
rect 29181 784 29233 836
rect 30429 784 30481 836
rect 31677 784 31729 836
rect 32925 784 32977 836
rect 34173 784 34225 836
rect 35421 784 35473 836
rect 36669 784 36721 836
rect 37917 784 37969 836
rect 39165 784 39217 836
rect 40413 784 40465 836
rect 1610 581 1662 633
rect 2858 581 2910 633
rect 4106 581 4158 633
rect 5354 581 5406 633
rect 6602 581 6654 633
rect 7850 581 7902 633
rect 9098 581 9150 633
rect 10346 581 10398 633
rect 11594 581 11646 633
rect 12842 581 12894 633
rect 14090 581 14142 633
rect 15338 581 15390 633
rect 16586 581 16638 633
rect 17834 581 17886 633
rect 19082 581 19134 633
rect 20330 581 20382 633
rect 21578 581 21630 633
rect 22826 581 22878 633
rect 24074 581 24126 633
rect 25322 581 25374 633
rect 26570 581 26622 633
rect 27818 581 27870 633
rect 29066 581 29118 633
rect 30314 581 30366 633
rect 31562 581 31614 633
rect 32810 581 32862 633
rect 34058 581 34110 633
rect 35306 581 35358 633
rect 36554 581 36606 633
rect 37802 581 37854 633
rect 39050 581 39102 633
rect 40298 581 40350 633
rect 1624 165 1676 217
rect 2872 165 2924 217
rect 4120 165 4172 217
rect 5368 165 5420 217
rect 6616 165 6668 217
rect 7864 165 7916 217
rect 9112 165 9164 217
rect 10360 165 10412 217
rect 11608 165 11660 217
rect 12856 165 12908 217
rect 14104 165 14156 217
rect 15352 165 15404 217
rect 16600 165 16652 217
rect 17848 165 17900 217
rect 19096 165 19148 217
rect 20344 165 20396 217
rect 21592 165 21644 217
rect 22840 165 22892 217
rect 24088 165 24140 217
rect 25336 165 25388 217
rect 26584 165 26636 217
rect 27832 165 27884 217
rect 29080 165 29132 217
rect 30328 165 30380 217
rect 31576 165 31628 217
rect 32824 165 32876 217
rect 34072 165 34124 217
rect 35320 165 35372 217
rect 36568 165 36620 217
rect 37816 165 37868 217
rect 39064 165 39116 217
rect 40312 165 40364 217
<< metal2 >>
rect 1613 1606 1669 1615
rect 1613 1541 1669 1550
rect 2861 1606 2917 1615
rect 2861 1541 2917 1550
rect 4109 1606 4165 1615
rect 4109 1541 4165 1550
rect 5357 1606 5413 1615
rect 5357 1541 5413 1550
rect 6605 1606 6661 1615
rect 6605 1541 6661 1550
rect 7853 1606 7909 1615
rect 7853 1541 7909 1550
rect 9101 1606 9157 1615
rect 9101 1541 9157 1550
rect 10349 1606 10405 1615
rect 10349 1541 10405 1550
rect 11597 1606 11653 1615
rect 11597 1541 11653 1550
rect 12845 1606 12901 1615
rect 12845 1541 12901 1550
rect 14093 1606 14149 1615
rect 14093 1541 14149 1550
rect 15341 1606 15397 1615
rect 15341 1541 15397 1550
rect 16589 1606 16645 1615
rect 16589 1541 16645 1550
rect 17837 1606 17893 1615
rect 17837 1541 17893 1550
rect 19085 1606 19141 1615
rect 19085 1541 19141 1550
rect 20333 1606 20389 1615
rect 20333 1541 20389 1550
rect 21581 1606 21637 1615
rect 21581 1541 21637 1550
rect 22829 1606 22885 1615
rect 22829 1541 22885 1550
rect 24077 1606 24133 1615
rect 24077 1541 24133 1550
rect 25325 1606 25381 1615
rect 25325 1541 25381 1550
rect 26573 1606 26629 1615
rect 26573 1541 26629 1550
rect 27821 1606 27877 1615
rect 27821 1541 27877 1550
rect 29069 1606 29125 1615
rect 29069 1541 29125 1550
rect 30317 1606 30373 1615
rect 30317 1541 30373 1550
rect 31565 1606 31621 1615
rect 31565 1541 31621 1550
rect 32813 1606 32869 1615
rect 32813 1541 32869 1550
rect 34061 1606 34117 1615
rect 34061 1541 34117 1550
rect 35309 1606 35365 1615
rect 35309 1541 35365 1550
rect 36557 1606 36613 1615
rect 36557 1541 36613 1550
rect 37805 1606 37861 1615
rect 37805 1541 37861 1550
rect 39053 1606 39109 1615
rect 39053 1541 39109 1550
rect 40301 1606 40357 1615
rect 40301 1541 40357 1550
rect 1602 1169 1658 1178
rect 1602 1104 1658 1113
rect 2850 1169 2906 1178
rect 2850 1104 2906 1113
rect 4098 1169 4154 1178
rect 4098 1104 4154 1113
rect 5346 1169 5402 1178
rect 5346 1104 5402 1113
rect 6594 1169 6650 1178
rect 6594 1104 6650 1113
rect 7842 1169 7898 1178
rect 7842 1104 7898 1113
rect 9090 1169 9146 1178
rect 9090 1104 9146 1113
rect 10338 1169 10394 1178
rect 10338 1104 10394 1113
rect 11586 1169 11642 1178
rect 11586 1104 11642 1113
rect 12834 1169 12890 1178
rect 12834 1104 12890 1113
rect 14082 1169 14138 1178
rect 14082 1104 14138 1113
rect 15330 1169 15386 1178
rect 15330 1104 15386 1113
rect 16578 1169 16634 1178
rect 16578 1104 16634 1113
rect 17826 1169 17882 1178
rect 17826 1104 17882 1113
rect 19074 1169 19130 1178
rect 19074 1104 19130 1113
rect 20322 1169 20378 1178
rect 20322 1104 20378 1113
rect 21570 1169 21626 1178
rect 21570 1104 21626 1113
rect 22818 1169 22874 1178
rect 22818 1104 22874 1113
rect 24066 1169 24122 1178
rect 24066 1104 24122 1113
rect 25314 1169 25370 1178
rect 25314 1104 25370 1113
rect 26562 1169 26618 1178
rect 26562 1104 26618 1113
rect 27810 1169 27866 1178
rect 27810 1104 27866 1113
rect 29058 1169 29114 1178
rect 29058 1104 29114 1113
rect 30306 1169 30362 1178
rect 30306 1104 30362 1113
rect 31554 1169 31610 1178
rect 31554 1104 31610 1113
rect 32802 1169 32858 1178
rect 32802 1104 32858 1113
rect 34050 1169 34106 1178
rect 34050 1104 34106 1113
rect 35298 1169 35354 1178
rect 35298 1104 35354 1113
rect 36546 1169 36602 1178
rect 36546 1104 36602 1113
rect 37794 1169 37850 1178
rect 37794 1104 37850 1113
rect 39042 1169 39098 1178
rect 39042 1104 39098 1113
rect 40290 1169 40346 1178
rect 40290 1104 40346 1113
rect 1723 837 1779 846
rect 1723 772 1779 781
rect 2971 837 3027 846
rect 2971 772 3027 781
rect 4219 837 4275 846
rect 4219 772 4275 781
rect 5467 837 5523 846
rect 5467 772 5523 781
rect 6715 837 6771 846
rect 6715 772 6771 781
rect 7963 837 8019 846
rect 7963 772 8019 781
rect 9211 837 9267 846
rect 9211 772 9267 781
rect 10459 837 10515 846
rect 10459 772 10515 781
rect 11707 837 11763 846
rect 11707 772 11763 781
rect 12955 837 13011 846
rect 12955 772 13011 781
rect 14203 837 14259 846
rect 14203 772 14259 781
rect 15451 837 15507 846
rect 15451 772 15507 781
rect 16699 837 16755 846
rect 16699 772 16755 781
rect 17947 837 18003 846
rect 17947 772 18003 781
rect 19195 837 19251 846
rect 19195 772 19251 781
rect 20443 837 20499 846
rect 20443 772 20499 781
rect 21691 837 21747 846
rect 21691 772 21747 781
rect 22939 837 22995 846
rect 22939 772 22995 781
rect 24187 837 24243 846
rect 24187 772 24243 781
rect 25435 837 25491 846
rect 25435 772 25491 781
rect 26683 837 26739 846
rect 26683 772 26739 781
rect 27931 837 27987 846
rect 27931 772 27987 781
rect 29179 837 29235 846
rect 29179 772 29235 781
rect 30427 837 30483 846
rect 30427 772 30483 781
rect 31675 837 31731 846
rect 31675 772 31731 781
rect 32923 837 32979 846
rect 32923 772 32979 781
rect 34171 837 34227 846
rect 34171 772 34227 781
rect 35419 837 35475 846
rect 35419 772 35475 781
rect 36667 837 36723 846
rect 36667 772 36723 781
rect 37915 837 37971 846
rect 37915 772 37971 781
rect 39163 837 39219 846
rect 39163 772 39219 781
rect 40411 837 40467 846
rect 40411 772 40467 781
rect 1608 635 1664 644
rect 1608 570 1664 579
rect 2856 635 2912 644
rect 2856 570 2912 579
rect 4104 635 4160 644
rect 4104 570 4160 579
rect 5352 635 5408 644
rect 5352 570 5408 579
rect 6600 635 6656 644
rect 6600 570 6656 579
rect 7848 635 7904 644
rect 7848 570 7904 579
rect 9096 635 9152 644
rect 9096 570 9152 579
rect 10344 635 10400 644
rect 10344 570 10400 579
rect 11592 635 11648 644
rect 11592 570 11648 579
rect 12840 635 12896 644
rect 12840 570 12896 579
rect 14088 635 14144 644
rect 14088 570 14144 579
rect 15336 635 15392 644
rect 15336 570 15392 579
rect 16584 635 16640 644
rect 16584 570 16640 579
rect 17832 635 17888 644
rect 17832 570 17888 579
rect 19080 635 19136 644
rect 19080 570 19136 579
rect 20328 635 20384 644
rect 20328 570 20384 579
rect 21576 635 21632 644
rect 21576 570 21632 579
rect 22824 635 22880 644
rect 22824 570 22880 579
rect 24072 635 24128 644
rect 24072 570 24128 579
rect 25320 635 25376 644
rect 25320 570 25376 579
rect 26568 635 26624 644
rect 26568 570 26624 579
rect 27816 635 27872 644
rect 27816 570 27872 579
rect 29064 635 29120 644
rect 29064 570 29120 579
rect 30312 635 30368 644
rect 30312 570 30368 579
rect 31560 635 31616 644
rect 31560 570 31616 579
rect 32808 635 32864 644
rect 32808 570 32864 579
rect 34056 635 34112 644
rect 34056 570 34112 579
rect 35304 635 35360 644
rect 35304 570 35360 579
rect 36552 635 36608 644
rect 36552 570 36608 579
rect 37800 635 37856 644
rect 37800 570 37856 579
rect 39048 635 39104 644
rect 39048 570 39104 579
rect 40296 635 40352 644
rect 40296 570 40352 579
rect 1622 219 1678 228
rect 1622 154 1678 163
rect 2870 219 2926 228
rect 2870 154 2926 163
rect 4118 219 4174 228
rect 4118 154 4174 163
rect 5366 219 5422 228
rect 5366 154 5422 163
rect 6614 219 6670 228
rect 6614 154 6670 163
rect 7862 219 7918 228
rect 7862 154 7918 163
rect 9110 219 9166 228
rect 9110 154 9166 163
rect 10358 219 10414 228
rect 10358 154 10414 163
rect 11606 219 11662 228
rect 11606 154 11662 163
rect 12854 219 12910 228
rect 12854 154 12910 163
rect 14102 219 14158 228
rect 14102 154 14158 163
rect 15350 219 15406 228
rect 15350 154 15406 163
rect 16598 219 16654 228
rect 16598 154 16654 163
rect 17846 219 17902 228
rect 17846 154 17902 163
rect 19094 219 19150 228
rect 19094 154 19150 163
rect 20342 219 20398 228
rect 20342 154 20398 163
rect 21590 219 21646 228
rect 21590 154 21646 163
rect 22838 219 22894 228
rect 22838 154 22894 163
rect 24086 219 24142 228
rect 24086 154 24142 163
rect 25334 219 25390 228
rect 25334 154 25390 163
rect 26582 219 26638 228
rect 26582 154 26638 163
rect 27830 219 27886 228
rect 27830 154 27886 163
rect 29078 219 29134 228
rect 29078 154 29134 163
rect 30326 219 30382 228
rect 30326 154 30382 163
rect 31574 219 31630 228
rect 31574 154 31630 163
rect 32822 219 32878 228
rect 32822 154 32878 163
rect 34070 219 34126 228
rect 34070 154 34126 163
rect 35318 219 35374 228
rect 35318 154 35374 163
rect 36566 219 36622 228
rect 36566 154 36622 163
rect 37814 219 37870 228
rect 37814 154 37870 163
rect 39062 219 39118 228
rect 39062 154 39118 163
rect 40310 219 40366 228
rect 40310 154 40366 163
<< via2 >>
rect 1613 1604 1669 1606
rect 1613 1552 1615 1604
rect 1615 1552 1667 1604
rect 1667 1552 1669 1604
rect 1613 1550 1669 1552
rect 2861 1604 2917 1606
rect 2861 1552 2863 1604
rect 2863 1552 2915 1604
rect 2915 1552 2917 1604
rect 2861 1550 2917 1552
rect 4109 1604 4165 1606
rect 4109 1552 4111 1604
rect 4111 1552 4163 1604
rect 4163 1552 4165 1604
rect 4109 1550 4165 1552
rect 5357 1604 5413 1606
rect 5357 1552 5359 1604
rect 5359 1552 5411 1604
rect 5411 1552 5413 1604
rect 5357 1550 5413 1552
rect 6605 1604 6661 1606
rect 6605 1552 6607 1604
rect 6607 1552 6659 1604
rect 6659 1552 6661 1604
rect 6605 1550 6661 1552
rect 7853 1604 7909 1606
rect 7853 1552 7855 1604
rect 7855 1552 7907 1604
rect 7907 1552 7909 1604
rect 7853 1550 7909 1552
rect 9101 1604 9157 1606
rect 9101 1552 9103 1604
rect 9103 1552 9155 1604
rect 9155 1552 9157 1604
rect 9101 1550 9157 1552
rect 10349 1604 10405 1606
rect 10349 1552 10351 1604
rect 10351 1552 10403 1604
rect 10403 1552 10405 1604
rect 10349 1550 10405 1552
rect 11597 1604 11653 1606
rect 11597 1552 11599 1604
rect 11599 1552 11651 1604
rect 11651 1552 11653 1604
rect 11597 1550 11653 1552
rect 12845 1604 12901 1606
rect 12845 1552 12847 1604
rect 12847 1552 12899 1604
rect 12899 1552 12901 1604
rect 12845 1550 12901 1552
rect 14093 1604 14149 1606
rect 14093 1552 14095 1604
rect 14095 1552 14147 1604
rect 14147 1552 14149 1604
rect 14093 1550 14149 1552
rect 15341 1604 15397 1606
rect 15341 1552 15343 1604
rect 15343 1552 15395 1604
rect 15395 1552 15397 1604
rect 15341 1550 15397 1552
rect 16589 1604 16645 1606
rect 16589 1552 16591 1604
rect 16591 1552 16643 1604
rect 16643 1552 16645 1604
rect 16589 1550 16645 1552
rect 17837 1604 17893 1606
rect 17837 1552 17839 1604
rect 17839 1552 17891 1604
rect 17891 1552 17893 1604
rect 17837 1550 17893 1552
rect 19085 1604 19141 1606
rect 19085 1552 19087 1604
rect 19087 1552 19139 1604
rect 19139 1552 19141 1604
rect 19085 1550 19141 1552
rect 20333 1604 20389 1606
rect 20333 1552 20335 1604
rect 20335 1552 20387 1604
rect 20387 1552 20389 1604
rect 20333 1550 20389 1552
rect 21581 1604 21637 1606
rect 21581 1552 21583 1604
rect 21583 1552 21635 1604
rect 21635 1552 21637 1604
rect 21581 1550 21637 1552
rect 22829 1604 22885 1606
rect 22829 1552 22831 1604
rect 22831 1552 22883 1604
rect 22883 1552 22885 1604
rect 22829 1550 22885 1552
rect 24077 1604 24133 1606
rect 24077 1552 24079 1604
rect 24079 1552 24131 1604
rect 24131 1552 24133 1604
rect 24077 1550 24133 1552
rect 25325 1604 25381 1606
rect 25325 1552 25327 1604
rect 25327 1552 25379 1604
rect 25379 1552 25381 1604
rect 25325 1550 25381 1552
rect 26573 1604 26629 1606
rect 26573 1552 26575 1604
rect 26575 1552 26627 1604
rect 26627 1552 26629 1604
rect 26573 1550 26629 1552
rect 27821 1604 27877 1606
rect 27821 1552 27823 1604
rect 27823 1552 27875 1604
rect 27875 1552 27877 1604
rect 27821 1550 27877 1552
rect 29069 1604 29125 1606
rect 29069 1552 29071 1604
rect 29071 1552 29123 1604
rect 29123 1552 29125 1604
rect 29069 1550 29125 1552
rect 30317 1604 30373 1606
rect 30317 1552 30319 1604
rect 30319 1552 30371 1604
rect 30371 1552 30373 1604
rect 30317 1550 30373 1552
rect 31565 1604 31621 1606
rect 31565 1552 31567 1604
rect 31567 1552 31619 1604
rect 31619 1552 31621 1604
rect 31565 1550 31621 1552
rect 32813 1604 32869 1606
rect 32813 1552 32815 1604
rect 32815 1552 32867 1604
rect 32867 1552 32869 1604
rect 32813 1550 32869 1552
rect 34061 1604 34117 1606
rect 34061 1552 34063 1604
rect 34063 1552 34115 1604
rect 34115 1552 34117 1604
rect 34061 1550 34117 1552
rect 35309 1604 35365 1606
rect 35309 1552 35311 1604
rect 35311 1552 35363 1604
rect 35363 1552 35365 1604
rect 35309 1550 35365 1552
rect 36557 1604 36613 1606
rect 36557 1552 36559 1604
rect 36559 1552 36611 1604
rect 36611 1552 36613 1604
rect 36557 1550 36613 1552
rect 37805 1604 37861 1606
rect 37805 1552 37807 1604
rect 37807 1552 37859 1604
rect 37859 1552 37861 1604
rect 37805 1550 37861 1552
rect 39053 1604 39109 1606
rect 39053 1552 39055 1604
rect 39055 1552 39107 1604
rect 39107 1552 39109 1604
rect 39053 1550 39109 1552
rect 40301 1604 40357 1606
rect 40301 1552 40303 1604
rect 40303 1552 40355 1604
rect 40355 1552 40357 1604
rect 40301 1550 40357 1552
rect 1602 1167 1658 1169
rect 1602 1115 1604 1167
rect 1604 1115 1656 1167
rect 1656 1115 1658 1167
rect 1602 1113 1658 1115
rect 2850 1167 2906 1169
rect 2850 1115 2852 1167
rect 2852 1115 2904 1167
rect 2904 1115 2906 1167
rect 2850 1113 2906 1115
rect 4098 1167 4154 1169
rect 4098 1115 4100 1167
rect 4100 1115 4152 1167
rect 4152 1115 4154 1167
rect 4098 1113 4154 1115
rect 5346 1167 5402 1169
rect 5346 1115 5348 1167
rect 5348 1115 5400 1167
rect 5400 1115 5402 1167
rect 5346 1113 5402 1115
rect 6594 1167 6650 1169
rect 6594 1115 6596 1167
rect 6596 1115 6648 1167
rect 6648 1115 6650 1167
rect 6594 1113 6650 1115
rect 7842 1167 7898 1169
rect 7842 1115 7844 1167
rect 7844 1115 7896 1167
rect 7896 1115 7898 1167
rect 7842 1113 7898 1115
rect 9090 1167 9146 1169
rect 9090 1115 9092 1167
rect 9092 1115 9144 1167
rect 9144 1115 9146 1167
rect 9090 1113 9146 1115
rect 10338 1167 10394 1169
rect 10338 1115 10340 1167
rect 10340 1115 10392 1167
rect 10392 1115 10394 1167
rect 10338 1113 10394 1115
rect 11586 1167 11642 1169
rect 11586 1115 11588 1167
rect 11588 1115 11640 1167
rect 11640 1115 11642 1167
rect 11586 1113 11642 1115
rect 12834 1167 12890 1169
rect 12834 1115 12836 1167
rect 12836 1115 12888 1167
rect 12888 1115 12890 1167
rect 12834 1113 12890 1115
rect 14082 1167 14138 1169
rect 14082 1115 14084 1167
rect 14084 1115 14136 1167
rect 14136 1115 14138 1167
rect 14082 1113 14138 1115
rect 15330 1167 15386 1169
rect 15330 1115 15332 1167
rect 15332 1115 15384 1167
rect 15384 1115 15386 1167
rect 15330 1113 15386 1115
rect 16578 1167 16634 1169
rect 16578 1115 16580 1167
rect 16580 1115 16632 1167
rect 16632 1115 16634 1167
rect 16578 1113 16634 1115
rect 17826 1167 17882 1169
rect 17826 1115 17828 1167
rect 17828 1115 17880 1167
rect 17880 1115 17882 1167
rect 17826 1113 17882 1115
rect 19074 1167 19130 1169
rect 19074 1115 19076 1167
rect 19076 1115 19128 1167
rect 19128 1115 19130 1167
rect 19074 1113 19130 1115
rect 20322 1167 20378 1169
rect 20322 1115 20324 1167
rect 20324 1115 20376 1167
rect 20376 1115 20378 1167
rect 20322 1113 20378 1115
rect 21570 1167 21626 1169
rect 21570 1115 21572 1167
rect 21572 1115 21624 1167
rect 21624 1115 21626 1167
rect 21570 1113 21626 1115
rect 22818 1167 22874 1169
rect 22818 1115 22820 1167
rect 22820 1115 22872 1167
rect 22872 1115 22874 1167
rect 22818 1113 22874 1115
rect 24066 1167 24122 1169
rect 24066 1115 24068 1167
rect 24068 1115 24120 1167
rect 24120 1115 24122 1167
rect 24066 1113 24122 1115
rect 25314 1167 25370 1169
rect 25314 1115 25316 1167
rect 25316 1115 25368 1167
rect 25368 1115 25370 1167
rect 25314 1113 25370 1115
rect 26562 1167 26618 1169
rect 26562 1115 26564 1167
rect 26564 1115 26616 1167
rect 26616 1115 26618 1167
rect 26562 1113 26618 1115
rect 27810 1167 27866 1169
rect 27810 1115 27812 1167
rect 27812 1115 27864 1167
rect 27864 1115 27866 1167
rect 27810 1113 27866 1115
rect 29058 1167 29114 1169
rect 29058 1115 29060 1167
rect 29060 1115 29112 1167
rect 29112 1115 29114 1167
rect 29058 1113 29114 1115
rect 30306 1167 30362 1169
rect 30306 1115 30308 1167
rect 30308 1115 30360 1167
rect 30360 1115 30362 1167
rect 30306 1113 30362 1115
rect 31554 1167 31610 1169
rect 31554 1115 31556 1167
rect 31556 1115 31608 1167
rect 31608 1115 31610 1167
rect 31554 1113 31610 1115
rect 32802 1167 32858 1169
rect 32802 1115 32804 1167
rect 32804 1115 32856 1167
rect 32856 1115 32858 1167
rect 32802 1113 32858 1115
rect 34050 1167 34106 1169
rect 34050 1115 34052 1167
rect 34052 1115 34104 1167
rect 34104 1115 34106 1167
rect 34050 1113 34106 1115
rect 35298 1167 35354 1169
rect 35298 1115 35300 1167
rect 35300 1115 35352 1167
rect 35352 1115 35354 1167
rect 35298 1113 35354 1115
rect 36546 1167 36602 1169
rect 36546 1115 36548 1167
rect 36548 1115 36600 1167
rect 36600 1115 36602 1167
rect 36546 1113 36602 1115
rect 37794 1167 37850 1169
rect 37794 1115 37796 1167
rect 37796 1115 37848 1167
rect 37848 1115 37850 1167
rect 37794 1113 37850 1115
rect 39042 1167 39098 1169
rect 39042 1115 39044 1167
rect 39044 1115 39096 1167
rect 39096 1115 39098 1167
rect 39042 1113 39098 1115
rect 40290 1167 40346 1169
rect 40290 1115 40292 1167
rect 40292 1115 40344 1167
rect 40344 1115 40346 1167
rect 40290 1113 40346 1115
rect 1723 836 1779 837
rect 1723 784 1725 836
rect 1725 784 1777 836
rect 1777 784 1779 836
rect 1723 781 1779 784
rect 2971 836 3027 837
rect 2971 784 2973 836
rect 2973 784 3025 836
rect 3025 784 3027 836
rect 2971 781 3027 784
rect 4219 836 4275 837
rect 4219 784 4221 836
rect 4221 784 4273 836
rect 4273 784 4275 836
rect 4219 781 4275 784
rect 5467 836 5523 837
rect 5467 784 5469 836
rect 5469 784 5521 836
rect 5521 784 5523 836
rect 5467 781 5523 784
rect 6715 836 6771 837
rect 6715 784 6717 836
rect 6717 784 6769 836
rect 6769 784 6771 836
rect 6715 781 6771 784
rect 7963 836 8019 837
rect 7963 784 7965 836
rect 7965 784 8017 836
rect 8017 784 8019 836
rect 7963 781 8019 784
rect 9211 836 9267 837
rect 9211 784 9213 836
rect 9213 784 9265 836
rect 9265 784 9267 836
rect 9211 781 9267 784
rect 10459 836 10515 837
rect 10459 784 10461 836
rect 10461 784 10513 836
rect 10513 784 10515 836
rect 10459 781 10515 784
rect 11707 836 11763 837
rect 11707 784 11709 836
rect 11709 784 11761 836
rect 11761 784 11763 836
rect 11707 781 11763 784
rect 12955 836 13011 837
rect 12955 784 12957 836
rect 12957 784 13009 836
rect 13009 784 13011 836
rect 12955 781 13011 784
rect 14203 836 14259 837
rect 14203 784 14205 836
rect 14205 784 14257 836
rect 14257 784 14259 836
rect 14203 781 14259 784
rect 15451 836 15507 837
rect 15451 784 15453 836
rect 15453 784 15505 836
rect 15505 784 15507 836
rect 15451 781 15507 784
rect 16699 836 16755 837
rect 16699 784 16701 836
rect 16701 784 16753 836
rect 16753 784 16755 836
rect 16699 781 16755 784
rect 17947 836 18003 837
rect 17947 784 17949 836
rect 17949 784 18001 836
rect 18001 784 18003 836
rect 17947 781 18003 784
rect 19195 836 19251 837
rect 19195 784 19197 836
rect 19197 784 19249 836
rect 19249 784 19251 836
rect 19195 781 19251 784
rect 20443 836 20499 837
rect 20443 784 20445 836
rect 20445 784 20497 836
rect 20497 784 20499 836
rect 20443 781 20499 784
rect 21691 836 21747 837
rect 21691 784 21693 836
rect 21693 784 21745 836
rect 21745 784 21747 836
rect 21691 781 21747 784
rect 22939 836 22995 837
rect 22939 784 22941 836
rect 22941 784 22993 836
rect 22993 784 22995 836
rect 22939 781 22995 784
rect 24187 836 24243 837
rect 24187 784 24189 836
rect 24189 784 24241 836
rect 24241 784 24243 836
rect 24187 781 24243 784
rect 25435 836 25491 837
rect 25435 784 25437 836
rect 25437 784 25489 836
rect 25489 784 25491 836
rect 25435 781 25491 784
rect 26683 836 26739 837
rect 26683 784 26685 836
rect 26685 784 26737 836
rect 26737 784 26739 836
rect 26683 781 26739 784
rect 27931 836 27987 837
rect 27931 784 27933 836
rect 27933 784 27985 836
rect 27985 784 27987 836
rect 27931 781 27987 784
rect 29179 836 29235 837
rect 29179 784 29181 836
rect 29181 784 29233 836
rect 29233 784 29235 836
rect 29179 781 29235 784
rect 30427 836 30483 837
rect 30427 784 30429 836
rect 30429 784 30481 836
rect 30481 784 30483 836
rect 30427 781 30483 784
rect 31675 836 31731 837
rect 31675 784 31677 836
rect 31677 784 31729 836
rect 31729 784 31731 836
rect 31675 781 31731 784
rect 32923 836 32979 837
rect 32923 784 32925 836
rect 32925 784 32977 836
rect 32977 784 32979 836
rect 32923 781 32979 784
rect 34171 836 34227 837
rect 34171 784 34173 836
rect 34173 784 34225 836
rect 34225 784 34227 836
rect 34171 781 34227 784
rect 35419 836 35475 837
rect 35419 784 35421 836
rect 35421 784 35473 836
rect 35473 784 35475 836
rect 35419 781 35475 784
rect 36667 836 36723 837
rect 36667 784 36669 836
rect 36669 784 36721 836
rect 36721 784 36723 836
rect 36667 781 36723 784
rect 37915 836 37971 837
rect 37915 784 37917 836
rect 37917 784 37969 836
rect 37969 784 37971 836
rect 37915 781 37971 784
rect 39163 836 39219 837
rect 39163 784 39165 836
rect 39165 784 39217 836
rect 39217 784 39219 836
rect 39163 781 39219 784
rect 40411 836 40467 837
rect 40411 784 40413 836
rect 40413 784 40465 836
rect 40465 784 40467 836
rect 40411 781 40467 784
rect 1608 633 1664 635
rect 1608 581 1610 633
rect 1610 581 1662 633
rect 1662 581 1664 633
rect 1608 579 1664 581
rect 2856 633 2912 635
rect 2856 581 2858 633
rect 2858 581 2910 633
rect 2910 581 2912 633
rect 2856 579 2912 581
rect 4104 633 4160 635
rect 4104 581 4106 633
rect 4106 581 4158 633
rect 4158 581 4160 633
rect 4104 579 4160 581
rect 5352 633 5408 635
rect 5352 581 5354 633
rect 5354 581 5406 633
rect 5406 581 5408 633
rect 5352 579 5408 581
rect 6600 633 6656 635
rect 6600 581 6602 633
rect 6602 581 6654 633
rect 6654 581 6656 633
rect 6600 579 6656 581
rect 7848 633 7904 635
rect 7848 581 7850 633
rect 7850 581 7902 633
rect 7902 581 7904 633
rect 7848 579 7904 581
rect 9096 633 9152 635
rect 9096 581 9098 633
rect 9098 581 9150 633
rect 9150 581 9152 633
rect 9096 579 9152 581
rect 10344 633 10400 635
rect 10344 581 10346 633
rect 10346 581 10398 633
rect 10398 581 10400 633
rect 10344 579 10400 581
rect 11592 633 11648 635
rect 11592 581 11594 633
rect 11594 581 11646 633
rect 11646 581 11648 633
rect 11592 579 11648 581
rect 12840 633 12896 635
rect 12840 581 12842 633
rect 12842 581 12894 633
rect 12894 581 12896 633
rect 12840 579 12896 581
rect 14088 633 14144 635
rect 14088 581 14090 633
rect 14090 581 14142 633
rect 14142 581 14144 633
rect 14088 579 14144 581
rect 15336 633 15392 635
rect 15336 581 15338 633
rect 15338 581 15390 633
rect 15390 581 15392 633
rect 15336 579 15392 581
rect 16584 633 16640 635
rect 16584 581 16586 633
rect 16586 581 16638 633
rect 16638 581 16640 633
rect 16584 579 16640 581
rect 17832 633 17888 635
rect 17832 581 17834 633
rect 17834 581 17886 633
rect 17886 581 17888 633
rect 17832 579 17888 581
rect 19080 633 19136 635
rect 19080 581 19082 633
rect 19082 581 19134 633
rect 19134 581 19136 633
rect 19080 579 19136 581
rect 20328 633 20384 635
rect 20328 581 20330 633
rect 20330 581 20382 633
rect 20382 581 20384 633
rect 20328 579 20384 581
rect 21576 633 21632 635
rect 21576 581 21578 633
rect 21578 581 21630 633
rect 21630 581 21632 633
rect 21576 579 21632 581
rect 22824 633 22880 635
rect 22824 581 22826 633
rect 22826 581 22878 633
rect 22878 581 22880 633
rect 22824 579 22880 581
rect 24072 633 24128 635
rect 24072 581 24074 633
rect 24074 581 24126 633
rect 24126 581 24128 633
rect 24072 579 24128 581
rect 25320 633 25376 635
rect 25320 581 25322 633
rect 25322 581 25374 633
rect 25374 581 25376 633
rect 25320 579 25376 581
rect 26568 633 26624 635
rect 26568 581 26570 633
rect 26570 581 26622 633
rect 26622 581 26624 633
rect 26568 579 26624 581
rect 27816 633 27872 635
rect 27816 581 27818 633
rect 27818 581 27870 633
rect 27870 581 27872 633
rect 27816 579 27872 581
rect 29064 633 29120 635
rect 29064 581 29066 633
rect 29066 581 29118 633
rect 29118 581 29120 633
rect 29064 579 29120 581
rect 30312 633 30368 635
rect 30312 581 30314 633
rect 30314 581 30366 633
rect 30366 581 30368 633
rect 30312 579 30368 581
rect 31560 633 31616 635
rect 31560 581 31562 633
rect 31562 581 31614 633
rect 31614 581 31616 633
rect 31560 579 31616 581
rect 32808 633 32864 635
rect 32808 581 32810 633
rect 32810 581 32862 633
rect 32862 581 32864 633
rect 32808 579 32864 581
rect 34056 633 34112 635
rect 34056 581 34058 633
rect 34058 581 34110 633
rect 34110 581 34112 633
rect 34056 579 34112 581
rect 35304 633 35360 635
rect 35304 581 35306 633
rect 35306 581 35358 633
rect 35358 581 35360 633
rect 35304 579 35360 581
rect 36552 633 36608 635
rect 36552 581 36554 633
rect 36554 581 36606 633
rect 36606 581 36608 633
rect 36552 579 36608 581
rect 37800 633 37856 635
rect 37800 581 37802 633
rect 37802 581 37854 633
rect 37854 581 37856 633
rect 37800 579 37856 581
rect 39048 633 39104 635
rect 39048 581 39050 633
rect 39050 581 39102 633
rect 39102 581 39104 633
rect 39048 579 39104 581
rect 40296 633 40352 635
rect 40296 581 40298 633
rect 40298 581 40350 633
rect 40350 581 40352 633
rect 40296 579 40352 581
rect 1622 217 1678 219
rect 1622 165 1624 217
rect 1624 165 1676 217
rect 1676 165 1678 217
rect 1622 163 1678 165
rect 2870 217 2926 219
rect 2870 165 2872 217
rect 2872 165 2924 217
rect 2924 165 2926 217
rect 2870 163 2926 165
rect 4118 217 4174 219
rect 4118 165 4120 217
rect 4120 165 4172 217
rect 4172 165 4174 217
rect 4118 163 4174 165
rect 5366 217 5422 219
rect 5366 165 5368 217
rect 5368 165 5420 217
rect 5420 165 5422 217
rect 5366 163 5422 165
rect 6614 217 6670 219
rect 6614 165 6616 217
rect 6616 165 6668 217
rect 6668 165 6670 217
rect 6614 163 6670 165
rect 7862 217 7918 219
rect 7862 165 7864 217
rect 7864 165 7916 217
rect 7916 165 7918 217
rect 7862 163 7918 165
rect 9110 217 9166 219
rect 9110 165 9112 217
rect 9112 165 9164 217
rect 9164 165 9166 217
rect 9110 163 9166 165
rect 10358 217 10414 219
rect 10358 165 10360 217
rect 10360 165 10412 217
rect 10412 165 10414 217
rect 10358 163 10414 165
rect 11606 217 11662 219
rect 11606 165 11608 217
rect 11608 165 11660 217
rect 11660 165 11662 217
rect 11606 163 11662 165
rect 12854 217 12910 219
rect 12854 165 12856 217
rect 12856 165 12908 217
rect 12908 165 12910 217
rect 12854 163 12910 165
rect 14102 217 14158 219
rect 14102 165 14104 217
rect 14104 165 14156 217
rect 14156 165 14158 217
rect 14102 163 14158 165
rect 15350 217 15406 219
rect 15350 165 15352 217
rect 15352 165 15404 217
rect 15404 165 15406 217
rect 15350 163 15406 165
rect 16598 217 16654 219
rect 16598 165 16600 217
rect 16600 165 16652 217
rect 16652 165 16654 217
rect 16598 163 16654 165
rect 17846 217 17902 219
rect 17846 165 17848 217
rect 17848 165 17900 217
rect 17900 165 17902 217
rect 17846 163 17902 165
rect 19094 217 19150 219
rect 19094 165 19096 217
rect 19096 165 19148 217
rect 19148 165 19150 217
rect 19094 163 19150 165
rect 20342 217 20398 219
rect 20342 165 20344 217
rect 20344 165 20396 217
rect 20396 165 20398 217
rect 20342 163 20398 165
rect 21590 217 21646 219
rect 21590 165 21592 217
rect 21592 165 21644 217
rect 21644 165 21646 217
rect 21590 163 21646 165
rect 22838 217 22894 219
rect 22838 165 22840 217
rect 22840 165 22892 217
rect 22892 165 22894 217
rect 22838 163 22894 165
rect 24086 217 24142 219
rect 24086 165 24088 217
rect 24088 165 24140 217
rect 24140 165 24142 217
rect 24086 163 24142 165
rect 25334 217 25390 219
rect 25334 165 25336 217
rect 25336 165 25388 217
rect 25388 165 25390 217
rect 25334 163 25390 165
rect 26582 217 26638 219
rect 26582 165 26584 217
rect 26584 165 26636 217
rect 26636 165 26638 217
rect 26582 163 26638 165
rect 27830 217 27886 219
rect 27830 165 27832 217
rect 27832 165 27884 217
rect 27884 165 27886 217
rect 27830 163 27886 165
rect 29078 217 29134 219
rect 29078 165 29080 217
rect 29080 165 29132 217
rect 29132 165 29134 217
rect 29078 163 29134 165
rect 30326 217 30382 219
rect 30326 165 30328 217
rect 30328 165 30380 217
rect 30380 165 30382 217
rect 30326 163 30382 165
rect 31574 217 31630 219
rect 31574 165 31576 217
rect 31576 165 31628 217
rect 31628 165 31630 217
rect 31574 163 31630 165
rect 32822 217 32878 219
rect 32822 165 32824 217
rect 32824 165 32876 217
rect 32876 165 32878 217
rect 32822 163 32878 165
rect 34070 217 34126 219
rect 34070 165 34072 217
rect 34072 165 34124 217
rect 34124 165 34126 217
rect 34070 163 34126 165
rect 35318 217 35374 219
rect 35318 165 35320 217
rect 35320 165 35372 217
rect 35372 165 35374 217
rect 35318 163 35374 165
rect 36566 217 36622 219
rect 36566 165 36568 217
rect 36568 165 36620 217
rect 36620 165 36622 217
rect 36566 163 36622 165
rect 37814 217 37870 219
rect 37814 165 37816 217
rect 37816 165 37868 217
rect 37868 165 37870 217
rect 37814 163 37870 165
rect 39062 217 39118 219
rect 39062 165 39064 217
rect 39064 165 39116 217
rect 39116 165 39118 217
rect 39062 163 39118 165
rect 40310 217 40366 219
rect 40310 165 40312 217
rect 40312 165 40364 217
rect 40364 165 40366 217
rect 40310 163 40366 165
<< metal3 >>
rect 1592 1606 1690 1627
rect 1592 1550 1613 1606
rect 1669 1550 1690 1606
rect 1592 1529 1690 1550
rect 2840 1606 2938 1627
rect 2840 1550 2861 1606
rect 2917 1550 2938 1606
rect 2840 1529 2938 1550
rect 4088 1606 4186 1627
rect 4088 1550 4109 1606
rect 4165 1550 4186 1606
rect 4088 1529 4186 1550
rect 5336 1606 5434 1627
rect 5336 1550 5357 1606
rect 5413 1550 5434 1606
rect 5336 1529 5434 1550
rect 6584 1606 6682 1627
rect 6584 1550 6605 1606
rect 6661 1550 6682 1606
rect 6584 1529 6682 1550
rect 7832 1606 7930 1627
rect 7832 1550 7853 1606
rect 7909 1550 7930 1606
rect 7832 1529 7930 1550
rect 9080 1606 9178 1627
rect 9080 1550 9101 1606
rect 9157 1550 9178 1606
rect 9080 1529 9178 1550
rect 10328 1606 10426 1627
rect 10328 1550 10349 1606
rect 10405 1550 10426 1606
rect 10328 1529 10426 1550
rect 11576 1606 11674 1627
rect 11576 1550 11597 1606
rect 11653 1550 11674 1606
rect 11576 1529 11674 1550
rect 12824 1606 12922 1627
rect 12824 1550 12845 1606
rect 12901 1550 12922 1606
rect 12824 1529 12922 1550
rect 14072 1606 14170 1627
rect 14072 1550 14093 1606
rect 14149 1550 14170 1606
rect 14072 1529 14170 1550
rect 15320 1606 15418 1627
rect 15320 1550 15341 1606
rect 15397 1550 15418 1606
rect 15320 1529 15418 1550
rect 16568 1606 16666 1627
rect 16568 1550 16589 1606
rect 16645 1550 16666 1606
rect 16568 1529 16666 1550
rect 17816 1606 17914 1627
rect 17816 1550 17837 1606
rect 17893 1550 17914 1606
rect 17816 1529 17914 1550
rect 19064 1606 19162 1627
rect 19064 1550 19085 1606
rect 19141 1550 19162 1606
rect 19064 1529 19162 1550
rect 20312 1606 20410 1627
rect 20312 1550 20333 1606
rect 20389 1550 20410 1606
rect 20312 1529 20410 1550
rect 21560 1606 21658 1627
rect 21560 1550 21581 1606
rect 21637 1550 21658 1606
rect 21560 1529 21658 1550
rect 22808 1606 22906 1627
rect 22808 1550 22829 1606
rect 22885 1550 22906 1606
rect 22808 1529 22906 1550
rect 24056 1606 24154 1627
rect 24056 1550 24077 1606
rect 24133 1550 24154 1606
rect 24056 1529 24154 1550
rect 25304 1606 25402 1627
rect 25304 1550 25325 1606
rect 25381 1550 25402 1606
rect 25304 1529 25402 1550
rect 26552 1606 26650 1627
rect 26552 1550 26573 1606
rect 26629 1550 26650 1606
rect 26552 1529 26650 1550
rect 27800 1606 27898 1627
rect 27800 1550 27821 1606
rect 27877 1550 27898 1606
rect 27800 1529 27898 1550
rect 29048 1606 29146 1627
rect 29048 1550 29069 1606
rect 29125 1550 29146 1606
rect 29048 1529 29146 1550
rect 30296 1606 30394 1627
rect 30296 1550 30317 1606
rect 30373 1550 30394 1606
rect 30296 1529 30394 1550
rect 31544 1606 31642 1627
rect 31544 1550 31565 1606
rect 31621 1550 31642 1606
rect 31544 1529 31642 1550
rect 32792 1606 32890 1627
rect 32792 1550 32813 1606
rect 32869 1550 32890 1606
rect 32792 1529 32890 1550
rect 34040 1606 34138 1627
rect 34040 1550 34061 1606
rect 34117 1550 34138 1606
rect 34040 1529 34138 1550
rect 35288 1606 35386 1627
rect 35288 1550 35309 1606
rect 35365 1550 35386 1606
rect 35288 1529 35386 1550
rect 36536 1606 36634 1627
rect 36536 1550 36557 1606
rect 36613 1550 36634 1606
rect 36536 1529 36634 1550
rect 37784 1606 37882 1627
rect 37784 1550 37805 1606
rect 37861 1550 37882 1606
rect 37784 1529 37882 1550
rect 39032 1606 39130 1627
rect 39032 1550 39053 1606
rect 39109 1550 39130 1606
rect 39032 1529 39130 1550
rect 40280 1606 40378 1627
rect 40280 1550 40301 1606
rect 40357 1550 40378 1606
rect 40280 1529 40378 1550
rect 1581 1169 1679 1190
rect 1581 1113 1602 1169
rect 1658 1113 1679 1169
rect 1581 1092 1679 1113
rect 2829 1169 2927 1190
rect 2829 1113 2850 1169
rect 2906 1113 2927 1169
rect 2829 1092 2927 1113
rect 4077 1169 4175 1190
rect 4077 1113 4098 1169
rect 4154 1113 4175 1169
rect 4077 1092 4175 1113
rect 5325 1169 5423 1190
rect 5325 1113 5346 1169
rect 5402 1113 5423 1169
rect 5325 1092 5423 1113
rect 6573 1169 6671 1190
rect 6573 1113 6594 1169
rect 6650 1113 6671 1169
rect 6573 1092 6671 1113
rect 7821 1169 7919 1190
rect 7821 1113 7842 1169
rect 7898 1113 7919 1169
rect 7821 1092 7919 1113
rect 9069 1169 9167 1190
rect 9069 1113 9090 1169
rect 9146 1113 9167 1169
rect 9069 1092 9167 1113
rect 10317 1169 10415 1190
rect 10317 1113 10338 1169
rect 10394 1113 10415 1169
rect 10317 1092 10415 1113
rect 11565 1169 11663 1190
rect 11565 1113 11586 1169
rect 11642 1113 11663 1169
rect 11565 1092 11663 1113
rect 12813 1169 12911 1190
rect 12813 1113 12834 1169
rect 12890 1113 12911 1169
rect 12813 1092 12911 1113
rect 14061 1169 14159 1190
rect 14061 1113 14082 1169
rect 14138 1113 14159 1169
rect 14061 1092 14159 1113
rect 15309 1169 15407 1190
rect 15309 1113 15330 1169
rect 15386 1113 15407 1169
rect 15309 1092 15407 1113
rect 16557 1169 16655 1190
rect 16557 1113 16578 1169
rect 16634 1113 16655 1169
rect 16557 1092 16655 1113
rect 17805 1169 17903 1190
rect 17805 1113 17826 1169
rect 17882 1113 17903 1169
rect 17805 1092 17903 1113
rect 19053 1169 19151 1190
rect 19053 1113 19074 1169
rect 19130 1113 19151 1169
rect 19053 1092 19151 1113
rect 20301 1169 20399 1190
rect 20301 1113 20322 1169
rect 20378 1113 20399 1169
rect 20301 1092 20399 1113
rect 21549 1169 21647 1190
rect 21549 1113 21570 1169
rect 21626 1113 21647 1169
rect 21549 1092 21647 1113
rect 22797 1169 22895 1190
rect 22797 1113 22818 1169
rect 22874 1113 22895 1169
rect 22797 1092 22895 1113
rect 24045 1169 24143 1190
rect 24045 1113 24066 1169
rect 24122 1113 24143 1169
rect 24045 1092 24143 1113
rect 25293 1169 25391 1190
rect 25293 1113 25314 1169
rect 25370 1113 25391 1169
rect 25293 1092 25391 1113
rect 26541 1169 26639 1190
rect 26541 1113 26562 1169
rect 26618 1113 26639 1169
rect 26541 1092 26639 1113
rect 27789 1169 27887 1190
rect 27789 1113 27810 1169
rect 27866 1113 27887 1169
rect 27789 1092 27887 1113
rect 29037 1169 29135 1190
rect 29037 1113 29058 1169
rect 29114 1113 29135 1169
rect 29037 1092 29135 1113
rect 30285 1169 30383 1190
rect 30285 1113 30306 1169
rect 30362 1113 30383 1169
rect 30285 1092 30383 1113
rect 31533 1169 31631 1190
rect 31533 1113 31554 1169
rect 31610 1113 31631 1169
rect 31533 1092 31631 1113
rect 32781 1169 32879 1190
rect 32781 1113 32802 1169
rect 32858 1113 32879 1169
rect 32781 1092 32879 1113
rect 34029 1169 34127 1190
rect 34029 1113 34050 1169
rect 34106 1113 34127 1169
rect 34029 1092 34127 1113
rect 35277 1169 35375 1190
rect 35277 1113 35298 1169
rect 35354 1113 35375 1169
rect 35277 1092 35375 1113
rect 36525 1169 36623 1190
rect 36525 1113 36546 1169
rect 36602 1113 36623 1169
rect 36525 1092 36623 1113
rect 37773 1169 37871 1190
rect 37773 1113 37794 1169
rect 37850 1113 37871 1169
rect 37773 1092 37871 1113
rect 39021 1169 39119 1190
rect 39021 1113 39042 1169
rect 39098 1113 39119 1169
rect 39021 1092 39119 1113
rect 40269 1169 40367 1190
rect 40269 1113 40290 1169
rect 40346 1113 40367 1169
rect 40269 1092 40367 1113
rect 1702 837 1800 858
rect 1702 781 1723 837
rect 1779 781 1800 837
rect 1702 760 1800 781
rect 2950 837 3048 858
rect 2950 781 2971 837
rect 3027 781 3048 837
rect 2950 760 3048 781
rect 4198 837 4296 858
rect 4198 781 4219 837
rect 4275 781 4296 837
rect 4198 760 4296 781
rect 5446 837 5544 858
rect 5446 781 5467 837
rect 5523 781 5544 837
rect 5446 760 5544 781
rect 6694 837 6792 858
rect 6694 781 6715 837
rect 6771 781 6792 837
rect 6694 760 6792 781
rect 7942 837 8040 858
rect 7942 781 7963 837
rect 8019 781 8040 837
rect 7942 760 8040 781
rect 9190 837 9288 858
rect 9190 781 9211 837
rect 9267 781 9288 837
rect 9190 760 9288 781
rect 10438 837 10536 858
rect 10438 781 10459 837
rect 10515 781 10536 837
rect 10438 760 10536 781
rect 11686 837 11784 858
rect 11686 781 11707 837
rect 11763 781 11784 837
rect 11686 760 11784 781
rect 12934 837 13032 858
rect 12934 781 12955 837
rect 13011 781 13032 837
rect 12934 760 13032 781
rect 14182 837 14280 858
rect 14182 781 14203 837
rect 14259 781 14280 837
rect 14182 760 14280 781
rect 15430 837 15528 858
rect 15430 781 15451 837
rect 15507 781 15528 837
rect 15430 760 15528 781
rect 16678 837 16776 858
rect 16678 781 16699 837
rect 16755 781 16776 837
rect 16678 760 16776 781
rect 17926 837 18024 858
rect 17926 781 17947 837
rect 18003 781 18024 837
rect 17926 760 18024 781
rect 19174 837 19272 858
rect 19174 781 19195 837
rect 19251 781 19272 837
rect 19174 760 19272 781
rect 20422 837 20520 858
rect 20422 781 20443 837
rect 20499 781 20520 837
rect 20422 760 20520 781
rect 21670 837 21768 858
rect 21670 781 21691 837
rect 21747 781 21768 837
rect 21670 760 21768 781
rect 22918 837 23016 858
rect 22918 781 22939 837
rect 22995 781 23016 837
rect 22918 760 23016 781
rect 24166 837 24264 858
rect 24166 781 24187 837
rect 24243 781 24264 837
rect 24166 760 24264 781
rect 25414 837 25512 858
rect 25414 781 25435 837
rect 25491 781 25512 837
rect 25414 760 25512 781
rect 26662 837 26760 858
rect 26662 781 26683 837
rect 26739 781 26760 837
rect 26662 760 26760 781
rect 27910 837 28008 858
rect 27910 781 27931 837
rect 27987 781 28008 837
rect 27910 760 28008 781
rect 29158 837 29256 858
rect 29158 781 29179 837
rect 29235 781 29256 837
rect 29158 760 29256 781
rect 30406 837 30504 858
rect 30406 781 30427 837
rect 30483 781 30504 837
rect 30406 760 30504 781
rect 31654 837 31752 858
rect 31654 781 31675 837
rect 31731 781 31752 837
rect 31654 760 31752 781
rect 32902 837 33000 858
rect 32902 781 32923 837
rect 32979 781 33000 837
rect 32902 760 33000 781
rect 34150 837 34248 858
rect 34150 781 34171 837
rect 34227 781 34248 837
rect 34150 760 34248 781
rect 35398 837 35496 858
rect 35398 781 35419 837
rect 35475 781 35496 837
rect 35398 760 35496 781
rect 36646 837 36744 858
rect 36646 781 36667 837
rect 36723 781 36744 837
rect 36646 760 36744 781
rect 37894 837 37992 858
rect 37894 781 37915 837
rect 37971 781 37992 837
rect 37894 760 37992 781
rect 39142 837 39240 858
rect 39142 781 39163 837
rect 39219 781 39240 837
rect 39142 760 39240 781
rect 40390 837 40488 858
rect 40390 781 40411 837
rect 40467 781 40488 837
rect 40390 760 40488 781
rect 1587 635 1685 656
rect 1587 579 1608 635
rect 1664 579 1685 635
rect 1587 558 1685 579
rect 2835 635 2933 656
rect 2835 579 2856 635
rect 2912 579 2933 635
rect 2835 558 2933 579
rect 4083 635 4181 656
rect 4083 579 4104 635
rect 4160 579 4181 635
rect 4083 558 4181 579
rect 5331 635 5429 656
rect 5331 579 5352 635
rect 5408 579 5429 635
rect 5331 558 5429 579
rect 6579 635 6677 656
rect 6579 579 6600 635
rect 6656 579 6677 635
rect 6579 558 6677 579
rect 7827 635 7925 656
rect 7827 579 7848 635
rect 7904 579 7925 635
rect 7827 558 7925 579
rect 9075 635 9173 656
rect 9075 579 9096 635
rect 9152 579 9173 635
rect 9075 558 9173 579
rect 10323 635 10421 656
rect 10323 579 10344 635
rect 10400 579 10421 635
rect 10323 558 10421 579
rect 11571 635 11669 656
rect 11571 579 11592 635
rect 11648 579 11669 635
rect 11571 558 11669 579
rect 12819 635 12917 656
rect 12819 579 12840 635
rect 12896 579 12917 635
rect 12819 558 12917 579
rect 14067 635 14165 656
rect 14067 579 14088 635
rect 14144 579 14165 635
rect 14067 558 14165 579
rect 15315 635 15413 656
rect 15315 579 15336 635
rect 15392 579 15413 635
rect 15315 558 15413 579
rect 16563 635 16661 656
rect 16563 579 16584 635
rect 16640 579 16661 635
rect 16563 558 16661 579
rect 17811 635 17909 656
rect 17811 579 17832 635
rect 17888 579 17909 635
rect 17811 558 17909 579
rect 19059 635 19157 656
rect 19059 579 19080 635
rect 19136 579 19157 635
rect 19059 558 19157 579
rect 20307 635 20405 656
rect 20307 579 20328 635
rect 20384 579 20405 635
rect 20307 558 20405 579
rect 21555 635 21653 656
rect 21555 579 21576 635
rect 21632 579 21653 635
rect 21555 558 21653 579
rect 22803 635 22901 656
rect 22803 579 22824 635
rect 22880 579 22901 635
rect 22803 558 22901 579
rect 24051 635 24149 656
rect 24051 579 24072 635
rect 24128 579 24149 635
rect 24051 558 24149 579
rect 25299 635 25397 656
rect 25299 579 25320 635
rect 25376 579 25397 635
rect 25299 558 25397 579
rect 26547 635 26645 656
rect 26547 579 26568 635
rect 26624 579 26645 635
rect 26547 558 26645 579
rect 27795 635 27893 656
rect 27795 579 27816 635
rect 27872 579 27893 635
rect 27795 558 27893 579
rect 29043 635 29141 656
rect 29043 579 29064 635
rect 29120 579 29141 635
rect 29043 558 29141 579
rect 30291 635 30389 656
rect 30291 579 30312 635
rect 30368 579 30389 635
rect 30291 558 30389 579
rect 31539 635 31637 656
rect 31539 579 31560 635
rect 31616 579 31637 635
rect 31539 558 31637 579
rect 32787 635 32885 656
rect 32787 579 32808 635
rect 32864 579 32885 635
rect 32787 558 32885 579
rect 34035 635 34133 656
rect 34035 579 34056 635
rect 34112 579 34133 635
rect 34035 558 34133 579
rect 35283 635 35381 656
rect 35283 579 35304 635
rect 35360 579 35381 635
rect 35283 558 35381 579
rect 36531 635 36629 656
rect 36531 579 36552 635
rect 36608 579 36629 635
rect 36531 558 36629 579
rect 37779 635 37877 656
rect 37779 579 37800 635
rect 37856 579 37877 635
rect 37779 558 37877 579
rect 39027 635 39125 656
rect 39027 579 39048 635
rect 39104 579 39125 635
rect 39027 558 39125 579
rect 40275 635 40373 656
rect 40275 579 40296 635
rect 40352 579 40373 635
rect 40275 558 40373 579
rect 1601 219 1699 240
rect 1601 163 1622 219
rect 1678 163 1699 219
rect 1601 142 1699 163
rect 2849 219 2947 240
rect 2849 163 2870 219
rect 2926 163 2947 219
rect 2849 142 2947 163
rect 4097 219 4195 240
rect 4097 163 4118 219
rect 4174 163 4195 219
rect 4097 142 4195 163
rect 5345 219 5443 240
rect 5345 163 5366 219
rect 5422 163 5443 219
rect 5345 142 5443 163
rect 6593 219 6691 240
rect 6593 163 6614 219
rect 6670 163 6691 219
rect 6593 142 6691 163
rect 7841 219 7939 240
rect 7841 163 7862 219
rect 7918 163 7939 219
rect 7841 142 7939 163
rect 9089 219 9187 240
rect 9089 163 9110 219
rect 9166 163 9187 219
rect 9089 142 9187 163
rect 10337 219 10435 240
rect 10337 163 10358 219
rect 10414 163 10435 219
rect 10337 142 10435 163
rect 11585 219 11683 240
rect 11585 163 11606 219
rect 11662 163 11683 219
rect 11585 142 11683 163
rect 12833 219 12931 240
rect 12833 163 12854 219
rect 12910 163 12931 219
rect 12833 142 12931 163
rect 14081 219 14179 240
rect 14081 163 14102 219
rect 14158 163 14179 219
rect 14081 142 14179 163
rect 15329 219 15427 240
rect 15329 163 15350 219
rect 15406 163 15427 219
rect 15329 142 15427 163
rect 16577 219 16675 240
rect 16577 163 16598 219
rect 16654 163 16675 219
rect 16577 142 16675 163
rect 17825 219 17923 240
rect 17825 163 17846 219
rect 17902 163 17923 219
rect 17825 142 17923 163
rect 19073 219 19171 240
rect 19073 163 19094 219
rect 19150 163 19171 219
rect 19073 142 19171 163
rect 20321 219 20419 240
rect 20321 163 20342 219
rect 20398 163 20419 219
rect 20321 142 20419 163
rect 21569 219 21667 240
rect 21569 163 21590 219
rect 21646 163 21667 219
rect 21569 142 21667 163
rect 22817 219 22915 240
rect 22817 163 22838 219
rect 22894 163 22915 219
rect 22817 142 22915 163
rect 24065 219 24163 240
rect 24065 163 24086 219
rect 24142 163 24163 219
rect 24065 142 24163 163
rect 25313 219 25411 240
rect 25313 163 25334 219
rect 25390 163 25411 219
rect 25313 142 25411 163
rect 26561 219 26659 240
rect 26561 163 26582 219
rect 26638 163 26659 219
rect 26561 142 26659 163
rect 27809 219 27907 240
rect 27809 163 27830 219
rect 27886 163 27907 219
rect 27809 142 27907 163
rect 29057 219 29155 240
rect 29057 163 29078 219
rect 29134 163 29155 219
rect 29057 142 29155 163
rect 30305 219 30403 240
rect 30305 163 30326 219
rect 30382 163 30403 219
rect 30305 142 30403 163
rect 31553 219 31651 240
rect 31553 163 31574 219
rect 31630 163 31651 219
rect 31553 142 31651 163
rect 32801 219 32899 240
rect 32801 163 32822 219
rect 32878 163 32899 219
rect 32801 142 32899 163
rect 34049 219 34147 240
rect 34049 163 34070 219
rect 34126 163 34147 219
rect 34049 142 34147 163
rect 35297 219 35395 240
rect 35297 163 35318 219
rect 35374 163 35395 219
rect 35297 142 35395 163
rect 36545 219 36643 240
rect 36545 163 36566 219
rect 36622 163 36643 219
rect 36545 142 36643 163
rect 37793 219 37891 240
rect 37793 163 37814 219
rect 37870 163 37891 219
rect 37793 142 37891 163
rect 39041 219 39139 240
rect 39041 163 39062 219
rect 39118 163 39139 219
rect 39041 142 39139 163
rect 40289 219 40387 240
rect 40289 163 40310 219
rect 40366 163 40387 219
rect 40289 142 40387 163
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1694700623
transform 1 0 2622 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1694700623
transform 1 0 1374 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1694700623
transform 1 0 6366 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1694700623
transform 1 0 5118 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1694700623
transform 1 0 3870 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1694700623
transform 1 0 8862 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1694700623
transform 1 0 7614 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1694700623
transform 1 0 18846 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_8
timestamp 1694700623
transform 1 0 17598 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_9
timestamp 1694700623
transform 1 0 16350 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_10
timestamp 1694700623
transform 1 0 15102 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_11
timestamp 1694700623
transform 1 0 13854 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_12
timestamp 1694700623
transform 1 0 12606 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_13
timestamp 1694700623
transform 1 0 11358 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_14
timestamp 1694700623
transform 1 0 10110 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_15
timestamp 1694700623
transform 1 0 25086 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_16
timestamp 1694700623
transform 1 0 23838 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_17
timestamp 1694700623
transform 1 0 22590 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_18
timestamp 1694700623
transform 1 0 28830 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_19
timestamp 1694700623
transform 1 0 27582 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_20
timestamp 1694700623
transform 1 0 26334 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_21
timestamp 1694700623
transform 1 0 40062 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_22
timestamp 1694700623
transform 1 0 38814 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_23
timestamp 1694700623
transform 1 0 37566 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_24
timestamp 1694700623
transform 1 0 36318 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_25
timestamp 1694700623
transform 1 0 35070 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_26
timestamp 1694700623
transform 1 0 33822 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_27
timestamp 1694700623
transform 1 0 32574 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_28
timestamp 1694700623
transform 1 0 31326 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_29
timestamp 1694700623
transform 1 0 30078 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_30
timestamp 1694700623
transform 1 0 21342 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver  sky130_fd_bd_sram__openram_write_driver_31
timestamp 1694700623
transform 1 0 20094 0 1 0
box -376 4 880 2011
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_0
timestamp 1694700623
transform 1 0 7965 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_1
timestamp 1694700623
transform 1 0 7850 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_2
timestamp 1694700623
transform 1 0 7844 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_3
timestamp 1694700623
transform 1 0 7864 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_4
timestamp 1694700623
transform 1 0 6607 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_5
timestamp 1694700623
transform 1 0 6717 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_6
timestamp 1694700623
transform 1 0 6602 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_7
timestamp 1694700623
transform 1 0 6596 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_8
timestamp 1694700623
transform 1 0 6616 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_9
timestamp 1694700623
transform 1 0 5359 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_10
timestamp 1694700623
transform 1 0 5469 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_11
timestamp 1694700623
transform 1 0 5354 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_12
timestamp 1694700623
transform 1 0 5348 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_13
timestamp 1694700623
transform 1 0 5368 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_14
timestamp 1694700623
transform 1 0 4111 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_15
timestamp 1694700623
transform 1 0 4221 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_16
timestamp 1694700623
transform 1 0 4106 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_17
timestamp 1694700623
transform 1 0 4100 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_18
timestamp 1694700623
transform 1 0 4120 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_19
timestamp 1694700623
transform 1 0 2863 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_20
timestamp 1694700623
transform 1 0 2973 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_21
timestamp 1694700623
transform 1 0 2858 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_22
timestamp 1694700623
transform 1 0 2852 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_23
timestamp 1694700623
transform 1 0 2872 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_24
timestamp 1694700623
transform 1 0 1615 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_25
timestamp 1694700623
transform 1 0 1725 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_26
timestamp 1694700623
transform 1 0 1610 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_27
timestamp 1694700623
transform 1 0 1604 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_28
timestamp 1694700623
transform 1 0 1624 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_29
timestamp 1694700623
transform 1 0 10351 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_30
timestamp 1694700623
transform 1 0 10461 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_31
timestamp 1694700623
transform 1 0 10346 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_32
timestamp 1694700623
transform 1 0 10340 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_33
timestamp 1694700623
transform 1 0 10360 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_34
timestamp 1694700623
transform 1 0 9103 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_35
timestamp 1694700623
transform 1 0 9213 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_36
timestamp 1694700623
transform 1 0 9098 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_37
timestamp 1694700623
transform 1 0 9092 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_38
timestamp 1694700623
transform 1 0 9112 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_39
timestamp 1694700623
transform 1 0 7855 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_40
timestamp 1694700623
transform 1 0 19082 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_41
timestamp 1694700623
transform 1 0 19076 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_42
timestamp 1694700623
transform 1 0 19096 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_43
timestamp 1694700623
transform 1 0 17839 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_44
timestamp 1694700623
transform 1 0 17949 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_45
timestamp 1694700623
transform 1 0 17834 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_46
timestamp 1694700623
transform 1 0 17828 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_47
timestamp 1694700623
transform 1 0 17848 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_48
timestamp 1694700623
transform 1 0 16591 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_49
timestamp 1694700623
transform 1 0 16701 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_50
timestamp 1694700623
transform 1 0 16586 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_51
timestamp 1694700623
transform 1 0 16580 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_52
timestamp 1694700623
transform 1 0 16600 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_53
timestamp 1694700623
transform 1 0 15343 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_54
timestamp 1694700623
transform 1 0 15453 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_55
timestamp 1694700623
transform 1 0 15338 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_56
timestamp 1694700623
transform 1 0 15332 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_57
timestamp 1694700623
transform 1 0 15352 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_58
timestamp 1694700623
transform 1 0 14095 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_59
timestamp 1694700623
transform 1 0 14205 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_60
timestamp 1694700623
transform 1 0 14090 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_61
timestamp 1694700623
transform 1 0 14084 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_62
timestamp 1694700623
transform 1 0 14104 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_63
timestamp 1694700623
transform 1 0 12847 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_64
timestamp 1694700623
transform 1 0 12957 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_65
timestamp 1694700623
transform 1 0 12842 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_66
timestamp 1694700623
transform 1 0 12836 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_67
timestamp 1694700623
transform 1 0 12856 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_68
timestamp 1694700623
transform 1 0 11599 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_69
timestamp 1694700623
transform 1 0 11709 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_70
timestamp 1694700623
transform 1 0 11594 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_71
timestamp 1694700623
transform 1 0 11588 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_72
timestamp 1694700623
transform 1 0 11608 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_73
timestamp 1694700623
transform 1 0 19197 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_74
timestamp 1694700623
transform 1 0 20335 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_75
timestamp 1694700623
transform 1 0 20445 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_76
timestamp 1694700623
transform 1 0 20330 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_77
timestamp 1694700623
transform 1 0 20324 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_78
timestamp 1694700623
transform 1 0 20344 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_79
timestamp 1694700623
transform 1 0 19087 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_80
timestamp 1694700623
transform 1 0 30308 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_81
timestamp 1694700623
transform 1 0 30328 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_82
timestamp 1694700623
transform 1 0 29071 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_83
timestamp 1694700623
transform 1 0 29181 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_84
timestamp 1694700623
transform 1 0 29066 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_85
timestamp 1694700623
transform 1 0 29060 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_86
timestamp 1694700623
transform 1 0 29080 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_87
timestamp 1694700623
transform 1 0 27823 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_88
timestamp 1694700623
transform 1 0 27933 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_89
timestamp 1694700623
transform 1 0 27818 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_90
timestamp 1694700623
transform 1 0 27812 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_91
timestamp 1694700623
transform 1 0 27832 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_92
timestamp 1694700623
transform 1 0 26575 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_93
timestamp 1694700623
transform 1 0 26685 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_94
timestamp 1694700623
transform 1 0 26570 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_95
timestamp 1694700623
transform 1 0 26564 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_96
timestamp 1694700623
transform 1 0 26584 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_97
timestamp 1694700623
transform 1 0 25327 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_98
timestamp 1694700623
transform 1 0 25437 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_99
timestamp 1694700623
transform 1 0 25322 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_100
timestamp 1694700623
transform 1 0 25316 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_101
timestamp 1694700623
transform 1 0 25336 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_102
timestamp 1694700623
transform 1 0 24079 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_103
timestamp 1694700623
transform 1 0 24189 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_104
timestamp 1694700623
transform 1 0 24074 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_105
timestamp 1694700623
transform 1 0 24068 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_106
timestamp 1694700623
transform 1 0 24088 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_107
timestamp 1694700623
transform 1 0 22831 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_108
timestamp 1694700623
transform 1 0 22941 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_109
timestamp 1694700623
transform 1 0 22826 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_110
timestamp 1694700623
transform 1 0 22820 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_111
timestamp 1694700623
transform 1 0 22840 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_112
timestamp 1694700623
transform 1 0 21583 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_113
timestamp 1694700623
transform 1 0 21693 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_114
timestamp 1694700623
transform 1 0 21578 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_115
timestamp 1694700623
transform 1 0 21572 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_116
timestamp 1694700623
transform 1 0 21592 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_117
timestamp 1694700623
transform 1 0 30319 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_118
timestamp 1694700623
transform 1 0 30429 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_119
timestamp 1694700623
transform 1 0 30314 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_120
timestamp 1694700623
transform 1 0 40303 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_121
timestamp 1694700623
transform 1 0 40413 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_122
timestamp 1694700623
transform 1 0 40298 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_123
timestamp 1694700623
transform 1 0 40292 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_124
timestamp 1694700623
transform 1 0 40312 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_125
timestamp 1694700623
transform 1 0 39055 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_126
timestamp 1694700623
transform 1 0 39165 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_127
timestamp 1694700623
transform 1 0 39050 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_128
timestamp 1694700623
transform 1 0 39044 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_129
timestamp 1694700623
transform 1 0 39064 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_130
timestamp 1694700623
transform 1 0 37807 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_131
timestamp 1694700623
transform 1 0 37917 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_132
timestamp 1694700623
transform 1 0 37802 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_133
timestamp 1694700623
transform 1 0 37796 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_134
timestamp 1694700623
transform 1 0 37816 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_135
timestamp 1694700623
transform 1 0 36559 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_136
timestamp 1694700623
transform 1 0 36669 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_137
timestamp 1694700623
transform 1 0 36554 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_138
timestamp 1694700623
transform 1 0 36548 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_139
timestamp 1694700623
transform 1 0 36568 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_140
timestamp 1694700623
transform 1 0 35311 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_141
timestamp 1694700623
transform 1 0 35421 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_142
timestamp 1694700623
transform 1 0 35306 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_143
timestamp 1694700623
transform 1 0 35300 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_144
timestamp 1694700623
transform 1 0 35320 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_145
timestamp 1694700623
transform 1 0 34063 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_146
timestamp 1694700623
transform 1 0 34173 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_147
timestamp 1694700623
transform 1 0 34058 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_148
timestamp 1694700623
transform 1 0 34052 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_149
timestamp 1694700623
transform 1 0 34072 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_150
timestamp 1694700623
transform 1 0 32815 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_151
timestamp 1694700623
transform 1 0 32925 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_152
timestamp 1694700623
transform 1 0 32810 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_153
timestamp 1694700623
transform 1 0 32804 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_154
timestamp 1694700623
transform 1 0 32824 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_155
timestamp 1694700623
transform 1 0 31567 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_156
timestamp 1694700623
transform 1 0 31677 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_157
timestamp 1694700623
transform 1 0 31562 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_158
timestamp 1694700623
transform 1 0 31556 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_21  sky130_sram_1kbyte_1rw1r_32x256_8_contact_21_159
timestamp 1694700623
transform 1 0 31576 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_0
timestamp 1694700623
transform 1 0 7958 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_1
timestamp 1694700623
transform 1 0 7843 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_2
timestamp 1694700623
transform 1 0 7837 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_3
timestamp 1694700623
transform 1 0 7857 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_4
timestamp 1694700623
transform 1 0 6600 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_5
timestamp 1694700623
transform 1 0 6710 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_6
timestamp 1694700623
transform 1 0 6595 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_7
timestamp 1694700623
transform 1 0 6589 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_8
timestamp 1694700623
transform 1 0 6609 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_9
timestamp 1694700623
transform 1 0 5352 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_10
timestamp 1694700623
transform 1 0 5462 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_11
timestamp 1694700623
transform 1 0 5347 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_12
timestamp 1694700623
transform 1 0 5341 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_13
timestamp 1694700623
transform 1 0 5361 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_14
timestamp 1694700623
transform 1 0 4104 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_15
timestamp 1694700623
transform 1 0 4214 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_16
timestamp 1694700623
transform 1 0 4099 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_17
timestamp 1694700623
transform 1 0 4093 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_18
timestamp 1694700623
transform 1 0 4113 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_19
timestamp 1694700623
transform 1 0 2856 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_20
timestamp 1694700623
transform 1 0 2966 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_21
timestamp 1694700623
transform 1 0 2851 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_22
timestamp 1694700623
transform 1 0 2845 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_23
timestamp 1694700623
transform 1 0 2865 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_24
timestamp 1694700623
transform 1 0 1608 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_25
timestamp 1694700623
transform 1 0 1718 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_26
timestamp 1694700623
transform 1 0 1603 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_27
timestamp 1694700623
transform 1 0 1597 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_28
timestamp 1694700623
transform 1 0 1617 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_29
timestamp 1694700623
transform 1 0 10344 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_30
timestamp 1694700623
transform 1 0 10454 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_31
timestamp 1694700623
transform 1 0 10339 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_32
timestamp 1694700623
transform 1 0 10333 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_33
timestamp 1694700623
transform 1 0 10353 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_34
timestamp 1694700623
transform 1 0 9096 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_35
timestamp 1694700623
transform 1 0 9206 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_36
timestamp 1694700623
transform 1 0 9091 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_37
timestamp 1694700623
transform 1 0 9085 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_38
timestamp 1694700623
transform 1 0 9105 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_39
timestamp 1694700623
transform 1 0 7848 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_40
timestamp 1694700623
transform 1 0 19069 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_41
timestamp 1694700623
transform 1 0 19089 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_42
timestamp 1694700623
transform 1 0 17832 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_43
timestamp 1694700623
transform 1 0 17942 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_44
timestamp 1694700623
transform 1 0 17827 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_45
timestamp 1694700623
transform 1 0 17821 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_46
timestamp 1694700623
transform 1 0 17841 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_47
timestamp 1694700623
transform 1 0 16584 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_48
timestamp 1694700623
transform 1 0 16694 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_49
timestamp 1694700623
transform 1 0 16579 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_50
timestamp 1694700623
transform 1 0 16573 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_51
timestamp 1694700623
transform 1 0 16593 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_52
timestamp 1694700623
transform 1 0 15336 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_53
timestamp 1694700623
transform 1 0 15446 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_54
timestamp 1694700623
transform 1 0 15331 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_55
timestamp 1694700623
transform 1 0 15325 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_56
timestamp 1694700623
transform 1 0 15345 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_57
timestamp 1694700623
transform 1 0 14088 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_58
timestamp 1694700623
transform 1 0 14198 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_59
timestamp 1694700623
transform 1 0 14083 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_60
timestamp 1694700623
transform 1 0 14077 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_61
timestamp 1694700623
transform 1 0 14097 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_62
timestamp 1694700623
transform 1 0 12840 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_63
timestamp 1694700623
transform 1 0 12950 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_64
timestamp 1694700623
transform 1 0 12835 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_65
timestamp 1694700623
transform 1 0 12829 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_66
timestamp 1694700623
transform 1 0 12849 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_67
timestamp 1694700623
transform 1 0 11592 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_68
timestamp 1694700623
transform 1 0 11702 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_69
timestamp 1694700623
transform 1 0 11587 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_70
timestamp 1694700623
transform 1 0 11581 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_71
timestamp 1694700623
transform 1 0 11601 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_72
timestamp 1694700623
transform 1 0 19075 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_73
timestamp 1694700623
transform 1 0 20328 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_74
timestamp 1694700623
transform 1 0 20438 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_75
timestamp 1694700623
transform 1 0 20323 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_76
timestamp 1694700623
transform 1 0 20317 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_77
timestamp 1694700623
transform 1 0 20337 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_78
timestamp 1694700623
transform 1 0 19080 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_79
timestamp 1694700623
transform 1 0 19190 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_80
timestamp 1694700623
transform 1 0 30301 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_81
timestamp 1694700623
transform 1 0 30321 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_82
timestamp 1694700623
transform 1 0 29064 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_83
timestamp 1694700623
transform 1 0 29174 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_84
timestamp 1694700623
transform 1 0 29059 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_85
timestamp 1694700623
transform 1 0 29053 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_86
timestamp 1694700623
transform 1 0 29073 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_87
timestamp 1694700623
transform 1 0 27816 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_88
timestamp 1694700623
transform 1 0 27926 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_89
timestamp 1694700623
transform 1 0 27811 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_90
timestamp 1694700623
transform 1 0 27805 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_91
timestamp 1694700623
transform 1 0 27825 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_92
timestamp 1694700623
transform 1 0 26568 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_93
timestamp 1694700623
transform 1 0 26678 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_94
timestamp 1694700623
transform 1 0 26563 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_95
timestamp 1694700623
transform 1 0 26557 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_96
timestamp 1694700623
transform 1 0 26577 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_97
timestamp 1694700623
transform 1 0 25320 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_98
timestamp 1694700623
transform 1 0 25430 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_99
timestamp 1694700623
transform 1 0 25315 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_100
timestamp 1694700623
transform 1 0 25309 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_101
timestamp 1694700623
transform 1 0 25329 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_102
timestamp 1694700623
transform 1 0 24072 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_103
timestamp 1694700623
transform 1 0 24182 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_104
timestamp 1694700623
transform 1 0 24067 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_105
timestamp 1694700623
transform 1 0 24061 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_106
timestamp 1694700623
transform 1 0 24081 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_107
timestamp 1694700623
transform 1 0 22824 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_108
timestamp 1694700623
transform 1 0 22934 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_109
timestamp 1694700623
transform 1 0 22819 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_110
timestamp 1694700623
transform 1 0 22813 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_111
timestamp 1694700623
transform 1 0 22833 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_112
timestamp 1694700623
transform 1 0 21576 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_113
timestamp 1694700623
transform 1 0 21686 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_114
timestamp 1694700623
transform 1 0 21571 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_115
timestamp 1694700623
transform 1 0 21565 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_116
timestamp 1694700623
transform 1 0 21585 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_117
timestamp 1694700623
transform 1 0 30312 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_118
timestamp 1694700623
transform 1 0 30422 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_119
timestamp 1694700623
transform 1 0 30307 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_120
timestamp 1694700623
transform 1 0 40296 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_121
timestamp 1694700623
transform 1 0 40406 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_122
timestamp 1694700623
transform 1 0 40291 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_123
timestamp 1694700623
transform 1 0 40285 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_124
timestamp 1694700623
transform 1 0 40305 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_125
timestamp 1694700623
transform 1 0 39048 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_126
timestamp 1694700623
transform 1 0 39158 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_127
timestamp 1694700623
transform 1 0 39043 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_128
timestamp 1694700623
transform 1 0 39037 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_129
timestamp 1694700623
transform 1 0 39057 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_130
timestamp 1694700623
transform 1 0 37800 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_131
timestamp 1694700623
transform 1 0 37910 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_132
timestamp 1694700623
transform 1 0 37795 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_133
timestamp 1694700623
transform 1 0 37789 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_134
timestamp 1694700623
transform 1 0 37809 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_135
timestamp 1694700623
transform 1 0 36552 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_136
timestamp 1694700623
transform 1 0 36662 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_137
timestamp 1694700623
transform 1 0 36547 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_138
timestamp 1694700623
transform 1 0 36541 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_139
timestamp 1694700623
transform 1 0 36561 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_140
timestamp 1694700623
transform 1 0 35304 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_141
timestamp 1694700623
transform 1 0 35414 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_142
timestamp 1694700623
transform 1 0 35299 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_143
timestamp 1694700623
transform 1 0 35293 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_144
timestamp 1694700623
transform 1 0 35313 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_145
timestamp 1694700623
transform 1 0 34056 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_146
timestamp 1694700623
transform 1 0 34166 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_147
timestamp 1694700623
transform 1 0 34051 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_148
timestamp 1694700623
transform 1 0 34045 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_149
timestamp 1694700623
transform 1 0 34065 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_150
timestamp 1694700623
transform 1 0 32808 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_151
timestamp 1694700623
transform 1 0 32918 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_152
timestamp 1694700623
transform 1 0 32803 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_153
timestamp 1694700623
transform 1 0 32797 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_154
timestamp 1694700623
transform 1 0 32817 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_155
timestamp 1694700623
transform 1 0 31560 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_156
timestamp 1694700623
transform 1 0 31670 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_157
timestamp 1694700623
transform 1 0 31555 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_158
timestamp 1694700623
transform 1 0 31549 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_22  sky130_sram_1kbyte_1rw1r_32x256_8_contact_22_159
timestamp 1694700623
transform 1 0 31569 0 1 154
box 0 0 1 1
<< labels >>
rlabel metal3 s 40269 1092 40367 1190 4 vdd
port 1 nsew
rlabel metal3 s 21549 1092 21647 1190 4 vdd
port 1 nsew
rlabel metal3 s 31533 1092 31631 1190 4 vdd
port 1 nsew
rlabel metal3 s 26541 1092 26639 1190 4 vdd
port 1 nsew
rlabel metal3 s 30285 1092 30383 1190 4 vdd
port 1 nsew
rlabel metal3 s 27789 1092 27887 1190 4 vdd
port 1 nsew
rlabel metal3 s 24045 1092 24143 1190 4 vdd
port 1 nsew
rlabel metal3 s 36525 1092 36623 1190 4 vdd
port 1 nsew
rlabel metal3 s 37773 1092 37871 1190 4 vdd
port 1 nsew
rlabel metal3 s 39021 1092 39119 1190 4 vdd
port 1 nsew
rlabel metal3 s 34029 1092 34127 1190 4 vdd
port 1 nsew
rlabel metal3 s 25293 1092 25391 1190 4 vdd
port 1 nsew
rlabel metal3 s 29037 1092 29135 1190 4 vdd
port 1 nsew
rlabel metal3 s 22797 1092 22895 1190 4 vdd
port 1 nsew
rlabel metal3 s 35277 1092 35375 1190 4 vdd
port 1 nsew
rlabel metal3 s 32781 1092 32879 1190 4 vdd
port 1 nsew
rlabel metal3 s 27800 1529 27898 1627 4 gnd
port 2 nsew
rlabel metal3 s 26552 1529 26650 1627 4 gnd
port 2 nsew
rlabel metal3 s 39142 760 39240 858 4 gnd
port 2 nsew
rlabel metal3 s 40390 760 40488 858 4 gnd
port 2 nsew
rlabel metal3 s 34040 1529 34138 1627 4 gnd
port 2 nsew
rlabel metal3 s 31654 760 31752 858 4 gnd
port 2 nsew
rlabel metal3 s 34150 760 34248 858 4 gnd
port 2 nsew
rlabel metal3 s 32792 1529 32890 1627 4 gnd
port 2 nsew
rlabel metal3 s 30406 760 30504 858 4 gnd
port 2 nsew
rlabel metal3 s 27795 558 27893 656 4 gnd
port 2 nsew
rlabel metal3 s 21555 558 21653 656 4 gnd
port 2 nsew
rlabel metal3 s 30291 558 30389 656 4 gnd
port 2 nsew
rlabel metal3 s 24056 1529 24154 1627 4 gnd
port 2 nsew
rlabel metal3 s 29158 760 29256 858 4 gnd
port 2 nsew
rlabel metal3 s 37779 558 37877 656 4 gnd
port 2 nsew
rlabel metal3 s 22918 760 23016 858 4 gnd
port 2 nsew
rlabel metal3 s 22803 558 22901 656 4 gnd
port 2 nsew
rlabel metal3 s 21670 760 21768 858 4 gnd
port 2 nsew
rlabel metal3 s 40275 558 40373 656 4 gnd
port 2 nsew
rlabel metal3 s 27910 760 28008 858 4 gnd
port 2 nsew
rlabel metal3 s 26662 760 26760 858 4 gnd
port 2 nsew
rlabel metal3 s 29048 1529 29146 1627 4 gnd
port 2 nsew
rlabel metal3 s 25414 760 25512 858 4 gnd
port 2 nsew
rlabel metal3 s 30296 1529 30394 1627 4 gnd
port 2 nsew
rlabel metal3 s 32787 558 32885 656 4 gnd
port 2 nsew
rlabel metal3 s 29043 558 29141 656 4 gnd
port 2 nsew
rlabel metal3 s 31544 1529 31642 1627 4 gnd
port 2 nsew
rlabel metal3 s 31539 558 31637 656 4 gnd
port 2 nsew
rlabel metal3 s 36531 558 36629 656 4 gnd
port 2 nsew
rlabel metal3 s 37784 1529 37882 1627 4 gnd
port 2 nsew
rlabel metal3 s 39027 558 39125 656 4 gnd
port 2 nsew
rlabel metal3 s 40280 1529 40378 1627 4 gnd
port 2 nsew
rlabel metal3 s 22808 1529 22906 1627 4 gnd
port 2 nsew
rlabel metal3 s 37894 760 37992 858 4 gnd
port 2 nsew
rlabel metal3 s 35283 558 35381 656 4 gnd
port 2 nsew
rlabel metal3 s 24166 760 24264 858 4 gnd
port 2 nsew
rlabel metal3 s 35398 760 35496 858 4 gnd
port 2 nsew
rlabel metal3 s 39032 1529 39130 1627 4 gnd
port 2 nsew
rlabel metal3 s 32902 760 33000 858 4 gnd
port 2 nsew
rlabel metal3 s 35288 1529 35386 1627 4 gnd
port 2 nsew
rlabel metal3 s 24051 558 24149 656 4 gnd
port 2 nsew
rlabel metal3 s 25304 1529 25402 1627 4 gnd
port 2 nsew
rlabel metal3 s 34035 558 34133 656 4 gnd
port 2 nsew
rlabel metal3 s 21560 1529 21658 1627 4 gnd
port 2 nsew
rlabel metal3 s 36536 1529 36634 1627 4 gnd
port 2 nsew
rlabel metal3 s 25299 558 25397 656 4 gnd
port 2 nsew
rlabel metal3 s 26547 558 26645 656 4 gnd
port 2 nsew
rlabel metal3 s 36646 760 36744 858 4 gnd
port 2 nsew
rlabel metal3 s 11686 760 11784 858 4 gnd
port 2 nsew
rlabel metal3 s 15320 1529 15418 1627 4 gnd
port 2 nsew
rlabel metal3 s 7942 760 8040 858 4 gnd
port 2 nsew
rlabel metal3 s 19053 1092 19151 1190 4 vdd
port 1 nsew
rlabel metal3 s 20301 1092 20399 1190 4 vdd
port 1 nsew
rlabel metal3 s 6579 558 6677 656 4 gnd
port 2 nsew
rlabel metal3 s 5446 760 5544 858 4 gnd
port 2 nsew
rlabel metal3 s 19064 1529 19162 1627 4 gnd
port 2 nsew
rlabel metal3 s 5325 1092 5423 1190 4 vdd
port 1 nsew
rlabel metal3 s 6694 760 6792 858 4 gnd
port 2 nsew
rlabel metal3 s 20312 1529 20410 1627 4 gnd
port 2 nsew
rlabel metal3 s 20422 760 20520 858 4 gnd
port 2 nsew
rlabel metal3 s 10323 558 10421 656 4 gnd
port 2 nsew
rlabel metal3 s 20307 558 20405 656 4 gnd
port 2 nsew
rlabel metal3 s 14072 1529 14170 1627 4 gnd
port 2 nsew
rlabel metal3 s 19059 558 19157 656 4 gnd
port 2 nsew
rlabel metal3 s 6573 1092 6671 1190 4 vdd
port 1 nsew
rlabel metal3 s 9069 1092 9167 1190 4 vdd
port 1 nsew
rlabel metal3 s 4198 760 4296 858 4 gnd
port 2 nsew
rlabel metal3 s 5331 558 5429 656 4 gnd
port 2 nsew
rlabel metal3 s 12819 558 12917 656 4 gnd
port 2 nsew
rlabel metal3 s 10317 1092 10415 1190 4 vdd
port 1 nsew
rlabel metal3 s 1702 760 1800 858 4 gnd
port 2 nsew
rlabel metal3 s 9075 558 9173 656 4 gnd
port 2 nsew
rlabel metal3 s 11571 558 11669 656 4 gnd
port 2 nsew
rlabel metal3 s 4077 1092 4175 1190 4 vdd
port 1 nsew
rlabel metal3 s 4083 558 4181 656 4 gnd
port 2 nsew
rlabel metal3 s 12824 1529 12922 1627 4 gnd
port 2 nsew
rlabel metal3 s 1581 1092 1679 1190 4 vdd
port 1 nsew
rlabel metal3 s 7832 1529 7930 1627 4 gnd
port 2 nsew
rlabel metal3 s 17805 1092 17903 1190 4 vdd
port 1 nsew
rlabel metal3 s 6584 1529 6682 1627 4 gnd
port 2 nsew
rlabel metal3 s 1587 558 1685 656 4 gnd
port 2 nsew
rlabel metal3 s 17811 558 17909 656 4 gnd
port 2 nsew
rlabel metal3 s 5336 1529 5434 1627 4 gnd
port 2 nsew
rlabel metal3 s 2840 1529 2938 1627 4 gnd
port 2 nsew
rlabel metal3 s 9190 760 9288 858 4 gnd
port 2 nsew
rlabel metal3 s 7827 558 7925 656 4 gnd
port 2 nsew
rlabel metal3 s 14061 1092 14159 1190 4 vdd
port 1 nsew
rlabel metal3 s 16678 760 16776 858 4 gnd
port 2 nsew
rlabel metal3 s 17926 760 18024 858 4 gnd
port 2 nsew
rlabel metal3 s 4088 1529 4186 1627 4 gnd
port 2 nsew
rlabel metal3 s 1592 1529 1690 1627 4 gnd
port 2 nsew
rlabel metal3 s 10328 1529 10426 1627 4 gnd
port 2 nsew
rlabel metal3 s 12813 1092 12911 1190 4 vdd
port 1 nsew
rlabel metal3 s 17816 1529 17914 1627 4 gnd
port 2 nsew
rlabel metal3 s 2829 1092 2927 1190 4 vdd
port 1 nsew
rlabel metal3 s 14067 558 14165 656 4 gnd
port 2 nsew
rlabel metal3 s 19174 760 19272 858 4 gnd
port 2 nsew
rlabel metal3 s 15309 1092 15407 1190 4 vdd
port 1 nsew
rlabel metal3 s 15315 558 15413 656 4 gnd
port 2 nsew
rlabel metal3 s 15430 760 15528 858 4 gnd
port 2 nsew
rlabel metal3 s 16557 1092 16655 1190 4 vdd
port 1 nsew
rlabel metal3 s 11565 1092 11663 1190 4 vdd
port 1 nsew
rlabel metal3 s 11576 1529 11674 1627 4 gnd
port 2 nsew
rlabel metal3 s 12934 760 13032 858 4 gnd
port 2 nsew
rlabel metal3 s 10438 760 10536 858 4 gnd
port 2 nsew
rlabel metal3 s 16568 1529 16666 1627 4 gnd
port 2 nsew
rlabel metal3 s 9080 1529 9178 1627 4 gnd
port 2 nsew
rlabel metal3 s 2950 760 3048 858 4 gnd
port 2 nsew
rlabel metal3 s 14182 760 14280 858 4 gnd
port 2 nsew
rlabel metal3 s 7821 1092 7919 1190 4 vdd
port 1 nsew
rlabel metal3 s 16563 558 16661 656 4 gnd
port 2 nsew
rlabel metal3 s 2835 558 2933 656 4 gnd
port 2 nsew
rlabel metal3 s 4097 142 4195 240 4 vdd
port 1 nsew
rlabel metal3 s 1601 142 1699 240 4 vdd
port 1 nsew
rlabel metal3 s 14081 142 14179 240 4 vdd
port 1 nsew
rlabel metal3 s 20321 142 20419 240 4 vdd
port 1 nsew
rlabel metal3 s 7841 142 7939 240 4 vdd
port 1 nsew
rlabel metal3 s 12833 142 12931 240 4 vdd
port 1 nsew
rlabel metal3 s 2849 142 2947 240 4 vdd
port 1 nsew
rlabel metal3 s 10337 142 10435 240 4 vdd
port 1 nsew
rlabel metal3 s 11585 142 11683 240 4 vdd
port 1 nsew
rlabel metal3 s 17825 142 17923 240 4 vdd
port 1 nsew
rlabel metal3 s 9089 142 9187 240 4 vdd
port 1 nsew
rlabel metal3 s 19073 142 19171 240 4 vdd
port 1 nsew
rlabel metal3 s 6593 142 6691 240 4 vdd
port 1 nsew
rlabel metal3 s 5345 142 5443 240 4 vdd
port 1 nsew
rlabel metal3 s 16577 142 16675 240 4 vdd
port 1 nsew
rlabel metal3 s 15329 142 15427 240 4 vdd
port 1 nsew
rlabel metal3 s 22817 142 22915 240 4 vdd
port 1 nsew
rlabel metal3 s 27809 142 27907 240 4 vdd
port 1 nsew
rlabel metal3 s 24065 142 24163 240 4 vdd
port 1 nsew
rlabel metal3 s 31553 142 31651 240 4 vdd
port 1 nsew
rlabel metal3 s 32801 142 32899 240 4 vdd
port 1 nsew
rlabel metal3 s 30305 142 30403 240 4 vdd
port 1 nsew
rlabel metal3 s 40289 142 40387 240 4 vdd
port 1 nsew
rlabel metal3 s 39041 142 39139 240 4 vdd
port 1 nsew
rlabel metal3 s 35297 142 35395 240 4 vdd
port 1 nsew
rlabel metal3 s 25313 142 25411 240 4 vdd
port 1 nsew
rlabel metal3 s 37793 142 37891 240 4 vdd
port 1 nsew
rlabel metal3 s 26561 142 26659 240 4 vdd
port 1 nsew
rlabel metal3 s 21569 142 21667 240 4 vdd
port 1 nsew
rlabel metal3 s 34049 142 34147 240 4 vdd
port 1 nsew
rlabel metal3 s 29057 142 29155 240 4 vdd
port 1 nsew
rlabel metal3 s 36545 142 36643 240 4 vdd
port 1 nsew
rlabel metal1 s 1629 4 1689 60 4 data_0
port 3 nsew
rlabel metal1 s 1500 1959 1530 2011 4 bl_0
port 4 nsew
rlabel metal1 s 1702 1959 1732 2011 4 br_0
port 5 nsew
rlabel metal1 s 2877 4 2937 60 4 data_1
port 6 nsew
rlabel metal1 s 2748 1959 2778 2011 4 bl_1
port 7 nsew
rlabel metal1 s 2950 1959 2980 2011 4 br_1
port 8 nsew
rlabel metal1 s 4125 4 4185 60 4 data_2
port 9 nsew
rlabel metal1 s 3996 1959 4026 2011 4 bl_2
port 10 nsew
rlabel metal1 s 4198 1959 4228 2011 4 br_2
port 11 nsew
rlabel metal1 s 5373 4 5433 60 4 data_3
port 12 nsew
rlabel metal1 s 5244 1959 5274 2011 4 bl_3
port 13 nsew
rlabel metal1 s 5446 1959 5476 2011 4 br_3
port 14 nsew
rlabel metal1 s 6621 4 6681 60 4 data_4
port 15 nsew
rlabel metal1 s 6492 1959 6522 2011 4 bl_4
port 16 nsew
rlabel metal1 s 6694 1959 6724 2011 4 br_4
port 17 nsew
rlabel metal1 s 7869 4 7929 60 4 data_5
port 18 nsew
rlabel metal1 s 7740 1959 7770 2011 4 bl_5
port 19 nsew
rlabel metal1 s 7942 1959 7972 2011 4 br_5
port 20 nsew
rlabel metal1 s 9117 4 9177 60 4 data_6
port 21 nsew
rlabel metal1 s 8988 1959 9018 2011 4 bl_6
port 22 nsew
rlabel metal1 s 9190 1959 9220 2011 4 br_6
port 23 nsew
rlabel metal1 s 10365 4 10425 60 4 data_7
port 24 nsew
rlabel metal1 s 10236 1959 10266 2011 4 bl_7
port 25 nsew
rlabel metal1 s 10438 1959 10468 2011 4 br_7
port 26 nsew
rlabel metal1 s 11613 4 11673 60 4 data_8
port 27 nsew
rlabel metal1 s 11484 1959 11514 2011 4 bl_8
port 28 nsew
rlabel metal1 s 11686 1959 11716 2011 4 br_8
port 29 nsew
rlabel metal1 s 12861 4 12921 60 4 data_9
port 30 nsew
rlabel metal1 s 12732 1959 12762 2011 4 bl_9
port 31 nsew
rlabel metal1 s 12934 1959 12964 2011 4 br_9
port 32 nsew
rlabel metal1 s 14109 4 14169 60 4 data_10
port 33 nsew
rlabel metal1 s 13980 1959 14010 2011 4 bl_10
port 34 nsew
rlabel metal1 s 14182 1959 14212 2011 4 br_10
port 35 nsew
rlabel metal1 s 15357 4 15417 60 4 data_11
port 36 nsew
rlabel metal1 s 15228 1959 15258 2011 4 bl_11
port 37 nsew
rlabel metal1 s 15430 1959 15460 2011 4 br_11
port 38 nsew
rlabel metal1 s 16605 4 16665 60 4 data_12
port 39 nsew
rlabel metal1 s 16476 1959 16506 2011 4 bl_12
port 40 nsew
rlabel metal1 s 16678 1959 16708 2011 4 br_12
port 41 nsew
rlabel metal1 s 17853 4 17913 60 4 data_13
port 42 nsew
rlabel metal1 s 17724 1959 17754 2011 4 bl_13
port 43 nsew
rlabel metal1 s 17926 1959 17956 2011 4 br_13
port 44 nsew
rlabel metal1 s 19101 4 19161 60 4 data_14
port 45 nsew
rlabel metal1 s 18972 1959 19002 2011 4 bl_14
port 46 nsew
rlabel metal1 s 19174 1959 19204 2011 4 br_14
port 47 nsew
rlabel metal1 s 20349 4 20409 60 4 data_15
port 48 nsew
rlabel metal1 s 20220 1959 20250 2011 4 bl_15
port 49 nsew
rlabel metal1 s 20422 1959 20452 2011 4 br_15
port 50 nsew
rlabel metal1 s 21597 4 21657 60 4 data_16
port 51 nsew
rlabel metal1 s 21468 1959 21498 2011 4 bl_16
port 52 nsew
rlabel metal1 s 21670 1959 21700 2011 4 br_16
port 53 nsew
rlabel metal1 s 22845 4 22905 60 4 data_17
port 54 nsew
rlabel metal1 s 22716 1959 22746 2011 4 bl_17
port 55 nsew
rlabel metal1 s 22918 1959 22948 2011 4 br_17
port 56 nsew
rlabel metal1 s 24093 4 24153 60 4 data_18
port 57 nsew
rlabel metal1 s 23964 1959 23994 2011 4 bl_18
port 58 nsew
rlabel metal1 s 24166 1959 24196 2011 4 br_18
port 59 nsew
rlabel metal1 s 25341 4 25401 60 4 data_19
port 60 nsew
rlabel metal1 s 25212 1959 25242 2011 4 bl_19
port 61 nsew
rlabel metal1 s 25414 1959 25444 2011 4 br_19
port 62 nsew
rlabel metal1 s 26589 4 26649 60 4 data_20
port 63 nsew
rlabel metal1 s 26460 1959 26490 2011 4 bl_20
port 64 nsew
rlabel metal1 s 26662 1959 26692 2011 4 br_20
port 65 nsew
rlabel metal1 s 27837 4 27897 60 4 data_21
port 66 nsew
rlabel metal1 s 27708 1959 27738 2011 4 bl_21
port 67 nsew
rlabel metal1 s 27910 1959 27940 2011 4 br_21
port 68 nsew
rlabel metal1 s 29085 4 29145 60 4 data_22
port 69 nsew
rlabel metal1 s 28956 1959 28986 2011 4 bl_22
port 70 nsew
rlabel metal1 s 29158 1959 29188 2011 4 br_22
port 71 nsew
rlabel metal1 s 30333 4 30393 60 4 data_23
port 72 nsew
rlabel metal1 s 30204 1959 30234 2011 4 bl_23
port 73 nsew
rlabel metal1 s 30406 1959 30436 2011 4 br_23
port 74 nsew
rlabel metal1 s 31581 4 31641 60 4 data_24
port 75 nsew
rlabel metal1 s 31452 1959 31482 2011 4 bl_24
port 76 nsew
rlabel metal1 s 31654 1959 31684 2011 4 br_24
port 77 nsew
rlabel metal1 s 32829 4 32889 60 4 data_25
port 78 nsew
rlabel metal1 s 32700 1959 32730 2011 4 bl_25
port 79 nsew
rlabel metal1 s 32902 1959 32932 2011 4 br_25
port 80 nsew
rlabel metal1 s 34077 4 34137 60 4 data_26
port 81 nsew
rlabel metal1 s 33948 1959 33978 2011 4 bl_26
port 82 nsew
rlabel metal1 s 34150 1959 34180 2011 4 br_26
port 83 nsew
rlabel metal1 s 35325 4 35385 60 4 data_27
port 84 nsew
rlabel metal1 s 35196 1959 35226 2011 4 bl_27
port 85 nsew
rlabel metal1 s 35398 1959 35428 2011 4 br_27
port 86 nsew
rlabel metal1 s 36573 4 36633 60 4 data_28
port 87 nsew
rlabel metal1 s 36444 1959 36474 2011 4 bl_28
port 88 nsew
rlabel metal1 s 36646 1959 36676 2011 4 br_28
port 89 nsew
rlabel metal1 s 37821 4 37881 60 4 data_29
port 90 nsew
rlabel metal1 s 37692 1959 37722 2011 4 bl_29
port 91 nsew
rlabel metal1 s 37894 1959 37924 2011 4 br_29
port 92 nsew
rlabel metal1 s 39069 4 39129 60 4 data_30
port 93 nsew
rlabel metal1 s 38940 1959 38970 2011 4 bl_30
port 94 nsew
rlabel metal1 s 39142 1959 39172 2011 4 br_30
port 95 nsew
rlabel metal1 s 40317 4 40377 60 4 data_31
port 96 nsew
rlabel metal1 s 40188 1959 40218 2011 4 bl_31
port 97 nsew
rlabel metal1 s 40390 1959 40420 2011 4 br_31
port 98 nsew
rlabel metal1 s 1473 94 10833 128 4 en_0
port 99 nsew
rlabel metal1 s 11457 94 20817 128 4 en_1
port 100 nsew
rlabel metal1 s 21441 94 30801 128 4 en_2
port 101 nsew
rlabel metal1 s 31425 94 40785 128 4 en_3
port 102 nsew
<< properties >>
string FIXED_BBOX 0 0 40562 2011
string GDS_END 1195608
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 1113880
<< end >>
