magic
tech sky130B
timestamp 1694700623
<< properties >>
string GDS_END 15503532
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15500328
<< end >>
