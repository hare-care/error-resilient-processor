magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< locali >>
rect 167 752 179 786
rect 213 752 251 786
rect 285 752 323 786
rect 357 752 369 786
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 454 672 488 674
rect 454 600 488 638
rect 454 528 488 566
rect 454 456 488 494
rect 454 384 488 422
rect 454 312 488 350
rect 454 240 488 278
rect 454 168 488 206
rect 454 132 488 134
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
<< viali >>
rect 179 752 213 786
rect 251 752 285 786
rect 323 752 357 786
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 454 638 488 672
rect 454 566 488 600
rect 454 494 488 528
rect 454 422 488 456
rect 454 350 488 384
rect 454 278 488 312
rect 454 206 488 240
rect 454 134 488 168
rect 179 20 213 54
rect 251 20 285 54
rect 323 20 357 54
<< obsli1 >>
rect 159 98 193 708
rect 251 98 285 708
rect 343 98 377 708
<< metal1 >>
rect 167 786 369 806
rect 167 752 179 786
rect 213 752 251 786
rect 285 752 323 786
rect 357 752 369 786
rect 167 740 369 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 442 672 500 684
rect 442 638 454 672
rect 488 638 500 672
rect 442 600 500 638
rect 442 566 454 600
rect 488 566 500 600
rect 442 528 500 566
rect 442 494 454 528
rect 488 494 500 528
rect 442 456 500 494
rect 442 422 454 456
rect 488 422 500 456
rect 442 384 500 422
rect 442 350 454 384
rect 488 350 500 384
rect 442 312 500 350
rect 442 278 454 312
rect 488 278 500 312
rect 442 240 500 278
rect 442 206 454 240
rect 488 206 500 240
rect 442 168 500 206
rect 442 134 454 168
rect 488 134 500 168
rect 442 122 500 134
rect 167 54 369 66
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
rect 167 0 369 20
<< obsm1 >>
rect 150 122 202 684
rect 242 122 294 684
rect 334 122 386 684
<< metal2 >>
rect 10 428 526 684
rect 10 122 526 378
<< labels >>
rlabel viali s 454 638 488 672 6 BULK
port 1 nsew
rlabel viali s 454 566 488 600 6 BULK
port 1 nsew
rlabel viali s 454 494 488 528 6 BULK
port 1 nsew
rlabel viali s 454 422 488 456 6 BULK
port 1 nsew
rlabel viali s 454 350 488 384 6 BULK
port 1 nsew
rlabel viali s 454 278 488 312 6 BULK
port 1 nsew
rlabel viali s 454 206 488 240 6 BULK
port 1 nsew
rlabel viali s 454 134 488 168 6 BULK
port 1 nsew
rlabel viali s 48 638 82 672 6 BULK
port 1 nsew
rlabel viali s 48 566 82 600 6 BULK
port 1 nsew
rlabel viali s 48 494 82 528 6 BULK
port 1 nsew
rlabel viali s 48 422 82 456 6 BULK
port 1 nsew
rlabel viali s 48 350 82 384 6 BULK
port 1 nsew
rlabel viali s 48 278 82 312 6 BULK
port 1 nsew
rlabel viali s 48 206 82 240 6 BULK
port 1 nsew
rlabel viali s 48 134 82 168 6 BULK
port 1 nsew
rlabel locali s 454 132 488 674 6 BULK
port 1 nsew
rlabel locali s 48 132 82 674 6 BULK
port 1 nsew
rlabel metal1 s 442 122 500 684 6 BULK
port 1 nsew
rlabel metal1 s 36 122 94 684 6 BULK
port 1 nsew
rlabel metal2 s 10 428 526 684 6 DRAIN
port 2 nsew
rlabel viali s 323 752 357 786 6 GATE
port 3 nsew
rlabel viali s 323 20 357 54 6 GATE
port 3 nsew
rlabel viali s 251 752 285 786 6 GATE
port 3 nsew
rlabel viali s 251 20 285 54 6 GATE
port 3 nsew
rlabel viali s 179 752 213 786 6 GATE
port 3 nsew
rlabel viali s 179 20 213 54 6 GATE
port 3 nsew
rlabel locali s 167 752 369 786 6 GATE
port 3 nsew
rlabel locali s 167 20 369 54 6 GATE
port 3 nsew
rlabel metal1 s 167 740 369 806 6 GATE
port 3 nsew
rlabel metal1 s 167 0 369 66 6 GATE
port 3 nsew
rlabel metal2 s 10 122 526 378 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 536 806
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9273642
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9262726
<< end >>
