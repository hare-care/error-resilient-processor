magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< locali >>
rect 0 1396 1940 1432
rect 1510 909 1544 925
rect 1509 875 1510 892
rect 1509 859 1544 875
rect 1509 726 1543 859
rect 1268 705 1302 721
rect 1509 705 1653 726
rect 1400 692 1653 705
rect 1768 692 1887 726
rect 1400 671 1543 692
rect 1268 655 1302 671
rect 1853 522 1887 692
rect 1853 472 1887 488
rect 0 -20 1940 16
<< viali >>
rect 1510 875 1544 909
rect 1268 671 1302 705
rect 1853 488 1887 522
<< metal1 >>
rect 1494 866 1500 918
rect 1552 866 1559 918
rect 1253 662 1259 714
rect 1311 662 1317 714
rect 1838 479 1844 531
rect 1896 479 1902 531
<< via1 >>
rect 1500 909 1552 918
rect 1500 875 1510 909
rect 1510 875 1544 909
rect 1544 875 1552 909
rect 1500 866 1552 875
rect 1259 705 1311 714
rect 1259 671 1268 705
rect 1268 671 1302 705
rect 1302 671 1311 705
rect 1259 662 1311 671
rect 1844 522 1896 531
rect 1844 488 1853 522
rect 1853 488 1887 522
rect 1887 488 1896 522
rect 1844 479 1896 488
<< metal2 >>
rect 1500 918 1552 924
rect 1500 860 1552 866
rect 369 692 423 756
rect 1259 714 1311 720
rect 1259 661 1311 662
rect 1115 609 1311 661
rect 137 538 203 590
rect 1844 531 1896 537
rect 1844 473 1896 479
use contact_7  contact_7_0
timestamp 1694700623
transform 1 0 1498 0 1 859
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1694700623
transform 1 0 1841 0 1 472
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1694700623
transform 1 0 1256 0 1 655
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1694700623
transform 1 0 1494 0 1 860
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1694700623
transform 1 0 1838 0 1 473
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1694700623
transform 1 0 1253 0 1 656
box 0 0 1 1
use dff  dff_0
timestamp 1694700623
transform 1 0 0 0 1 0
box -8 -43 1176 1467
use pinv_1  pinv_1_0
timestamp 1694700623
transform 1 0 1204 0 1 0
box -36 -17 404 1471
use pinv_2  pinv_2_0
timestamp 1694700623
transform 1 0 1572 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 970 1414 970 1414 4 vdd
port 5 nsew
rlabel locali s 970 -2 970 -2 4 gnd
port 6 nsew
rlabel metal2 s 170 564 170 564 4 D
port 1 nsew
rlabel metal2 s 1870 505 1870 505 4 Q
port 2 nsew
rlabel metal2 s 1526 892 1526 892 4 Qb
port 3 nsew
rlabel metal2 s 396 724 396 724 4 clk
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1940 1414
string GDS_END 4235272
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4233162
<< end >>
