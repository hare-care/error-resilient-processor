magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 604 203
rect 1 67 827 157
rect 29 21 827 67
rect 29 -17 63 21
<< scnmos >>
rect 79 93 109 177
rect 188 47 218 177
rect 296 47 326 177
rect 396 47 426 177
rect 496 47 526 177
rect 684 47 714 131
<< scpmoshvt >>
rect 79 413 109 497
rect 188 297 218 497
rect 296 297 326 497
rect 396 297 426 497
rect 496 297 526 497
rect 684 413 714 497
<< ndiff >>
rect 27 139 79 177
rect 27 105 35 139
rect 69 105 79 139
rect 27 93 79 105
rect 109 93 188 177
rect 124 59 132 93
rect 166 59 188 93
rect 124 47 188 59
rect 218 47 296 177
rect 326 47 396 177
rect 426 47 496 177
rect 526 161 578 177
rect 526 127 536 161
rect 570 127 578 161
rect 526 93 578 127
rect 526 59 536 93
rect 570 59 578 93
rect 526 47 578 59
rect 632 93 684 131
rect 632 59 640 93
rect 674 59 684 93
rect 632 47 684 59
rect 714 93 801 131
rect 714 59 743 93
rect 777 59 801 93
rect 714 47 801 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 413 79 451
rect 109 485 188 497
rect 109 451 135 485
rect 169 451 188 485
rect 109 413 188 451
rect 124 401 188 413
rect 124 367 135 401
rect 169 367 188 401
rect 124 297 188 367
rect 218 485 296 497
rect 218 451 240 485
rect 274 451 296 485
rect 218 417 296 451
rect 218 383 240 417
rect 274 383 296 417
rect 218 349 296 383
rect 218 315 240 349
rect 274 315 296 349
rect 218 297 296 315
rect 326 485 396 497
rect 326 451 344 485
rect 378 451 396 485
rect 326 417 396 451
rect 326 383 344 417
rect 378 383 396 417
rect 326 297 396 383
rect 426 485 496 497
rect 426 451 444 485
rect 478 451 496 485
rect 426 417 496 451
rect 426 383 444 417
rect 478 383 496 417
rect 426 349 496 383
rect 426 315 444 349
rect 478 315 496 349
rect 426 297 496 315
rect 526 485 578 497
rect 526 451 536 485
rect 570 451 578 485
rect 526 297 578 451
rect 632 485 684 497
rect 632 451 640 485
rect 674 451 684 485
rect 632 413 684 451
rect 714 485 801 497
rect 714 451 743 485
rect 777 451 801 485
rect 714 413 801 451
<< ndiffc >>
rect 35 105 69 139
rect 132 59 166 93
rect 536 127 570 161
rect 536 59 570 93
rect 640 59 674 93
rect 743 59 777 93
<< pdiffc >>
rect 35 451 69 485
rect 135 451 169 485
rect 135 367 169 401
rect 240 451 274 485
rect 240 383 274 417
rect 240 315 274 349
rect 344 451 378 485
rect 344 383 378 417
rect 444 451 478 485
rect 444 383 478 417
rect 444 315 478 349
rect 536 451 570 485
rect 640 451 674 485
rect 743 451 777 485
<< poly >>
rect 79 497 109 523
rect 188 497 218 523
rect 296 497 326 523
rect 396 497 426 523
rect 496 497 526 523
rect 684 497 714 523
rect 79 265 109 413
rect 188 265 218 297
rect 296 265 326 297
rect 396 265 426 297
rect 496 265 526 297
rect 79 249 146 265
rect 79 215 102 249
rect 136 215 146 249
rect 79 199 146 215
rect 188 249 254 265
rect 188 215 210 249
rect 244 215 254 249
rect 188 199 254 215
rect 296 249 354 265
rect 296 215 310 249
rect 344 215 354 249
rect 296 199 354 215
rect 396 249 450 265
rect 396 215 406 249
rect 440 215 450 249
rect 396 199 450 215
rect 496 249 618 265
rect 496 215 568 249
rect 602 215 618 249
rect 496 199 618 215
rect 684 264 714 413
rect 684 248 738 264
rect 684 214 694 248
rect 728 214 738 248
rect 79 177 109 199
rect 188 177 218 199
rect 296 177 326 199
rect 396 177 426 199
rect 496 177 526 199
rect 684 198 738 214
rect 79 67 109 93
rect 684 131 714 198
rect 188 21 218 47
rect 296 21 326 47
rect 396 21 426 47
rect 496 21 526 47
rect 684 21 714 47
<< polycont >>
rect 102 215 136 249
rect 210 215 244 249
rect 310 215 344 249
rect 406 215 440 249
rect 568 215 602 249
rect 694 214 728 248
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 413 85 451
rect 119 485 185 527
rect 119 451 135 485
rect 169 451 185 485
rect 17 181 52 413
rect 119 401 185 451
rect 119 367 135 401
rect 169 367 185 401
rect 224 485 290 493
rect 224 451 240 485
rect 274 451 290 485
rect 224 417 290 451
rect 224 383 240 417
rect 274 383 290 417
rect 224 349 290 383
rect 328 485 394 527
rect 328 451 344 485
rect 378 451 394 485
rect 328 417 394 451
rect 328 383 344 417
rect 378 383 394 417
rect 328 367 394 383
rect 428 485 494 493
rect 428 451 444 485
rect 478 451 494 485
rect 428 417 494 451
rect 536 485 690 527
rect 570 451 640 485
rect 674 451 690 485
rect 536 435 690 451
rect 727 485 811 493
rect 727 451 743 485
rect 777 451 811 485
rect 428 383 444 417
rect 478 383 494 417
rect 727 401 811 451
rect 86 249 156 331
rect 224 315 240 349
rect 274 333 290 349
rect 428 349 494 383
rect 428 333 444 349
rect 274 315 444 333
rect 478 333 494 349
rect 568 367 811 401
rect 478 315 534 333
rect 224 299 534 315
rect 86 215 102 249
rect 136 215 156 249
rect 194 249 264 265
rect 194 215 210 249
rect 244 215 264 249
rect 300 249 344 265
rect 300 215 310 249
rect 17 143 254 181
rect 300 147 344 215
rect 394 249 450 265
rect 394 215 406 249
rect 440 215 450 249
rect 17 139 85 143
rect 17 105 35 139
rect 69 105 85 139
rect 216 111 254 143
rect 394 111 450 215
rect 17 97 85 105
rect 119 93 180 109
rect 119 59 132 93
rect 166 59 180 93
rect 216 73 450 111
rect 484 165 534 299
rect 568 249 618 367
rect 602 215 618 249
rect 568 199 618 215
rect 678 248 728 323
rect 678 214 694 248
rect 484 161 586 165
rect 484 127 536 161
rect 570 127 586 161
rect 678 145 728 214
rect 484 93 586 127
rect 762 109 811 367
rect 119 17 180 59
rect 484 59 536 93
rect 570 59 586 93
rect 484 51 586 59
rect 620 93 690 109
rect 620 59 640 93
rect 674 59 690 93
rect 620 17 690 59
rect 724 93 811 109
rect 724 59 743 93
rect 777 59 811 93
rect 724 51 811 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 678 289 712 323 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 490 289 524 323 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 490 153 524 187 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 B_N
port 2 nsew signal input
flabel locali s 490 85 524 119 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4bb_1
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1933288
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1926132
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
