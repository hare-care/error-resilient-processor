magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 5 217 267 283
rect 5 43 467 217
rect -26 -43 506 43
<< locali >>
rect 23 435 110 751
rect 23 99 73 435
rect 293 293 359 652
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 146 735 257 751
rect 146 701 148 735
rect 182 701 220 735
rect 254 701 257 735
rect 146 435 257 701
rect 135 257 201 349
rect 395 257 445 601
rect 135 223 445 257
rect 109 113 359 187
rect 143 79 181 113
rect 215 79 253 113
rect 287 79 325 113
rect 395 99 445 223
rect 109 73 359 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 148 701 182 735
rect 220 701 254 735
rect 109 79 143 113
rect 181 79 215 113
rect 253 79 287 113
rect 325 79 359 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 148 735
rect 182 701 220 735
rect 254 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 109 113
rect 143 79 181 113
rect 215 79 253 113
rect 287 79 325 113
rect 359 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel locali s 293 293 359 652 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 480 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 480 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 506 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 5 43 467 217 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 5 217 267 283 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 480 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 546 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 480 763 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 23 99 73 435 6 X
port 6 nsew signal output
rlabel locali s 23 435 110 751 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 480 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 821242
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 813686
<< end >>
