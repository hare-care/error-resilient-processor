magic
tech sky130B
timestamp 1694700623
<< properties >>
string GDS_END 31290980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31290592
<< end >>
