magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -83 34302 16087 35388
rect -83 33688 1503 34302
rect 13394 33688 16087 34302
rect -83 33639 16087 33688
rect -83 33296 16088 33639
rect -83 28931 1277 33296
rect 15726 28931 16088 33296
rect -83 28569 16088 28931
rect 9208 27669 16088 27670
rect -83 25726 16088 27669
rect 9388 18442 16134 18626
rect 12530 18340 16134 18442
rect -83 17957 559 18073
rect -83 17290 1195 17957
rect -24 17249 1195 17290
rect -24 17141 1684 17249
rect -24 16925 1699 17141
rect -24 16709 906 16925
rect 15848 16462 16134 18340
rect 9388 16226 16134 16462
rect -143 15554 4963 15840
rect -143 12061 143 15554
rect 15848 14348 16134 16226
rect 12530 14246 16134 14348
rect 9388 14112 16134 14246
rect 15825 12802 16134 14112
rect 14067 12632 16134 12802
rect -143 11797 762 12061
rect -143 11747 2707 11797
rect -143 11629 2092 11747
rect -143 11197 143 11629
rect -143 10911 4703 11197
rect 15825 10003 16134 12632
rect 14067 9717 16134 10003
rect 9783 6446 16090 6804
rect 11655 6075 16090 6446
rect 12966 5550 16090 6075
rect 2257 3424 10099 4209
rect 0 2152 1591 2424
rect 0 1458 272 2152
rect -83 726 332 1458
rect 0 293 272 726
rect 0 272 699 293
rect 1319 272 1591 2152
rect 0 0 1591 272
rect 2257 34 10099 293
rect 12966 4209 16090 4662
rect 11657 3424 16090 4209
rect 11657 34 12298 293
rect 12806 34 13078 427
rect 0 -220 699 0
rect 2257 -220 23593 34
rect 0 -270 23593 -220
rect 0 -407 12298 -270
<< pwell >>
rect -58 27730 16058 28506
rect -43 25456 8049 25664
rect 13382 25456 16058 25664
rect -43 24620 16058 25456
rect -43 20303 1147 24620
rect 15573 20303 16058 24620
rect -43 19986 16058 20303
rect -43 18844 1043 19986
rect 7877 19757 16058 19986
rect 10576 19497 16058 19757
rect 15354 19190 16058 19497
rect 7877 18844 16058 19190
rect -43 18788 16058 18844
rect -43 18645 9168 18788
rect -43 18584 9318 18645
rect -43 18180 1860 18584
rect 699 2424 2257 4351
rect 699 2092 1319 2152
rect 332 332 1319 2092
rect 699 272 1319 332
rect 1591 0 2257 2424
rect 10099 34 11657 4351
rect 699 -220 2257 0
rect 12849 -383 13241 -270
rect 13322 -383 13642 -270
<< locali >>
rect 66 2305 1525 2358
rect 66 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1525 2305
rect 66 2218 1525 2271
rect 66 2035 206 2218
rect 66 2001 119 2035
rect 153 2001 206 2035
rect 66 1963 206 2001
rect 66 1929 119 1963
rect 153 1929 206 1963
rect 66 1891 206 1929
rect 66 1857 119 1891
rect 153 1857 206 1891
rect 66 1819 206 1857
rect 66 1785 119 1819
rect 153 1785 206 1819
rect 66 1747 206 1785
rect 66 1713 119 1747
rect 153 1713 206 1747
rect 66 1675 206 1713
rect 66 1641 119 1675
rect 153 1641 206 1675
rect 66 1603 206 1641
rect 66 1569 119 1603
rect 153 1569 206 1603
rect 66 1531 206 1569
rect 66 1497 119 1531
rect 153 1497 206 1531
rect 66 1459 206 1497
rect 66 1425 119 1459
rect 153 1425 206 1459
rect 66 1387 206 1425
rect 66 1353 119 1387
rect 153 1353 206 1387
rect 66 1315 206 1353
rect 66 1281 119 1315
rect 153 1281 206 1315
rect 66 1243 206 1281
rect 66 1209 119 1243
rect 153 1209 206 1243
rect 66 1171 206 1209
rect 66 1137 119 1171
rect 153 1137 206 1171
rect 66 1099 206 1137
rect 66 1065 119 1099
rect 153 1065 206 1099
rect 66 1027 206 1065
rect 66 993 119 1027
rect 153 993 206 1027
rect 66 955 206 993
rect 66 921 119 955
rect 153 921 206 955
rect 66 883 206 921
rect 66 849 119 883
rect 153 849 206 883
rect 66 811 206 849
rect 66 777 119 811
rect 153 777 206 811
rect 66 739 206 777
rect 66 705 119 739
rect 153 705 206 739
rect 66 667 206 705
rect 66 633 119 667
rect 153 633 206 667
rect 66 595 206 633
rect 66 561 119 595
rect 153 561 206 595
rect 66 523 206 561
rect 66 489 119 523
rect 153 489 206 523
rect 66 451 206 489
rect 66 417 119 451
rect 153 417 206 451
rect 66 379 206 417
rect 66 345 119 379
rect 153 345 206 379
rect 358 2003 1233 2066
rect 358 1969 454 2003
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 1969 1233 2003
rect 358 1924 1233 1969
rect 358 1803 498 1924
rect 358 1769 395 1803
rect 429 1769 498 1803
rect 662 1847 927 1867
rect 662 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 927 1847
rect 662 1785 927 1813
rect 1093 1803 1233 1924
rect 358 1731 498 1769
rect 1093 1769 1146 1803
rect 1180 1769 1233 1803
rect 358 1697 395 1731
rect 429 1697 498 1731
rect 358 1659 498 1697
rect 358 1625 395 1659
rect 429 1625 498 1659
rect 358 1587 498 1625
rect 358 1553 395 1587
rect 429 1553 498 1587
rect 358 1515 498 1553
rect 358 1481 395 1515
rect 429 1481 498 1515
rect 358 1443 498 1481
rect 358 1409 395 1443
rect 429 1409 498 1443
rect 358 1371 498 1409
rect 358 1337 395 1371
rect 429 1337 498 1371
rect 358 1299 498 1337
rect 358 1265 395 1299
rect 429 1265 498 1299
rect 358 1227 498 1265
rect 358 1193 395 1227
rect 429 1193 498 1227
rect 358 1155 498 1193
rect 358 1121 395 1155
rect 429 1121 498 1155
rect 358 1083 498 1121
rect 358 1049 395 1083
rect 429 1049 498 1083
rect 358 1011 498 1049
rect 358 977 395 1011
rect 429 977 498 1011
rect 358 939 498 977
rect 358 905 395 939
rect 429 905 498 939
rect 358 867 498 905
rect 358 833 395 867
rect 429 833 498 867
rect 358 795 498 833
rect 358 761 395 795
rect 429 761 498 795
rect 358 723 498 761
rect 358 689 395 723
rect 429 689 498 723
rect 358 651 498 689
rect 593 1583 701 1751
rect 593 1549 621 1583
rect 655 1549 701 1583
rect 593 1511 701 1549
rect 593 1477 621 1511
rect 655 1477 701 1511
rect 593 1439 701 1477
rect 593 1405 621 1439
rect 655 1405 701 1439
rect 593 1367 701 1405
rect 593 1333 621 1367
rect 655 1333 701 1367
rect 593 1295 701 1333
rect 593 1261 621 1295
rect 655 1261 701 1295
rect 593 1223 701 1261
rect 593 1189 621 1223
rect 655 1189 701 1223
rect 593 1151 701 1189
rect 593 1117 621 1151
rect 655 1117 701 1151
rect 593 1079 701 1117
rect 593 1045 621 1079
rect 655 1045 701 1079
rect 593 1007 701 1045
rect 593 973 621 1007
rect 655 973 701 1007
rect 593 935 701 973
rect 593 901 621 935
rect 655 901 701 935
rect 593 863 701 901
rect 593 829 621 863
rect 655 829 701 863
rect 593 791 701 829
rect 593 757 621 791
rect 655 757 701 791
rect 593 672 701 757
rect 888 1583 996 1751
rect 888 1549 915 1583
rect 949 1549 996 1583
rect 888 1511 996 1549
rect 888 1477 915 1511
rect 949 1477 996 1511
rect 888 1439 996 1477
rect 888 1405 915 1439
rect 949 1405 996 1439
rect 888 1367 996 1405
rect 888 1333 915 1367
rect 949 1333 996 1367
rect 888 1295 996 1333
rect 888 1261 915 1295
rect 949 1261 996 1295
rect 888 1223 996 1261
rect 888 1189 915 1223
rect 949 1189 996 1223
rect 888 1151 996 1189
rect 888 1117 915 1151
rect 949 1117 996 1151
rect 888 1079 996 1117
rect 888 1045 915 1079
rect 949 1045 996 1079
rect 888 1007 996 1045
rect 888 973 915 1007
rect 949 973 996 1007
rect 888 935 996 973
rect 888 901 915 935
rect 949 901 996 935
rect 888 863 996 901
rect 888 829 915 863
rect 949 829 996 863
rect 888 791 996 829
rect 888 757 915 791
rect 949 757 996 791
rect 888 672 996 757
rect 1093 1731 1233 1769
rect 1093 1697 1146 1731
rect 1180 1697 1233 1731
rect 1093 1659 1233 1697
rect 1093 1625 1146 1659
rect 1180 1625 1233 1659
rect 1093 1587 1233 1625
rect 1093 1553 1146 1587
rect 1180 1553 1233 1587
rect 1093 1515 1233 1553
rect 1093 1481 1146 1515
rect 1180 1481 1233 1515
rect 1093 1443 1233 1481
rect 1093 1409 1146 1443
rect 1180 1409 1233 1443
rect 1093 1371 1233 1409
rect 1093 1337 1146 1371
rect 1180 1337 1233 1371
rect 1093 1299 1233 1337
rect 1093 1265 1146 1299
rect 1180 1265 1233 1299
rect 1093 1227 1233 1265
rect 1093 1193 1146 1227
rect 1180 1193 1233 1227
rect 1093 1155 1233 1193
rect 1093 1121 1146 1155
rect 1180 1121 1233 1155
rect 1093 1083 1233 1121
rect 1093 1049 1146 1083
rect 1180 1049 1233 1083
rect 1093 1011 1233 1049
rect 1093 977 1146 1011
rect 1180 977 1233 1011
rect 1093 939 1233 977
rect 1093 905 1146 939
rect 1180 905 1233 939
rect 1093 867 1233 905
rect 1093 833 1146 867
rect 1180 833 1233 867
rect 1093 795 1233 833
rect 1093 761 1146 795
rect 1180 761 1233 795
rect 1093 723 1233 761
rect 1093 689 1146 723
rect 1180 689 1233 723
rect 358 617 395 651
rect 429 617 498 651
rect 358 579 498 617
rect 358 545 395 579
rect 429 545 498 579
rect 358 507 498 545
rect 358 473 395 507
rect 429 498 498 507
rect 1093 651 1233 689
rect 1093 617 1146 651
rect 1180 617 1233 651
rect 1093 579 1233 617
rect 1093 545 1146 579
rect 1180 545 1233 579
rect 1093 507 1233 545
rect 1093 498 1146 507
rect 429 473 1146 498
rect 1180 473 1233 507
rect 358 435 1233 473
rect 358 401 395 435
rect 429 401 1146 435
rect 1180 401 1233 435
rect 358 358 1233 401
rect 1385 2035 1525 2218
rect 1385 2001 1438 2035
rect 1472 2001 1525 2035
rect 1385 1963 1525 2001
rect 1385 1929 1438 1963
rect 1472 1929 1525 1963
rect 1385 1891 1525 1929
rect 1385 1857 1438 1891
rect 1472 1857 1525 1891
rect 1385 1819 1525 1857
rect 1385 1785 1438 1819
rect 1472 1785 1525 1819
rect 1385 1747 1525 1785
rect 1385 1713 1438 1747
rect 1472 1713 1525 1747
rect 1385 1675 1525 1713
rect 1385 1641 1438 1675
rect 1472 1641 1525 1675
rect 1385 1603 1525 1641
rect 1385 1569 1438 1603
rect 1472 1569 1525 1603
rect 1385 1531 1525 1569
rect 1385 1497 1438 1531
rect 1472 1497 1525 1531
rect 1385 1459 1525 1497
rect 1385 1425 1438 1459
rect 1472 1425 1525 1459
rect 1385 1387 1525 1425
rect 1385 1353 1438 1387
rect 1472 1353 1525 1387
rect 1385 1315 1525 1353
rect 1385 1281 1438 1315
rect 1472 1281 1525 1315
rect 1385 1243 1525 1281
rect 1385 1209 1438 1243
rect 1472 1209 1525 1243
rect 1385 1171 1525 1209
rect 1385 1137 1438 1171
rect 1472 1137 1525 1171
rect 1385 1099 1525 1137
rect 1385 1065 1438 1099
rect 1472 1065 1525 1099
rect 1385 1027 1525 1065
rect 1385 993 1438 1027
rect 1472 993 1525 1027
rect 1385 955 1525 993
rect 1385 921 1438 955
rect 1472 921 1525 955
rect 1385 883 1525 921
rect 1385 849 1438 883
rect 1472 849 1525 883
rect 1385 811 1525 849
rect 1385 777 1438 811
rect 1472 777 1525 811
rect 1385 739 1525 777
rect 1385 705 1438 739
rect 1472 705 1525 739
rect 1385 667 1525 705
rect 1385 633 1438 667
rect 1472 633 1525 667
rect 1385 595 1525 633
rect 1385 561 1438 595
rect 1472 561 1525 595
rect 1385 523 1525 561
rect 1385 489 1438 523
rect 1472 489 1525 523
rect 1385 451 1525 489
rect 1385 417 1438 451
rect 1472 417 1525 451
rect 1385 379 1525 417
rect 66 307 206 345
rect 66 273 119 307
rect 153 273 206 307
rect 66 206 206 273
rect 1385 345 1438 379
rect 1472 345 1525 379
rect 1385 307 1525 345
rect 1385 273 1438 307
rect 1472 273 1525 307
rect 1385 206 1525 273
rect 66 142 1525 206
rect 66 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1525 142
rect 66 66 1525 108
<< viali >>
rect 307 2271 341 2305
rect 379 2271 413 2305
rect 451 2271 485 2305
rect 523 2271 557 2305
rect 595 2271 629 2305
rect 959 2271 993 2305
rect 1031 2271 1065 2305
rect 1103 2271 1137 2305
rect 1175 2271 1209 2305
rect 1247 2271 1281 2305
rect 119 2001 153 2035
rect 119 1929 153 1963
rect 119 1857 153 1891
rect 119 1785 153 1819
rect 119 1713 153 1747
rect 119 1641 153 1675
rect 119 1569 153 1603
rect 119 1497 153 1531
rect 119 1425 153 1459
rect 119 1353 153 1387
rect 119 1281 153 1315
rect 119 1209 153 1243
rect 119 1137 153 1171
rect 119 1065 153 1099
rect 119 993 153 1027
rect 119 921 153 955
rect 119 849 153 883
rect 119 777 153 811
rect 119 705 153 739
rect 119 633 153 667
rect 119 561 153 595
rect 119 489 153 523
rect 119 417 153 451
rect 119 345 153 379
rect 454 1969 488 2003
rect 526 1969 560 2003
rect 598 1969 632 2003
rect 928 1969 962 2003
rect 1000 1969 1034 2003
rect 1072 1969 1106 2003
rect 395 1769 429 1803
rect 725 1813 759 1847
rect 797 1813 831 1847
rect 1146 1769 1180 1803
rect 395 1697 429 1731
rect 395 1625 429 1659
rect 395 1553 429 1587
rect 395 1481 429 1515
rect 395 1409 429 1443
rect 395 1337 429 1371
rect 395 1265 429 1299
rect 395 1193 429 1227
rect 395 1121 429 1155
rect 395 1049 429 1083
rect 395 977 429 1011
rect 395 905 429 939
rect 395 833 429 867
rect 395 761 429 795
rect 395 689 429 723
rect 621 1549 655 1583
rect 621 1477 655 1511
rect 621 1405 655 1439
rect 621 1333 655 1367
rect 621 1261 655 1295
rect 621 1189 655 1223
rect 621 1117 655 1151
rect 621 1045 655 1079
rect 621 973 655 1007
rect 621 901 655 935
rect 621 829 655 863
rect 621 757 655 791
rect 915 1549 949 1583
rect 915 1477 949 1511
rect 915 1405 949 1439
rect 915 1333 949 1367
rect 915 1261 949 1295
rect 915 1189 949 1223
rect 915 1117 949 1151
rect 915 1045 949 1079
rect 915 973 949 1007
rect 915 901 949 935
rect 915 829 949 863
rect 915 757 949 791
rect 1146 1697 1180 1731
rect 1146 1625 1180 1659
rect 1146 1553 1180 1587
rect 1146 1481 1180 1515
rect 1146 1409 1180 1443
rect 1146 1337 1180 1371
rect 1146 1265 1180 1299
rect 1146 1193 1180 1227
rect 1146 1121 1180 1155
rect 1146 1049 1180 1083
rect 1146 977 1180 1011
rect 1146 905 1180 939
rect 1146 833 1180 867
rect 1146 761 1180 795
rect 1146 689 1180 723
rect 395 617 429 651
rect 395 545 429 579
rect 395 473 429 507
rect 1146 617 1180 651
rect 1146 545 1180 579
rect 1146 473 1180 507
rect 395 401 429 435
rect 1146 401 1180 435
rect 1438 2001 1472 2035
rect 1438 1929 1472 1963
rect 1438 1857 1472 1891
rect 1438 1785 1472 1819
rect 1438 1713 1472 1747
rect 1438 1641 1472 1675
rect 1438 1569 1472 1603
rect 1438 1497 1472 1531
rect 1438 1425 1472 1459
rect 1438 1353 1472 1387
rect 1438 1281 1472 1315
rect 1438 1209 1472 1243
rect 1438 1137 1472 1171
rect 1438 1065 1472 1099
rect 1438 993 1472 1027
rect 1438 921 1472 955
rect 1438 849 1472 883
rect 1438 777 1472 811
rect 1438 705 1472 739
rect 1438 633 1472 667
rect 1438 561 1472 595
rect 1438 489 1472 523
rect 1438 417 1472 451
rect 119 273 153 307
rect 1438 345 1472 379
rect 1438 273 1472 307
rect 1118 108 1152 142
rect 1190 108 1224 142
rect 1262 108 1296 142
<< obsli1 >>
rect -32 39532 16032 42134
rect -32 2358 23971 39532
rect -32 2239 66 2358
rect 0 1392 66 2239
rect 206 2066 1385 2218
rect -17 792 66 1392
rect 0 66 66 792
rect 206 358 358 2066
rect 498 1867 1093 1924
rect 498 1785 662 1867
rect 927 1785 1093 1867
rect 498 1751 1093 1785
rect 498 672 593 1751
rect 701 672 888 1751
rect 996 672 1093 1751
rect 498 498 1093 672
rect 1233 358 1385 2066
rect 206 206 1385 358
rect 1525 66 23971 2358
rect 0 0 23971 66
rect 122 -194 2260 0
rect 141 -300 175 -194
rect 297 -278 332 -194
rect 518 -269 552 -194
rect 694 -239 728 -194
rect 870 -269 904 -194
rect 1046 -239 1080 -194
rect 1222 -269 1256 -194
rect 1346 -269 1380 -194
rect 1522 -241 1556 -194
rect 1698 -269 1732 -194
rect 1874 -241 1908 -194
rect 2050 -269 2084 -194
rect 2226 -241 2260 -194
rect 2350 -269 2384 0
rect 2407 -23 2609 0
rect 2702 -23 2736 0
rect 2878 -23 2912 0
rect 3054 -23 3088 0
rect 3230 -23 3264 0
rect 3406 -23 3440 0
rect 3582 -23 3616 0
rect 3758 -23 3792 0
rect 3934 -23 3968 0
rect 4110 -23 4144 0
rect 4286 -23 4320 0
rect 4462 -23 4496 0
rect 4638 -23 4672 0
rect 4814 -23 4848 0
rect 4990 -23 5024 0
rect 5166 -23 5200 0
rect 5342 -23 5376 0
rect 5518 -23 5552 0
rect 5694 -23 5728 0
rect 5870 -23 5904 0
rect 5993 -10 6099 0
rect 5994 -23 6028 -10
rect 6170 -23 6204 0
rect 6294 -23 6328 0
rect 6470 -23 6504 0
rect 6646 -23 6680 0
rect 6822 -23 6857 0
rect 7598 -23 7632 0
rect 7774 -23 7808 0
rect 7950 -23 7984 0
rect 8126 -23 8160 0
rect 8250 -23 8284 0
rect 8426 -23 8460 0
rect 8602 -23 8636 0
rect 9058 -23 9092 0
rect 9234 -23 9268 0
rect 9410 -23 9444 0
rect 9522 -23 11631 0
rect 11694 -23 11728 0
rect 11804 -23 12014 0
rect 12156 -23 12190 0
rect 13658 -19 14136 0
rect 14463 -19 14867 0
rect 13946 -23 14136 -19
rect 23346 -23 23536 0
rect 2407 -213 23536 -23
rect 2526 -241 2560 -213
rect 2702 -269 2736 -213
rect 2878 -241 2912 -213
rect 3054 -269 3088 -213
rect 3230 -241 3264 -213
rect 3406 -269 3440 -213
rect 3582 -241 3616 -213
rect 3758 -269 3792 -213
rect 3934 -241 3968 -213
rect 4110 -269 4144 -213
rect 4286 -241 4320 -213
rect 4462 -269 4496 -213
rect 4638 -241 4672 -213
rect 4814 -269 4848 -213
rect 4990 -241 5024 -213
rect 5166 -269 5200 -213
rect 5342 -241 5376 -213
rect 5518 -269 5552 -213
rect 5694 -241 5728 -213
rect 5870 -269 5904 -213
rect 5994 -241 6028 -213
rect 6170 -269 6204 -213
rect 6294 -269 6328 -213
rect 6470 -241 6504 -213
rect 6646 -269 6680 -213
rect 6822 -241 6856 -213
rect 7598 -269 7632 -213
rect 7774 -241 7808 -213
rect 7950 -269 7984 -213
rect 8126 -241 8160 -213
rect 8250 -269 8284 -213
rect 8426 -239 8460 -213
rect 8602 -269 8636 -213
rect 9058 -241 9092 -213
rect 9234 -269 9268 -213
rect 9410 -239 9444 -213
rect 9586 -269 9620 -213
rect 9699 -269 9733 -213
rect 9875 -241 9909 -213
rect 10051 -269 10085 -213
rect 10227 -241 10261 -213
rect 10403 -269 10437 -213
rect 10528 -241 10562 -213
rect 10704 -269 10738 -213
rect 10880 -241 10914 -213
rect 11056 -269 11090 -213
rect 11166 -269 11200 -213
rect 11342 -241 11376 -213
rect 11518 -269 11552 -213
rect 11694 -241 11728 -213
rect 11804 -269 11838 -213
rect 11980 -241 12014 -213
rect 12156 -269 12190 -213
rect 297 -300 331 -278
rect 510 -341 12198 -307
rect 12875 -357 13215 -213
rect 13359 -361 13393 -213
rect 13465 -361 13499 -213
rect 13571 -361 13605 -213
<< metal1 >>
tri 66 2216 208 2358 se
rect 208 2305 669 2358
rect 208 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 669 2305
rect 208 2218 669 2271
rect 208 2216 286 2218
tri 286 2216 288 2218 nw
rect 66 2035 206 2216
tri 206 2136 286 2216 nw
rect 66 2001 119 2035
rect 153 2001 206 2035
rect 66 1963 206 2001
rect 66 1929 119 1963
rect 153 1929 206 1963
rect 66 1891 206 1929
rect 66 1857 119 1891
rect 153 1857 206 1891
rect 66 1819 206 1857
rect 66 1785 119 1819
rect 153 1785 206 1819
rect 66 1747 206 1785
rect 66 1713 119 1747
rect 153 1713 206 1747
rect 66 1675 206 1713
rect 66 1641 119 1675
rect 153 1641 206 1675
rect 66 1603 206 1641
rect 66 1569 119 1603
rect 153 1569 206 1603
rect 66 1531 206 1569
rect 66 1497 119 1531
rect 153 1497 206 1531
rect 66 1459 206 1497
rect 66 1425 119 1459
rect 153 1425 206 1459
rect 66 1387 206 1425
rect 66 1353 119 1387
rect 153 1353 206 1387
rect 66 1315 206 1353
rect 66 1281 119 1315
rect 153 1281 206 1315
rect 66 1243 206 1281
rect 66 1209 119 1243
rect 153 1209 206 1243
rect 66 1171 206 1209
rect 66 1137 119 1171
rect 153 1137 206 1171
rect 66 1099 206 1137
rect 66 1065 119 1099
rect 153 1065 206 1099
rect 66 1027 206 1065
rect 66 993 119 1027
rect 153 993 206 1027
rect 66 955 206 993
rect 66 921 119 955
rect 153 921 206 955
rect 66 883 206 921
rect 66 849 119 883
rect 153 849 206 883
rect 66 811 206 849
rect 66 777 119 811
rect 153 777 206 811
rect 66 739 206 777
rect 66 705 119 739
rect 153 705 206 739
rect 66 667 206 705
rect 66 633 119 667
rect 153 633 206 667
rect 66 595 206 633
rect 66 561 119 595
rect 153 561 206 595
rect 66 523 206 561
rect 66 489 119 523
rect 153 489 206 523
rect 66 451 206 489
rect 66 417 119 451
rect 153 417 206 451
rect 66 379 206 417
rect 66 345 119 379
rect 153 345 206 379
rect 66 307 206 345
rect 66 273 119 307
rect 153 273 206 307
rect 66 69 206 273
tri 358 2000 424 2066 se
rect 424 2003 669 2066
rect 424 2000 454 2003
rect 358 1969 454 2000
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 669 2003
rect 358 1901 669 1969
rect 358 1803 536 1901
tri 536 1826 611 1901 nw
rect 703 1847 852 2359
rect 886 2305 1383 2358
rect 886 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1383 2305
rect 886 2218 1383 2271
tri 1289 2216 1291 2218 ne
rect 1291 2216 1383 2218
tri 1383 2216 1525 2358 sw
tri 1291 2136 1371 2216 ne
rect 1371 2136 1525 2216
tri 1371 2124 1383 2136 ne
rect 1383 2124 1525 2136
tri 1383 2122 1385 2124 ne
rect 886 2003 1167 2066
rect 886 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 2000 1167 2003
tri 1167 2000 1233 2066 sw
rect 1106 1969 1233 2000
rect 886 1901 1233 1969
rect 358 1769 395 1803
rect 429 1769 536 1803
rect 703 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 852 1847
tri 1012 1826 1087 1901 ne
rect 1087 1826 1233 1901
tri 1087 1820 1093 1826 ne
rect 703 1791 852 1813
rect 1093 1803 1233 1826
rect 358 1731 536 1769
rect 1093 1769 1146 1803
rect 1180 1769 1233 1803
rect 358 1697 395 1731
rect 429 1697 536 1731
rect 358 1659 536 1697
rect 358 1625 395 1659
rect 429 1625 536 1659
rect 358 1587 536 1625
rect 358 1553 395 1587
rect 429 1553 536 1587
rect 358 1515 536 1553
rect 358 1481 395 1515
rect 429 1481 536 1515
rect 358 1443 536 1481
rect 358 1409 395 1443
rect 429 1409 536 1443
rect 358 1371 536 1409
rect 358 1337 395 1371
rect 429 1337 536 1371
rect 358 1299 536 1337
rect 358 1265 395 1299
rect 429 1265 536 1299
rect 358 1227 536 1265
rect 358 1193 395 1227
rect 429 1193 536 1227
rect 358 1155 536 1193
rect 358 1121 395 1155
rect 429 1121 536 1155
rect 358 1083 536 1121
rect 358 1049 395 1083
rect 429 1049 536 1083
rect 358 1011 536 1049
rect 358 977 395 1011
rect 429 977 536 1011
rect 358 939 536 977
rect 358 905 395 939
rect 429 905 536 939
rect 358 867 536 905
rect 358 833 395 867
rect 429 833 536 867
rect 358 795 536 833
rect 358 761 395 795
rect 429 761 536 795
rect 358 723 536 761
rect 358 689 395 723
rect 429 689 536 723
rect 358 651 536 689
rect 358 617 395 651
rect 429 617 536 651
rect 358 579 536 617
rect 358 545 395 579
rect 429 545 536 579
rect 358 507 536 545
rect 358 473 395 507
rect 429 473 536 507
rect 358 435 536 473
rect 358 401 395 435
rect 429 401 536 435
rect 358 69 536 401
rect 572 1583 772 1709
rect 572 1549 621 1583
rect 655 1549 772 1583
rect 572 1511 772 1549
rect 572 1477 621 1511
rect 655 1477 772 1511
rect 572 1439 772 1477
rect 572 1405 621 1439
rect 655 1405 772 1439
rect 572 1367 772 1405
rect 572 1333 621 1367
rect 655 1333 772 1367
rect 572 1295 772 1333
rect 572 1261 621 1295
rect 655 1261 772 1295
rect 572 1223 772 1261
rect 572 1189 621 1223
rect 655 1189 772 1223
rect 572 1151 772 1189
rect 572 1117 621 1151
rect 655 1117 772 1151
rect 572 1079 772 1117
rect 572 1045 621 1079
rect 655 1045 772 1079
rect 572 1007 772 1045
rect 572 973 621 1007
rect 655 973 772 1007
rect 572 935 772 973
rect 572 901 621 935
rect 655 901 772 935
rect 572 863 772 901
rect 572 829 621 863
rect 655 829 772 863
rect 572 791 772 829
rect 572 757 621 791
rect 655 757 772 791
rect 66 66 203 69
rect 358 66 533 69
rect 572 66 772 757
rect 831 1583 1031 1752
rect 831 1549 915 1583
rect 949 1549 1031 1583
rect 831 1511 1031 1549
rect 831 1477 915 1511
rect 949 1477 1031 1511
rect 831 1439 1031 1477
rect 831 1405 915 1439
rect 949 1405 1031 1439
rect 831 1367 1031 1405
rect 831 1333 915 1367
rect 949 1333 1031 1367
rect 831 1295 1031 1333
rect 831 1261 915 1295
rect 949 1261 1031 1295
rect 831 1223 1031 1261
rect 831 1189 915 1223
rect 949 1189 1031 1223
rect 831 1151 1031 1189
rect 831 1117 915 1151
rect 949 1117 1031 1151
rect 831 1079 1031 1117
rect 831 1045 915 1079
rect 949 1045 1031 1079
rect 831 1007 1031 1045
rect 831 973 915 1007
rect 949 973 1031 1007
rect 831 935 1031 973
rect 831 901 915 935
rect 949 901 1031 935
rect 831 863 1031 901
rect 831 829 915 863
rect 949 829 1031 863
rect 831 791 1031 829
rect 831 757 915 791
rect 949 757 1031 791
rect 831 66 1031 757
rect 1093 1731 1233 1769
rect 1093 1697 1146 1731
rect 1180 1697 1233 1731
rect 1093 1659 1233 1697
rect 1093 1625 1146 1659
rect 1180 1625 1233 1659
rect 1093 1587 1233 1625
rect 1093 1553 1146 1587
rect 1180 1553 1233 1587
rect 1093 1515 1233 1553
rect 1093 1481 1146 1515
rect 1180 1481 1233 1515
rect 1093 1443 1233 1481
rect 1093 1409 1146 1443
rect 1180 1409 1233 1443
rect 1093 1371 1233 1409
rect 1093 1337 1146 1371
rect 1180 1337 1233 1371
rect 1093 1299 1233 1337
rect 1093 1265 1146 1299
rect 1180 1265 1233 1299
rect 1093 1227 1233 1265
rect 1093 1193 1146 1227
rect 1180 1193 1233 1227
rect 1093 1155 1233 1193
rect 1093 1121 1146 1155
rect 1180 1121 1233 1155
rect 1093 1083 1233 1121
rect 1093 1049 1146 1083
rect 1180 1049 1233 1083
rect 1093 1011 1233 1049
rect 1093 977 1146 1011
rect 1180 977 1233 1011
rect 1093 939 1233 977
rect 1093 905 1146 939
rect 1180 905 1233 939
rect 1093 867 1233 905
rect 1093 833 1146 867
rect 1180 833 1233 867
rect 1093 795 1233 833
rect 1093 761 1146 795
rect 1180 761 1233 795
rect 1093 723 1233 761
rect 1093 689 1146 723
rect 1180 689 1233 723
rect 1093 651 1233 689
rect 1093 617 1146 651
rect 1180 617 1233 651
rect 1093 579 1233 617
rect 1093 545 1146 579
rect 1180 545 1233 579
rect 1093 507 1233 545
rect 1093 473 1146 507
rect 1180 473 1233 507
rect 1093 435 1233 473
rect 1093 401 1146 435
rect 1180 401 1233 435
rect 1093 358 1233 401
rect 1385 2035 1525 2124
rect 1385 2001 1438 2035
rect 1472 2001 1525 2035
rect 1385 1963 1525 2001
rect 1385 1929 1438 1963
rect 1472 1929 1525 1963
rect 1385 1891 1525 1929
rect 1385 1857 1438 1891
rect 1472 1857 1525 1891
rect 1385 1819 1525 1857
rect 1385 1785 1438 1819
rect 1472 1785 1525 1819
rect 1385 1747 1525 1785
rect 1385 1713 1438 1747
rect 1472 1713 1525 1747
rect 1385 1675 1525 1713
rect 1385 1641 1438 1675
rect 1472 1641 1525 1675
rect 1385 1603 1525 1641
rect 1385 1569 1438 1603
rect 1472 1569 1525 1603
rect 1385 1531 1525 1569
rect 1385 1497 1438 1531
rect 1472 1497 1525 1531
rect 1385 1459 1525 1497
rect 1385 1425 1438 1459
rect 1472 1425 1525 1459
rect 1385 1387 1525 1425
rect 1385 1353 1438 1387
rect 1472 1353 1525 1387
rect 1385 1315 1525 1353
rect 1385 1281 1438 1315
rect 1472 1281 1525 1315
rect 1385 1243 1525 1281
rect 1385 1209 1438 1243
rect 1472 1209 1525 1243
rect 1385 1171 1525 1209
rect 1385 1137 1438 1171
rect 1472 1137 1525 1171
rect 1385 1099 1525 1137
rect 1385 1065 1438 1099
rect 1472 1065 1525 1099
rect 1385 1027 1525 1065
rect 1385 993 1438 1027
rect 1472 993 1525 1027
rect 1385 955 1525 993
rect 1385 921 1438 955
rect 1472 921 1525 955
rect 1385 883 1525 921
rect 1385 849 1438 883
rect 1472 849 1525 883
rect 1385 811 1525 849
rect 1385 777 1438 811
rect 1472 777 1525 811
rect 1385 739 1525 777
rect 1385 705 1438 739
rect 1472 705 1525 739
rect 1385 667 1525 705
rect 1385 633 1438 667
rect 1472 633 1525 667
rect 1385 595 1525 633
rect 1385 561 1438 595
rect 1472 561 1525 595
rect 1385 523 1525 561
rect 1385 489 1438 523
rect 1472 489 1525 523
rect 1385 451 1525 489
rect 1385 417 1438 451
rect 1472 417 1525 451
rect 1385 379 1525 417
rect 1385 345 1438 379
rect 1472 345 1525 379
rect 1385 307 1525 345
tri 1289 206 1385 302 se
rect 1385 273 1438 307
rect 1472 273 1525 307
rect 1385 208 1525 273
rect 1385 206 1386 208
rect 1070 142 1386 206
rect 1070 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1386 142
rect 1070 69 1386 108
tri 1386 69 1525 208 nw
rect 1070 66 1383 69
tri 1383 66 1386 69 nw
<< obsm1 >>
rect -29 39538 16029 42193
rect -29 2359 23983 39538
rect -29 2358 703 2359
rect -29 824 66 2358
tri 66 2216 208 2358 nw
rect 669 2218 703 2358
tri 286 2216 288 2218 se
rect 288 2216 703 2218
tri 206 2136 286 2216 se
rect 286 2136 703 2216
rect 206 2066 703 2136
rect 0 66 66 824
rect 206 69 358 2066
tri 358 2000 424 2066 nw
rect 669 1901 703 2066
tri 536 1826 611 1901 se
rect 611 1826 703 1901
rect 852 2358 23983 2359
rect 852 2218 886 2358
rect 852 2216 1289 2218
tri 1289 2216 1291 2218 sw
tri 1383 2216 1525 2358 ne
rect 852 2136 1291 2216
tri 1291 2136 1371 2216 sw
rect 852 2124 1371 2136
tri 1371 2124 1383 2136 sw
rect 852 2122 1383 2124
tri 1383 2122 1385 2124 sw
rect 852 2066 1385 2122
rect 852 1901 886 2066
tri 1167 2000 1233 2066 ne
rect 536 1791 703 1826
rect 852 1826 1012 1901
tri 1012 1826 1087 1901 sw
rect 852 1820 1087 1826
tri 1087 1820 1093 1826 sw
rect 852 1791 1093 1820
rect 536 1752 1093 1791
rect 536 1709 831 1752
rect 536 69 572 1709
rect 203 66 358 69
rect 533 66 572 69
rect 772 66 831 1709
rect 1031 358 1093 1752
rect 1233 358 1385 2066
rect 1031 302 1385 358
rect 1031 206 1289 302
tri 1289 206 1385 302 nw
rect 1031 66 1070 206
tri 1386 69 1525 208 se
rect 1525 69 23983 2358
tri 1383 66 1386 69 se
rect 1386 66 23983 69
rect 0 0 23983 66
rect 52 -26 104 0
tri 181 -48 209 -20 se
rect 209 -40 255 0
rect 209 -48 247 -40
tri 247 -48 255 -40 nw
tri 135 -94 181 -48 se
rect 135 -293 181 -94
tri 181 -114 247 -48 nw
rect 292 -122 338 0
tri 338 -122 413 -47 sw
rect 428 -51 474 0
rect 725 -16 11313 0
tri 474 -51 508 -17 sw
rect 725 -51 1771 -16
rect 2407 -23 2686 -16
tri 2686 -23 2693 -16 sw
rect 4099 -23 11313 -16
rect 11336 -23 11382 0
rect 11807 -23 12070 0
tri 12070 -23 12093 0 sw
rect 12736 -23 12976 0
tri 13106 -21 13127 0 ne
rect 13127 -23 13155 0
tri 13359 -23 13366 -16 se
rect 13366 -23 13419 0
rect 13471 -23 13499 0
tri 13600 -23 13623 0 ne
rect 13623 -23 13643 0
tri 13643 -23 13666 0 sw
tri 13885 -23 13908 0 se
rect 13908 -23 14136 0
rect 15240 -23 17187 0
tri 23285 -23 23308 0 se
rect 23308 -23 23536 0
rect 2407 -51 23536 -23
rect 428 -97 23536 -51
rect 292 -150 413 -122
tri 413 -150 441 -122 sw
rect 725 -150 1771 -97
rect 2407 -150 23536 -97
rect 292 -213 23536 -150
rect 292 -353 17187 -213
tri 3331 -603 3581 -353 se
rect 3581 -603 17187 -353
rect 3331 -1384 17187 -603
rect 3331 -1391 17180 -1384
tri 17180 -1391 17187 -1384 nw
rect 3331 -1398 17173 -1391
tri 17173 -1398 17180 -1391 nw
rect 3331 -1405 17166 -1398
tri 17166 -1405 17173 -1398 nw
rect 3331 -1412 17159 -1405
tri 17159 -1412 17166 -1405 nw
rect 3331 -1419 17152 -1412
tri 17152 -1419 17159 -1412 nw
rect 3331 -1426 17145 -1419
tri 17145 -1426 17152 -1419 nw
rect 3331 -1433 17138 -1426
tri 17138 -1433 17145 -1426 nw
rect 3331 -1440 17131 -1433
tri 17131 -1440 17138 -1433 nw
rect 3331 -1447 17124 -1440
tri 17124 -1447 17131 -1440 nw
rect 3331 -1454 17117 -1447
tri 17117 -1454 17124 -1447 nw
rect 3331 -1461 17110 -1454
tri 17110 -1461 17117 -1454 nw
rect 3331 -1468 17103 -1461
tri 17103 -1468 17110 -1461 nw
rect 3331 -1475 17096 -1468
tri 17096 -1475 17103 -1468 nw
rect 3331 -1482 17089 -1475
tri 17089 -1482 17096 -1475 nw
rect 3331 -1489 17082 -1482
tri 17082 -1489 17089 -1482 nw
rect 3331 -1496 17075 -1489
tri 17075 -1496 17082 -1489 nw
rect 3331 -1503 17068 -1496
tri 17068 -1503 17075 -1496 nw
rect 3331 -1510 17061 -1503
tri 17061 -1510 17068 -1503 nw
rect 3331 -1517 17054 -1510
tri 17054 -1517 17061 -1510 nw
rect 3331 -1524 17047 -1517
tri 17047 -1524 17054 -1517 nw
rect 3331 -1531 17040 -1524
tri 17040 -1531 17047 -1524 nw
rect 3331 -1538 17033 -1531
tri 17033 -1538 17040 -1531 nw
rect 3331 -1545 17026 -1538
tri 17026 -1545 17033 -1538 nw
rect 3331 -1552 17019 -1545
tri 17019 -1552 17026 -1545 nw
rect 3331 -1559 17012 -1552
tri 17012 -1559 17019 -1552 nw
rect 3331 -1566 17005 -1559
tri 17005 -1566 17012 -1559 nw
rect 3331 -1573 16998 -1566
tri 16998 -1573 17005 -1566 nw
rect 3331 -1580 16991 -1573
tri 16991 -1580 16998 -1573 nw
rect 3331 -1587 16984 -1580
tri 16984 -1587 16991 -1580 nw
rect 3331 -1594 16977 -1587
tri 16977 -1594 16984 -1587 nw
rect 3331 -1601 16970 -1594
tri 16970 -1601 16977 -1594 nw
rect 3331 -1608 16963 -1601
tri 16963 -1608 16970 -1601 nw
rect 3331 -1615 16956 -1608
tri 16956 -1615 16963 -1608 nw
rect 3331 -1622 16949 -1615
tri 16949 -1622 16956 -1615 nw
rect 3331 -1629 16942 -1622
tri 16942 -1629 16949 -1622 nw
rect 3331 -1636 16935 -1629
tri 16935 -1636 16942 -1629 nw
rect 3331 -1643 16928 -1636
tri 16928 -1643 16935 -1636 nw
rect 3331 -1650 16921 -1643
tri 16921 -1650 16928 -1643 nw
rect 3331 -1657 16914 -1650
tri 16914 -1657 16921 -1650 nw
rect 3331 -1664 16907 -1657
tri 16907 -1664 16914 -1657 nw
rect 3331 -1671 16900 -1664
tri 16900 -1671 16907 -1664 nw
rect 3331 -1678 16893 -1671
tri 16893 -1678 16900 -1671 nw
rect 3331 -1685 16886 -1678
tri 16886 -1685 16893 -1678 nw
rect 3331 -1692 16879 -1685
tri 16879 -1692 16886 -1685 nw
rect 3331 -1699 16872 -1692
tri 16872 -1699 16879 -1692 nw
rect 3331 -1706 16865 -1699
tri 16865 -1706 16872 -1699 nw
rect 3331 -1707 16858 -1706
tri 3331 -2107 3731 -1707 ne
rect 3731 -1713 16858 -1707
tri 16858 -1713 16865 -1706 nw
rect 3731 -1720 16851 -1713
tri 16851 -1720 16858 -1713 nw
rect 3731 -1727 16844 -1720
tri 16844 -1727 16851 -1720 nw
rect 3731 -1734 16837 -1727
tri 16837 -1734 16844 -1727 nw
rect 3731 -1741 16830 -1734
tri 16830 -1741 16837 -1734 nw
rect 3731 -1748 16823 -1741
tri 16823 -1748 16830 -1741 nw
rect 3731 -1755 16816 -1748
tri 16816 -1755 16823 -1748 nw
rect 3731 -1762 16809 -1755
tri 16809 -1762 16816 -1755 nw
rect 3731 -1769 16802 -1762
tri 16802 -1769 16809 -1762 nw
rect 3731 -1776 16795 -1769
tri 16795 -1776 16802 -1769 nw
rect 3731 -1778 16793 -1776
tri 16793 -1778 16795 -1776 nw
rect 3731 -1785 16786 -1778
tri 16786 -1785 16793 -1778 nw
rect 3731 -1792 16779 -1785
tri 16779 -1792 16786 -1785 nw
rect 3731 -1799 16772 -1792
tri 16772 -1799 16779 -1792 nw
rect 3731 -1806 16765 -1799
tri 16765 -1806 16772 -1799 nw
rect 3731 -1813 16758 -1806
tri 16758 -1813 16765 -1806 nw
rect 3731 -1820 16751 -1813
tri 16751 -1820 16758 -1813 nw
rect 3731 -1827 16744 -1820
tri 16744 -1827 16751 -1820 nw
rect 3731 -1834 16737 -1827
tri 16737 -1834 16744 -1827 nw
rect 3731 -1841 16730 -1834
tri 16730 -1841 16737 -1834 nw
rect 3731 -1848 16723 -1841
tri 16723 -1848 16730 -1841 nw
rect 3731 -1855 16716 -1848
tri 16716 -1855 16723 -1848 nw
rect 3731 -1862 16709 -1855
tri 16709 -1862 16716 -1855 nw
rect 3731 -1869 16702 -1862
tri 16702 -1869 16709 -1862 nw
rect 3731 -1876 16695 -1869
tri 16695 -1876 16702 -1869 nw
rect 3731 -1883 16688 -1876
tri 16688 -1883 16695 -1876 nw
rect 3731 -1890 16681 -1883
tri 16681 -1890 16688 -1883 nw
rect 3731 -1897 16674 -1890
tri 16674 -1897 16681 -1890 nw
rect 3731 -1904 16667 -1897
tri 16667 -1904 16674 -1897 nw
rect 3731 -1911 16660 -1904
tri 16660 -1911 16667 -1904 nw
rect 3731 -1918 16653 -1911
tri 16653 -1918 16660 -1911 nw
rect 3731 -1925 16646 -1918
tri 16646 -1925 16653 -1918 nw
rect 3731 -1932 16639 -1925
tri 16639 -1932 16646 -1925 nw
rect 3731 -1939 16632 -1932
tri 16632 -1939 16639 -1932 nw
rect 3731 -1946 16625 -1939
tri 16625 -1946 16632 -1939 nw
rect 3731 -1953 16618 -1946
tri 16618 -1953 16625 -1946 nw
rect 3731 -1960 16611 -1953
tri 16611 -1960 16618 -1953 nw
rect 3731 -1967 16604 -1960
tri 16604 -1967 16611 -1960 nw
rect 3731 -1974 16597 -1967
tri 16597 -1974 16604 -1967 nw
rect 3731 -1981 16590 -1974
tri 16590 -1981 16597 -1974 nw
rect 3731 -1988 16583 -1981
tri 16583 -1988 16590 -1981 nw
rect 3731 -1995 16576 -1988
tri 16576 -1995 16583 -1988 nw
rect 3731 -2002 16569 -1995
tri 16569 -2002 16576 -1995 nw
rect 3731 -2009 16562 -2002
tri 16562 -2009 16569 -2002 nw
rect 3731 -2016 16555 -2009
tri 16555 -2016 16562 -2009 nw
rect 3731 -2023 16548 -2016
tri 16548 -2023 16555 -2016 nw
rect 3731 -2030 16541 -2023
tri 16541 -2030 16548 -2023 nw
rect 3731 -2037 16534 -2030
tri 16534 -2037 16541 -2030 nw
rect 3731 -2044 16527 -2037
tri 16527 -2044 16534 -2037 nw
rect 3731 -2051 16520 -2044
tri 16520 -2051 16527 -2044 nw
rect 3731 -2058 16513 -2051
tri 16513 -2058 16520 -2051 nw
rect 3731 -2065 16506 -2058
tri 16506 -2065 16513 -2058 nw
rect 3731 -2072 16499 -2065
tri 16499 -2072 16506 -2065 nw
rect 3731 -2079 16492 -2072
tri 16492 -2079 16499 -2072 nw
rect 3731 -2086 16485 -2079
tri 16485 -2086 16492 -2079 nw
rect 3731 -2093 16478 -2086
tri 16478 -2093 16485 -2086 nw
rect 3731 -2100 16471 -2093
tri 16471 -2100 16478 -2093 nw
rect 3731 -2107 16464 -2100
tri 16464 -2107 16471 -2100 nw
rect 4185 -2114 16457 -2107
tri 16457 -2114 16464 -2107 nw
rect 4185 -2121 16450 -2114
tri 16450 -2121 16457 -2114 nw
rect 4185 -2128 16443 -2121
tri 16443 -2128 16450 -2121 nw
rect 4185 -2135 16436 -2128
tri 16436 -2135 16443 -2128 nw
rect 4185 -2142 16429 -2135
tri 16429 -2142 16436 -2135 nw
rect 4185 -2149 16422 -2142
tri 16422 -2149 16429 -2142 nw
rect 4185 -2156 16415 -2149
tri 16415 -2156 16422 -2149 nw
rect 4185 -2163 16408 -2156
tri 16408 -2163 16415 -2156 nw
rect 4185 -2170 16401 -2163
tri 16401 -2170 16408 -2163 nw
rect 4185 -2177 16394 -2170
tri 16394 -2177 16401 -2170 nw
rect 4185 -2184 16387 -2177
tri 16387 -2184 16394 -2177 nw
<< metal2 >>
rect 10887 725 14858 781
rect 100 4 4099 290
rect 99 0 4155 4
rect 99 -7 4185 0
rect 6888 -7 8888 58
rect 10707 -7 10819 0
rect 10943 -7 14940 725
rect 99 -407 4879 -7
rect 5320 -23 5372 -7
rect 5698 -407 5750 -7
rect 6150 -407 6202 -7
rect 6363 -407 6415 -7
rect 7092 -407 7144 -97
rect 7678 -407 7730 -7
rect 9049 -407 9101 -7
rect 9499 -407 14858 -7
rect 15256 -407 15384 0
rect 15522 -407 15574 -170
rect 15741 -407 15781 -164
rect 15943 -407 15983 0
rect 19478 -407 24258 4725
<< obsm2 >>
rect 42 39593 15983 42193
rect 42 39586 17187 39593
rect 0 38608 17187 39586
rect 0 8833 24258 38608
rect -2195 7903 24258 8833
rect 0 4781 24258 7903
rect 0 781 19422 4781
rect 0 725 10887 781
rect 14858 725 19422 781
rect 0 290 10943 725
rect 0 4 100 290
rect 4099 58 10943 290
rect 4099 4 6888 58
rect 0 0 99 4
rect 4155 0 6888 4
rect 52 -213 99 0
rect 4185 -7 6888 0
rect 8888 0 10943 58
rect 8888 -7 10707 0
rect 10819 -7 10943 0
rect 14940 0 19422 725
tri 52 -259 98 -213 ne
rect 98 -407 99 -213
rect 4879 -23 5253 -7
rect 4879 -352 5579 -23
rect 5179 -407 5579 -352
tri 5798 -56 5817 -37 se
rect 5817 -56 5877 -7
tri 5877 -56 5926 -7 sw
rect 5798 -108 5926 -56
rect 5954 -107 6082 -7
tri 6455 -33 6471 -17 se
rect 6471 -33 6523 -7
rect 6455 -55 6523 -33
tri 6523 -55 6561 -17 sw
rect 6455 -107 6583 -55
rect 6680 -353 6934 -7
tri 7072 -27 7092 -7 ne
rect 7092 -45 7146 -7
tri 7146 -45 7184 -7 sw
tri 7496 -45 7534 -7 se
rect 7534 -45 7624 -7
rect 7092 -97 7220 -45
rect 7496 -97 7624 -45
tri 7144 -137 7184 -97 nw
tri 7885 -70 7948 -7 se
rect 7948 -70 8006 -7
tri 8350 -62 8405 -7 se
rect 8405 -62 8424 -7
tri 8424 -62 8479 -7 nw
rect 7878 -122 8006 -70
tri 8276 -136 8350 -62 se
tri 8350 -136 8424 -62 nw
tri 7730 -180 7769 -141 sw
tri 8232 -180 8276 -136 se
rect 8276 -180 8306 -136
tri 8306 -180 8350 -136 nw
rect 7730 -232 8254 -180
tri 8254 -232 8306 -180 nw
tri 7730 -271 7769 -232 nw
tri 9441 -70 9475 -36 se
rect 9475 -70 9499 -7
rect 9354 -122 9499 -70
rect 14858 -23 14940 -7
rect 14858 -407 14979 -23
rect 15025 -295 15179 -239
tri 15384 -82 15466 0 nw
rect 15478 -170 15642 -114
tri 15741 -164 15742 -163 se
rect 15742 -164 15782 0
tri 15482 -210 15522 -170 ne
tri 15574 -232 15636 -170 nw
rect 15781 -181 15782 -164
tri 15781 -182 15782 -181 nw
rect 15822 -295 15874 0
rect 98 -502 4204 -407
tri 4204 -502 4299 -407 sw
tri 10619 -502 10714 -407 se
rect 10714 -502 14940 -407
rect 98 -512 14940 -502
tri 98 -1512 1098 -512 ne
rect 1098 -1512 13940 -512
tri 13940 -1512 14940 -512 nw
<< metal3 >>
rect 99 1453 4900 4843
rect 5200 2078 7376 4037
rect 20 862 4959 1453
rect 20 0 98 862
rect 0 -407 98 0
rect 99 0 4959 862
rect 5179 0 7379 2078
rect 7676 2069 9851 4573
rect 7596 339 9851 2069
rect 10078 1453 14940 4843
rect 7578 0 9851 339
rect 10071 138 14940 1453
rect 15716 138 15782 218
rect 15848 138 15914 218
rect 10071 0 16779 138
rect 99 -7 16779 0
rect 99 -407 9778 -7
rect 9851 -407 16779 -7
rect 16978 -407 19178 1859
rect 19478 -407 33800 2730
rect 100 -1896 4900 -407
rect 5200 -502 9851 -458
rect 5190 -1506 9852 -502
rect 5200 -1898 9851 -1506
rect 10151 -1902 14940 -407
<< obsm3 >>
rect 62 39593 15914 42193
rect -2195 7903 -179 8833
rect 0 4843 33800 39593
rect 0 1453 99 4843
rect 4900 4573 10078 4843
rect 4900 4037 7676 4573
rect 4900 2078 5200 4037
rect 7376 2078 7676 4037
rect 4900 1453 5179 2078
rect 0 0 20 1453
rect 98 -407 99 862
rect 4959 0 5179 1453
rect 7379 2069 7676 2078
rect 7379 339 7596 2069
rect 9851 1453 10078 4573
rect 14940 2810 33800 4843
rect 14940 1939 19398 2810
rect 7379 0 7578 339
rect 9851 0 10071 1453
rect 14940 218 16898 1939
rect 14940 138 15636 218
rect 16859 138 16898 218
rect 9778 -407 9851 -7
rect 19258 138 19398 1939
rect 98 -1566 100 -407
rect 5200 -458 7376 -407
rect 7676 -458 9851 -407
<< metal4 >>
rect 0 40800 254 42193
rect 0 39593 287 40800
rect 14746 39593 15000 40000
rect 0 34750 9641 39593
rect 14746 34750 15294 39593
rect 15746 34750 16000 42193
rect 25649 34750 33800 39593
rect 0 19800 254 21193
rect 0 18593 529 19800
rect 0 14540 9543 18593
rect -540 14516 12540 14540
rect -540 -516 -516 14516
rect 574 14280 12540 14516
rect -280 14000 12540 14280
rect -280 13600 9543 14000
rect -280 13540 254 13600
rect 12000 13540 12540 14000
rect 14746 13540 15000 19000
rect 15746 13600 16000 21193
rect 25177 13600 33800 18593
rect -280 13474 522 13540
rect 9418 13474 16000 13540
rect -280 13414 254 13474
rect 12000 13414 12540 13474
rect 14746 13414 15000 13474
rect -280 13300 7288 13414
rect 7752 13300 16000 13414
rect -280 12818 16000 13300
rect -280 12462 9543 12818
rect 12000 12462 12540 12818
rect 14746 12462 15000 12818
rect 15746 12462 16000 12818
rect -280 11866 10429 12462
rect 10893 11866 16000 12462
rect 25177 12410 33800 13300
rect -280 11806 9543 11866
rect 12000 11806 12540 11866
rect 14746 11806 15000 11866
rect 15746 11806 16000 11866
rect -280 11740 16000 11806
rect -280 11347 9543 11740
rect 12000 11347 12540 11740
rect 14746 11347 15000 11740
rect -280 11281 15000 11347
rect -280 11240 9543 11281
rect -280 11221 4310 11240
rect 12000 11221 12540 11281
rect 14746 11240 15000 11281
rect -280 10940 15000 11221
rect 15746 10940 16000 11740
rect 25177 11240 33800 12130
rect -280 10874 33800 10940
rect -280 10814 15000 10874
rect 15746 10814 16000 10874
rect -280 10218 33800 10814
rect -280 9862 15000 10218
rect 15746 9862 16000 10218
rect 25177 9922 33800 10158
rect -280 9266 33800 9862
rect -280 9206 295 9266
rect 12000 9206 12540 9266
rect 14746 9206 15000 9247
rect 15746 9206 16000 9260
rect -280 9140 33800 9206
rect -280 9117 295 9140
rect -280 8840 254 9117
rect -280 7910 9450 8840
rect -280 7867 254 7910
rect -280 7630 277 7867
rect -280 6940 9543 7630
rect -280 6897 254 6940
rect -280 6660 320 6897
rect -280 5970 9543 6660
rect -280 5967 320 5970
rect -280 5690 254 5967
rect -280 4760 9543 5690
rect -280 4757 305 4760
rect -280 4480 254 4757
rect -280 3550 9543 4480
rect -280 3507 254 3550
rect -280 3270 757 3507
rect -280 2580 9543 3270
rect -280 2577 757 2580
rect -280 2300 254 2577
rect -280 1370 9543 2300
rect -280 1207 470 1370
rect -280 1090 254 1207
rect -280 0 9543 1090
rect 9547 0 9613 4715
rect 9673 0 10269 4175
rect 10329 0 10565 4311
rect 10625 0 11221 5382
rect 11281 0 11347 5435
rect 12000 254 12540 9140
rect 14746 3550 15000 9140
rect 15746 5970 16000 9140
rect 25177 7910 33800 8840
rect 25177 6940 33800 7630
rect 25177 5970 33800 6660
rect 15794 5690 16000 5870
rect 14807 2707 15000 3550
rect 14746 371 15000 2707
rect 15746 2600 16000 5690
rect 25177 4760 33800 5690
rect 24241 3550 33800 4480
rect 15794 2580 16000 2600
rect 24241 2580 33800 3270
rect 15746 1370 16000 2300
rect 25177 1370 33800 2300
rect 15746 371 16000 1090
rect 11647 20 12540 254
rect 11647 0 12280 20
rect -280 -280 12280 0
rect 12516 -516 12540 20
rect 12817 0 13707 254
rect 14007 0 19000 371
rect 25177 0 33800 1090
rect 35157 0 40000 254
rect -540 -540 12540 -516
<< obsm4 >>
rect 334 40800 15666 42193
rect 334 40000 15746 40800
rect 334 39993 14746 40000
rect 287 39593 14746 39993
rect 15000 39593 15746 40000
rect 9641 34750 14746 39593
rect 15294 34750 15746 39593
rect 16000 39593 40000 40800
rect 16000 34750 25649 39593
rect 33800 34750 40000 39593
rect 0 21193 40000 34750
rect 254 19800 15746 21193
rect 529 19000 15746 19800
rect 529 18593 14746 19000
rect 9543 14540 14746 18593
rect -2195 7903 -540 8833
rect 9543 13600 12000 14000
rect 334 13540 12000 13600
rect 12540 13540 14746 14540
rect 15000 13600 15746 19000
rect 16000 18593 40000 21193
rect 16000 13600 25177 18593
rect 33800 13600 40000 18593
rect 15000 13540 40000 13600
rect 522 13474 9418 13540
rect 16000 13474 40000 13540
rect 254 13414 12000 13474
rect 12540 13414 14746 13474
rect 15000 13414 40000 13474
rect 7288 13300 7752 13414
rect 16000 13300 40000 13414
rect 9543 12462 12000 12818
rect 12540 12462 14746 12818
rect 15000 12462 15746 12818
rect 10429 11866 10893 12462
rect 16000 12410 25177 13300
rect 33800 12410 40000 13300
rect 16000 12130 40000 12410
rect 9543 11806 12000 11866
rect 12540 11806 14746 11866
rect 15000 11806 15746 11866
rect 9543 11347 12000 11740
rect 12540 11347 14746 11740
rect 9543 11240 12000 11281
rect 4310 11221 12000 11240
rect 12540 11240 14746 11281
rect 15000 11240 15746 11740
rect 12540 11221 15746 11240
rect 15000 10940 15746 11221
rect 16000 11240 25177 12130
rect 33800 11240 40000 12130
rect 16000 10940 40000 11240
rect 33800 10874 40000 10940
rect 15000 10814 15746 10874
rect 16000 10814 40000 10874
rect 33800 10218 40000 10814
rect 15000 9862 15746 10218
rect 16000 10158 40000 10218
rect 16000 9922 25177 10158
rect 33800 9922 40000 10158
rect 16000 9862 40000 9922
rect 33800 9266 40000 9862
rect 334 9240 12000 9266
rect 295 9206 12000 9240
rect 12540 9260 40000 9266
rect 12540 9247 15746 9260
rect 12540 9206 14746 9247
rect 15000 9206 15746 9247
rect 16000 9206 40000 9260
rect 33800 9140 40000 9206
rect 334 9060 12000 9140
rect 254 8840 12000 9060
rect 9450 7910 12000 8840
rect 334 7830 12000 7910
rect 277 7630 12000 7830
rect 9543 6940 12000 7630
rect 334 6860 12000 6940
rect 320 6660 12000 6860
rect 9543 5970 12000 6660
rect 320 5967 12000 5970
rect 254 5950 12000 5967
rect 273 5890 12000 5950
rect 254 5690 12000 5890
rect 9543 5435 12000 5690
rect 9543 5382 11281 5435
rect 9543 4760 10625 5382
rect 334 4715 10625 4760
rect 334 4680 9547 4715
rect 254 4480 9547 4680
rect 9543 3550 9547 4480
rect 273 3507 9547 3550
rect 757 3270 9547 3507
rect 9543 2580 9547 3270
rect 757 2577 9547 2580
rect 273 2520 9547 2577
rect 254 2300 9547 2520
rect 9543 1370 9547 2300
rect 470 1207 9547 1370
rect 254 1090 9547 1207
rect 9543 0 9547 1090
rect 9613 4311 10625 4715
rect 9613 4175 10329 4311
rect 9613 0 9673 4175
rect 10269 0 10329 4175
rect 10565 0 10625 4311
rect 11221 0 11281 5382
rect 11347 254 12000 5435
rect 12540 3550 14746 9140
rect 15000 5970 15746 9140
rect 16000 8840 40000 9140
rect 16000 7910 25177 8840
rect 33800 7910 40000 8840
rect 16000 7630 40000 7910
rect 16000 6940 25177 7630
rect 33800 6940 40000 7630
rect 16000 6660 40000 6940
rect 16000 5970 25177 6660
rect 33800 5970 40000 6660
rect 15000 5870 40000 5970
rect 15000 5690 15794 5870
rect 16000 5690 40000 5870
rect 12540 2707 14807 3550
rect 12540 371 14746 2707
rect 15000 2600 15746 5690
rect 16000 4760 25177 5690
rect 33800 4760 40000 5690
rect 16000 4480 40000 4760
rect 16000 3550 24241 4480
rect 33800 3550 40000 4480
rect 16000 3270 40000 3550
rect 15000 2580 15794 2600
rect 16000 2580 24241 3270
rect 33800 2580 40000 3270
rect 15000 2300 40000 2580
rect 15000 1370 15746 2300
rect 16000 1370 25177 2300
rect 33800 1370 40000 2300
rect 15000 1090 40000 1370
rect 15000 371 15746 1090
rect 16000 371 25177 1090
rect 12540 254 14007 371
rect 11347 0 11647 254
rect 12540 0 12817 254
rect 13707 0 14007 254
rect 19000 251 25177 371
rect 19000 0 25097 251
rect 33800 334 40000 1090
rect 33800 251 35077 334
rect 13012 -174 13463 -108
rect 15029 -174 15633 -108
rect 12540 -300 15180 -234
<< via4 >>
rect -516 14280 574 14516
rect -516 -280 -280 14280
rect 12280 -280 12516 20
rect -516 -516 12516 -280
<< metal5 >>
rect 0 39593 254 40000
rect 0 35595 4000 39593
rect 14746 35595 15000 40000
rect 0 35157 15000 35595
rect 0 34750 14760 35157
rect 2240 33426 14760 34750
rect 2054 33189 14760 33426
rect 1410 32782 14760 33189
rect 0 19797 254 21190
rect 1410 20617 22978 32782
rect 2054 20505 14760 20617
rect 2054 19973 12934 20505
rect 0 18590 529 19797
rect 0 14540 9543 18590
rect -540 14516 12540 14540
rect -540 8833 -516 14516
rect 334 14280 12540 14516
rect -280 8833 12540 14280
rect -540 7903 12540 8833
rect -540 -516 -516 7903
rect -280 0 12540 7903
rect 14746 3570 15000 18997
rect 15746 13600 16000 20617
rect 25177 13600 33800 18590
rect 15746 5990 16000 13540
rect 25177 12430 33800 13280
rect 25177 11260 33800 12110
rect 25177 9140 33800 10940
rect 25177 7930 33800 8820
rect 25177 6960 33800 7610
rect 25177 5990 33800 6640
rect 15794 5670 16000 5850
rect 14807 2687 15000 3570
rect 14746 371 15000 2687
rect 15746 2620 16000 5670
rect 25177 4780 33800 5670
rect 25177 3570 33800 4460
rect 15794 2600 16000 2620
rect 24241 2600 33800 3250
rect 15746 1390 16000 2280
rect 25177 1390 33800 2280
rect 15746 371 16000 1070
rect 12837 0 13687 254
rect 14007 0 18997 371
rect 25177 20 33800 1070
rect -280 -234 12280 0
rect 12516 -234 12540 0
rect -280 -280 12540 -234
rect 731 -300 12540 -280
rect 12516 -516 12540 -300
rect -540 -540 12540 -516
<< obsm5 >>
rect 0 40800 16000 42193
rect 0 40000 40000 40800
rect 254 39593 14746 40000
rect 4000 35595 14746 39593
rect 15000 35157 40000 40000
rect 0 33426 2240 34750
rect 0 33189 2054 33426
rect 0 21190 1410 33189
rect 14760 32782 40000 35157
rect 254 20617 1410 21190
rect 22978 20617 40000 32782
rect 254 19973 2054 20617
rect 14760 20505 15746 20617
rect 12934 19973 15746 20505
rect 254 19797 15746 19973
rect 529 18997 15746 19797
rect 529 18910 14746 18997
rect 574 18729 14746 18910
rect 529 18629 14746 18729
rect 574 18590 14746 18629
rect 9543 14540 14746 18590
rect 12540 3570 14746 14540
rect 15000 13600 15746 18997
rect 16000 18590 40000 20617
rect 16000 13600 25177 18590
rect 33800 13600 40000 18590
rect 15000 13540 40000 13600
rect 15000 5990 15746 13540
rect 16000 13280 40000 13540
rect 16000 12430 25177 13280
rect 33800 12430 40000 13280
rect 16000 12110 40000 12430
rect 16000 11260 25177 12110
rect 33800 11260 40000 12110
rect 16000 10940 40000 11260
rect 16000 9140 25177 10940
rect 33800 9140 40000 10940
rect 16000 8820 40000 9140
rect 16000 7930 25177 8820
rect 33800 7930 40000 8820
rect 16000 7610 40000 7930
rect 16000 6960 25177 7610
rect 33800 6960 40000 7610
rect 16000 6640 40000 6960
rect 16000 5990 25177 6640
rect 33800 5990 40000 6640
rect 15000 5850 40000 5990
rect 15000 5670 15794 5850
rect 16000 5670 40000 5850
rect 12540 2687 14807 3570
rect 12540 371 14746 2687
rect 15000 2620 15746 5670
rect 16000 4780 25177 5670
rect 33800 4780 40000 5670
rect 16000 4460 40000 4780
rect 16000 3570 25177 4460
rect 33800 3570 40000 4460
rect 16000 3250 40000 3570
rect 15000 2600 15794 2620
rect 16000 2600 24241 3250
rect 33800 2600 40000 3250
rect 15000 2280 40000 2600
rect 15000 1390 15746 2280
rect 16000 1390 25177 2280
rect 33800 1390 40000 2280
rect 15000 1070 40000 1390
rect 15000 371 15746 1070
rect 16000 371 25177 1070
rect 12540 254 14007 371
rect 12540 20 12837 254
rect 13687 20 14007 254
rect 18997 20 25177 371
rect 33800 20 40000 1070
rect 19317 0 40000 20
<< labels >>
rlabel metal3 s 4944 0 9944 16470 6 P_CORE
port 1 nsew
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 2 nsew
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 2 nsew
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 2 nsew
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 2 nsew
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 2 nsew
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 2 nsew
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 2 nsew
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 2 nsew
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 2 nsew
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 2 nsew
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 2 nsew
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 2 nsew
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 3 nsew
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 3 nsew
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 3 nsew
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 3 nsew
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 4 nsew
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 4 nsew
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 5 nsew
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 5 nsew
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 6 nsew
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 6 nsew
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 6 nsew
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 6 nsew
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 7 nsew
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 7 nsew
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 7 nsew
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 7 nsew
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 7 nsew
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 7 nsew
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 7 nsew
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 7 nsew
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 8 nsew
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 8 nsew
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 8 nsew
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 8 nsew
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 9 nsew
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 9 nsew
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 9 nsew
rlabel metal4 s 126 38320 128 38322 6 VSSIO
port 9 nsew
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 9 nsew
rlabel metal4 s 14872 38320 14874 38322 6 VSSIO
port 9 nsew
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 9 nsew
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 9 nsew
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 9 nsew
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 9 nsew
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 10 nsew
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 10 nsew
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 10 nsew
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 10 nsew
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 11 nsew
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 11 nsew
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 11 nsew
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 11 nsew
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 12 nsew
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 12 nsew
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 12 nsew
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 12 nsew
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 13 nsew
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 13 nsew
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 13 nsew
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 13 nsew
rlabel metal5 s 1410 21024 13578 33189 6 P_PAD
port 14 nsew
rlabel metal3 s 4944 0 9944 16470 6 P_CORE
port 15 nsew
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 16 nsew
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 16 nsew
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 16 nsew
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 16 nsew
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 16 nsew
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 16 nsew
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 16 nsew
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 16 nsew
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 16 nsew
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 16 nsew
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 16 nsew
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 16 nsew
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 17 nsew
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 17 nsew
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 17 nsew
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 17 nsew
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 18 nsew
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 18 nsew
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 19 nsew
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 19 nsew
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 20 nsew
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 20 nsew
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 20 nsew
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 20 nsew
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 21 nsew
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 21 nsew
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 21 nsew
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 21 nsew
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 21 nsew
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 21 nsew
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 21 nsew
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 21 nsew
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 22 nsew
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 22 nsew
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 22 nsew
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 22 nsew
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 23 nsew
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 23 nsew
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 23 nsew
rlabel metal4 s 126 38320 128 38322 6 VSSIO
port 23 nsew
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 23 nsew
rlabel metal4 s 14872 38320 14874 38322 6 VSSIO
port 23 nsew
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 23 nsew
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 23 nsew
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 23 nsew
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 23 nsew
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 24 nsew
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 24 nsew
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 24 nsew
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 24 nsew
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 25 nsew
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 25 nsew
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 25 nsew
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 25 nsew
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 26 nsew
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 26 nsew
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 26 nsew
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 26 nsew
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 27 nsew
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 27 nsew
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 27 nsew
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 27 nsew
rlabel metal5 s 1410 21024 13578 33189 6 P_PAD
port 28 nsew
rlabel metal3 s 4944 0 9944 16470 6 P_CORE
port 29 nsew
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 30 nsew
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 30 nsew
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 30 nsew
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 30 nsew
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 30 nsew
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 30 nsew
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 30 nsew
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 30 nsew
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 30 nsew
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 30 nsew
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 30 nsew
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 30 nsew
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 31 nsew
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 31 nsew
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 31 nsew
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 31 nsew
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 32 nsew
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 32 nsew
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 33 nsew
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 33 nsew
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 34 nsew
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 34 nsew
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 34 nsew
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 34 nsew
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 35 nsew
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 35 nsew
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 35 nsew
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 35 nsew
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 35 nsew
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 35 nsew
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 35 nsew
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 35 nsew
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 36 nsew
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 36 nsew
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 36 nsew
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 36 nsew
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 37 nsew
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 37 nsew
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 37 nsew
rlabel metal4 s 126 38320 128 38322 6 VSSIO
port 37 nsew
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 37 nsew
rlabel metal4 s 14872 38320 14874 38322 6 VSSIO
port 37 nsew
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 37 nsew
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 37 nsew
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 37 nsew
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 37 nsew
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 38 nsew
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 38 nsew
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 38 nsew
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 38 nsew
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 39 nsew
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 39 nsew
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 39 nsew
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 39 nsew
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 40 nsew
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 40 nsew
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 40 nsew
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 40 nsew
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 41 nsew
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 41 nsew
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 41 nsew
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 41 nsew
rlabel metal5 s 1410 21024 13578 33189 6 P_PAD
port 42 nsew
rlabel metal5 s -540 -540 12540 14540 6 PAD
port 43 nsew
rlabel via4 s -516 -516 12516 -280 8 PAD
port 43 nsew
rlabel via4 s 12280 -280 12516 14280 6 PAD
port 43 nsew
rlabel via4 s -516 -280 -280 14280 4 PAD
port 43 nsew
rlabel via4 s -516 14280 12516 14516 6 PAD
port 43 nsew
rlabel metal4 s -540 -540 12540 0 8 PAD
port 43 nsew
rlabel metal4 s 12000 0 12540 14000 6 PAD
port 43 nsew
rlabel metal4 s -540 0 0 14000 4 PAD
port 43 nsew
rlabel metal4 s -540 14000 12540 14540 6 PAD
port 43 nsew
rlabel metal4 s 0 10218 200 10814 6 AMUXBUS_A
port 44 nsew signal bidirectional
rlabel metal4 s 0 9266 200 9862 6 AMUXBUS_B
port 45 nsew signal bidirectional
rlabel metal5 s 0 9140 200 10940 6 VSSA
port 46 nsew ground bidirectional
rlabel metal4 s 0 10874 200 10940 6 VSSA
port 46 nsew ground bidirectional
rlabel metal4 s 0 9140 200 9206 6 VSSA
port 46 nsew ground bidirectional
rlabel metal5 s 0 6960 200 7610 6 VSSA
port 46 nsew ground bidirectional
rlabel metal4 s 0 6940 200 7630 6 VSSA
port 46 nsew ground bidirectional
rlabel metal5 s 0 2600 200 3250 6 VDDA
port 47 nsew power bidirectional
rlabel metal4 s 0 2580 200 3270 6 VDDA
port 47 nsew power bidirectional
rlabel metal5 s 0 5990 200 6640 6 VSWITCH
port 48 nsew power bidirectional
rlabel metal4 s 0 5970 200 6660 6 VSWITCH
port 48 nsew power bidirectional
rlabel metal5 s 0 12430 200 13280 6 VDDIO_Q
port 49 nsew power bidirectional
rlabel metal4 s 0 12410 200 13300 6 VDDIO_Q
port 49 nsew power bidirectional
rlabel metal5 s 0 20 200 1070 6 VCCHIB
port 50 nsew power bidirectional
rlabel metal4 s 0 0 200 1090 6 VCCHIB
port 50 nsew power bidirectional
rlabel metal5 s 0 13600 200 18590 6 VDDIO
port 51 nsew power bidirectional
rlabel metal4 s 0 13600 200 18593 6 VDDIO
port 51 nsew power bidirectional
rlabel metal5 s 0 3570 200 4460 6 VDDIO
port 51 nsew power bidirectional
rlabel metal4 s 0 3550 200 4480 6 VDDIO
port 51 nsew power bidirectional
rlabel metal5 s 0 1390 200 2280 6 VCCD
port 52 nsew power bidirectional
rlabel metal4 s 0 1370 200 2300 6 VCCD
port 52 nsew power bidirectional
rlabel metal5 s 0 4780 200 5670 6 VSSIO
port 53 nsew ground bidirectional
rlabel metal4 s 0 4760 200 5690 6 VSSIO
port 53 nsew ground bidirectional
rlabel metal5 s 0 34750 200 39593 6 VSSIO
port 53 nsew ground bidirectional
rlabel metal5 s 0 7930 200 8820 6 VSSD
port 54 nsew ground bidirectional
rlabel metal4 s 0 7910 200 8840 6 VSSD
port 54 nsew ground bidirectional
rlabel metal5 s 0 11260 200 12110 6 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 0 11240 200 12130 6 VSSIO_Q
port 55 nsew ground bidirectional
rlabel metal4 s 0 10218 1000 10814 6 AMUXBUS_A
port 56 nsew signal bidirectional
rlabel metal4 s 0 9266 1000 9862 6 AMUXBUS_B
port 57 nsew signal bidirectional
rlabel metal5 s 0 9140 1000 10940 6 VSSA
port 58 nsew ground bidirectional
rlabel metal4 s 0 10874 1000 10940 6 VSSA
port 58 nsew ground bidirectional
rlabel metal4 s 0 9140 1000 9206 6 VSSA
port 58 nsew ground bidirectional
rlabel metal5 s 0 6960 1000 7610 6 VSSA
port 58 nsew ground bidirectional
rlabel metal4 s 0 6940 1000 7630 6 VSSA
port 58 nsew ground bidirectional
rlabel metal5 s 0 2600 1000 3250 6 VDDA
port 59 nsew power bidirectional
rlabel metal4 s 0 2580 1000 3270 6 VDDA
port 59 nsew power bidirectional
rlabel metal5 s 0 5990 1000 6640 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal4 s 0 5970 1000 6660 6 VSWITCH
port 60 nsew power bidirectional
rlabel metal5 s 0 12430 1000 13280 6 VDDIO_Q
port 61 nsew power bidirectional
rlabel metal4 s 0 12410 1000 13300 6 VDDIO_Q
port 61 nsew power bidirectional
rlabel metal5 s 0 20 1000 1070 6 VCCHIB
port 62 nsew power bidirectional
rlabel metal4 s 0 0 1000 1090 6 VCCHIB
port 62 nsew power bidirectional
rlabel metal5 s 0 13600 1000 18590 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 0 13600 1000 18593 6 VDDIO
port 63 nsew power bidirectional
rlabel metal5 s 0 3570 1000 4460 6 VDDIO
port 63 nsew power bidirectional
rlabel metal4 s 0 3550 1000 4480 6 VDDIO
port 63 nsew power bidirectional
rlabel metal5 s 0 1390 1000 2280 6 VCCD
port 64 nsew power bidirectional
rlabel metal4 s 0 1370 1000 2300 6 VCCD
port 64 nsew power bidirectional
rlabel metal5 s 0 4780 1000 5670 6 VSSIO
port 65 nsew ground bidirectional
rlabel metal4 s 0 4760 1000 5690 6 VSSIO
port 65 nsew ground bidirectional
rlabel metal5 s 0 34750 1000 39593 6 VSSIO
port 65 nsew ground bidirectional
rlabel metal5 s 0 7930 1000 8820 6 VSSD
port 66 nsew ground bidirectional
rlabel metal4 s 0 7910 1000 8840 6 VSSD
port 66 nsew ground bidirectional
rlabel metal5 s 0 11260 1000 12110 6 VSSIO_Q
port 67 nsew ground bidirectional
rlabel metal4 s 0 11240 1000 12130 6 VSSIO_Q
port 67 nsew ground bidirectional
rlabel metal4 s 0 10218 2000 10814 6 AMUXBUS_A
port 68 nsew signal bidirectional
rlabel metal4 s 0 9266 2000 9862 6 AMUXBUS_B
port 69 nsew signal bidirectional
rlabel metal5 s 0 9140 2000 10940 6 VSSA
port 70 nsew ground bidirectional
rlabel metal4 s 0 10874 2000 10940 6 VSSA
port 70 nsew ground bidirectional
rlabel metal4 s 0 9140 2000 9206 6 VSSA
port 70 nsew ground bidirectional
rlabel metal5 s 0 6960 2000 7610 6 VSSA
port 70 nsew ground bidirectional
rlabel metal4 s 0 6940 2000 7630 6 VSSA
port 70 nsew ground bidirectional
rlabel metal5 s 0 2600 2000 3250 6 VDDA
port 71 nsew power bidirectional
rlabel metal4 s 0 2580 2000 3270 6 VDDA
port 71 nsew power bidirectional
rlabel metal5 s 0 5990 2000 6640 6 VSWITCH
port 72 nsew power bidirectional
rlabel metal4 s 0 5970 2000 6660 6 VSWITCH
port 72 nsew power bidirectional
rlabel metal5 s 0 12430 2000 13280 6 VDDIO_Q
port 73 nsew power bidirectional
rlabel metal4 s 0 12410 2000 13300 6 VDDIO_Q
port 73 nsew power bidirectional
rlabel metal5 s 0 20 2000 1070 6 VCCHIB
port 74 nsew power bidirectional
rlabel metal4 s 0 0 2000 1090 6 VCCHIB
port 74 nsew power bidirectional
rlabel metal5 s 0 13600 2000 18590 6 VDDIO
port 75 nsew power bidirectional
rlabel metal4 s 0 13600 2000 18593 6 VDDIO
port 75 nsew power bidirectional
rlabel metal5 s 0 3570 2000 4460 6 VDDIO
port 75 nsew power bidirectional
rlabel metal4 s 0 3550 2000 4480 6 VDDIO
port 75 nsew power bidirectional
rlabel metal5 s 0 1390 2000 2280 6 VCCD
port 76 nsew power bidirectional
rlabel metal4 s 0 1370 2000 2300 6 VCCD
port 76 nsew power bidirectional
rlabel metal5 s 0 4780 2000 5670 6 VSSIO
port 77 nsew ground bidirectional
rlabel metal4 s 0 4760 2000 5690 6 VSSIO
port 77 nsew ground bidirectional
rlabel metal5 s 0 34750 2000 39593 6 VSSIO
port 77 nsew ground bidirectional
rlabel metal5 s 0 7930 2000 8820 6 VSSD
port 78 nsew ground bidirectional
rlabel metal4 s 0 7910 2000 8840 6 VSSD
port 78 nsew ground bidirectional
rlabel metal5 s 0 11260 2000 12110 6 VSSIO_Q
port 79 nsew ground bidirectional
rlabel metal4 s 0 11240 2000 12130 6 VSSIO_Q
port 79 nsew ground bidirectional
rlabel metal4 s 0 10218 4000 10814 6 AMUXBUS_A
port 80 nsew signal bidirectional
rlabel metal4 s 0 9266 4000 9862 6 AMUXBUS_B
port 81 nsew signal bidirectional
rlabel metal5 s 0 9140 4000 10940 6 VSSA
port 82 nsew ground bidirectional
rlabel metal4 s 0 10874 4000 10940 6 VSSA
port 82 nsew ground bidirectional
rlabel metal4 s 0 9140 4000 9206 6 VSSA
port 82 nsew ground bidirectional
rlabel metal5 s 0 6960 4000 7610 6 VSSA
port 82 nsew ground bidirectional
rlabel metal4 s 0 6940 4000 7630 6 VSSA
port 82 nsew ground bidirectional
rlabel metal5 s 0 2600 4000 3250 6 VDDA
port 83 nsew power bidirectional
rlabel metal4 s 0 2580 4000 3270 6 VDDA
port 83 nsew power bidirectional
rlabel metal5 s 0 5990 4000 6640 6 VSWITCH
port 84 nsew power bidirectional
rlabel metal4 s 0 5970 4000 6660 6 VSWITCH
port 84 nsew power bidirectional
rlabel metal5 s 0 12430 4000 13280 6 VDDIO_Q
port 85 nsew power bidirectional
rlabel metal4 s 0 12410 4000 13300 6 VDDIO_Q
port 85 nsew power bidirectional
rlabel metal5 s 0 20 4000 1070 6 VCCHIB
port 86 nsew power bidirectional
rlabel metal4 s 0 0 4000 1090 6 VCCHIB
port 86 nsew power bidirectional
rlabel metal5 s 0 13600 4000 18590 6 VDDIO
port 87 nsew power bidirectional
rlabel metal4 s 0 13600 4000 18593 6 VDDIO
port 87 nsew power bidirectional
rlabel metal5 s 0 3570 4000 4460 6 VDDIO
port 87 nsew power bidirectional
rlabel metal4 s 0 3550 4000 4480 6 VDDIO
port 87 nsew power bidirectional
rlabel metal5 s 0 1390 4000 2280 6 VCCD
port 88 nsew power bidirectional
rlabel metal4 s 0 1370 4000 2300 6 VCCD
port 88 nsew power bidirectional
rlabel metal5 s 0 4780 4000 5670 6 VSSIO
port 89 nsew ground bidirectional
rlabel metal4 s 0 4760 4000 5690 6 VSSIO
port 89 nsew ground bidirectional
rlabel metal5 s 0 34750 4000 39593 6 VSSIO
port 89 nsew ground bidirectional
rlabel metal5 s 0 7930 4000 8820 6 VSSD
port 90 nsew ground bidirectional
rlabel metal4 s 0 7910 4000 8840 6 VSSD
port 90 nsew ground bidirectional
rlabel metal5 s 0 11260 4000 12110 6 VSSIO_Q
port 91 nsew ground bidirectional
rlabel metal4 s 0 11240 4000 12130 6 VSSIO_Q
port 91 nsew ground bidirectional
rlabel metal4 s 0 10218 4000 10814 6 AMUXBUS_A
port 92 nsew signal bidirectional
rlabel metal4 s 0 9266 4000 9862 6 AMUXBUS_B
port 93 nsew signal bidirectional
rlabel metal5 s 0 9140 4000 10940 6 VSSA
port 94 nsew ground bidirectional
rlabel metal4 s 0 10874 4000 10940 6 VSSA
port 94 nsew ground bidirectional
rlabel metal4 s 0 9140 4000 9206 6 VSSA
port 94 nsew ground bidirectional
rlabel metal5 s 0 6960 4000 7610 6 VSSA
port 94 nsew ground bidirectional
rlabel metal4 s 0 6940 4000 7630 6 VSSA
port 94 nsew ground bidirectional
rlabel metal5 s 0 2600 4000 3250 6 VDDA
port 95 nsew power bidirectional
rlabel metal4 s 0 2580 4000 3270 6 VDDA
port 95 nsew power bidirectional
rlabel metal5 s 0 5990 4000 6640 6 VSWITCH
port 96 nsew power bidirectional
rlabel metal4 s 0 3550 4000 4480 6 VSWITCH
port 96 nsew power bidirectional
rlabel metal4 s 0 5970 4000 6660 6 VSWITCH
port 96 nsew power bidirectional
rlabel via3 s 256 3616 3754 4418 6 VSWITCH
port 96 nsew power bidirectional
rlabel via3 s 218 6016 3748 6606 6 VSWITCH
port 96 nsew power bidirectional
rlabel metal3 s 198 3576 3800 6640 6 VSWITCH
port 96 nsew power bidirectional
rlabel metal5 s 0 12430 4000 13280 6 VDDIO_Q
port 97 nsew power bidirectional
rlabel metal4 s 0 12410 4000 13300 6 VDDIO_Q
port 97 nsew power bidirectional
rlabel metal5 s 0 20 4000 2280 6 VCCHIB
port 98 nsew power bidirectional
rlabel metal4 s 0 0 4000 1090 6 VCCHIB
port 98 nsew power bidirectional
rlabel metal5 s 0 13600 4000 18590 6 VDDIO
port 99 nsew power bidirectional
rlabel metal4 s 0 13600 4000 18593 6 VDDIO
port 99 nsew power bidirectional
rlabel metal5 s 0 3570 4000 4460 6 VDDIO
port 99 nsew power bidirectional
rlabel metal4 s 0 1370 4000 2300 6 VCCD
port 100 nsew power bidirectional
rlabel metal5 s 0 4780 4000 5670 6 VSSIO
port 101 nsew ground bidirectional
rlabel metal4 s 0 4760 4000 5690 6 VSSIO
port 101 nsew ground bidirectional
rlabel metal5 s 0 34750 4000 39593 6 VSSIO
port 101 nsew ground bidirectional
rlabel metal5 s 0 7930 4000 8820 6 VSSD
port 102 nsew ground bidirectional
rlabel metal4 s 0 7910 4000 8840 6 VSSD
port 102 nsew ground bidirectional
rlabel metal5 s 0 11260 4000 12110 6 VSSIO_Q
port 103 nsew ground bidirectional
rlabel metal4 s 0 11240 4000 12130 6 VSSIO_Q
port 103 nsew ground bidirectional
rlabel metal4 s 0 11425 4582 12021 6 AMUXBUS_A
port 104 nsew signal bidirectional
rlabel metal4 s 10625 0 11221 5382 6 AMUXBUS_A
port 104 nsew signal bidirectional
rlabel metal4 s 0 10473 4187 11069 6 AMUXBUS_B
port 105 nsew signal bidirectional
rlabel metal4 s 9673 0 10269 4175 6 AMUXBUS_B
port 105 nsew signal bidirectional
rlabel metal5 s 0 10347 4631 12147 6 VSSA
port 106 nsew ground bidirectional
rlabel metal5 s 0 8167 267 8817 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 0 10347 3915 10413 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 0 8147 267 8837 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 0 11129 4310 11365 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 0 12081 4635 12147 6 VSSA
port 106 nsew ground bidirectional
rlabel metal5 s 7368 0 8017 254 6 VSSA
port 106 nsew ground bidirectional
rlabel metal5 s 9547 0 11347 5431 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 11281 0 11347 5435 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 10329 0 10565 4311 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 7347 0 8037 254 6 VSSA
port 106 nsew ground bidirectional
rlabel metal4 s 9547 0 9613 4715 6 VSSA
port 106 nsew ground bidirectional
rlabel metal5 s 0 3807 294 4457 6 VDDA
port 107 nsew power bidirectional
rlabel metal4 s 0 3787 294 4477 6 VDDA
port 107 nsew power bidirectional
rlabel metal5 s 3007 0 3657 251 6 VDDA
port 107 nsew power bidirectional
rlabel metal4 s 2987 0 3677 251 6 VDDA
port 107 nsew power bidirectional
rlabel metal5 s 0 7197 277 7847 6 VSWITCH
port 108 nsew power bidirectional
rlabel metal4 s 0 7177 277 7867 6 VSWITCH
port 108 nsew power bidirectional
rlabel metal5 s 6397 0 7047 254 6 VSWITCH
port 108 nsew power bidirectional
rlabel metal4 s 6377 0 7067 254 6 VSWITCH
port 108 nsew power bidirectional
rlabel metal5 s 0 13637 296 14487 6 VDDIO_Q
port 109 nsew power bidirectional
rlabel metal4 s 0 13617 296 14507 6 VDDIO_Q
port 109 nsew power bidirectional
rlabel metal5 s 12837 0 13687 254 6 VDDIO_Q
port 109 nsew power bidirectional
rlabel metal4 s 12817 0 13707 254 6 VDDIO_Q
port 109 nsew power bidirectional
rlabel metal5 s 0 1227 470 2277 6 VCCHIB
port 110 nsew power bidirectional
rlabel metal4 s 0 1207 470 2297 6 VCCHIB
port 110 nsew power bidirectional
rlabel metal5 s 427 0 1477 254 6 VCCHIB
port 110 nsew power bidirectional
rlabel metal4 s 407 0 1497 254 6 VCCHIB
port 110 nsew power bidirectional
rlabel metal5 s 0 14807 529 19797 6 VDDIO
port 111 nsew power bidirectional
rlabel metal5 s 0 4777 305 5667 6 VDDIO
port 111 nsew power bidirectional
rlabel metal4 s 0 4757 305 5687 6 VDDIO
port 111 nsew power bidirectional
rlabel metal4 s 0 14807 529 19800 6 VDDIO
port 111 nsew power bidirectional
rlabel metal5 s 3977 0 4867 254 6 VDDIO
port 111 nsew power bidirectional
rlabel metal5 s 14007 0 18997 371 6 VDDIO
port 111 nsew power bidirectional
rlabel metal4 s 14007 0 19000 371 6 VDDIO
port 111 nsew power bidirectional
rlabel metal4 s 3957 0 4887 254 6 VDDIO
port 111 nsew power bidirectional
rlabel metal5 s 0 2597 757 3487 6 VCCD
port 112 nsew power bidirectional
rlabel metal4 s 0 2577 757 3507 6 VCCD
port 112 nsew power bidirectional
rlabel metal5 s 1797 0 2687 254 6 VCCD
port 112 nsew power bidirectional
rlabel metal4 s 1777 0 2707 254 6 VCCD
port 112 nsew power bidirectional
rlabel metal5 s 0 5987 320 6877 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal4 s 0 5967 320 6897 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal4 s 0 35957 287 40800 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal5 s 5187 0 6077 254 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal4 s 5167 0 6097 254 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal4 s 35157 0 40000 254 6 VSSIO
port 113 nsew ground bidirectional
rlabel metal5 s 0 9137 295 10027 6 VSSD
port 114 nsew ground bidirectional
rlabel metal4 s 0 9117 295 10047 6 VSSD
port 114 nsew ground bidirectional
rlabel metal5 s 8337 0 9227 254 6 VSSD
port 114 nsew ground bidirectional
rlabel metal4 s 8317 0 9247 254 6 VSSD
port 114 nsew ground bidirectional
rlabel metal5 s 0 12467 325 13317 6 VSSIO_Q
port 115 nsew ground bidirectional
rlabel metal4 s 0 12447 325 13337 6 VSSIO_Q
port 115 nsew ground bidirectional
rlabel metal5 s 11667 0 12517 254 6 VSSIO_Q
port 115 nsew ground bidirectional
rlabel metal4 s 11647 0 12537 254 6 VSSIO_Q
port 115 nsew ground bidirectional
rlabel metal4 s 0 10218 1000 10814 6 AMUXBUS_A
port 116 nsew signal bidirectional
rlabel metal4 s 0 9266 1000 9862 6 AMUXBUS_B
port 117 nsew signal bidirectional
rlabel metal5 s 0 9140 1000 10940 6 VSSA
port 118 nsew ground bidirectional
rlabel metal4 s 0 10874 1000 10940 6 VSSA
port 118 nsew ground bidirectional
rlabel metal4 s 0 9140 1000 9206 6 VSSA
port 118 nsew ground bidirectional
rlabel metal5 s 0 6960 1000 7610 6 VSSA
port 118 nsew ground bidirectional
rlabel metal4 s 0 6940 1000 7630 6 VSSA
port 118 nsew ground bidirectional
rlabel metal5 s 0 2600 1000 3250 6 VDDA
port 119 nsew power bidirectional
rlabel metal4 s 0 2580 1000 3270 6 VDDA
port 119 nsew power bidirectional
rlabel metal5 s 0 5990 1000 6640 6 VSWITCH
port 120 nsew power bidirectional
rlabel metal4 s 0 5970 1000 6660 6 VSWITCH
port 120 nsew power bidirectional
rlabel metal5 s 0 12430 1000 13280 6 VDDIO_Q
port 121 nsew power bidirectional
rlabel metal4 s 0 12410 1000 13300 6 VDDIO_Q
port 121 nsew power bidirectional
rlabel metal5 s 0 20 1000 1070 6 VCCHIB
port 122 nsew power bidirectional
rlabel metal4 s 0 0 1000 1090 6 VCCHIB
port 122 nsew power bidirectional
rlabel metal5 s 0 13600 1000 18590 6 VDDIO
port 123 nsew power bidirectional
rlabel metal4 s 0 13600 1000 18593 6 VDDIO
port 123 nsew power bidirectional
rlabel metal5 s 0 3570 1000 4460 6 VDDIO
port 123 nsew power bidirectional
rlabel metal4 s 0 3550 1000 4480 6 VDDIO
port 123 nsew power bidirectional
rlabel metal5 s 0 4780 1000 5670 6 VSSIO
port 124 nsew ground bidirectional
rlabel metal4 s 0 4760 1000 5690 6 VSSIO
port 124 nsew ground bidirectional
rlabel metal5 s 0 34750 1000 39593 6 VSSIO
port 124 nsew ground bidirectional
rlabel metal5 s 0 11260 1000 12110 6 VSSIO_Q
port 125 nsew ground bidirectional
rlabel metal4 s 0 11240 1000 12130 6 VSSIO_Q
port 125 nsew ground bidirectional
rlabel metal4 s 0 10218 1000 10814 6 AMUXBUS_A
port 126 nsew signal bidirectional
rlabel metal4 s 0 9266 1000 9862 6 AMUXBUS_B
port 127 nsew signal bidirectional
rlabel metal5 s 0 5990 1000 6640 6 VSWITCH
port 128 nsew power bidirectional
rlabel metal4 s 0 5970 1000 6660 6 VSWITCH
port 128 nsew power bidirectional
rlabel metal5 s 0 12430 1000 13280 6 VDDIO_Q
port 129 nsew power bidirectional
rlabel metal4 s 0 12410 1000 13300 6 VDDIO_Q
port 129 nsew power bidirectional
rlabel metal5 s 0 20 1000 1070 6 VCCHIB
port 130 nsew power bidirectional
rlabel metal4 s 0 0 1000 1090 6 VCCHIB
port 130 nsew power bidirectional
rlabel metal4 s 0 3550 1000 4480 6 VDDIO
port 131 nsew power bidirectional
rlabel metal5 s 0 13600 1000 18590 6 VDDIO
port 131 nsew power bidirectional
rlabel metal4 s 0 13600 1000 18593 6 VDDIO
port 131 nsew power bidirectional
rlabel metal5 s 0 3570 1000 4460 6 VDDIO
port 131 nsew power bidirectional
rlabel metal5 s 0 1390 1000 2280 6 VCCD
port 132 nsew power bidirectional
rlabel metal4 s 0 1370 1000 2300 6 VCCD
port 132 nsew power bidirectional
rlabel metal5 s 0 4780 1000 5670 6 VSSIO
port 133 nsew ground bidirectional
rlabel metal4 s 0 4760 1000 5690 6 VSSIO
port 133 nsew ground bidirectional
rlabel metal5 s 0 34750 1000 39593 6 VSSIO
port 133 nsew ground bidirectional
rlabel metal5 s 0 7930 1000 8820 6 VSSD
port 134 nsew ground bidirectional
rlabel metal4 s 0 7910 1000 8840 6 VSSD
port 134 nsew ground bidirectional
rlabel metal5 s 0 11260 1000 12110 6 VSSIO_Q
port 135 nsew ground bidirectional
rlabel metal4 s 0 11240 1000 12130 6 VSSIO_Q
port 135 nsew ground bidirectional
rlabel metal4 s 0 10218 7288 10814 6 AMUXBUS_A
port 136 nsew signal bidirectional
rlabel metal4 s 7752 10218 16000 10814 6 AMUXBUS_A
port 136 nsew signal bidirectional
rlabel metal4 s 0 9266 10429 9862 6 AMUXBUS_B
port 137 nsew signal bidirectional
rlabel metal4 s 10893 9266 16000 9862 6 AMUXBUS_B
port 137 nsew signal bidirectional
rlabel metal1 s 12486 -407 12538 -146 8 ANALOG_EN
port 138 nsew signal input
rlabel metal3 s 9173 -407 9239 6954 6 ANALOG_POL
port 139 nsew signal input
rlabel metal2 s 6150 -407 6202 46 8 ANALOG_SEL
port 140 nsew signal input
rlabel metal2 s 5698 -407 5750 407 8 DM[2]
port 141 nsew signal input
rlabel metal2 s 13367 -407 13419 -168 8 DM[1]
port 142 nsew signal input
rlabel metal2 s 9971 -407 10023 -298 8 DM[0]
port 143 nsew signal input
rlabel metal2 s 7092 -407 7144 -97 8 ENABLE_H
port 144 nsew signal input
rlabel metal2 s 7678 -407 7730 211 8 ENABLE_INP_H
port 145 nsew signal input
rlabel metal2 s 2551 -407 2603 663 6 ENABLE_VDDA_H
port 146 nsew signal input
rlabel metal3 s 15716 -407 15782 36548 6 ENABLE_VDDIO
port 147 nsew signal input
rlabel metal2 s 3262 -407 3314 57 8 ENABLE_VSWITCH_H
port 148 nsew signal input
rlabel metal2 s 6363 -407 6415 261 8 HLD_H_N
port 149 nsew signal input
rlabel metal2 s 5320 -407 5372 134 8 HLD_OVR
port 150 nsew signal input
rlabel metal2 s 1084 -407 1130 488 6 IB_MODE_SEL
port 151 nsew signal input
rlabel metal3 s 15848 -407 15914 37505 6 IN
port 152 nsew signal output
rlabel metal3 s 80 -407 204 35290 6 IN_H
port 153 nsew signal output
rlabel metal2 s 9049 -407 9101 611 6 INP_DIS
port 154 nsew signal input
rlabel metal2 s 675 -407 721 488 6 OE_N
port 155 nsew signal input
rlabel metal2 s 4471 -407 4523 878 6 OUT
port 156 nsew signal input
rlabel metal5 s 2240 20505 14760 32995 6 PAD
port 157 nsew signal bidirectional
rlabel metal2 s 15256 -407 15384 4 8 PAD_A_ESD_0_H
port 158 nsew signal bidirectional
rlabel metal2 s 13655 -407 13785 47 8 PAD_A_ESD_1_H
port 159 nsew signal bidirectional
rlabel metal3 s 12564 -407 12778 1534 6 PAD_A_NOESD_H
port 160 nsew signal bidirectional
rlabel metal2 s 15522 -407 15574 -170 8 SLOW
port 161 nsew signal input
rlabel metal2 s 15741 -407 15781 -164 8 TIE_HI_ESD
port 162 nsew signal output
rlabel metal2 s 15943 -407 15983 35167 6 TIE_LO_ESD
port 163 nsew signal output
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 164 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 164 nsew power bidirectional
rlabel metal5 s 15746 1390 16000 2280 6 VCCD
port 164 nsew power bidirectional
rlabel metal4 s 15746 1370 16000 2300 6 VCCD
port 164 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 165 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 165 nsew power bidirectional
rlabel metal5 s 15746 20 16000 1070 6 VCCHIB
port 165 nsew power bidirectional
rlabel metal4 s 15746 0 16000 1090 6 VCCHIB
port 165 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 166 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 166 nsew power bidirectional
rlabel metal5 s 15794 2600 16000 3250 6 VDDA
port 166 nsew power bidirectional
rlabel metal4 s 15794 2580 16000 3270 6 VDDA
port 166 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 167 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 167 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 167 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 167 nsew power bidirectional
rlabel metal5 s 15746 13600 16000 18590 6 VDDIO
port 167 nsew power bidirectional
rlabel metal5 s 15746 3570 16000 4460 6 VDDIO
port 167 nsew power bidirectional
rlabel metal4 s 15746 3550 16000 4480 6 VDDIO
port 167 nsew power bidirectional
rlabel metal4 s 15746 13600 16000 18593 6 VDDIO
port 167 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 168 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 168 nsew power bidirectional
rlabel metal5 s 15746 12430 16000 13280 6 VDDIO_Q
port 168 nsew power bidirectional
rlabel metal4 s 15746 12410 16000 13300 6 VDDIO_Q
port 168 nsew power bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 169 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 0 9140 522 9206 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 0 10874 522 10940 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 169 nsew ground bidirectional
rlabel metal5 s 15746 9140 16000 10940 6 VSSA
port 169 nsew ground bidirectional
rlabel metal5 s 15746 6961 16000 7610 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 15746 9922 16000 10158 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 9418 10874 16000 10940 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 9418 9140 16000 9206 6 VSSA
port 169 nsew ground bidirectional
rlabel metal4 s 15746 6940 16000 7630 6 VSSA
port 169 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 170 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 170 nsew ground bidirectional
rlabel metal5 s 15746 7930 16000 8820 6 VSSD
port 170 nsew ground bidirectional
rlabel metal4 s 15746 7910 16000 8840 6 VSSD
port 170 nsew ground bidirectional
rlabel metal4 s 0 34750 162 39593 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal4 s 15794 34750 16000 39593 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal5 s 15746 4780 16000 5670 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal4 s 15746 4760 16000 5690 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal4 s 15746 34750 16000 39593 6 VSSIO
port 171 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 172 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 172 nsew ground bidirectional
rlabel metal5 s 15746 11260 16000 12110 6 VSSIO_Q
port 172 nsew ground bidirectional
rlabel metal4 s 15746 11240 16000 12130 6 VSSIO_Q
port 172 nsew ground bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 173 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 173 nsew power bidirectional
rlabel metal5 s 15746 5990 16000 6640 6 VSWITCH
port 173 nsew power bidirectional
rlabel metal4 s 15746 5970 16000 6660 6 VSWITCH
port 173 nsew power bidirectional
rlabel metal2 s 1226 -407 1278 -97 8 VTRIP_SEL
port 174 nsew signal input
rlabel metal4 s 0 12818 7288 13414 6 AMUXBUS_A
port 175 nsew signal bidirectional
rlabel metal4 s 7752 12818 16000 13414 6 AMUXBUS_A
port 175 nsew signal bidirectional
rlabel metal4 s 0 11866 10429 12462 6 AMUXBUS_B
port 176 nsew signal bidirectional
rlabel metal4 s 10893 11866 16000 12462 6 AMUXBUS_B
port 176 nsew signal bidirectional
rlabel metal2 s 10141 0 10197 480 6 ANALOG_EN
port 177 nsew signal input
rlabel metal2 s 8853 0 8909 480 6 ANALOG_POL
port 178 nsew signal input
rlabel metal2 s 5817 0 5873 480 6 ANALOG_SEL
port 179 nsew signal input
rlabel metal2 s 5173 0 5229 480 6 DM[2]
port 180 nsew signal input
rlabel metal2 s 11337 0 11393 480 6 DM[1]
port 181 nsew signal input
rlabel metal2 s 9497 0 9553 480 6 DM[0]
port 182 nsew signal input
rlabel metal2 s 7013 0 7069 480 6 ENABLE_H
port 183 nsew signal input
rlabel metal2 s 7657 0 7713 480 6 ENABLE_INP_H
port 184 nsew signal input
rlabel metal2 s 2689 0 2745 480 6 ENABLE_VDDA_H
port 185 nsew signal input
rlabel metal2 s 13821 0 13877 480 6 ENABLE_VDDIO
port 186 nsew signal input
rlabel metal2 s 3333 0 3389 480 6 ENABLE_VSWITCH_H
port 187 nsew signal input
rlabel metal2 s 6369 0 6425 480 6 HLD_H_N
port 188 nsew signal input
rlabel metal2 s 4529 0 4585 480 6 HLD_OVR
port 189 nsew signal input
rlabel metal2 s 1493 0 1549 480 6 IB_MODE_SEL
port 190 nsew signal input
rlabel metal2 s 15017 0 15073 480 6 IN
port 191 nsew signal output
rlabel metal2 s 297 0 353 480 6 IN_H
port 192 nsew signal output
rlabel metal2 s 8301 0 8357 480 6 INP_DIS
port 193 nsew signal input
rlabel metal2 s 849 0 905 480 6 OE_N
port 194 nsew signal input
rlabel metal2 s 3977 0 4033 480 6 OUT
port 195 nsew signal input
rlabel metal5 s 2240 23105 14760 35595 6 PAD
port 196 nsew signal bidirectional
rlabel metal2 s 12533 0 12589 480 6 PAD_A_ESD_0_H
port 197 nsew signal bidirectional
rlabel metal2 s 11981 0 12037 480 6 PAD_A_ESD_1_H
port 198 nsew signal bidirectional
rlabel metal2 s 10693 0 10749 480 6 PAD_A_NOESD_H
port 199 nsew signal bidirectional
rlabel metal2 s 13177 0 13233 480 6 SLOW
port 200 nsew signal input
rlabel metal2 s 14373 0 14429 480 6 TIE_HI_ESD
port 201 nsew signal output
rlabel metal2 s 15661 0 15717 480 6 TIE_LO_ESD
port 202 nsew signal output
rlabel metal5 s 0 3990 254 4880 6 VCCD
port 203 nsew power bidirectional
rlabel metal4 s 0 3970 254 4900 6 VCCD
port 203 nsew power bidirectional
rlabel metal5 s 15746 3990 16000 4880 6 VCCD
port 203 nsew power bidirectional
rlabel metal4 s 15746 3970 16000 4900 6 VCCD
port 203 nsew power bidirectional
rlabel metal5 s 0 2620 254 3670 6 VCCHIB
port 204 nsew power bidirectional
rlabel metal4 s 0 2600 254 3690 6 VCCHIB
port 204 nsew power bidirectional
rlabel metal5 s 15746 2620 16000 3670 6 VCCHIB
port 204 nsew power bidirectional
rlabel metal4 s 15746 2600 16000 3690 6 VCCHIB
port 204 nsew power bidirectional
rlabel metal5 s 0 5200 193 5850 6 VDDA
port 205 nsew power bidirectional
rlabel metal4 s 0 5180 193 5870 6 VDDA
port 205 nsew power bidirectional
rlabel metal5 s 15794 5200 16000 5850 6 VDDA
port 205 nsew power bidirectional
rlabel metal4 s 15794 5180 16000 5870 6 VDDA
port 205 nsew power bidirectional
rlabel metal5 s 0 16200 254 21190 6 VDDIO
port 206 nsew power bidirectional
rlabel metal5 s 0 6170 254 7060 6 VDDIO
port 206 nsew power bidirectional
rlabel metal4 s 0 6150 254 7080 6 VDDIO
port 206 nsew power bidirectional
rlabel metal4 s 0 16200 254 21193 6 VDDIO
port 206 nsew power bidirectional
rlabel metal5 s 15746 16200 16000 21190 6 VDDIO
port 206 nsew power bidirectional
rlabel metal5 s 15746 6170 16000 7060 6 VDDIO
port 206 nsew power bidirectional
rlabel metal4 s 15746 6150 16000 7080 6 VDDIO
port 206 nsew power bidirectional
rlabel metal4 s 15746 16200 16000 21193 6 VDDIO
port 206 nsew power bidirectional
rlabel metal5 s 0 15030 254 15880 6 VDDIO_Q
port 207 nsew power bidirectional
rlabel metal4 s 0 15010 254 15900 6 VDDIO_Q
port 207 nsew power bidirectional
rlabel metal5 s 15746 15030 16000 15880 6 VDDIO_Q
port 207 nsew power bidirectional
rlabel metal4 s 15746 15010 16000 15900 6 VDDIO_Q
port 207 nsew power bidirectional
rlabel metal5 s 0 11740 254 13540 6 VSSA
port 208 nsew ground bidirectional
rlabel metal5 s 0 9561 254 10210 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 0 11740 522 11806 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 0 12522 254 12758 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 0 13474 522 13540 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 0 9540 254 10230 6 VSSA
port 208 nsew ground bidirectional
rlabel metal5 s 15746 11740 16000 13540 6 VSSA
port 208 nsew ground bidirectional
rlabel metal5 s 15746 9561 16000 10210 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 15746 12522 16000 12758 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 9418 13474 16000 13540 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 9418 11740 16000 11806 6 VSSA
port 208 nsew ground bidirectional
rlabel metal4 s 15746 9540 16000 10230 6 VSSA
port 208 nsew ground bidirectional
rlabel metal5 s 0 10530 254 11420 6 VSSD
port 209 nsew ground bidirectional
rlabel metal4 s 0 10510 254 11440 6 VSSD
port 209 nsew ground bidirectional
rlabel metal5 s 15746 10530 16000 11420 6 VSSD
port 209 nsew ground bidirectional
rlabel metal4 s 15746 10510 16000 11440 6 VSSD
port 209 nsew ground bidirectional
rlabel metal4 s 0 37350 254 42193 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal5 s 0 7380 254 8270 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal4 s 0 7360 254 8290 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal4 s 15746 37350 16000 42193 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal5 s 15746 7380 16000 8270 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal4 s 15746 7360 16000 8290 6 VSSIO
port 210 nsew ground bidirectional
rlabel metal5 s 0 13860 254 14710 6 VSSIO_Q
port 211 nsew ground bidirectional
rlabel metal4 s 0 13840 254 14730 6 VSSIO_Q
port 211 nsew ground bidirectional
rlabel metal5 s 15746 13860 16000 14710 6 VSSIO_Q
port 211 nsew ground bidirectional
rlabel metal4 s 15746 13840 16000 14730 6 VSSIO_Q
port 211 nsew ground bidirectional
rlabel metal5 s 0 8590 254 9240 6 VSWITCH
port 212 nsew power bidirectional
rlabel metal4 s 0 8570 254 9260 6 VSWITCH
port 212 nsew power bidirectional
rlabel metal5 s 15746 8590 16000 9240 6 VSWITCH
port 212 nsew power bidirectional
rlabel metal4 s 15746 8570 16000 9260 6 VSWITCH
port 212 nsew power bidirectional
rlabel metal2 s 2137 0 2193 480 6 VTRIP_SEL
port 213 nsew signal input
rlabel metal4 s 0 10218 33800 10814 6 AMUXBUS_A
port 214 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 214 nsew signal bidirectional
rlabel metal4 s 0 9266 33800 9862 6 AMUXBUS_B
port 215 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 215 nsew signal bidirectional
rlabel metal2 s 19478 -407 24258 4725 6 DRN_HVC
port 216 nsew power bidirectional
rlabel metal3 s 16978 -407 19178 1859 6 DRN_HVC
port 216 nsew power bidirectional
rlabel metal3 s 0 -407 14279 2730 6 P_CORE
port 217 nsew power bidirectional
rlabel metal3 s 19478 -407 33800 2730 6 P_CORE
port 217 nsew power bidirectional
rlabel metal5 s 10810 20617 22978 32782 6 P_PAD
port 218 nsew power bidirectional
rlabel metal2 s 9499 -407 14279 4 8 SRC_BDY_HVC
port 219 nsew ground bidirectional
rlabel metal3 s 14579 -407 16779 138 8 SRC_BDY_HVC
port 219 nsew ground bidirectional
rlabel metal5 s 25177 9140 33800 10940 6 VSSA
port 220 nsew ground bidirectional
rlabel metal5 s 25177 6960 33800 7610 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 25177 9922 33800 10158 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 10874 33800 10940 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 9140 33800 9206 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 25177 6940 33800 7630 6 VSSA
port 220 nsew ground bidirectional
rlabel metal5 s 0 9140 9448 10940 6 VSSA
port 220 nsew ground bidirectional
rlabel metal5 s 0 6960 9543 7610 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 9922 9448 10158 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 220 nsew ground bidirectional
rlabel metal4 s 0 6940 9543 7630 6 VSSA
port 220 nsew ground bidirectional
rlabel metal5 s 24241 2600 33800 3250 6 VDDA
port 221 nsew power bidirectional
rlabel metal4 s 24241 2580 33800 3270 6 VDDA
port 221 nsew power bidirectional
rlabel metal5 s 0 2600 9543 3250 6 VDDA
port 221 nsew power bidirectional
rlabel metal4 s 0 2580 9543 3270 6 VDDA
port 221 nsew power bidirectional
rlabel metal5 s 25177 5990 33800 6640 6 VSWITCH
port 222 nsew power bidirectional
rlabel metal4 s 25177 5970 33800 6660 6 VSWITCH
port 222 nsew power bidirectional
rlabel metal5 s 0 5990 9543 6640 6 VSWITCH
port 222 nsew power bidirectional
rlabel metal4 s 0 5970 9543 6660 6 VSWITCH
port 222 nsew power bidirectional
rlabel metal5 s 25177 12430 33800 13280 6 VDDIO_Q
port 223 nsew power bidirectional
rlabel metal4 s 25177 12410 33800 13300 6 VDDIO_Q
port 223 nsew power bidirectional
rlabel metal5 s 0 12430 9543 13280 6 VDDIO_Q
port 223 nsew power bidirectional
rlabel metal4 s 0 12410 9543 13300 6 VDDIO_Q
port 223 nsew power bidirectional
rlabel metal5 s 25177 20 33800 1070 6 VCCHIB
port 224 nsew power bidirectional
rlabel metal4 s 25177 0 33800 1090 6 VCCHIB
port 224 nsew power bidirectional
rlabel metal5 s 0 20 9543 1070 6 VCCHIB
port 224 nsew power bidirectional
rlabel metal4 s 0 0 9543 1090 6 VCCHIB
port 224 nsew power bidirectional
rlabel metal5 s 25177 13600 33800 18590 6 VDDIO
port 225 nsew power bidirectional
rlabel metal5 s 25177 3570 33800 4460 6 VDDIO
port 225 nsew power bidirectional
rlabel metal4 s 24241 3550 33800 4480 6 VDDIO
port 225 nsew power bidirectional
rlabel metal4 s 25177 13600 33800 18593 6 VDDIO
port 225 nsew power bidirectional
rlabel metal5 s 0 13600 9543 18590 6 VDDIO
port 225 nsew power bidirectional
rlabel metal5 s 0 3570 9543 4460 6 VDDIO
port 225 nsew power bidirectional
rlabel metal4 s 0 3550 9543 4480 6 VDDIO
port 225 nsew power bidirectional
rlabel metal4 s 0 13600 9543 18593 6 VDDIO
port 225 nsew power bidirectional
rlabel metal5 s 25177 1390 33800 2280 6 VCCD
port 226 nsew power bidirectional
rlabel metal4 s 25177 1370 33800 2300 6 VCCD
port 226 nsew power bidirectional
rlabel metal5 s 0 1390 9543 2280 6 VCCD
port 226 nsew power bidirectional
rlabel metal4 s 0 1370 9543 2300 6 VCCD
port 226 nsew power bidirectional
rlabel metal4 s 25649 34750 33800 39593 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 33672 37913 33674 37915 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal5 s 25177 4780 33800 5670 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 25177 4760 33800 5690 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 33546 34750 33800 39593 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 0 34750 9641 39593 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal5 s 0 4780 9543 5670 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal4 s 0 4760 9543 5690 6 VSSIO
port 227 nsew ground bidirectional
rlabel metal5 s 25177 7930 33800 8820 6 VSSD
port 228 nsew ground bidirectional
rlabel metal4 s 25177 7910 33800 8840 6 VSSD
port 228 nsew ground bidirectional
rlabel metal5 s 0 7930 9543 8820 6 VSSD
port 228 nsew ground bidirectional
rlabel metal4 s 0 7910 9450 8840 6 VSSD
port 228 nsew ground bidirectional
rlabel metal5 s 25177 11260 33800 12110 6 VSSIO_Q
port 229 nsew ground bidirectional
rlabel metal4 s 25177 11240 33800 12130 6 VSSIO_Q
port 229 nsew ground bidirectional
rlabel metal5 s 0 11260 9543 12110 6 VSSIO_Q
port 229 nsew ground bidirectional
rlabel metal4 s 0 11240 9543 12130 6 VSSIO_Q
port 229 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 230 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 230 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 231 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 231 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 232 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 1859 6 DRN_HVC
port 232 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 233 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 138 8 SRC_BDY_HVC
port 233 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VCCD_PAD
port 234 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 235 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 235 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 235 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 235 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 235 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 236 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 236 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 236 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 236 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 237 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 237 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 237 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 237 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 238 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 238 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 238 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 238 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 239 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 239 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 239 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 239 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 240 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 240 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 240 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 240 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 240 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 240 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 240 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 240 nsew power bidirectional
rlabel metal3 s 10078 -407 14858 1373 6 VCCD
port 241 nsew power bidirectional
rlabel metal3 s 99 -407 4879 1373 6 VCCD
port 241 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 241 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 241 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 241 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 241 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 242 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 243 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 243 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 243 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 243 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 244 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 244 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 244 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 244 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 245 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 245 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 246 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 246 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VCCD_PAD
port 247 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 248 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 248 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 248 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 248 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 248 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 249 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 249 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 249 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 249 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 250 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 250 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 250 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 250 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 251 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 251 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 251 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 251 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 252 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 252 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 252 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 252 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 253 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 253 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 253 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 253 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 253 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 253 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 253 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 253 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 1373 6 VCCD
port 254 nsew power bidirectional
rlabel metal3 s 100 -7 4900 1373 6 VCCD
port 254 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 254 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 254 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 254 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 254 nsew power bidirectional
rlabel metal4 s 14845 34750 15294 39586 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 255 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 256 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 256 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 256 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 256 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 257 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 257 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 257 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 257 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 258 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 259 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VCCD_PAD
port 260 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 261 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 261 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 261 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 261 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 261 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 262 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 262 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 262 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 262 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 263 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 263 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 263 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 263 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 264 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 264 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 264 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 264 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 265 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 265 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 265 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 265 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 266 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 266 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 266 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 266 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 266 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 266 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 266 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 266 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 267 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 267 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 267 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 267 nsew power bidirectional
rlabel metal4 s 14845 34750 15294 39593 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 268 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 269 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 269 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 269 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 269 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 270 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 270 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 270 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 270 nsew ground bidirectional
rlabel metal3 s 100 -1566 4900 9469 6 VCCD1
port 271 nsew power bidirectional
rlabel metal3 s 10151 -1542 14940 16886 6 VCCD1
port 271 nsew power bidirectional
rlabel metal3 s 5190 -1506 9852 -502 8 VSSD1
port 272 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 273 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 273 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 274 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 274 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VCCD_PAD
port 275 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 276 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 276 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 276 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 276 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 276 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 277 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 277 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 277 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 277 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 278 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 278 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 278 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 278 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 279 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 279 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 279 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 279 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 280 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 280 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 280 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 280 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 281 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 281 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 281 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 281 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 281 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 281 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 281 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 281 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 1373 6 VCCD
port 282 nsew power bidirectional
rlabel metal3 s 100 -7 4900 1373 6 VCCD
port 282 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 282 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 282 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 282 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 282 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal4 s 0 34750 141 39593 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 283 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 284 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 284 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 284 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 284 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 285 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 285 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 285 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 285 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 286 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 286 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 287 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 287 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 288 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 289 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 290 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 291 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 292 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VCCD_PAD
port 293 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 294 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 294 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 294 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 294 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 294 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 295 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 295 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 295 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 295 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 296 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 296 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 296 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 296 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 297 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 297 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 297 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 297 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 298 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 298 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 298 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 298 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 299 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 299 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 299 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 299 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 299 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 299 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 299 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 299 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 1373 6 VCCD
port 300 nsew power bidirectional
rlabel metal3 s 100 -7 4900 1373 6 VCCD
port 300 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 300 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 300 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 300 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 300 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 301 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 302 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 302 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 302 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 302 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 303 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 303 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 303 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 303 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 304 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 304 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 305 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 305 nsew signal bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VDDA_PAD
port 306 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 307 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 307 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 307 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 307 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 307 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 2585 6 VDDA
port 308 nsew power bidirectional
rlabel metal3 s 99 -407 4879 2585 6 VDDA
port 308 nsew power bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 308 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 308 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 308 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 308 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 309 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 309 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 309 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 309 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 310 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 310 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 310 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 310 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 311 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 311 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 311 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 311 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 312 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 312 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 312 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 312 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 312 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 312 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 312 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 312 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 313 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 313 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 313 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 313 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 14872 37913 14874 37915 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 314 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 315 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 315 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 315 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 315 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 316 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 316 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 316 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 316 nsew ground bidirectional
rlabel metal4 s 14746 10218 15000 10814 6 AMUXBUS_A
port 317 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 317 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9922 6 AMUXBUS_B
port 318 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 318 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 319 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 1859 6 DRN_HVC
port 319 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 320 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 138 8 SRC_BDY_HVC
port 320 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VDDA_PAD
port 321 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 322 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 322 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 322 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 0 10814 15000 11214 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 14746 9140 15000 9206 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 322 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 322 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 2985 6 VDDA
port 323 nsew power bidirectional
rlabel metal3 s 99 -407 4879 2985 6 VDDA
port 323 nsew power bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 323 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 323 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 323 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 323 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 324 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 324 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 324 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 324 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 325 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 325 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 325 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 325 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 326 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 326 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 326 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 326 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 327 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 327 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 327 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 327 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 327 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 327 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 327 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 327 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 328 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 328 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 328 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 328 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39993 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39993 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 14872 37913 14874 37915 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 329 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 330 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 330 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 330 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 330 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 331 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 331 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 331 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 331 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 332 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 332 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 333 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 333 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 334 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 335 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 336 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 337 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 338 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VDDA_PAD
port 339 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 340 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 340 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 340 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 340 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 340 nsew ground bidirectional
rlabel metal3 s 10151 -7 14940 2585 6 VDDA
port 341 nsew power bidirectional
rlabel metal3 s 100 -7 4900 2585 6 VDDA
port 341 nsew power bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 341 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 341 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 341 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 341 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 342 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 342 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 342 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 342 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 343 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 343 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 343 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 343 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 344 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 344 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 344 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 344 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 345 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 345 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 345 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 345 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 345 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 345 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 345 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 345 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 346 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 346 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 346 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 346 nsew power bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 347 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 348 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 348 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 348 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 348 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 349 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 349 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 349 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 349 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 350 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 350 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 351 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 351 nsew signal bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VDDIO_PAD
port 352 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 353 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 353 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 353 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 353 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 353 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 354 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 354 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 354 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 354 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 355 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 355 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 355 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 355 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 356 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 356 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 356 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 356 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 357 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 357 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 357 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 357 nsew power bidirectional
rlabel metal3 s 10078 -407 14858 3553 6 VDDIO
port 358 nsew power bidirectional
rlabel metal3 s 99 -407 4879 3553 6 VDDIO
port 358 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 358 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 358 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 358 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 358 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 358 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 358 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 358 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 358 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 359 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 359 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 359 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 359 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 360 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 361 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 361 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 361 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 361 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 362 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 362 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 362 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 362 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 363 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 363 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 364 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 364 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 365 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 1859 6 DRN_HVC
port 365 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 366 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 138 8 SRC_BDY_HVC
port 366 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VDDIO_PAD
port 367 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 368 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 368 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 368 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 368 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 368 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 369 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 369 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 369 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 369 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 370 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 370 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 370 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 370 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 371 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 371 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 371 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 371 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 372 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 372 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 372 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 372 nsew power bidirectional
rlabel metal3 s 10078 -407 14858 3553 6 VDDIO
port 373 nsew power bidirectional
rlabel metal3 s 99 -407 4879 3553 6 VDDIO
port 373 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 373 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 373 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 373 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 373 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 373 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 373 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 373 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 373 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 374 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 374 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 374 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 374 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 375 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 376 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 376 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 376 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 376 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 377 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 377 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 377 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 377 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 378 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 378 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 379 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 379 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 380 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 381 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 382 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 383 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 384 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VDDIO_PAD
port 385 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 386 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 386 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 386 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 386 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 386 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 387 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 387 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 387 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 387 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 388 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 388 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 388 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 388 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 389 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 389 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 389 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 389 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 390 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 390 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 390 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 390 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 3553 6 VDDIO
port 391 nsew power bidirectional
rlabel metal3 s 100 -7 4900 3553 6 VDDIO
port 391 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 391 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 391 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 391 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 391 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 391 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 391 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 391 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 391 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 392 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 392 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 392 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 392 nsew power bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 393 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 394 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 394 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 394 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 394 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 395 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 395 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 395 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 395 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 396 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 396 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 397 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 397 nsew signal bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VSSA_PAD
port 398 nsew ground bidirectional
rlabel metal3 s 99 -407 4879 6096 6 VSSA
port 399 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 6945 6 VSSA
port 399 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 399 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 399 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 399 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 14746 10874 15000 10940 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 14746 9140 15000 9206 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 399 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 399 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 400 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 400 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 400 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 400 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 401 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 401 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 401 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 401 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 402 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 402 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 402 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 402 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 403 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 403 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 403 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 403 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 404 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 404 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 404 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 404 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 404 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 404 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 404 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 404 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 405 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 405 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 405 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 405 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 406 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 407 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 407 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 407 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 407 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 408 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 408 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 408 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 408 nsew ground bidirectional
rlabel metal4 s 14872 37913 14874 37915 6 VSSIO
port 409 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 410 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 410 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 411 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 411 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 412 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 2069 6 DRN_HVC
port 412 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 413 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 2078 6 SRC_BDY_HVC
port 413 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VSSA_PAD
port 414 nsew ground bidirectional
rlabel metal3 s 99 -407 4879 6096 6 VSSA
port 415 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 6945 6 VSSA
port 415 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 415 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 415 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 415 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 14746 10874 15000 10940 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 14746 9140 15000 9206 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 415 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 415 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 416 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 416 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 416 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 416 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 417 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 417 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 417 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 417 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 418 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 418 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 418 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 418 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 419 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 419 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 419 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 419 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 420 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 420 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 420 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 420 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 420 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 420 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 420 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 420 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 421 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 421 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 421 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 421 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 422 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 423 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 423 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 423 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 423 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 424 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 424 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 424 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 424 nsew ground bidirectional
rlabel metal4 s 14872 37913 14874 37915 6 VSSIO
port 425 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 426 nsew signal bidirectional
rlabel metal4 s 14746 10218 15000 10814 6 AMUXBUS_A
port 426 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 427 nsew signal bidirectional
rlabel metal4 s 14746 9266 15000 9862 6 AMUXBUS_B
port 427 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 428 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 429 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 430 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 431 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 432 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSA_PAD
port 433 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 14746 9140 15000 9206 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 14746 10874 15000 10940 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 434 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 434 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 434 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 434 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 434 nsew ground bidirectional
rlabel metal3 s 100 -7 4900 6945 6 VSSA
port 434 nsew ground bidirectional
rlabel metal3 s 10151 -7 14940 6945 6 VSSA
port 434 nsew ground bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 435 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 435 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 435 nsew power bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 435 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 436 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 436 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 436 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 436 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 437 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 437 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 437 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 437 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 438 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 438 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 438 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 438 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 439 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 439 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 439 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 439 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 439 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 439 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 439 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 439 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 440 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 440 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 440 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 440 nsew power bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 441 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 442 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 442 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 442 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 442 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 443 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 443 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 443 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 443 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 444 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 444 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 445 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 445 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 446 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 2069 6 DRN_HVC
port 446 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 447 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 2078 6 SRC_BDY_HVC
port 447 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VSSD_PAD
port 448 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 449 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 449 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 449 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 449 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 449 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 450 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 450 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 450 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 450 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 451 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 451 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 451 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 451 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 452 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 452 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 452 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 452 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 453 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 453 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 453 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 453 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 454 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 454 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 454 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 454 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 454 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 454 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 454 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 454 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 455 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 455 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 455 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 455 nsew power bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 456 nsew ground bidirectional
rlabel metal3 s 99 -407 4879 6096 6 VSSD
port 457 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 7913 6 VSSD
port 457 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 457 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 457 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 457 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 457 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 458 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 458 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 458 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 458 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 459 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 459 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 460 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 460 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSD_PAD
port 461 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 462 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 462 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 462 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 462 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 462 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 463 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 463 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 463 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 463 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 464 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 464 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 464 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 464 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 465 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 465 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 465 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 465 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 466 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 466 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 466 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 466 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 467 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 467 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 467 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 467 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 467 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 467 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 467 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 467 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 468 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 468 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 468 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 468 nsew power bidirectional
rlabel metal4 s 14845 34750 15294 39586 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 469 nsew ground bidirectional
rlabel metal3 s 10151 -7 14940 7913 6 VSSD
port 470 nsew ground bidirectional
rlabel metal3 s 100 -7 4900 7913 6 VSSD
port 470 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 470 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 470 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 470 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 470 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 471 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 471 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 471 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 471 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 472 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 473 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSD_PAD
port 474 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 475 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 475 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 475 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 475 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 475 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 476 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 476 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 476 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 476 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 477 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 477 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 477 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 477 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 478 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 478 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 478 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 478 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 479 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 479 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 479 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 479 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 480 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 480 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 480 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 480 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 480 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 480 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 480 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 480 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 481 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 481 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 481 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 481 nsew power bidirectional
rlabel metal4 s 14845 34750 15294 39593 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 482 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 483 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 483 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 483 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 483 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 484 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 484 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 484 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 484 nsew ground bidirectional
rlabel metal3 s 100 -1896 4900 5280 6 VSSD1
port 485 nsew ground bidirectional
rlabel metal3 s 10151 -1902 14940 5424 6 VSSD1
port 485 nsew ground bidirectional
rlabel metal3 s 5200 -1898 9851 -458 8 VCCD1
port 486 nsew power bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 487 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 487 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 488 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 488 nsew signal bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSD_PAD
port 489 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 490 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 490 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 490 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 490 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 490 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 491 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 491 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 491 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 491 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 492 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 492 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 492 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 492 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 493 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 493 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 493 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 493 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 494 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 494 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 494 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 494 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 495 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 495 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 495 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 495 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 495 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 495 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 495 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 495 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 496 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 496 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 496 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 496 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal4 s 0 34750 141 39593 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 497 nsew ground bidirectional
rlabel metal3 s 10151 -7 14940 7913 6 VSSD
port 498 nsew ground bidirectional
rlabel metal3 s 100 -7 4900 7913 6 VSSD
port 498 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 498 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 498 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 498 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 498 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 499 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 499 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 499 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 499 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 500 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 500 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 501 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 501 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 502 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 503 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 504 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 505 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 506 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSD_PAD
port 507 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 508 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 508 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 508 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 508 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 508 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 509 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 509 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 509 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 509 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 510 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 510 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 510 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 510 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 511 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 511 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 511 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 511 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 512 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 512 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 512 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 512 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 513 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 513 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 513 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 513 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 513 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 513 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 513 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 513 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 514 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 514 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 514 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 514 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39593 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39593 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 515 nsew ground bidirectional
rlabel metal3 s 10151 -7 14940 7913 6 VSSD
port 516 nsew ground bidirectional
rlabel metal3 s 100 -7 4900 7913 6 VSSD
port 516 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 516 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 516 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 516 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 516 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 517 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 517 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 517 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 517 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 518 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 518 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 519 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 519 nsew signal bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VSSIO_PAD
port 520 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 521 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 521 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 521 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 521 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 521 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 522 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 522 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 522 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 522 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 523 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 523 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 523 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 523 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 524 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 524 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 524 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 524 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 525 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 525 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 525 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 525 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 526 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 526 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 526 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 526 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 526 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 526 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 526 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 526 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 527 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 527 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 527 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 527 nsew power bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal4 s 14850 34750 15000 39593 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal3 s 99 -407 4879 4763 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 4763 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 528 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 529 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 529 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 529 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 529 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 530 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 530 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 530 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 530 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 531 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 531 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 532 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 532 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 533 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 2069 6 DRN_HVC
port 533 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 534 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 2078 6 SRC_BDY_HVC
port 534 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VSSIO_PAD
port 535 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 536 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 536 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 536 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 536 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 536 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 537 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 537 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 537 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 537 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 538 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 538 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 538 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 538 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 539 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 539 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 539 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 539 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 540 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 540 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 540 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 540 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 541 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 541 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 541 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 541 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 541 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 541 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 541 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 541 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 542 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 542 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 542 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 542 nsew power bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal4 s 14850 34750 15000 39593 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal3 s 99 -407 4879 4763 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 4763 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 543 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 544 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 544 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 544 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 544 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 545 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 545 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 545 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 545 nsew ground bidirectional
rlabel metal4 s 0 10218 15000 10814 6 AMUXBUS_A
port 546 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 546 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9862 6 AMUXBUS_B
port 547 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 547 nsew signal bidirectional
rlabel metal3 s 5200 -7 7376 4037 6 DRN_LVC1
port 548 nsew power bidirectional
rlabel metal3 s 7676 -7 9851 4573 6 DRN_LVC2
port 549 nsew power bidirectional
rlabel metal2 s 100 -7 4099 290 6 SRC_BDY_LVC1
port 550 nsew ground bidirectional
rlabel metal2 s 10943 -7 14940 725 6 SRC_BDY_LVC2
port 551 nsew ground bidirectional
rlabel metal2 s 6888 -7 8888 58 6 BDY2_B2B
port 552 nsew ground bidirectional
rlabel metal5 s 2054 19973 12934 33426 6 VSSIO_PAD
port 553 nsew ground bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 554 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 554 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 554 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 10874 15000 10940 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 9140 15000 9206 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 554 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 554 nsew ground bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 555 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 555 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 555 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 555 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 556 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 556 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 556 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 556 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 557 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 557 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 557 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 557 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 558 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 558 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 558 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 558 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 559 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 559 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 559 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 559 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 559 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 559 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 559 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 559 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 560 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 560 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 560 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 560 nsew power bidirectional
rlabel metal3 s 10151 -7 14940 4763 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal3 s 100 -7 4900 4763 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 561 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 562 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 562 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 562 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 562 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 563 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 563 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 563 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 563 nsew ground bidirectional
rlabel metal1 s 703 1791 852 2359 6 GATE
port 564 nsew
rlabel viali s 797 1813 831 1847 6 GATE
port 564 nsew
rlabel viali s 725 1813 759 1847 6 GATE
port 564 nsew
rlabel locali s 662 1785 927 1867 6 GATE
port 564 nsew
rlabel metal1 s 1070 66 1383 69 6 NWELLRING
port 565 nsew
rlabel metal1 s 66 66 203 69 6 NWELLRING
port 565 nsew
rlabel metal1 s 1070 69 1386 206 6 NWELLRING
port 565 nsew
rlabel metal1 s 1385 206 1386 208 6 NWELLRING
port 565 nsew
rlabel metal1 s 1385 208 1525 2124 6 NWELLRING
port 565 nsew
rlabel metal1 s 1383 2124 1525 2136 6 NWELLRING
port 565 nsew
rlabel metal1 s 1371 2136 1525 2216 6 NWELLRING
port 565 nsew
rlabel metal1 s 66 69 206 2216 6 NWELLRING
port 565 nsew
rlabel metal1 s 1291 2216 1383 2218 6 NWELLRING
port 565 nsew
rlabel metal1 s 208 2216 286 2218 6 NWELLRING
port 565 nsew
rlabel metal1 s 886 2218 1383 2358 6 NWELLRING
port 565 nsew
rlabel metal1 s 208 2218 669 2358 6 NWELLRING
port 565 nsew
rlabel viali s 1262 108 1296 142 6 NWELLRING
port 565 nsew
rlabel viali s 1190 108 1224 142 6 NWELLRING
port 565 nsew
rlabel viali s 1118 108 1152 142 6 NWELLRING
port 565 nsew
rlabel viali s 1438 273 1472 307 6 NWELLRING
port 565 nsew
rlabel viali s 1438 345 1472 379 6 NWELLRING
port 565 nsew
rlabel viali s 1438 417 1472 451 6 NWELLRING
port 565 nsew
rlabel viali s 1438 489 1472 523 6 NWELLRING
port 565 nsew
rlabel viali s 1438 561 1472 595 6 NWELLRING
port 565 nsew
rlabel viali s 1438 633 1472 667 6 NWELLRING
port 565 nsew
rlabel viali s 1438 705 1472 739 6 NWELLRING
port 565 nsew
rlabel viali s 1438 777 1472 811 6 NWELLRING
port 565 nsew
rlabel viali s 1438 849 1472 883 6 NWELLRING
port 565 nsew
rlabel viali s 1438 921 1472 955 6 NWELLRING
port 565 nsew
rlabel viali s 1438 993 1472 1027 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1065 1472 1099 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1137 1472 1171 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1209 1472 1243 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1281 1472 1315 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1353 1472 1387 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1425 1472 1459 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1497 1472 1531 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1569 1472 1603 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1641 1472 1675 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1713 1472 1747 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1785 1472 1819 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1857 1472 1891 6 NWELLRING
port 565 nsew
rlabel viali s 1438 1929 1472 1963 6 NWELLRING
port 565 nsew
rlabel viali s 1438 2001 1472 2035 6 NWELLRING
port 565 nsew
rlabel viali s 119 273 153 307 6 NWELLRING
port 565 nsew
rlabel viali s 119 345 153 379 6 NWELLRING
port 565 nsew
rlabel viali s 119 417 153 451 6 NWELLRING
port 565 nsew
rlabel viali s 119 489 153 523 6 NWELLRING
port 565 nsew
rlabel viali s 119 561 153 595 6 NWELLRING
port 565 nsew
rlabel viali s 119 633 153 667 6 NWELLRING
port 565 nsew
rlabel viali s 119 705 153 739 6 NWELLRING
port 565 nsew
rlabel viali s 119 777 153 811 6 NWELLRING
port 565 nsew
rlabel viali s 119 849 153 883 6 NWELLRING
port 565 nsew
rlabel viali s 119 921 153 955 6 NWELLRING
port 565 nsew
rlabel viali s 119 993 153 1027 6 NWELLRING
port 565 nsew
rlabel viali s 119 1065 153 1099 6 NWELLRING
port 565 nsew
rlabel viali s 119 1137 153 1171 6 NWELLRING
port 565 nsew
rlabel viali s 119 1209 153 1243 6 NWELLRING
port 565 nsew
rlabel viali s 119 1281 153 1315 6 NWELLRING
port 565 nsew
rlabel viali s 119 1353 153 1387 6 NWELLRING
port 565 nsew
rlabel viali s 119 1425 153 1459 6 NWELLRING
port 565 nsew
rlabel viali s 119 1497 153 1531 6 NWELLRING
port 565 nsew
rlabel viali s 119 1569 153 1603 6 NWELLRING
port 565 nsew
rlabel viali s 119 1641 153 1675 6 NWELLRING
port 565 nsew
rlabel viali s 119 1713 153 1747 6 NWELLRING
port 565 nsew
rlabel viali s 119 1785 153 1819 6 NWELLRING
port 565 nsew
rlabel viali s 119 1857 153 1891 6 NWELLRING
port 565 nsew
rlabel viali s 119 1929 153 1963 6 NWELLRING
port 565 nsew
rlabel viali s 119 2001 153 2035 6 NWELLRING
port 565 nsew
rlabel viali s 1247 2271 1281 2305 6 NWELLRING
port 565 nsew
rlabel viali s 1175 2271 1209 2305 6 NWELLRING
port 565 nsew
rlabel viali s 1103 2271 1137 2305 6 NWELLRING
port 565 nsew
rlabel viali s 1031 2271 1065 2305 6 NWELLRING
port 565 nsew
rlabel viali s 959 2271 993 2305 6 NWELLRING
port 565 nsew
rlabel viali s 595 2271 629 2305 6 NWELLRING
port 565 nsew
rlabel viali s 523 2271 557 2305 6 NWELLRING
port 565 nsew
rlabel viali s 451 2271 485 2305 6 NWELLRING
port 565 nsew
rlabel viali s 379 2271 413 2305 6 NWELLRING
port 565 nsew
rlabel viali s 307 2271 341 2305 6 NWELLRING
port 565 nsew
rlabel locali s 66 66 1525 206 6 NWELLRING
port 565 nsew
rlabel locali s 1385 206 1525 2218 6 NWELLRING
port 565 nsew
rlabel locali s 66 206 206 2218 6 NWELLRING
port 565 nsew
rlabel locali s 66 2218 1525 2358 6 NWELLRING
port 565 nsew
rlabel nwell s 0 0 1591 272 6 NWELLRING
port 565 nsew
rlabel nwell s 1319 272 1591 2152 6 NWELLRING
port 565 nsew
rlabel nwell s 0 272 272 2152 6 NWELLRING
port 565 nsew
rlabel nwell s 0 2152 1591 2424 6 NWELLRING
port 565 nsew
rlabel metal1 s 572 66 772 1709 6 VGND
port 566 nsew ground default
rlabel viali s 621 757 655 791 6 VGND
port 566 nsew ground default
rlabel viali s 621 829 655 863 6 VGND
port 566 nsew ground default
rlabel viali s 621 901 655 935 6 VGND
port 566 nsew ground default
rlabel viali s 621 973 655 1007 6 VGND
port 566 nsew ground default
rlabel viali s 621 1045 655 1079 6 VGND
port 566 nsew ground default
rlabel viali s 621 1117 655 1151 6 VGND
port 566 nsew ground default
rlabel viali s 621 1189 655 1223 6 VGND
port 566 nsew ground default
rlabel viali s 621 1261 655 1295 6 VGND
port 566 nsew ground default
rlabel viali s 621 1333 655 1367 6 VGND
port 566 nsew ground default
rlabel viali s 621 1405 655 1439 6 VGND
port 566 nsew ground default
rlabel viali s 621 1477 655 1511 6 VGND
port 566 nsew ground default
rlabel viali s 621 1549 655 1583 6 VGND
port 566 nsew ground default
rlabel locali s 593 672 701 1751 6 VGND
port 566 nsew ground default
rlabel metal1 s 358 66 533 69 6 NBODY
port 567 nsew
rlabel metal1 s 1093 358 1233 1826 6 NBODY
port 567 nsew
rlabel metal1 s 1087 1826 1233 1901 6 NBODY
port 567 nsew
rlabel metal1 s 358 69 536 1901 6 NBODY
port 567 nsew
rlabel metal1 s 886 1901 1233 2000 6 NBODY
port 567 nsew
rlabel metal1 s 886 2000 1167 2066 6 NBODY
port 567 nsew
rlabel metal1 s 358 1901 669 2000 6 NBODY
port 567 nsew
rlabel metal1 s 424 2000 669 2066 6 NBODY
port 567 nsew
rlabel viali s 1146 401 1180 435 6 NBODY
port 567 nsew
rlabel viali s 395 401 429 435 6 NBODY
port 567 nsew
rlabel viali s 1146 473 1180 507 6 NBODY
port 567 nsew
rlabel viali s 1146 545 1180 579 6 NBODY
port 567 nsew
rlabel viali s 1146 617 1180 651 6 NBODY
port 567 nsew
rlabel viali s 1146 689 1180 723 6 NBODY
port 567 nsew
rlabel viali s 1146 761 1180 795 6 NBODY
port 567 nsew
rlabel viali s 1146 833 1180 867 6 NBODY
port 567 nsew
rlabel viali s 1146 905 1180 939 6 NBODY
port 567 nsew
rlabel viali s 1146 977 1180 1011 6 NBODY
port 567 nsew
rlabel viali s 1146 1049 1180 1083 6 NBODY
port 567 nsew
rlabel viali s 1146 1121 1180 1155 6 NBODY
port 567 nsew
rlabel viali s 1146 1193 1180 1227 6 NBODY
port 567 nsew
rlabel viali s 1146 1265 1180 1299 6 NBODY
port 567 nsew
rlabel viali s 1146 1337 1180 1371 6 NBODY
port 567 nsew
rlabel viali s 1146 1409 1180 1443 6 NBODY
port 567 nsew
rlabel viali s 1146 1481 1180 1515 6 NBODY
port 567 nsew
rlabel viali s 1146 1553 1180 1587 6 NBODY
port 567 nsew
rlabel viali s 1146 1625 1180 1659 6 NBODY
port 567 nsew
rlabel viali s 1146 1697 1180 1731 6 NBODY
port 567 nsew
rlabel viali s 1146 1769 1180 1803 6 NBODY
port 567 nsew
rlabel viali s 395 473 429 507 6 NBODY
port 567 nsew
rlabel viali s 395 545 429 579 6 NBODY
port 567 nsew
rlabel viali s 395 617 429 651 6 NBODY
port 567 nsew
rlabel viali s 395 689 429 723 6 NBODY
port 567 nsew
rlabel viali s 395 761 429 795 6 NBODY
port 567 nsew
rlabel viali s 395 833 429 867 6 NBODY
port 567 nsew
rlabel viali s 395 905 429 939 6 NBODY
port 567 nsew
rlabel viali s 395 977 429 1011 6 NBODY
port 567 nsew
rlabel viali s 395 1049 429 1083 6 NBODY
port 567 nsew
rlabel viali s 395 1121 429 1155 6 NBODY
port 567 nsew
rlabel viali s 395 1193 429 1227 6 NBODY
port 567 nsew
rlabel viali s 395 1265 429 1299 6 NBODY
port 567 nsew
rlabel viali s 395 1337 429 1371 6 NBODY
port 567 nsew
rlabel viali s 395 1409 429 1443 6 NBODY
port 567 nsew
rlabel viali s 395 1481 429 1515 6 NBODY
port 567 nsew
rlabel viali s 395 1553 429 1587 6 NBODY
port 567 nsew
rlabel viali s 395 1625 429 1659 6 NBODY
port 567 nsew
rlabel viali s 395 1697 429 1731 6 NBODY
port 567 nsew
rlabel viali s 395 1769 429 1803 6 NBODY
port 567 nsew
rlabel viali s 1072 1969 1106 2003 6 NBODY
port 567 nsew
rlabel viali s 1000 1969 1034 2003 6 NBODY
port 567 nsew
rlabel viali s 928 1969 962 2003 6 NBODY
port 567 nsew
rlabel viali s 598 1969 632 2003 6 NBODY
port 567 nsew
rlabel viali s 526 1969 560 2003 6 NBODY
port 567 nsew
rlabel viali s 454 1969 488 2003 6 NBODY
port 567 nsew
rlabel locali s 358 358 1233 498 6 NBODY
port 567 nsew
rlabel locali s 1093 498 1233 1924 6 NBODY
port 567 nsew
rlabel locali s 358 498 498 1924 6 NBODY
port 567 nsew
rlabel locali s 358 1924 1233 2066 6 NBODY
port 567 nsew
rlabel pwell s 332 332 1259 2092 6 NBODY
port 567 nsew
rlabel metal1 s 831 66 1031 1752 6 IN
port 568 nsew
rlabel viali s 915 757 949 791 6 IN
port 568 nsew
rlabel viali s 915 829 949 863 6 IN
port 568 nsew
rlabel viali s 915 901 949 935 6 IN
port 568 nsew
rlabel viali s 915 973 949 1007 6 IN
port 568 nsew
rlabel viali s 915 1045 949 1079 6 IN
port 568 nsew
rlabel viali s 915 1117 949 1151 6 IN
port 568 nsew
rlabel viali s 915 1189 949 1223 6 IN
port 568 nsew
rlabel viali s 915 1261 949 1295 6 IN
port 568 nsew
rlabel viali s 915 1333 949 1367 6 IN
port 568 nsew
rlabel viali s 915 1405 949 1439 6 IN
port 568 nsew
rlabel viali s 915 1477 949 1511 6 IN
port 568 nsew
rlabel viali s 915 1549 949 1583 6 IN
port 568 nsew
rlabel locali s 888 672 996 1751 6 IN
port 568 nsew
<< properties >>
string FIXED_BBOX 0 0 1591 2424
string LEFclass PAD
string LEFview TRUE
string GDS_END 4186318
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 4173684
<< end >>
