magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1165 157 1347 201
rect 1650 157 2205 203
rect 1 145 817 157
rect 1019 145 2205 157
rect 1 21 2205 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 453 47 483 131
rect 531 47 561 131
rect 627 47 657 131
rect 703 47 733 131
rect 901 47 931 119
rect 997 47 1027 119
rect 1095 47 1125 131
rect 1241 47 1271 175
rect 1342 47 1372 119
rect 1445 47 1475 119
rect 1540 47 1570 131
rect 1728 47 1758 177
rect 1812 47 1842 177
rect 2000 47 2030 131
rect 2097 47 2127 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 526 369 556 497
rect 610 369 640 497
rect 703 369 733 497
rect 900 413 930 497
rect 993 413 1023 497
rect 1089 413 1119 497
rect 1221 347 1251 497
rect 1316 413 1346 497
rect 1400 413 1430 497
rect 1517 413 1547 497
rect 1728 297 1758 497
rect 1812 297 1842 497
rect 2000 369 2030 497
rect 2097 297 2127 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 101 351 131
rect 299 67 307 101
rect 341 67 351 101
rect 299 47 351 67
rect 381 89 453 131
rect 381 55 407 89
rect 441 55 453 89
rect 381 47 453 55
rect 483 47 531 131
rect 561 89 627 131
rect 561 55 582 89
rect 616 55 627 89
rect 561 47 627 55
rect 657 47 703 131
rect 733 93 791 131
rect 1191 131 1241 175
rect 1045 119 1095 131
rect 733 59 749 93
rect 783 59 791 93
rect 733 47 791 59
rect 845 107 901 119
rect 845 73 853 107
rect 887 73 901 107
rect 845 47 901 73
rect 931 107 997 119
rect 931 73 953 107
rect 987 73 997 107
rect 931 47 997 73
rect 1027 47 1095 119
rect 1125 101 1241 131
rect 1125 67 1169 101
rect 1203 67 1241 101
rect 1125 47 1241 67
rect 1271 119 1321 175
rect 1676 162 1728 177
rect 1490 119 1540 131
rect 1271 107 1342 119
rect 1271 73 1287 107
rect 1321 73 1342 107
rect 1271 47 1342 73
rect 1372 107 1445 119
rect 1372 73 1399 107
rect 1433 73 1445 107
rect 1372 47 1445 73
rect 1475 47 1540 119
rect 1570 107 1622 131
rect 1570 73 1580 107
rect 1614 73 1622 107
rect 1570 47 1622 73
rect 1676 128 1684 162
rect 1718 128 1728 162
rect 1676 94 1728 128
rect 1676 60 1684 94
rect 1718 60 1728 94
rect 1676 47 1728 60
rect 1758 123 1812 177
rect 1758 89 1768 123
rect 1802 89 1812 123
rect 1758 47 1812 89
rect 1842 164 1894 177
rect 1842 130 1852 164
rect 1886 130 1894 164
rect 2045 161 2097 177
rect 2045 131 2053 161
rect 1842 96 1894 130
rect 1842 62 1852 96
rect 1886 62 1894 96
rect 1842 47 1894 62
rect 1948 119 2000 131
rect 1948 85 1956 119
rect 1990 85 2000 119
rect 1948 47 2000 85
rect 2030 127 2053 131
rect 2087 127 2097 161
rect 2030 93 2097 127
rect 2030 59 2053 93
rect 2087 59 2097 93
rect 2030 47 2097 59
rect 2127 143 2179 177
rect 2127 109 2137 143
rect 2171 109 2179 143
rect 2127 47 2179 109
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 452 351 497
rect 299 418 307 452
rect 341 418 351 452
rect 299 369 351 418
rect 381 483 435 497
rect 381 449 391 483
rect 425 449 435 483
rect 381 369 435 449
rect 465 369 526 497
rect 556 483 610 497
rect 556 449 566 483
rect 600 449 610 483
rect 556 369 610 449
rect 640 369 703 497
rect 733 483 790 497
rect 733 449 748 483
rect 782 449 790 483
rect 733 369 790 449
rect 848 472 900 497
rect 848 438 856 472
rect 890 438 900 472
rect 848 413 900 438
rect 930 472 993 497
rect 930 438 945 472
rect 979 438 993 472
rect 930 413 993 438
rect 1023 413 1089 497
rect 1119 485 1221 497
rect 1119 451 1177 485
rect 1211 451 1221 485
rect 1119 417 1221 451
rect 1119 413 1177 417
rect 1134 383 1177 413
rect 1211 383 1221 417
rect 1134 347 1221 383
rect 1251 477 1316 497
rect 1251 443 1261 477
rect 1295 443 1316 477
rect 1251 413 1316 443
rect 1346 467 1400 497
rect 1346 433 1356 467
rect 1390 433 1400 467
rect 1346 413 1400 433
rect 1430 413 1517 497
rect 1547 477 1622 497
rect 1547 443 1579 477
rect 1613 443 1622 477
rect 1547 413 1622 443
rect 1676 475 1728 497
rect 1676 441 1684 475
rect 1718 441 1728 475
rect 1251 347 1301 413
rect 1676 407 1728 441
rect 1676 373 1684 407
rect 1718 373 1728 407
rect 1676 297 1728 373
rect 1758 455 1812 497
rect 1758 421 1768 455
rect 1802 421 1812 455
rect 1758 375 1812 421
rect 1758 341 1768 375
rect 1802 341 1812 375
rect 1758 297 1812 341
rect 1842 477 1894 497
rect 1842 443 1852 477
rect 1886 443 1894 477
rect 1842 351 1894 443
rect 1948 485 2000 497
rect 1948 451 1956 485
rect 1990 451 2000 485
rect 1948 417 2000 451
rect 1948 383 1956 417
rect 1990 383 2000 417
rect 1948 369 2000 383
rect 2030 485 2097 497
rect 2030 451 2053 485
rect 2087 451 2097 485
rect 2030 417 2097 451
rect 2030 383 2053 417
rect 2087 383 2097 417
rect 2030 369 2097 383
rect 1842 317 1852 351
rect 1886 317 1894 351
rect 1842 297 1894 317
rect 2045 349 2097 369
rect 2045 315 2053 349
rect 2087 315 2097 349
rect 2045 297 2097 315
rect 2127 449 2179 497
rect 2127 415 2137 449
rect 2171 415 2179 449
rect 2127 381 2179 415
rect 2127 347 2137 381
rect 2171 347 2179 381
rect 2127 297 2179 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 67 341 101
rect 407 55 441 89
rect 582 55 616 89
rect 749 59 783 93
rect 853 73 887 107
rect 953 73 987 107
rect 1169 67 1203 101
rect 1287 73 1321 107
rect 1399 73 1433 107
rect 1580 73 1614 107
rect 1684 128 1718 162
rect 1684 60 1718 94
rect 1768 89 1802 123
rect 1852 130 1886 164
rect 1852 62 1886 96
rect 1956 85 1990 119
rect 2053 127 2087 161
rect 2053 59 2087 93
rect 2137 109 2171 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 418 341 452
rect 391 449 425 483
rect 566 449 600 483
rect 748 449 782 483
rect 856 438 890 472
rect 945 438 979 472
rect 1177 451 1211 485
rect 1177 383 1211 417
rect 1261 443 1295 477
rect 1356 433 1390 467
rect 1579 443 1613 477
rect 1684 441 1718 475
rect 1684 373 1718 407
rect 1768 421 1802 455
rect 1768 341 1802 375
rect 1852 443 1886 477
rect 1956 451 1990 485
rect 1956 383 1990 417
rect 2053 451 2087 485
rect 2053 383 2087 417
rect 1852 317 1886 351
rect 2053 315 2087 349
rect 2137 415 2171 449
rect 2137 347 2171 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 526 497 556 523
rect 610 497 640 523
rect 703 497 733 523
rect 900 497 930 523
rect 993 497 1023 523
rect 1089 497 1119 523
rect 1221 497 1251 523
rect 1316 497 1346 523
rect 1400 497 1430 523
rect 1517 497 1547 523
rect 1728 497 1758 523
rect 1812 497 1842 523
rect 2000 497 2030 523
rect 2097 497 2127 523
rect 900 375 930 413
rect 993 381 1023 413
rect 79 348 109 363
rect 47 318 109 348
rect 47 265 77 318
rect 163 274 193 363
rect 351 331 381 369
rect 435 331 465 369
rect 526 337 556 369
rect 610 337 640 369
rect 336 321 465 331
rect 336 287 352 321
rect 386 301 465 321
rect 511 321 565 337
rect 386 287 402 301
rect 336 277 402 287
rect 511 287 521 321
rect 555 287 565 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 193 274
rect 119 230 135 264
rect 169 230 193 264
rect 119 220 193 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 131 381 277
rect 511 271 565 287
rect 607 321 661 337
rect 607 287 617 321
rect 651 287 661 321
rect 607 271 661 287
rect 703 304 733 369
rect 885 365 951 375
rect 885 331 901 365
rect 935 331 951 365
rect 885 321 951 331
rect 993 365 1047 381
rect 993 331 1003 365
rect 1037 331 1047 365
rect 993 315 1047 331
rect 703 288 757 304
rect 423 225 489 235
rect 423 191 439 225
rect 473 191 489 225
rect 423 181 489 191
rect 453 131 483 181
rect 531 131 561 271
rect 703 254 713 288
rect 747 254 757 288
rect 993 279 1023 315
rect 703 238 757 254
rect 901 249 1023 279
rect 603 207 657 223
rect 603 173 613 207
rect 647 173 657 207
rect 603 157 657 173
rect 627 131 657 157
rect 703 131 733 238
rect 901 119 931 249
rect 1089 213 1119 413
rect 1221 309 1251 347
rect 1316 315 1346 413
rect 1400 375 1430 413
rect 1517 381 1547 413
rect 1399 365 1465 375
rect 1399 331 1415 365
rect 1449 331 1465 365
rect 1399 321 1465 331
rect 1517 365 1595 381
rect 1517 331 1551 365
rect 1585 331 1595 365
rect 1517 315 1595 331
rect 1161 299 1251 309
rect 1161 265 1177 299
rect 1211 265 1251 299
rect 1161 255 1251 265
rect 1221 220 1251 255
rect 1303 299 1357 315
rect 1303 265 1313 299
rect 1347 279 1357 299
rect 1347 265 1475 279
rect 1303 249 1475 265
rect 973 191 1027 207
rect 973 157 983 191
rect 1017 157 1027 191
rect 1089 203 1169 213
rect 1089 183 1119 203
rect 973 141 1027 157
rect 997 119 1027 141
rect 1095 169 1119 183
rect 1153 169 1169 203
rect 1221 190 1271 220
rect 1241 175 1271 190
rect 1342 191 1403 207
rect 1095 159 1169 169
rect 1095 131 1125 159
rect 1342 157 1359 191
rect 1393 157 1403 191
rect 1342 141 1403 157
rect 1342 119 1372 141
rect 1445 119 1475 249
rect 1540 131 1570 315
rect 2000 333 2030 369
rect 1989 303 2030 333
rect 1728 265 1758 297
rect 1812 265 1842 297
rect 1989 265 2019 303
rect 2097 265 2127 297
rect 1619 249 1758 265
rect 1619 215 1629 249
rect 1663 215 1758 249
rect 1619 199 1758 215
rect 1800 249 2019 265
rect 1800 215 1810 249
rect 1844 215 2019 249
rect 1800 199 2019 215
rect 2068 249 2127 265
rect 2068 215 2078 249
rect 2112 215 2127 249
rect 2068 199 2127 215
rect 1728 177 1758 199
rect 1812 177 1842 199
rect 1989 176 2019 199
rect 2097 177 2127 199
rect 1989 146 2030 176
rect 2000 131 2030 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 453 21 483 47
rect 531 21 561 47
rect 627 21 657 47
rect 703 21 733 47
rect 901 21 931 47
rect 997 21 1027 47
rect 1095 21 1125 47
rect 1241 21 1271 47
rect 1342 21 1372 47
rect 1445 21 1475 47
rect 1540 21 1570 47
rect 1728 21 1758 47
rect 1812 21 1842 47
rect 2000 21 2030 47
rect 2097 21 2127 47
<< polycont >>
rect 352 287 386 321
rect 521 287 555 321
rect 33 215 67 249
rect 135 230 169 264
rect 617 287 651 321
rect 901 331 935 365
rect 1003 331 1037 365
rect 439 191 473 225
rect 713 254 747 288
rect 613 173 647 207
rect 1415 331 1449 365
rect 1551 331 1585 365
rect 1177 265 1211 299
rect 1313 265 1347 299
rect 983 157 1017 191
rect 1119 169 1153 203
rect 1359 157 1393 191
rect 1629 215 1663 249
rect 1810 215 1844 249
rect 2078 215 2112 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 203 409 237 443
rect 69 391 169 393
rect 69 375 129 391
rect 35 359 129 375
rect 123 357 129 359
rect 163 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 194 169 230
rect 123 161 162 194
rect 35 127 162 161
rect 203 187 237 375
rect 35 119 69 127
rect 203 119 237 153
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 284 452 341 489
rect 284 418 307 452
rect 375 483 441 527
rect 748 483 782 527
rect 375 449 391 483
rect 425 449 441 483
rect 535 449 566 483
rect 600 449 714 483
rect 284 415 341 418
rect 284 372 646 415
rect 284 117 318 372
rect 352 321 386 337
rect 352 176 386 287
rect 420 225 454 372
rect 612 337 646 372
rect 680 399 714 449
rect 748 433 782 449
rect 833 472 890 488
rect 1177 485 1211 527
rect 833 438 856 472
rect 929 438 945 472
rect 979 438 1143 472
rect 833 414 890 438
rect 833 399 867 414
rect 680 365 867 399
rect 987 391 1075 402
rect 488 321 555 337
rect 488 287 521 321
rect 488 271 555 287
rect 612 321 651 337
rect 612 287 617 321
rect 612 271 651 287
rect 703 288 799 331
rect 703 254 713 288
rect 747 254 799 288
rect 420 191 439 225
rect 473 191 489 225
rect 613 207 647 223
rect 703 211 799 254
rect 352 175 388 176
rect 352 174 389 175
rect 352 172 390 174
rect 833 177 867 365
rect 352 171 391 172
rect 352 170 392 171
rect 352 168 393 170
rect 352 167 394 168
rect 352 164 395 167
rect 352 162 398 164
rect 352 157 402 162
rect 613 157 647 173
rect 352 150 647 157
rect 358 147 647 150
rect 361 145 647 147
rect 364 143 647 145
rect 366 141 647 143
rect 368 138 647 141
rect 372 131 647 138
rect 375 123 647 131
rect 681 143 867 177
rect 284 101 341 117
rect 103 17 169 59
rect 284 67 307 101
rect 284 51 341 67
rect 391 55 407 89
rect 441 55 457 89
rect 491 61 526 123
rect 681 89 715 143
rect 560 55 582 89
rect 616 55 715 89
rect 749 93 789 109
rect 783 59 789 93
rect 833 107 867 143
rect 901 365 949 381
rect 935 331 949 365
rect 987 365 1033 391
rect 987 331 1003 365
rect 1067 357 1075 391
rect 1037 331 1075 357
rect 901 207 949 331
rect 1109 315 1143 438
rect 1177 417 1211 451
rect 1177 367 1211 383
rect 1245 477 1295 493
rect 1245 443 1261 477
rect 1553 477 1614 527
rect 1245 427 1295 443
rect 1340 433 1356 467
rect 1390 433 1517 467
rect 1109 299 1211 315
rect 1109 297 1177 299
rect 1051 265 1177 297
rect 1051 263 1211 265
rect 901 191 1017 207
rect 901 187 983 191
rect 901 153 949 187
rect 983 153 1017 157
rect 901 141 1017 153
rect 1051 107 1085 263
rect 1177 249 1211 263
rect 1119 213 1153 219
rect 1245 213 1279 427
rect 1313 391 1351 393
rect 1313 357 1315 391
rect 1349 357 1351 391
rect 1313 299 1351 357
rect 1347 265 1351 299
rect 1313 249 1351 265
rect 1385 365 1449 381
rect 1385 331 1415 365
rect 1385 315 1449 331
rect 1119 203 1279 213
rect 1385 207 1423 315
rect 1483 281 1517 433
rect 1553 443 1579 477
rect 1613 443 1614 477
rect 1553 427 1614 443
rect 1676 475 1734 491
rect 1676 441 1684 475
rect 1718 441 1734 475
rect 1676 407 1734 441
rect 1676 381 1684 407
rect 1551 373 1684 381
rect 1718 373 1734 407
rect 1551 365 1734 373
rect 1585 331 1734 365
rect 1551 315 1734 331
rect 1768 455 1802 527
rect 1768 375 1802 421
rect 1768 325 1802 341
rect 1840 477 1906 493
rect 2042 485 2103 527
rect 1840 443 1852 477
rect 1886 443 1906 477
rect 1840 351 1906 443
rect 1153 169 1279 203
rect 1119 153 1279 169
rect 833 73 853 107
rect 887 73 903 107
rect 937 73 953 107
rect 987 73 1085 107
rect 1135 101 1209 117
rect 391 17 457 55
rect 749 17 789 59
rect 1135 67 1169 101
rect 1203 67 1209 101
rect 1245 107 1279 153
rect 1313 191 1423 207
rect 1313 187 1359 191
rect 1313 153 1317 187
rect 1351 157 1359 187
rect 1393 157 1423 191
rect 1351 153 1423 157
rect 1313 141 1423 153
rect 1457 265 1517 281
rect 1697 265 1734 315
rect 1840 317 1852 351
rect 1886 317 1906 351
rect 1940 451 1956 485
rect 1990 451 2006 485
rect 1940 417 2006 451
rect 1940 383 1956 417
rect 1990 383 2006 417
rect 1940 337 2006 383
rect 1840 308 1906 317
rect 1840 301 1922 308
rect 1871 286 1922 301
rect 1457 249 1663 265
rect 1457 215 1629 249
rect 1457 199 1663 215
rect 1697 249 1844 265
rect 1697 215 1810 249
rect 1697 199 1844 215
rect 1457 107 1491 199
rect 1697 165 1734 199
rect 1878 165 1922 286
rect 1668 162 1734 165
rect 1668 128 1684 162
rect 1718 128 1734 162
rect 1836 164 1922 165
rect 1245 73 1287 107
rect 1321 73 1337 107
rect 1383 73 1399 107
rect 1433 73 1491 107
rect 1540 107 1614 123
rect 1540 73 1580 107
rect 1135 17 1209 67
rect 1540 17 1614 73
rect 1668 94 1734 128
rect 1668 60 1684 94
rect 1718 60 1734 94
rect 1768 123 1802 139
rect 1768 17 1802 89
rect 1836 130 1852 164
rect 1886 158 1922 164
rect 1956 265 2006 337
rect 2042 451 2053 485
rect 2087 451 2103 485
rect 2042 417 2103 451
rect 2042 383 2053 417
rect 2087 383 2103 417
rect 2042 349 2103 383
rect 2042 315 2053 349
rect 2087 315 2103 349
rect 2042 299 2103 315
rect 2137 449 2188 465
rect 2171 415 2188 449
rect 2137 381 2188 415
rect 2171 347 2188 381
rect 2137 289 2188 347
rect 1956 249 2112 265
rect 1956 215 2078 249
rect 1956 199 2112 215
rect 1886 145 1912 158
rect 1886 130 1906 145
rect 1836 96 1906 130
rect 1956 124 1990 199
rect 1836 62 1852 96
rect 1886 62 1906 96
rect 1940 119 1990 124
rect 1940 85 1956 119
rect 1940 69 1990 85
rect 2037 127 2053 161
rect 2087 127 2103 161
rect 2146 159 2188 289
rect 2037 93 2103 127
rect 1836 61 1906 62
rect 2037 59 2053 93
rect 2087 59 2103 93
rect 2037 17 2103 59
rect 2137 143 2188 159
rect 2171 109 2188 143
rect 2137 53 2188 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 129 357 163 391
rect 203 153 237 187
rect 1033 365 1067 391
rect 1033 357 1037 365
rect 1037 357 1067 365
rect 949 153 983 187
rect 1315 357 1349 391
rect 1317 153 1351 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 1021 391 1079 397
rect 1021 388 1033 391
rect 163 360 1033 388
rect 163 357 175 360
rect 117 351 175 357
rect 1021 357 1033 360
rect 1067 388 1079 391
rect 1303 391 1361 397
rect 1303 388 1315 391
rect 1067 360 1315 388
rect 1067 357 1079 360
rect 1021 351 1079 357
rect 1303 357 1315 360
rect 1349 357 1361 391
rect 1303 351 1361 357
rect 191 187 249 193
rect 191 153 203 187
rect 237 184 249 187
rect 937 187 995 193
rect 937 184 949 187
rect 237 156 949 184
rect 237 153 249 156
rect 191 147 249 153
rect 937 153 949 156
rect 983 184 995 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 983 156 1317 184
rect 983 153 995 156
rect 937 147 995 153
rect 1305 153 1317 156
rect 1351 153 1363 187
rect 1305 147 1363 153
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 763 221 797 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel locali s 2143 289 2177 323 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 491 85 525 119 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1867 85 1901 119 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 sdfxbp_1
rlabel metal1 s 0 -48 2208 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2208 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_END 343100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 326098
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.040 0.000 
<< end >>
