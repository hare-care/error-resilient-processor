magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 2274 897
<< pwell >>
rect 1928 281 2186 283
rect 1604 269 2186 281
rect 32 242 610 269
rect 1040 242 2186 269
rect 32 43 2186 242
rect -26 -43 2234 43
<< locali >>
rect 119 307 185 425
rect 295 307 361 425
rect 864 293 930 395
rect 1839 625 1912 689
rect 1862 405 1912 625
rect 1862 345 1928 405
rect 2118 379 2191 747
rect 2137 243 2191 379
rect 2118 103 2191 243
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 58 757 858 763
rect 58 729 364 757
rect 58 695 76 729
rect 110 695 148 729
rect 182 695 220 729
rect 254 695 292 729
rect 326 723 364 729
rect 398 723 436 757
rect 470 723 508 757
rect 542 723 591 757
rect 625 723 663 757
rect 697 729 858 757
rect 697 723 735 729
rect 326 695 397 723
rect 58 689 397 695
rect 725 695 735 723
rect 769 695 807 729
rect 841 695 858 729
rect 1329 757 2084 763
rect 1329 743 1831 757
rect 1329 729 1479 743
rect 725 689 858 695
rect 58 459 124 689
rect 431 645 691 689
rect 370 459 429 611
rect 395 273 429 459
rect 526 377 592 611
rect 647 463 691 645
rect 792 497 858 689
rect 896 677 1295 711
rect 1329 695 1335 729
rect 1369 695 1407 729
rect 1441 709 1479 729
rect 1513 709 1551 743
rect 1585 729 1831 743
rect 1585 709 1623 729
rect 1441 695 1623 709
rect 1657 695 1695 729
rect 1729 723 1831 729
rect 1865 723 1903 757
rect 1937 729 2084 757
rect 1937 723 1975 729
rect 1729 695 1805 723
rect 1329 689 1805 695
rect 1946 695 1975 723
rect 2009 695 2047 729
rect 2081 695 2084 729
rect 1946 689 2084 695
rect 896 463 930 677
rect 647 429 930 463
rect 964 601 1227 643
rect 511 311 613 377
rect 58 239 429 273
rect 58 168 124 239
rect 214 125 280 205
rect 370 168 429 239
rect 526 168 592 311
rect 647 216 686 429
rect 636 141 686 216
rect 720 259 786 393
rect 964 259 1006 601
rect 720 225 1006 259
rect 146 119 348 125
rect 146 85 158 119
rect 192 85 230 119
rect 264 85 302 119
rect 336 85 348 119
rect 146 73 348 85
rect 423 107 565 134
rect 720 107 754 225
rect 423 73 754 107
rect 788 125 858 191
rect 956 141 1006 225
rect 1067 466 1124 532
rect 1261 519 1295 677
rect 1219 485 1295 519
rect 1067 273 1101 466
rect 1219 389 1253 485
rect 1356 466 1422 689
rect 1524 417 1578 532
rect 1622 445 1688 689
rect 1135 323 1253 389
rect 1295 375 1578 417
rect 1295 307 1361 375
rect 1524 365 1578 375
rect 1683 365 1749 411
rect 1417 273 1490 331
rect 1067 239 1490 273
rect 788 119 922 125
rect 788 85 791 119
rect 825 85 863 119
rect 897 107 922 119
rect 1067 107 1124 239
rect 1356 125 1422 205
rect 897 105 977 107
rect 897 85 935 105
rect 788 71 935 85
rect 969 71 977 105
rect 788 51 977 71
rect 1011 51 1124 107
rect 1158 119 1422 125
rect 1158 105 1310 119
rect 1158 71 1166 105
rect 1200 71 1238 105
rect 1272 85 1310 105
rect 1344 85 1382 119
rect 1416 85 1422 119
rect 1272 71 1422 85
rect 1456 134 1490 239
rect 1524 323 1749 365
rect 1524 168 1578 323
rect 1683 277 1749 323
rect 1783 311 1828 591
rect 1946 439 2012 689
rect 1981 311 2103 345
rect 1783 277 2103 311
rect 1783 243 1828 277
rect 1622 177 1828 243
rect 1456 71 1574 134
rect 1946 125 2012 243
rect 1608 119 2084 125
rect 1608 105 1900 119
rect 1608 71 1612 105
rect 1646 71 1684 105
rect 1718 71 1756 105
rect 1790 71 1828 105
rect 1862 85 1900 105
rect 1934 85 1972 119
rect 2006 85 2044 119
rect 2078 85 2084 119
rect 1862 71 2084 85
rect 1158 51 1422 71
rect 1608 51 2084 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 76 695 110 729
rect 148 695 182 729
rect 220 695 254 729
rect 292 695 326 729
rect 364 723 398 757
rect 436 723 470 757
rect 508 723 542 757
rect 591 723 625 757
rect 663 723 697 757
rect 735 695 769 729
rect 807 695 841 729
rect 1335 695 1369 729
rect 1407 695 1441 729
rect 1479 709 1513 743
rect 1551 709 1585 743
rect 1623 695 1657 729
rect 1695 695 1729 729
rect 1831 723 1865 757
rect 1903 723 1937 757
rect 1975 695 2009 729
rect 2047 695 2081 729
rect 158 85 192 119
rect 230 85 264 119
rect 302 85 336 119
rect 791 85 825 119
rect 863 85 897 119
rect 935 71 969 105
rect 1166 71 1200 105
rect 1238 71 1272 105
rect 1310 85 1344 119
rect 1382 85 1416 119
rect 1612 71 1646 105
rect 1684 71 1718 105
rect 1756 71 1790 105
rect 1828 71 1862 105
rect 1900 85 1934 119
rect 1972 85 2006 119
rect 2044 85 2078 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 831 2208 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2208 831
rect 0 791 2208 797
rect 0 757 2208 763
rect 0 729 364 757
rect 0 695 76 729
rect 110 695 148 729
rect 182 695 220 729
rect 254 695 292 729
rect 326 723 364 729
rect 398 723 436 757
rect 470 723 508 757
rect 542 723 591 757
rect 625 723 663 757
rect 697 743 1831 757
rect 697 729 1479 743
rect 697 723 735 729
rect 326 695 735 723
rect 769 695 807 729
rect 841 695 1335 729
rect 1369 695 1407 729
rect 1441 709 1479 729
rect 1513 709 1551 743
rect 1585 729 1831 743
rect 1585 709 1623 729
rect 1441 695 1623 709
rect 1657 695 1695 729
rect 1729 723 1831 729
rect 1865 723 1903 757
rect 1937 729 2208 757
rect 1937 723 1975 729
rect 1729 695 1975 723
rect 2009 695 2047 729
rect 2081 695 2208 729
rect 0 689 2208 695
rect 0 119 2208 125
rect 0 85 158 119
rect 192 85 230 119
rect 264 85 302 119
rect 336 85 791 119
rect 825 85 863 119
rect 897 105 1310 119
rect 897 85 935 105
rect 0 71 935 85
rect 969 71 1166 105
rect 1200 71 1238 105
rect 1272 85 1310 105
rect 1344 85 1382 119
rect 1416 105 1900 119
rect 1416 85 1612 105
rect 1272 71 1612 85
rect 1646 71 1684 105
rect 1718 71 1756 105
rect 1790 71 1828 105
rect 1862 85 1900 105
rect 1934 85 1972 119
rect 2006 85 2044 119
rect 2078 85 2208 119
rect 1862 71 2208 85
rect 0 51 2208 71
rect 0 17 2208 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -23 2208 -17
<< labels >>
rlabel locali s 1862 345 1928 405 6 CLK
port 1 nsew clock input
rlabel locali s 864 293 930 395 6 CLK
port 1 nsew clock input
rlabel locali s 1862 405 1912 625 6 CLK
port 1 nsew clock input
rlabel locali s 1839 625 1912 689 6 CLK
port 1 nsew clock input
rlabel locali s 295 307 361 425 6 GATE
port 2 nsew signal input
rlabel locali s 119 307 185 425 6 SCE
port 3 nsew signal input
rlabel metal1 s 0 51 2208 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 2208 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 2234 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 32 43 2186 242 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1040 242 2186 269 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 32 242 610 269 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1604 269 2186 281 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1928 281 2186 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 2208 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 2274 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 2208 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 2118 103 2191 243 6 GCLK
port 8 nsew signal output
rlabel locali s 2137 243 2191 379 6 GCLK
port 8 nsew signal output
rlabel locali s 2118 379 2191 747 6 GCLK
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 695048
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 672184
<< end >>
