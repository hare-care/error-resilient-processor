magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 7273 3544 11349 3740
rect 7273 408 7483 3544
rect 11159 408 11349 3544
rect 7273 218 11349 408
<< pwell >>
rect 7497 450 11145 3502
<< psubdiff >>
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
<< nsubdiff >>
rect 7319 3646 11313 3698
rect 7319 3612 7421 3646
rect 7455 3612 7489 3646
rect 7523 3612 7557 3646
rect 7591 3612 7625 3646
rect 7659 3612 7693 3646
rect 7727 3612 7761 3646
rect 7795 3612 7829 3646
rect 7863 3612 7897 3646
rect 7931 3612 7965 3646
rect 7999 3612 8033 3646
rect 8067 3612 8101 3646
rect 8135 3612 8169 3646
rect 8203 3612 8237 3646
rect 8271 3612 8305 3646
rect 8339 3612 8373 3646
rect 8407 3612 8441 3646
rect 8475 3612 8509 3646
rect 8543 3612 8577 3646
rect 8611 3612 8645 3646
rect 8679 3612 8713 3646
rect 8747 3612 8781 3646
rect 8815 3612 8849 3646
rect 8883 3612 8917 3646
rect 8951 3612 8985 3646
rect 9019 3612 9053 3646
rect 9087 3612 9121 3646
rect 9155 3612 9189 3646
rect 9223 3612 9257 3646
rect 9291 3612 9325 3646
rect 9359 3612 9393 3646
rect 9427 3612 9461 3646
rect 9495 3612 9529 3646
rect 9563 3612 9597 3646
rect 9631 3612 9665 3646
rect 9699 3612 9733 3646
rect 9767 3612 9801 3646
rect 9835 3612 9869 3646
rect 9903 3612 9937 3646
rect 9971 3612 10005 3646
rect 10039 3612 10073 3646
rect 10107 3612 10141 3646
rect 10175 3612 10209 3646
rect 10243 3612 10277 3646
rect 10311 3612 10345 3646
rect 10379 3612 10413 3646
rect 10447 3612 10481 3646
rect 10515 3612 10549 3646
rect 10583 3612 10617 3646
rect 10651 3612 10685 3646
rect 10719 3612 10753 3646
rect 10787 3612 10821 3646
rect 10855 3612 10889 3646
rect 10923 3612 10957 3646
rect 10991 3612 11025 3646
rect 11059 3612 11093 3646
rect 11127 3612 11161 3646
rect 11195 3612 11313 3646
rect 7319 3580 11313 3612
rect 7319 3557 7447 3580
rect 7319 3523 7353 3557
rect 7387 3523 7447 3557
rect 7319 3489 7447 3523
rect 7319 3455 7353 3489
rect 7387 3455 7447 3489
rect 11195 3557 11313 3580
rect 11195 3523 11255 3557
rect 11289 3523 11313 3557
rect 11195 3489 11313 3523
rect 7319 3421 7447 3455
rect 7319 3387 7353 3421
rect 7387 3387 7447 3421
rect 7319 3353 7447 3387
rect 7319 3319 7353 3353
rect 7387 3319 7447 3353
rect 7319 3285 7447 3319
rect 7319 3251 7353 3285
rect 7387 3251 7447 3285
rect 7319 3217 7447 3251
rect 7319 3183 7353 3217
rect 7387 3183 7447 3217
rect 7319 3149 7447 3183
rect 7319 3115 7353 3149
rect 7387 3115 7447 3149
rect 7319 3081 7447 3115
rect 7319 3047 7353 3081
rect 7387 3047 7447 3081
rect 7319 3013 7447 3047
rect 7319 2979 7353 3013
rect 7387 2979 7447 3013
rect 7319 2945 7447 2979
rect 7319 2911 7353 2945
rect 7387 2911 7447 2945
rect 7319 2877 7447 2911
rect 7319 2843 7353 2877
rect 7387 2843 7447 2877
rect 7319 2809 7447 2843
rect 7319 2775 7353 2809
rect 7387 2775 7447 2809
rect 7319 2741 7447 2775
rect 7319 2707 7353 2741
rect 7387 2707 7447 2741
rect 7319 2673 7447 2707
rect 7319 2639 7353 2673
rect 7387 2639 7447 2673
rect 7319 2605 7447 2639
rect 7319 2571 7353 2605
rect 7387 2571 7447 2605
rect 7319 2537 7447 2571
rect 7319 2503 7353 2537
rect 7387 2503 7447 2537
rect 7319 2469 7447 2503
rect 7319 2435 7353 2469
rect 7387 2435 7447 2469
rect 7319 2401 7447 2435
rect 7319 2367 7353 2401
rect 7387 2367 7447 2401
rect 7319 2333 7447 2367
rect 7319 2299 7353 2333
rect 7387 2299 7447 2333
rect 7319 2265 7447 2299
rect 7319 2231 7353 2265
rect 7387 2231 7447 2265
rect 7319 2197 7447 2231
rect 7319 2163 7353 2197
rect 7387 2163 7447 2197
rect 7319 2129 7447 2163
rect 7319 2095 7353 2129
rect 7387 2095 7447 2129
rect 7319 2061 7447 2095
rect 7319 2027 7353 2061
rect 7387 2027 7447 2061
rect 7319 1993 7447 2027
rect 7319 1959 7353 1993
rect 7387 1959 7447 1993
rect 7319 1925 7447 1959
rect 7319 1891 7353 1925
rect 7387 1891 7447 1925
rect 7319 1857 7447 1891
rect 7319 1823 7353 1857
rect 7387 1823 7447 1857
rect 7319 1789 7447 1823
rect 7319 1755 7353 1789
rect 7387 1755 7447 1789
rect 7319 1721 7447 1755
rect 7319 1687 7353 1721
rect 7387 1687 7447 1721
rect 7319 1653 7447 1687
rect 7319 1619 7353 1653
rect 7387 1619 7447 1653
rect 7319 1585 7447 1619
rect 7319 1551 7353 1585
rect 7387 1551 7447 1585
rect 7319 1517 7447 1551
rect 7319 1483 7353 1517
rect 7387 1483 7447 1517
rect 7319 1449 7447 1483
rect 7319 1415 7353 1449
rect 7387 1415 7447 1449
rect 7319 1381 7447 1415
rect 7319 1347 7353 1381
rect 7387 1347 7447 1381
rect 7319 1313 7447 1347
rect 7319 1279 7353 1313
rect 7387 1279 7447 1313
rect 7319 1245 7447 1279
rect 7319 1211 7353 1245
rect 7387 1211 7447 1245
rect 7319 1177 7447 1211
rect 7319 1143 7353 1177
rect 7387 1143 7447 1177
rect 7319 1109 7447 1143
rect 7319 1075 7353 1109
rect 7387 1075 7447 1109
rect 7319 1041 7447 1075
rect 7319 1007 7353 1041
rect 7387 1007 7447 1041
rect 7319 973 7447 1007
rect 7319 939 7353 973
rect 7387 939 7447 973
rect 7319 905 7447 939
rect 7319 871 7353 905
rect 7387 871 7447 905
rect 7319 837 7447 871
rect 7319 803 7353 837
rect 7387 803 7447 837
rect 7319 769 7447 803
rect 7319 735 7353 769
rect 7387 735 7447 769
rect 7319 701 7447 735
rect 7319 667 7353 701
rect 7387 667 7447 701
rect 7319 633 7447 667
rect 7319 599 7353 633
rect 7387 599 7447 633
rect 7319 565 7447 599
rect 7319 531 7353 565
rect 7387 531 7447 565
rect 7319 497 7447 531
rect 7319 463 7353 497
rect 7387 463 7447 497
rect 11195 3455 11255 3489
rect 11289 3455 11313 3489
rect 11195 3421 11313 3455
rect 11195 3387 11255 3421
rect 11289 3387 11313 3421
rect 11195 3353 11313 3387
rect 11195 3319 11255 3353
rect 11289 3319 11313 3353
rect 11195 3285 11313 3319
rect 11195 3251 11255 3285
rect 11289 3251 11313 3285
rect 11195 3217 11313 3251
rect 11195 3183 11255 3217
rect 11289 3183 11313 3217
rect 11195 3149 11313 3183
rect 11195 3115 11255 3149
rect 11289 3115 11313 3149
rect 11195 3081 11313 3115
rect 11195 3047 11255 3081
rect 11289 3047 11313 3081
rect 11195 3013 11313 3047
rect 11195 2979 11255 3013
rect 11289 2979 11313 3013
rect 11195 2945 11313 2979
rect 11195 2911 11255 2945
rect 11289 2911 11313 2945
rect 11195 2877 11313 2911
rect 11195 2843 11255 2877
rect 11289 2843 11313 2877
rect 11195 2809 11313 2843
rect 11195 2775 11255 2809
rect 11289 2775 11313 2809
rect 11195 2741 11313 2775
rect 11195 2707 11255 2741
rect 11289 2707 11313 2741
rect 11195 2673 11313 2707
rect 11195 2639 11255 2673
rect 11289 2639 11313 2673
rect 11195 2605 11313 2639
rect 11195 2571 11255 2605
rect 11289 2571 11313 2605
rect 11195 2537 11313 2571
rect 11195 2503 11255 2537
rect 11289 2503 11313 2537
rect 11195 2469 11313 2503
rect 11195 2435 11255 2469
rect 11289 2435 11313 2469
rect 11195 2401 11313 2435
rect 11195 2367 11255 2401
rect 11289 2367 11313 2401
rect 11195 2333 11313 2367
rect 11195 2299 11255 2333
rect 11289 2299 11313 2333
rect 11195 2265 11313 2299
rect 11195 2231 11255 2265
rect 11289 2231 11313 2265
rect 11195 2197 11313 2231
rect 11195 2163 11255 2197
rect 11289 2163 11313 2197
rect 11195 2129 11313 2163
rect 11195 2095 11255 2129
rect 11289 2095 11313 2129
rect 11195 2061 11313 2095
rect 11195 2027 11255 2061
rect 11289 2027 11313 2061
rect 11195 1993 11313 2027
rect 11195 1959 11255 1993
rect 11289 1959 11313 1993
rect 11195 1925 11313 1959
rect 11195 1891 11255 1925
rect 11289 1891 11313 1925
rect 11195 1857 11313 1891
rect 11195 1823 11255 1857
rect 11289 1823 11313 1857
rect 11195 1789 11313 1823
rect 11195 1755 11255 1789
rect 11289 1755 11313 1789
rect 11195 1721 11313 1755
rect 11195 1687 11255 1721
rect 11289 1687 11313 1721
rect 11195 1653 11313 1687
rect 11195 1619 11255 1653
rect 11289 1619 11313 1653
rect 11195 1585 11313 1619
rect 11195 1551 11255 1585
rect 11289 1551 11313 1585
rect 11195 1517 11313 1551
rect 11195 1483 11255 1517
rect 11289 1483 11313 1517
rect 11195 1449 11313 1483
rect 11195 1415 11255 1449
rect 11289 1415 11313 1449
rect 11195 1381 11313 1415
rect 11195 1347 11255 1381
rect 11289 1347 11313 1381
rect 11195 1313 11313 1347
rect 11195 1279 11255 1313
rect 11289 1279 11313 1313
rect 11195 1245 11313 1279
rect 11195 1211 11255 1245
rect 11289 1211 11313 1245
rect 11195 1177 11313 1211
rect 11195 1143 11255 1177
rect 11289 1143 11313 1177
rect 11195 1109 11313 1143
rect 11195 1075 11255 1109
rect 11289 1075 11313 1109
rect 11195 1041 11313 1075
rect 11195 1007 11255 1041
rect 11289 1007 11313 1041
rect 11195 973 11313 1007
rect 11195 939 11255 973
rect 11289 939 11313 973
rect 11195 905 11313 939
rect 11195 871 11255 905
rect 11289 871 11313 905
rect 11195 837 11313 871
rect 11195 803 11255 837
rect 11289 803 11313 837
rect 11195 769 11313 803
rect 11195 735 11255 769
rect 11289 735 11313 769
rect 11195 701 11313 735
rect 11195 667 11255 701
rect 11289 667 11313 701
rect 11195 633 11313 667
rect 11195 599 11255 633
rect 11289 599 11313 633
rect 11195 565 11313 599
rect 11195 531 11255 565
rect 11289 531 11313 565
rect 11195 497 11313 531
rect 7319 429 7447 463
rect 7319 395 7353 429
rect 7387 395 7447 429
rect 7319 372 7447 395
rect 11195 463 11255 497
rect 11289 463 11313 497
rect 11195 429 11313 463
rect 11195 395 11255 429
rect 11289 395 11313 429
rect 11195 372 11313 395
rect 7319 334 11313 372
rect 7319 300 7411 334
rect 7445 300 7479 334
rect 7513 300 7547 334
rect 7581 300 7615 334
rect 7649 300 7683 334
rect 7717 300 7751 334
rect 7785 300 7819 334
rect 7853 300 7887 334
rect 7921 300 7955 334
rect 7989 300 8023 334
rect 8057 300 8091 334
rect 8125 300 8159 334
rect 8193 300 8227 334
rect 8261 300 8295 334
rect 8329 300 8363 334
rect 8397 300 8431 334
rect 8465 300 8499 334
rect 8533 300 8567 334
rect 8601 300 8635 334
rect 8669 300 8703 334
rect 8737 300 8771 334
rect 8805 300 8839 334
rect 8873 300 8907 334
rect 8941 300 8975 334
rect 9009 300 9043 334
rect 9077 300 9111 334
rect 9145 300 9179 334
rect 9213 300 9247 334
rect 9281 300 9315 334
rect 9349 300 9383 334
rect 9417 300 9451 334
rect 9485 300 9519 334
rect 9553 300 9587 334
rect 9621 300 9655 334
rect 9689 300 9723 334
rect 9757 300 9791 334
rect 9825 300 9859 334
rect 9893 300 9927 334
rect 9961 300 9995 334
rect 10029 300 10063 334
rect 10097 300 10131 334
rect 10165 300 10199 334
rect 10233 300 10267 334
rect 10301 300 10335 334
rect 10369 300 10403 334
rect 10437 300 10471 334
rect 10505 300 10539 334
rect 10573 300 10607 334
rect 10641 300 10675 334
rect 10709 300 10743 334
rect 10777 300 10811 334
rect 10845 300 10879 334
rect 10913 300 10947 334
rect 10981 300 11015 334
rect 11049 300 11083 334
rect 11117 300 11151 334
rect 11185 300 11313 334
rect 7319 254 11313 300
<< psubdiffcont >>
rect 7554 531 7792 3421
rect 8378 531 8616 3421
rect 9202 531 9440 3421
rect 10026 531 10264 3421
rect 10850 531 11088 3421
<< nsubdiffcont >>
rect 7421 3612 7455 3646
rect 7489 3612 7523 3646
rect 7557 3612 7591 3646
rect 7625 3612 7659 3646
rect 7693 3612 7727 3646
rect 7761 3612 7795 3646
rect 7829 3612 7863 3646
rect 7897 3612 7931 3646
rect 7965 3612 7999 3646
rect 8033 3612 8067 3646
rect 8101 3612 8135 3646
rect 8169 3612 8203 3646
rect 8237 3612 8271 3646
rect 8305 3612 8339 3646
rect 8373 3612 8407 3646
rect 8441 3612 8475 3646
rect 8509 3612 8543 3646
rect 8577 3612 8611 3646
rect 8645 3612 8679 3646
rect 8713 3612 8747 3646
rect 8781 3612 8815 3646
rect 8849 3612 8883 3646
rect 8917 3612 8951 3646
rect 8985 3612 9019 3646
rect 9053 3612 9087 3646
rect 9121 3612 9155 3646
rect 9189 3612 9223 3646
rect 9257 3612 9291 3646
rect 9325 3612 9359 3646
rect 9393 3612 9427 3646
rect 9461 3612 9495 3646
rect 9529 3612 9563 3646
rect 9597 3612 9631 3646
rect 9665 3612 9699 3646
rect 9733 3612 9767 3646
rect 9801 3612 9835 3646
rect 9869 3612 9903 3646
rect 9937 3612 9971 3646
rect 10005 3612 10039 3646
rect 10073 3612 10107 3646
rect 10141 3612 10175 3646
rect 10209 3612 10243 3646
rect 10277 3612 10311 3646
rect 10345 3612 10379 3646
rect 10413 3612 10447 3646
rect 10481 3612 10515 3646
rect 10549 3612 10583 3646
rect 10617 3612 10651 3646
rect 10685 3612 10719 3646
rect 10753 3612 10787 3646
rect 10821 3612 10855 3646
rect 10889 3612 10923 3646
rect 10957 3612 10991 3646
rect 11025 3612 11059 3646
rect 11093 3612 11127 3646
rect 11161 3612 11195 3646
rect 7353 3523 7387 3557
rect 7353 3455 7387 3489
rect 11255 3523 11289 3557
rect 7353 3387 7387 3421
rect 7353 3319 7387 3353
rect 7353 3251 7387 3285
rect 7353 3183 7387 3217
rect 7353 3115 7387 3149
rect 7353 3047 7387 3081
rect 7353 2979 7387 3013
rect 7353 2911 7387 2945
rect 7353 2843 7387 2877
rect 7353 2775 7387 2809
rect 7353 2707 7387 2741
rect 7353 2639 7387 2673
rect 7353 2571 7387 2605
rect 7353 2503 7387 2537
rect 7353 2435 7387 2469
rect 7353 2367 7387 2401
rect 7353 2299 7387 2333
rect 7353 2231 7387 2265
rect 7353 2163 7387 2197
rect 7353 2095 7387 2129
rect 7353 2027 7387 2061
rect 7353 1959 7387 1993
rect 7353 1891 7387 1925
rect 7353 1823 7387 1857
rect 7353 1755 7387 1789
rect 7353 1687 7387 1721
rect 7353 1619 7387 1653
rect 7353 1551 7387 1585
rect 7353 1483 7387 1517
rect 7353 1415 7387 1449
rect 7353 1347 7387 1381
rect 7353 1279 7387 1313
rect 7353 1211 7387 1245
rect 7353 1143 7387 1177
rect 7353 1075 7387 1109
rect 7353 1007 7387 1041
rect 7353 939 7387 973
rect 7353 871 7387 905
rect 7353 803 7387 837
rect 7353 735 7387 769
rect 7353 667 7387 701
rect 7353 599 7387 633
rect 7353 531 7387 565
rect 7353 463 7387 497
rect 11255 3455 11289 3489
rect 11255 3387 11289 3421
rect 11255 3319 11289 3353
rect 11255 3251 11289 3285
rect 11255 3183 11289 3217
rect 11255 3115 11289 3149
rect 11255 3047 11289 3081
rect 11255 2979 11289 3013
rect 11255 2911 11289 2945
rect 11255 2843 11289 2877
rect 11255 2775 11289 2809
rect 11255 2707 11289 2741
rect 11255 2639 11289 2673
rect 11255 2571 11289 2605
rect 11255 2503 11289 2537
rect 11255 2435 11289 2469
rect 11255 2367 11289 2401
rect 11255 2299 11289 2333
rect 11255 2231 11289 2265
rect 11255 2163 11289 2197
rect 11255 2095 11289 2129
rect 11255 2027 11289 2061
rect 11255 1959 11289 1993
rect 11255 1891 11289 1925
rect 11255 1823 11289 1857
rect 11255 1755 11289 1789
rect 11255 1687 11289 1721
rect 11255 1619 11289 1653
rect 11255 1551 11289 1585
rect 11255 1483 11289 1517
rect 11255 1415 11289 1449
rect 11255 1347 11289 1381
rect 11255 1279 11289 1313
rect 11255 1211 11289 1245
rect 11255 1143 11289 1177
rect 11255 1075 11289 1109
rect 11255 1007 11289 1041
rect 11255 939 11289 973
rect 11255 871 11289 905
rect 11255 803 11289 837
rect 11255 735 11289 769
rect 11255 667 11289 701
rect 11255 599 11289 633
rect 11255 531 11289 565
rect 7353 395 7387 429
rect 11255 463 11289 497
rect 11255 395 11289 429
rect 7411 300 7445 334
rect 7479 300 7513 334
rect 7547 300 7581 334
rect 7615 300 7649 334
rect 7683 300 7717 334
rect 7751 300 7785 334
rect 7819 300 7853 334
rect 7887 300 7921 334
rect 7955 300 7989 334
rect 8023 300 8057 334
rect 8091 300 8125 334
rect 8159 300 8193 334
rect 8227 300 8261 334
rect 8295 300 8329 334
rect 8363 300 8397 334
rect 8431 300 8465 334
rect 8499 300 8533 334
rect 8567 300 8601 334
rect 8635 300 8669 334
rect 8703 300 8737 334
rect 8771 300 8805 334
rect 8839 300 8873 334
rect 8907 300 8941 334
rect 8975 300 9009 334
rect 9043 300 9077 334
rect 9111 300 9145 334
rect 9179 300 9213 334
rect 9247 300 9281 334
rect 9315 300 9349 334
rect 9383 300 9417 334
rect 9451 300 9485 334
rect 9519 300 9553 334
rect 9587 300 9621 334
rect 9655 300 9689 334
rect 9723 300 9757 334
rect 9791 300 9825 334
rect 9859 300 9893 334
rect 9927 300 9961 334
rect 9995 300 10029 334
rect 10063 300 10097 334
rect 10131 300 10165 334
rect 10199 300 10233 334
rect 10267 300 10301 334
rect 10335 300 10369 334
rect 10403 300 10437 334
rect 10471 300 10505 334
rect 10539 300 10573 334
rect 10607 300 10641 334
rect 10675 300 10709 334
rect 10743 300 10777 334
rect 10811 300 10845 334
rect 10879 300 10913 334
rect 10947 300 10981 334
rect 11015 300 11049 334
rect 11083 300 11117 334
rect 11151 300 11185 334
<< ndiode >>
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
<< ndiodec >>
rect 7966 531 8204 3421
rect 8790 531 9028 3421
rect 9614 531 9852 3421
rect 10438 531 10676 3421
<< locali >>
rect 7319 3664 11313 3698
rect 7319 3646 7428 3664
rect 7462 3646 7501 3664
rect 7535 3646 7574 3664
rect 7608 3646 7646 3664
rect 7680 3646 7718 3664
rect 7752 3646 7790 3664
rect 7824 3646 7862 3664
rect 7896 3646 7934 3664
rect 7968 3646 8006 3664
rect 8040 3646 8078 3664
rect 8112 3646 8150 3664
rect 8184 3646 8222 3664
rect 8256 3646 8294 3664
rect 8328 3646 8366 3664
rect 8400 3646 8438 3664
rect 8472 3646 8510 3664
rect 8544 3646 8582 3664
rect 8616 3646 8654 3664
rect 8688 3646 8726 3664
rect 8760 3646 8798 3664
rect 8832 3646 8870 3664
rect 8904 3646 8942 3664
rect 8976 3646 9014 3664
rect 9048 3646 9086 3664
rect 9120 3646 9158 3664
rect 9192 3646 9230 3664
rect 9264 3646 9302 3664
rect 9336 3646 9374 3664
rect 9408 3646 9446 3664
rect 9480 3646 9518 3664
rect 9552 3646 9590 3664
rect 9624 3646 9662 3664
rect 9696 3646 9734 3664
rect 9768 3646 9806 3664
rect 9840 3646 9878 3664
rect 9912 3646 9950 3664
rect 9984 3646 10022 3664
rect 10056 3646 10094 3664
rect 10128 3646 10166 3664
rect 10200 3646 10238 3664
rect 10272 3646 10310 3664
rect 10344 3646 10382 3664
rect 10416 3646 10454 3664
rect 10488 3646 10526 3664
rect 10560 3646 10598 3664
rect 10632 3646 10670 3664
rect 10704 3646 10742 3664
rect 10776 3646 10814 3664
rect 10848 3646 10886 3664
rect 10920 3646 10958 3664
rect 10992 3646 11030 3664
rect 11064 3646 11102 3664
rect 11136 3646 11174 3664
rect 7319 3612 7421 3646
rect 7462 3630 7489 3646
rect 7535 3630 7557 3646
rect 7608 3630 7625 3646
rect 7680 3630 7693 3646
rect 7752 3630 7761 3646
rect 7824 3630 7829 3646
rect 7896 3630 7897 3646
rect 7455 3612 7489 3630
rect 7523 3612 7557 3630
rect 7591 3612 7625 3630
rect 7659 3612 7693 3630
rect 7727 3612 7761 3630
rect 7795 3612 7829 3630
rect 7863 3612 7897 3630
rect 7931 3630 7934 3646
rect 7999 3630 8006 3646
rect 8067 3630 8078 3646
rect 8135 3630 8150 3646
rect 8203 3630 8222 3646
rect 8271 3630 8294 3646
rect 8339 3630 8366 3646
rect 8407 3630 8438 3646
rect 7931 3612 7965 3630
rect 7999 3612 8033 3630
rect 8067 3612 8101 3630
rect 8135 3612 8169 3630
rect 8203 3612 8237 3630
rect 8271 3612 8305 3630
rect 8339 3612 8373 3630
rect 8407 3612 8441 3630
rect 8475 3612 8509 3646
rect 8544 3630 8577 3646
rect 8616 3630 8645 3646
rect 8688 3630 8713 3646
rect 8760 3630 8781 3646
rect 8832 3630 8849 3646
rect 8904 3630 8917 3646
rect 8976 3630 8985 3646
rect 9048 3630 9053 3646
rect 9120 3630 9121 3646
rect 8543 3612 8577 3630
rect 8611 3612 8645 3630
rect 8679 3612 8713 3630
rect 8747 3612 8781 3630
rect 8815 3612 8849 3630
rect 8883 3612 8917 3630
rect 8951 3612 8985 3630
rect 9019 3612 9053 3630
rect 9087 3612 9121 3630
rect 9155 3630 9158 3646
rect 9223 3630 9230 3646
rect 9291 3630 9302 3646
rect 9359 3630 9374 3646
rect 9427 3630 9446 3646
rect 9495 3630 9518 3646
rect 9563 3630 9590 3646
rect 9631 3630 9662 3646
rect 9155 3612 9189 3630
rect 9223 3612 9257 3630
rect 9291 3612 9325 3630
rect 9359 3612 9393 3630
rect 9427 3612 9461 3630
rect 9495 3612 9529 3630
rect 9563 3612 9597 3630
rect 9631 3612 9665 3630
rect 9699 3612 9733 3646
rect 9768 3630 9801 3646
rect 9840 3630 9869 3646
rect 9912 3630 9937 3646
rect 9984 3630 10005 3646
rect 10056 3630 10073 3646
rect 10128 3630 10141 3646
rect 10200 3630 10209 3646
rect 10272 3630 10277 3646
rect 10344 3630 10345 3646
rect 9767 3612 9801 3630
rect 9835 3612 9869 3630
rect 9903 3612 9937 3630
rect 9971 3612 10005 3630
rect 10039 3612 10073 3630
rect 10107 3612 10141 3630
rect 10175 3612 10209 3630
rect 10243 3612 10277 3630
rect 10311 3612 10345 3630
rect 10379 3630 10382 3646
rect 10447 3630 10454 3646
rect 10515 3630 10526 3646
rect 10583 3630 10598 3646
rect 10651 3630 10670 3646
rect 10719 3630 10742 3646
rect 10787 3630 10814 3646
rect 10855 3630 10886 3646
rect 10379 3612 10413 3630
rect 10447 3612 10481 3630
rect 10515 3612 10549 3630
rect 10583 3612 10617 3630
rect 10651 3612 10685 3630
rect 10719 3612 10753 3630
rect 10787 3612 10821 3630
rect 10855 3612 10889 3630
rect 10923 3612 10957 3646
rect 10992 3630 11025 3646
rect 11064 3630 11093 3646
rect 11136 3630 11161 3646
rect 11208 3630 11313 3664
rect 10991 3612 11025 3630
rect 11059 3612 11093 3630
rect 11127 3612 11161 3630
rect 11195 3612 11313 3630
rect 7319 3580 11313 3612
rect 7319 3557 7411 3580
rect 7319 3536 7353 3557
rect 7319 3502 7350 3536
rect 7387 3523 7411 3557
rect 7384 3502 7411 3523
rect 7319 3489 7411 3502
rect 7319 3464 7353 3489
rect 7319 3430 7350 3464
rect 7387 3455 7411 3489
rect 11231 3557 11313 3580
rect 11231 3536 11255 3557
rect 11231 3502 11252 3536
rect 11289 3523 11313 3557
rect 11286 3502 11313 3523
rect 11231 3489 11313 3502
rect 7384 3430 7411 3455
rect 7319 3421 7411 3430
rect 7319 3392 7353 3421
rect 7319 3358 7350 3392
rect 7387 3387 7411 3421
rect 7384 3358 7411 3387
rect 7319 3353 7411 3358
rect 7319 3320 7353 3353
rect 7319 3286 7350 3320
rect 7387 3319 7411 3353
rect 7384 3286 7411 3319
rect 7319 3285 7411 3286
rect 7319 3251 7353 3285
rect 7387 3251 7411 3285
rect 7319 3248 7411 3251
rect 7319 3214 7350 3248
rect 7384 3217 7411 3248
rect 7319 3183 7353 3214
rect 7387 3183 7411 3217
rect 7319 3176 7411 3183
rect 7319 3142 7350 3176
rect 7384 3149 7411 3176
rect 7319 3115 7353 3142
rect 7387 3115 7411 3149
rect 7319 3104 7411 3115
rect 7319 3070 7350 3104
rect 7384 3081 7411 3104
rect 7319 3047 7353 3070
rect 7387 3047 7411 3081
rect 7319 3032 7411 3047
rect 7319 2998 7350 3032
rect 7384 3013 7411 3032
rect 7319 2979 7353 2998
rect 7387 2979 7411 3013
rect 7319 2960 7411 2979
rect 7319 2926 7350 2960
rect 7384 2945 7411 2960
rect 7319 2911 7353 2926
rect 7387 2911 7411 2945
rect 7319 2888 7411 2911
rect 7319 2854 7350 2888
rect 7384 2877 7411 2888
rect 7319 2843 7353 2854
rect 7387 2843 7411 2877
rect 7319 2816 7411 2843
rect 7319 2782 7350 2816
rect 7384 2809 7411 2816
rect 7319 2775 7353 2782
rect 7387 2775 7411 2809
rect 7319 2744 7411 2775
rect 7319 2710 7350 2744
rect 7384 2741 7411 2744
rect 7319 2707 7353 2710
rect 7387 2707 7411 2741
rect 7319 2673 7411 2707
rect 7319 2672 7353 2673
rect 7319 2638 7350 2672
rect 7387 2639 7411 2673
rect 7384 2638 7411 2639
rect 7319 2605 7411 2638
rect 7319 2600 7353 2605
rect 7319 2566 7350 2600
rect 7387 2571 7411 2605
rect 7384 2566 7411 2571
rect 7319 2537 7411 2566
rect 7319 2528 7353 2537
rect 7319 2494 7350 2528
rect 7387 2503 7411 2537
rect 7384 2494 7411 2503
rect 7319 2469 7411 2494
rect 7319 2456 7353 2469
rect 7319 2422 7350 2456
rect 7387 2435 7411 2469
rect 7384 2422 7411 2435
rect 7319 2401 7411 2422
rect 7319 2384 7353 2401
rect 7319 2350 7350 2384
rect 7387 2367 7411 2401
rect 7384 2350 7411 2367
rect 7319 2333 7411 2350
rect 7319 2312 7353 2333
rect 7319 2278 7350 2312
rect 7387 2299 7411 2333
rect 7384 2278 7411 2299
rect 7319 2265 7411 2278
rect 7319 2240 7353 2265
rect 7319 2206 7350 2240
rect 7387 2231 7411 2265
rect 7384 2206 7411 2231
rect 7319 2197 7411 2206
rect 7319 2168 7353 2197
rect 7319 2134 7350 2168
rect 7387 2163 7411 2197
rect 7384 2134 7411 2163
rect 7319 2129 7411 2134
rect 7319 2096 7353 2129
rect 7319 2062 7350 2096
rect 7387 2095 7411 2129
rect 7384 2062 7411 2095
rect 7319 2061 7411 2062
rect 7319 2027 7353 2061
rect 7387 2027 7411 2061
rect 7319 2024 7411 2027
rect 7319 1990 7350 2024
rect 7384 1993 7411 2024
rect 7319 1959 7353 1990
rect 7387 1959 7411 1993
rect 7319 1952 7411 1959
rect 7319 1918 7350 1952
rect 7384 1925 7411 1952
rect 7319 1891 7353 1918
rect 7387 1891 7411 1925
rect 7319 1880 7411 1891
rect 7319 1846 7350 1880
rect 7384 1857 7411 1880
rect 7319 1823 7353 1846
rect 7387 1823 7411 1857
rect 7319 1808 7411 1823
rect 7319 1774 7350 1808
rect 7384 1789 7411 1808
rect 7319 1755 7353 1774
rect 7387 1755 7411 1789
rect 7319 1736 7411 1755
rect 7319 1702 7350 1736
rect 7384 1721 7411 1736
rect 7319 1687 7353 1702
rect 7387 1687 7411 1721
rect 7319 1664 7411 1687
rect 7319 1630 7350 1664
rect 7384 1653 7411 1664
rect 7319 1619 7353 1630
rect 7387 1619 7411 1653
rect 7319 1592 7411 1619
rect 7319 1558 7350 1592
rect 7384 1585 7411 1592
rect 7319 1551 7353 1558
rect 7387 1551 7411 1585
rect 7319 1520 7411 1551
rect 7319 1486 7350 1520
rect 7384 1517 7411 1520
rect 7319 1483 7353 1486
rect 7387 1483 7411 1517
rect 7319 1449 7411 1483
rect 7319 1448 7353 1449
rect 7319 1414 7350 1448
rect 7387 1415 7411 1449
rect 7384 1414 7411 1415
rect 7319 1381 7411 1414
rect 7319 1376 7353 1381
rect 7319 1342 7350 1376
rect 7387 1347 7411 1381
rect 7384 1342 7411 1347
rect 7319 1313 7411 1342
rect 7319 1304 7353 1313
rect 7319 1270 7350 1304
rect 7387 1279 7411 1313
rect 7384 1270 7411 1279
rect 7319 1245 7411 1270
rect 7319 1232 7353 1245
rect 7319 1198 7350 1232
rect 7387 1211 7411 1245
rect 7384 1198 7411 1211
rect 7319 1177 7411 1198
rect 7319 1160 7353 1177
rect 7319 1126 7350 1160
rect 7387 1143 7411 1177
rect 7384 1126 7411 1143
rect 7319 1109 7411 1126
rect 7319 1088 7353 1109
rect 7319 1054 7350 1088
rect 7387 1075 7411 1109
rect 7384 1054 7411 1075
rect 7319 1041 7411 1054
rect 7319 1016 7353 1041
rect 7319 982 7350 1016
rect 7387 1007 7411 1041
rect 7384 982 7411 1007
rect 7319 973 7411 982
rect 7319 944 7353 973
rect 7319 910 7350 944
rect 7387 939 7411 973
rect 7384 910 7411 939
rect 7319 905 7411 910
rect 7319 872 7353 905
rect 7319 838 7350 872
rect 7387 871 7411 905
rect 7384 838 7411 871
rect 7319 837 7411 838
rect 7319 803 7353 837
rect 7387 803 7411 837
rect 7319 800 7411 803
rect 7319 766 7350 800
rect 7384 769 7411 800
rect 7319 735 7353 766
rect 7387 735 7411 769
rect 7319 728 7411 735
rect 7319 694 7350 728
rect 7384 701 7411 728
rect 7319 667 7353 694
rect 7387 667 7411 701
rect 7319 656 7411 667
rect 7319 622 7350 656
rect 7384 633 7411 656
rect 7319 599 7353 622
rect 7387 599 7411 633
rect 7319 565 7411 599
rect 7319 531 7353 565
rect 7387 531 7411 565
rect 7319 497 7411 531
rect 7319 463 7353 497
rect 7387 463 7411 497
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
rect 11231 3464 11255 3489
rect 11231 3430 11252 3464
rect 11289 3455 11313 3489
rect 11286 3430 11313 3455
rect 11231 3421 11313 3430
rect 11231 3392 11255 3421
rect 11231 3358 11252 3392
rect 11289 3387 11313 3421
rect 11286 3358 11313 3387
rect 11231 3353 11313 3358
rect 11231 3320 11255 3353
rect 11231 3286 11252 3320
rect 11289 3319 11313 3353
rect 11286 3286 11313 3319
rect 11231 3285 11313 3286
rect 11231 3251 11255 3285
rect 11289 3251 11313 3285
rect 11231 3248 11313 3251
rect 11231 3214 11252 3248
rect 11286 3217 11313 3248
rect 11231 3183 11255 3214
rect 11289 3183 11313 3217
rect 11231 3176 11313 3183
rect 11231 3142 11252 3176
rect 11286 3149 11313 3176
rect 11231 3115 11255 3142
rect 11289 3115 11313 3149
rect 11231 3104 11313 3115
rect 11231 3070 11252 3104
rect 11286 3081 11313 3104
rect 11231 3047 11255 3070
rect 11289 3047 11313 3081
rect 11231 3032 11313 3047
rect 11231 2998 11252 3032
rect 11286 3013 11313 3032
rect 11231 2979 11255 2998
rect 11289 2979 11313 3013
rect 11231 2960 11313 2979
rect 11231 2926 11252 2960
rect 11286 2945 11313 2960
rect 11231 2911 11255 2926
rect 11289 2911 11313 2945
rect 11231 2888 11313 2911
rect 11231 2854 11252 2888
rect 11286 2877 11313 2888
rect 11231 2843 11255 2854
rect 11289 2843 11313 2877
rect 11231 2816 11313 2843
rect 11231 2782 11252 2816
rect 11286 2809 11313 2816
rect 11231 2775 11255 2782
rect 11289 2775 11313 2809
rect 11231 2744 11313 2775
rect 11231 2710 11252 2744
rect 11286 2741 11313 2744
rect 11231 2707 11255 2710
rect 11289 2707 11313 2741
rect 11231 2673 11313 2707
rect 11231 2672 11255 2673
rect 11231 2638 11252 2672
rect 11289 2639 11313 2673
rect 11286 2638 11313 2639
rect 11231 2605 11313 2638
rect 11231 2600 11255 2605
rect 11231 2566 11252 2600
rect 11289 2571 11313 2605
rect 11286 2566 11313 2571
rect 11231 2537 11313 2566
rect 11231 2528 11255 2537
rect 11231 2494 11252 2528
rect 11289 2503 11313 2537
rect 11286 2494 11313 2503
rect 11231 2469 11313 2494
rect 11231 2456 11255 2469
rect 11231 2422 11252 2456
rect 11289 2435 11313 2469
rect 11286 2422 11313 2435
rect 11231 2401 11313 2422
rect 11231 2384 11255 2401
rect 11231 2350 11252 2384
rect 11289 2367 11313 2401
rect 11286 2350 11313 2367
rect 11231 2333 11313 2350
rect 11231 2312 11255 2333
rect 11231 2278 11252 2312
rect 11289 2299 11313 2333
rect 11286 2278 11313 2299
rect 11231 2265 11313 2278
rect 11231 2240 11255 2265
rect 11231 2206 11252 2240
rect 11289 2231 11313 2265
rect 11286 2206 11313 2231
rect 11231 2197 11313 2206
rect 11231 2168 11255 2197
rect 11231 2134 11252 2168
rect 11289 2163 11313 2197
rect 11286 2134 11313 2163
rect 11231 2129 11313 2134
rect 11231 2096 11255 2129
rect 11231 2062 11252 2096
rect 11289 2095 11313 2129
rect 11286 2062 11313 2095
rect 11231 2061 11313 2062
rect 11231 2027 11255 2061
rect 11289 2027 11313 2061
rect 11231 2024 11313 2027
rect 11231 1990 11252 2024
rect 11286 1993 11313 2024
rect 11231 1959 11255 1990
rect 11289 1959 11313 1993
rect 11231 1952 11313 1959
rect 11231 1918 11252 1952
rect 11286 1925 11313 1952
rect 11231 1891 11255 1918
rect 11289 1891 11313 1925
rect 11231 1880 11313 1891
rect 11231 1846 11252 1880
rect 11286 1857 11313 1880
rect 11231 1823 11255 1846
rect 11289 1823 11313 1857
rect 11231 1808 11313 1823
rect 11231 1774 11252 1808
rect 11286 1789 11313 1808
rect 11231 1755 11255 1774
rect 11289 1755 11313 1789
rect 11231 1736 11313 1755
rect 11231 1702 11252 1736
rect 11286 1721 11313 1736
rect 11231 1687 11255 1702
rect 11289 1687 11313 1721
rect 11231 1664 11313 1687
rect 11231 1630 11252 1664
rect 11286 1653 11313 1664
rect 11231 1619 11255 1630
rect 11289 1619 11313 1653
rect 11231 1592 11313 1619
rect 11231 1558 11252 1592
rect 11286 1585 11313 1592
rect 11231 1551 11255 1558
rect 11289 1551 11313 1585
rect 11231 1520 11313 1551
rect 11231 1486 11252 1520
rect 11286 1517 11313 1520
rect 11231 1483 11255 1486
rect 11289 1483 11313 1517
rect 11231 1449 11313 1483
rect 11231 1448 11255 1449
rect 11231 1414 11252 1448
rect 11289 1415 11313 1449
rect 11286 1414 11313 1415
rect 11231 1381 11313 1414
rect 11231 1376 11255 1381
rect 11231 1342 11252 1376
rect 11289 1347 11313 1381
rect 11286 1342 11313 1347
rect 11231 1313 11313 1342
rect 11231 1304 11255 1313
rect 11231 1270 11252 1304
rect 11289 1279 11313 1313
rect 11286 1270 11313 1279
rect 11231 1245 11313 1270
rect 11231 1232 11255 1245
rect 11231 1198 11252 1232
rect 11289 1211 11313 1245
rect 11286 1198 11313 1211
rect 11231 1177 11313 1198
rect 11231 1160 11255 1177
rect 11231 1126 11252 1160
rect 11289 1143 11313 1177
rect 11286 1126 11313 1143
rect 11231 1109 11313 1126
rect 11231 1088 11255 1109
rect 11231 1054 11252 1088
rect 11289 1075 11313 1109
rect 11286 1054 11313 1075
rect 11231 1041 11313 1054
rect 11231 1016 11255 1041
rect 11231 982 11252 1016
rect 11289 1007 11313 1041
rect 11286 982 11313 1007
rect 11231 973 11313 982
rect 11231 944 11255 973
rect 11231 910 11252 944
rect 11289 939 11313 973
rect 11286 910 11313 939
rect 11231 905 11313 910
rect 11231 872 11255 905
rect 11231 838 11252 872
rect 11289 871 11313 905
rect 11286 838 11313 871
rect 11231 837 11313 838
rect 11231 803 11255 837
rect 11289 803 11313 837
rect 11231 800 11313 803
rect 11231 766 11252 800
rect 11286 769 11313 800
rect 11231 735 11255 766
rect 11289 735 11313 769
rect 11231 728 11313 735
rect 11231 694 11252 728
rect 11286 701 11313 728
rect 11231 667 11255 694
rect 11289 667 11313 701
rect 11231 656 11313 667
rect 11231 622 11252 656
rect 11286 633 11313 656
rect 11231 599 11255 622
rect 11289 599 11313 633
rect 11231 565 11313 599
rect 11231 531 11255 565
rect 11289 531 11313 565
rect 11231 497 11313 531
rect 7319 429 7411 463
rect 7319 395 7353 429
rect 7387 395 7411 429
rect 7319 364 7411 395
rect 11231 463 11255 497
rect 11289 463 11313 497
rect 11231 429 11313 463
rect 11231 395 11255 429
rect 11289 395 11313 429
rect 11231 364 11313 395
rect 7319 334 11313 364
rect 7319 300 7411 334
rect 7445 300 7479 334
rect 7513 300 7547 334
rect 7581 300 7615 334
rect 7649 300 7683 334
rect 7717 300 7751 334
rect 7785 300 7819 334
rect 7853 300 7887 334
rect 7921 300 7955 334
rect 7989 300 8023 334
rect 8057 300 8091 334
rect 8125 300 8159 334
rect 8193 300 8227 334
rect 8261 300 8295 334
rect 8329 300 8363 334
rect 8397 300 8431 334
rect 8465 300 8499 334
rect 8533 300 8567 334
rect 8601 300 8635 334
rect 8669 300 8703 334
rect 8737 300 8771 334
rect 8805 300 8839 334
rect 8873 300 8907 334
rect 8941 300 8975 334
rect 9009 300 9043 334
rect 9077 300 9111 334
rect 9145 300 9179 334
rect 9213 300 9247 334
rect 9281 300 9315 334
rect 9349 300 9383 334
rect 9417 300 9451 334
rect 9485 300 9519 334
rect 9553 300 9587 334
rect 9621 300 9655 334
rect 9689 300 9723 334
rect 9757 300 9791 334
rect 9825 300 9859 334
rect 9893 300 9927 334
rect 9961 300 9995 334
rect 10029 300 10063 334
rect 10097 300 10131 334
rect 10165 300 10199 334
rect 10233 300 10267 334
rect 10301 300 10335 334
rect 10369 300 10403 334
rect 10437 300 10471 334
rect 10505 300 10539 334
rect 10573 300 10607 334
rect 10641 300 10675 334
rect 10709 300 10743 334
rect 10777 300 10811 334
rect 10845 300 10879 334
rect 10913 300 10947 334
rect 10981 300 11015 334
rect 11049 300 11083 334
rect 11117 300 11151 334
rect 11185 300 11313 334
rect 7319 254 11313 300
<< viali >>
rect 7428 3646 7462 3664
rect 7501 3646 7535 3664
rect 7574 3646 7608 3664
rect 7646 3646 7680 3664
rect 7718 3646 7752 3664
rect 7790 3646 7824 3664
rect 7862 3646 7896 3664
rect 7934 3646 7968 3664
rect 8006 3646 8040 3664
rect 8078 3646 8112 3664
rect 8150 3646 8184 3664
rect 8222 3646 8256 3664
rect 8294 3646 8328 3664
rect 8366 3646 8400 3664
rect 8438 3646 8472 3664
rect 8510 3646 8544 3664
rect 8582 3646 8616 3664
rect 8654 3646 8688 3664
rect 8726 3646 8760 3664
rect 8798 3646 8832 3664
rect 8870 3646 8904 3664
rect 8942 3646 8976 3664
rect 9014 3646 9048 3664
rect 9086 3646 9120 3664
rect 9158 3646 9192 3664
rect 9230 3646 9264 3664
rect 9302 3646 9336 3664
rect 9374 3646 9408 3664
rect 9446 3646 9480 3664
rect 9518 3646 9552 3664
rect 9590 3646 9624 3664
rect 9662 3646 9696 3664
rect 9734 3646 9768 3664
rect 9806 3646 9840 3664
rect 9878 3646 9912 3664
rect 9950 3646 9984 3664
rect 10022 3646 10056 3664
rect 10094 3646 10128 3664
rect 10166 3646 10200 3664
rect 10238 3646 10272 3664
rect 10310 3646 10344 3664
rect 10382 3646 10416 3664
rect 10454 3646 10488 3664
rect 10526 3646 10560 3664
rect 10598 3646 10632 3664
rect 10670 3646 10704 3664
rect 10742 3646 10776 3664
rect 10814 3646 10848 3664
rect 10886 3646 10920 3664
rect 10958 3646 10992 3664
rect 11030 3646 11064 3664
rect 11102 3646 11136 3664
rect 11174 3646 11208 3664
rect 7428 3630 7455 3646
rect 7455 3630 7462 3646
rect 7501 3630 7523 3646
rect 7523 3630 7535 3646
rect 7574 3630 7591 3646
rect 7591 3630 7608 3646
rect 7646 3630 7659 3646
rect 7659 3630 7680 3646
rect 7718 3630 7727 3646
rect 7727 3630 7752 3646
rect 7790 3630 7795 3646
rect 7795 3630 7824 3646
rect 7862 3630 7863 3646
rect 7863 3630 7896 3646
rect 7934 3630 7965 3646
rect 7965 3630 7968 3646
rect 8006 3630 8033 3646
rect 8033 3630 8040 3646
rect 8078 3630 8101 3646
rect 8101 3630 8112 3646
rect 8150 3630 8169 3646
rect 8169 3630 8184 3646
rect 8222 3630 8237 3646
rect 8237 3630 8256 3646
rect 8294 3630 8305 3646
rect 8305 3630 8328 3646
rect 8366 3630 8373 3646
rect 8373 3630 8400 3646
rect 8438 3630 8441 3646
rect 8441 3630 8472 3646
rect 8510 3630 8543 3646
rect 8543 3630 8544 3646
rect 8582 3630 8611 3646
rect 8611 3630 8616 3646
rect 8654 3630 8679 3646
rect 8679 3630 8688 3646
rect 8726 3630 8747 3646
rect 8747 3630 8760 3646
rect 8798 3630 8815 3646
rect 8815 3630 8832 3646
rect 8870 3630 8883 3646
rect 8883 3630 8904 3646
rect 8942 3630 8951 3646
rect 8951 3630 8976 3646
rect 9014 3630 9019 3646
rect 9019 3630 9048 3646
rect 9086 3630 9087 3646
rect 9087 3630 9120 3646
rect 9158 3630 9189 3646
rect 9189 3630 9192 3646
rect 9230 3630 9257 3646
rect 9257 3630 9264 3646
rect 9302 3630 9325 3646
rect 9325 3630 9336 3646
rect 9374 3630 9393 3646
rect 9393 3630 9408 3646
rect 9446 3630 9461 3646
rect 9461 3630 9480 3646
rect 9518 3630 9529 3646
rect 9529 3630 9552 3646
rect 9590 3630 9597 3646
rect 9597 3630 9624 3646
rect 9662 3630 9665 3646
rect 9665 3630 9696 3646
rect 9734 3630 9767 3646
rect 9767 3630 9768 3646
rect 9806 3630 9835 3646
rect 9835 3630 9840 3646
rect 9878 3630 9903 3646
rect 9903 3630 9912 3646
rect 9950 3630 9971 3646
rect 9971 3630 9984 3646
rect 10022 3630 10039 3646
rect 10039 3630 10056 3646
rect 10094 3630 10107 3646
rect 10107 3630 10128 3646
rect 10166 3630 10175 3646
rect 10175 3630 10200 3646
rect 10238 3630 10243 3646
rect 10243 3630 10272 3646
rect 10310 3630 10311 3646
rect 10311 3630 10344 3646
rect 10382 3630 10413 3646
rect 10413 3630 10416 3646
rect 10454 3630 10481 3646
rect 10481 3630 10488 3646
rect 10526 3630 10549 3646
rect 10549 3630 10560 3646
rect 10598 3630 10617 3646
rect 10617 3630 10632 3646
rect 10670 3630 10685 3646
rect 10685 3630 10704 3646
rect 10742 3630 10753 3646
rect 10753 3630 10776 3646
rect 10814 3630 10821 3646
rect 10821 3630 10848 3646
rect 10886 3630 10889 3646
rect 10889 3630 10920 3646
rect 10958 3630 10991 3646
rect 10991 3630 10992 3646
rect 11030 3630 11059 3646
rect 11059 3630 11064 3646
rect 11102 3630 11127 3646
rect 11127 3630 11136 3646
rect 11174 3630 11195 3646
rect 11195 3630 11208 3646
rect 7350 3523 7353 3536
rect 7353 3523 7384 3536
rect 7350 3502 7384 3523
rect 7350 3455 7353 3464
rect 7353 3455 7384 3464
rect 11252 3523 11255 3536
rect 11255 3523 11286 3536
rect 11252 3502 11286 3523
rect 7350 3430 7384 3455
rect 7350 3387 7353 3392
rect 7353 3387 7384 3392
rect 7350 3358 7384 3387
rect 7350 3319 7353 3320
rect 7353 3319 7384 3320
rect 7350 3286 7384 3319
rect 7350 3217 7384 3248
rect 7350 3214 7353 3217
rect 7353 3214 7384 3217
rect 7350 3149 7384 3176
rect 7350 3142 7353 3149
rect 7353 3142 7384 3149
rect 7350 3081 7384 3104
rect 7350 3070 7353 3081
rect 7353 3070 7384 3081
rect 7350 3013 7384 3032
rect 7350 2998 7353 3013
rect 7353 2998 7384 3013
rect 7350 2945 7384 2960
rect 7350 2926 7353 2945
rect 7353 2926 7384 2945
rect 7350 2877 7384 2888
rect 7350 2854 7353 2877
rect 7353 2854 7384 2877
rect 7350 2809 7384 2816
rect 7350 2782 7353 2809
rect 7353 2782 7384 2809
rect 7350 2741 7384 2744
rect 7350 2710 7353 2741
rect 7353 2710 7384 2741
rect 7350 2639 7353 2672
rect 7353 2639 7384 2672
rect 7350 2638 7384 2639
rect 7350 2571 7353 2600
rect 7353 2571 7384 2600
rect 7350 2566 7384 2571
rect 7350 2503 7353 2528
rect 7353 2503 7384 2528
rect 7350 2494 7384 2503
rect 7350 2435 7353 2456
rect 7353 2435 7384 2456
rect 7350 2422 7384 2435
rect 7350 2367 7353 2384
rect 7353 2367 7384 2384
rect 7350 2350 7384 2367
rect 7350 2299 7353 2312
rect 7353 2299 7384 2312
rect 7350 2278 7384 2299
rect 7350 2231 7353 2240
rect 7353 2231 7384 2240
rect 7350 2206 7384 2231
rect 7350 2163 7353 2168
rect 7353 2163 7384 2168
rect 7350 2134 7384 2163
rect 7350 2095 7353 2096
rect 7353 2095 7384 2096
rect 7350 2062 7384 2095
rect 7350 1993 7384 2024
rect 7350 1990 7353 1993
rect 7353 1990 7384 1993
rect 7350 1925 7384 1952
rect 7350 1918 7353 1925
rect 7353 1918 7384 1925
rect 7350 1857 7384 1880
rect 7350 1846 7353 1857
rect 7353 1846 7384 1857
rect 7350 1789 7384 1808
rect 7350 1774 7353 1789
rect 7353 1774 7384 1789
rect 7350 1721 7384 1736
rect 7350 1702 7353 1721
rect 7353 1702 7384 1721
rect 7350 1653 7384 1664
rect 7350 1630 7353 1653
rect 7353 1630 7384 1653
rect 7350 1585 7384 1592
rect 7350 1558 7353 1585
rect 7353 1558 7384 1585
rect 7350 1517 7384 1520
rect 7350 1486 7353 1517
rect 7353 1486 7384 1517
rect 7350 1415 7353 1448
rect 7353 1415 7384 1448
rect 7350 1414 7384 1415
rect 7350 1347 7353 1376
rect 7353 1347 7384 1376
rect 7350 1342 7384 1347
rect 7350 1279 7353 1304
rect 7353 1279 7384 1304
rect 7350 1270 7384 1279
rect 7350 1211 7353 1232
rect 7353 1211 7384 1232
rect 7350 1198 7384 1211
rect 7350 1143 7353 1160
rect 7353 1143 7384 1160
rect 7350 1126 7384 1143
rect 7350 1075 7353 1088
rect 7353 1075 7384 1088
rect 7350 1054 7384 1075
rect 7350 1007 7353 1016
rect 7353 1007 7384 1016
rect 7350 982 7384 1007
rect 7350 939 7353 944
rect 7353 939 7384 944
rect 7350 910 7384 939
rect 7350 871 7353 872
rect 7353 871 7384 872
rect 7350 838 7384 871
rect 7350 769 7384 800
rect 7350 766 7353 769
rect 7353 766 7384 769
rect 7350 701 7384 728
rect 7350 694 7353 701
rect 7353 694 7384 701
rect 7350 633 7384 656
rect 7350 622 7353 633
rect 7353 622 7384 633
rect 7584 3303 7618 3337
rect 7656 3303 7690 3337
rect 7728 3303 7762 3337
rect 7584 3207 7618 3241
rect 7656 3207 7690 3241
rect 7728 3207 7762 3241
rect 7584 3111 7618 3145
rect 7656 3111 7690 3145
rect 7728 3111 7762 3145
rect 7584 3015 7618 3049
rect 7656 3015 7690 3049
rect 7728 3015 7762 3049
rect 7584 2919 7618 2953
rect 7656 2919 7690 2953
rect 7728 2919 7762 2953
rect 7584 2823 7618 2857
rect 7656 2823 7690 2857
rect 7728 2823 7762 2857
rect 7584 2727 7618 2761
rect 7656 2727 7690 2761
rect 7728 2727 7762 2761
rect 7584 2631 7618 2665
rect 7656 2631 7690 2665
rect 7728 2631 7762 2665
rect 7584 2535 7618 2569
rect 7656 2535 7690 2569
rect 7728 2535 7762 2569
rect 7584 2439 7618 2473
rect 7656 2439 7690 2473
rect 7728 2439 7762 2473
rect 7584 2343 7618 2377
rect 7656 2343 7690 2377
rect 7728 2343 7762 2377
rect 7584 2247 7618 2281
rect 7656 2247 7690 2281
rect 7728 2247 7762 2281
rect 7584 2151 7618 2185
rect 7656 2151 7690 2185
rect 7728 2151 7762 2185
rect 7584 2055 7618 2089
rect 7656 2055 7690 2089
rect 7728 2055 7762 2089
rect 7584 1959 7618 1993
rect 7656 1959 7690 1993
rect 7728 1959 7762 1993
rect 7584 1863 7618 1897
rect 7656 1863 7690 1897
rect 7728 1863 7762 1897
rect 7584 1767 7618 1801
rect 7656 1767 7690 1801
rect 7728 1767 7762 1801
rect 7584 1671 7618 1705
rect 7656 1671 7690 1705
rect 7728 1671 7762 1705
rect 7584 1575 7618 1609
rect 7656 1575 7690 1609
rect 7728 1575 7762 1609
rect 7584 1479 7618 1513
rect 7656 1479 7690 1513
rect 7728 1479 7762 1513
rect 7584 1383 7618 1417
rect 7656 1383 7690 1417
rect 7728 1383 7762 1417
rect 7584 1287 7618 1321
rect 7656 1287 7690 1321
rect 7728 1287 7762 1321
rect 7584 1191 7618 1225
rect 7656 1191 7690 1225
rect 7728 1191 7762 1225
rect 7584 1095 7618 1129
rect 7656 1095 7690 1129
rect 7728 1095 7762 1129
rect 7584 999 7618 1033
rect 7656 999 7690 1033
rect 7728 999 7762 1033
rect 7584 903 7618 937
rect 7656 903 7690 937
rect 7728 903 7762 937
rect 7584 807 7618 841
rect 7656 807 7690 841
rect 7728 807 7762 841
rect 7584 711 7618 745
rect 7656 711 7690 745
rect 7728 711 7762 745
rect 7584 615 7618 649
rect 7656 615 7690 649
rect 7728 615 7762 649
rect 7996 3303 8030 3337
rect 8068 3303 8102 3337
rect 8140 3303 8174 3337
rect 7996 3207 8030 3241
rect 8068 3207 8102 3241
rect 8140 3207 8174 3241
rect 7996 3111 8030 3145
rect 8068 3111 8102 3145
rect 8140 3111 8174 3145
rect 7996 3015 8030 3049
rect 8068 3015 8102 3049
rect 8140 3015 8174 3049
rect 7996 2919 8030 2953
rect 8068 2919 8102 2953
rect 8140 2919 8174 2953
rect 7996 2823 8030 2857
rect 8068 2823 8102 2857
rect 8140 2823 8174 2857
rect 7996 2727 8030 2761
rect 8068 2727 8102 2761
rect 8140 2727 8174 2761
rect 7996 2631 8030 2665
rect 8068 2631 8102 2665
rect 8140 2631 8174 2665
rect 7996 2535 8030 2569
rect 8068 2535 8102 2569
rect 8140 2535 8174 2569
rect 7996 2439 8030 2473
rect 8068 2439 8102 2473
rect 8140 2439 8174 2473
rect 7996 2343 8030 2377
rect 8068 2343 8102 2377
rect 8140 2343 8174 2377
rect 7996 2247 8030 2281
rect 8068 2247 8102 2281
rect 8140 2247 8174 2281
rect 7996 2151 8030 2185
rect 8068 2151 8102 2185
rect 8140 2151 8174 2185
rect 7996 2055 8030 2089
rect 8068 2055 8102 2089
rect 8140 2055 8174 2089
rect 7996 1959 8030 1993
rect 8068 1959 8102 1993
rect 8140 1959 8174 1993
rect 7996 1863 8030 1897
rect 8068 1863 8102 1897
rect 8140 1863 8174 1897
rect 7996 1767 8030 1801
rect 8068 1767 8102 1801
rect 8140 1767 8174 1801
rect 7996 1671 8030 1705
rect 8068 1671 8102 1705
rect 8140 1671 8174 1705
rect 7996 1575 8030 1609
rect 8068 1575 8102 1609
rect 8140 1575 8174 1609
rect 7996 1479 8030 1513
rect 8068 1479 8102 1513
rect 8140 1479 8174 1513
rect 7996 1383 8030 1417
rect 8068 1383 8102 1417
rect 8140 1383 8174 1417
rect 7996 1287 8030 1321
rect 8068 1287 8102 1321
rect 8140 1287 8174 1321
rect 7996 1191 8030 1225
rect 8068 1191 8102 1225
rect 8140 1191 8174 1225
rect 7996 1095 8030 1129
rect 8068 1095 8102 1129
rect 8140 1095 8174 1129
rect 7996 999 8030 1033
rect 8068 999 8102 1033
rect 8140 999 8174 1033
rect 7996 903 8030 937
rect 8068 903 8102 937
rect 8140 903 8174 937
rect 7996 807 8030 841
rect 8068 807 8102 841
rect 8140 807 8174 841
rect 7996 711 8030 745
rect 8068 711 8102 745
rect 8140 711 8174 745
rect 7996 615 8030 649
rect 8068 615 8102 649
rect 8140 615 8174 649
rect 8408 3303 8442 3337
rect 8480 3303 8514 3337
rect 8552 3303 8586 3337
rect 8408 3207 8442 3241
rect 8480 3207 8514 3241
rect 8552 3207 8586 3241
rect 8408 3111 8442 3145
rect 8480 3111 8514 3145
rect 8552 3111 8586 3145
rect 8408 3015 8442 3049
rect 8480 3015 8514 3049
rect 8552 3015 8586 3049
rect 8408 2919 8442 2953
rect 8480 2919 8514 2953
rect 8552 2919 8586 2953
rect 8408 2823 8442 2857
rect 8480 2823 8514 2857
rect 8552 2823 8586 2857
rect 8408 2727 8442 2761
rect 8480 2727 8514 2761
rect 8552 2727 8586 2761
rect 8408 2631 8442 2665
rect 8480 2631 8514 2665
rect 8552 2631 8586 2665
rect 8408 2535 8442 2569
rect 8480 2535 8514 2569
rect 8552 2535 8586 2569
rect 8408 2439 8442 2473
rect 8480 2439 8514 2473
rect 8552 2439 8586 2473
rect 8408 2343 8442 2377
rect 8480 2343 8514 2377
rect 8552 2343 8586 2377
rect 8408 2247 8442 2281
rect 8480 2247 8514 2281
rect 8552 2247 8586 2281
rect 8408 2151 8442 2185
rect 8480 2151 8514 2185
rect 8552 2151 8586 2185
rect 8408 2055 8442 2089
rect 8480 2055 8514 2089
rect 8552 2055 8586 2089
rect 8408 1959 8442 1993
rect 8480 1959 8514 1993
rect 8552 1959 8586 1993
rect 8408 1863 8442 1897
rect 8480 1863 8514 1897
rect 8552 1863 8586 1897
rect 8408 1767 8442 1801
rect 8480 1767 8514 1801
rect 8552 1767 8586 1801
rect 8408 1671 8442 1705
rect 8480 1671 8514 1705
rect 8552 1671 8586 1705
rect 8408 1575 8442 1609
rect 8480 1575 8514 1609
rect 8552 1575 8586 1609
rect 8408 1479 8442 1513
rect 8480 1479 8514 1513
rect 8552 1479 8586 1513
rect 8408 1383 8442 1417
rect 8480 1383 8514 1417
rect 8552 1383 8586 1417
rect 8408 1287 8442 1321
rect 8480 1287 8514 1321
rect 8552 1287 8586 1321
rect 8408 1191 8442 1225
rect 8480 1191 8514 1225
rect 8552 1191 8586 1225
rect 8408 1095 8442 1129
rect 8480 1095 8514 1129
rect 8552 1095 8586 1129
rect 8408 999 8442 1033
rect 8480 999 8514 1033
rect 8552 999 8586 1033
rect 8408 903 8442 937
rect 8480 903 8514 937
rect 8552 903 8586 937
rect 8408 807 8442 841
rect 8480 807 8514 841
rect 8552 807 8586 841
rect 8408 711 8442 745
rect 8480 711 8514 745
rect 8552 711 8586 745
rect 8408 615 8442 649
rect 8480 615 8514 649
rect 8552 615 8586 649
rect 8820 3303 8854 3337
rect 8892 3303 8926 3337
rect 8964 3303 8998 3337
rect 8820 3207 8854 3241
rect 8892 3207 8926 3241
rect 8964 3207 8998 3241
rect 8820 3111 8854 3145
rect 8892 3111 8926 3145
rect 8964 3111 8998 3145
rect 8820 3015 8854 3049
rect 8892 3015 8926 3049
rect 8964 3015 8998 3049
rect 8820 2919 8854 2953
rect 8892 2919 8926 2953
rect 8964 2919 8998 2953
rect 8820 2823 8854 2857
rect 8892 2823 8926 2857
rect 8964 2823 8998 2857
rect 8820 2727 8854 2761
rect 8892 2727 8926 2761
rect 8964 2727 8998 2761
rect 8820 2631 8854 2665
rect 8892 2631 8926 2665
rect 8964 2631 8998 2665
rect 8820 2535 8854 2569
rect 8892 2535 8926 2569
rect 8964 2535 8998 2569
rect 8820 2439 8854 2473
rect 8892 2439 8926 2473
rect 8964 2439 8998 2473
rect 8820 2343 8854 2377
rect 8892 2343 8926 2377
rect 8964 2343 8998 2377
rect 8820 2247 8854 2281
rect 8892 2247 8926 2281
rect 8964 2247 8998 2281
rect 8820 2151 8854 2185
rect 8892 2151 8926 2185
rect 8964 2151 8998 2185
rect 8820 2055 8854 2089
rect 8892 2055 8926 2089
rect 8964 2055 8998 2089
rect 8820 1959 8854 1993
rect 8892 1959 8926 1993
rect 8964 1959 8998 1993
rect 8820 1863 8854 1897
rect 8892 1863 8926 1897
rect 8964 1863 8998 1897
rect 8820 1767 8854 1801
rect 8892 1767 8926 1801
rect 8964 1767 8998 1801
rect 8820 1671 8854 1705
rect 8892 1671 8926 1705
rect 8964 1671 8998 1705
rect 8820 1575 8854 1609
rect 8892 1575 8926 1609
rect 8964 1575 8998 1609
rect 8820 1479 8854 1513
rect 8892 1479 8926 1513
rect 8964 1479 8998 1513
rect 8820 1383 8854 1417
rect 8892 1383 8926 1417
rect 8964 1383 8998 1417
rect 8820 1287 8854 1321
rect 8892 1287 8926 1321
rect 8964 1287 8998 1321
rect 8820 1191 8854 1225
rect 8892 1191 8926 1225
rect 8964 1191 8998 1225
rect 8820 1095 8854 1129
rect 8892 1095 8926 1129
rect 8964 1095 8998 1129
rect 8820 999 8854 1033
rect 8892 999 8926 1033
rect 8964 999 8998 1033
rect 8820 903 8854 937
rect 8892 903 8926 937
rect 8964 903 8998 937
rect 8820 807 8854 841
rect 8892 807 8926 841
rect 8964 807 8998 841
rect 8820 711 8854 745
rect 8892 711 8926 745
rect 8964 711 8998 745
rect 8820 615 8854 649
rect 8892 615 8926 649
rect 8964 615 8998 649
rect 9232 3303 9266 3337
rect 9304 3303 9338 3337
rect 9376 3303 9410 3337
rect 9232 3207 9266 3241
rect 9304 3207 9338 3241
rect 9376 3207 9410 3241
rect 9232 3111 9266 3145
rect 9304 3111 9338 3145
rect 9376 3111 9410 3145
rect 9232 3015 9266 3049
rect 9304 3015 9338 3049
rect 9376 3015 9410 3049
rect 9232 2919 9266 2953
rect 9304 2919 9338 2953
rect 9376 2919 9410 2953
rect 9232 2823 9266 2857
rect 9304 2823 9338 2857
rect 9376 2823 9410 2857
rect 9232 2727 9266 2761
rect 9304 2727 9338 2761
rect 9376 2727 9410 2761
rect 9232 2631 9266 2665
rect 9304 2631 9338 2665
rect 9376 2631 9410 2665
rect 9232 2535 9266 2569
rect 9304 2535 9338 2569
rect 9376 2535 9410 2569
rect 9232 2439 9266 2473
rect 9304 2439 9338 2473
rect 9376 2439 9410 2473
rect 9232 2343 9266 2377
rect 9304 2343 9338 2377
rect 9376 2343 9410 2377
rect 9232 2247 9266 2281
rect 9304 2247 9338 2281
rect 9376 2247 9410 2281
rect 9232 2151 9266 2185
rect 9304 2151 9338 2185
rect 9376 2151 9410 2185
rect 9232 2055 9266 2089
rect 9304 2055 9338 2089
rect 9376 2055 9410 2089
rect 9232 1959 9266 1993
rect 9304 1959 9338 1993
rect 9376 1959 9410 1993
rect 9232 1863 9266 1897
rect 9304 1863 9338 1897
rect 9376 1863 9410 1897
rect 9232 1767 9266 1801
rect 9304 1767 9338 1801
rect 9376 1767 9410 1801
rect 9232 1671 9266 1705
rect 9304 1671 9338 1705
rect 9376 1671 9410 1705
rect 9232 1575 9266 1609
rect 9304 1575 9338 1609
rect 9376 1575 9410 1609
rect 9232 1479 9266 1513
rect 9304 1479 9338 1513
rect 9376 1479 9410 1513
rect 9232 1383 9266 1417
rect 9304 1383 9338 1417
rect 9376 1383 9410 1417
rect 9232 1287 9266 1321
rect 9304 1287 9338 1321
rect 9376 1287 9410 1321
rect 9232 1191 9266 1225
rect 9304 1191 9338 1225
rect 9376 1191 9410 1225
rect 9232 1095 9266 1129
rect 9304 1095 9338 1129
rect 9376 1095 9410 1129
rect 9232 999 9266 1033
rect 9304 999 9338 1033
rect 9376 999 9410 1033
rect 9232 903 9266 937
rect 9304 903 9338 937
rect 9376 903 9410 937
rect 9232 807 9266 841
rect 9304 807 9338 841
rect 9376 807 9410 841
rect 9232 711 9266 745
rect 9304 711 9338 745
rect 9376 711 9410 745
rect 9232 615 9266 649
rect 9304 615 9338 649
rect 9376 615 9410 649
rect 9644 3303 9678 3337
rect 9716 3303 9750 3337
rect 9788 3303 9822 3337
rect 9644 3207 9678 3241
rect 9716 3207 9750 3241
rect 9788 3207 9822 3241
rect 9644 3111 9678 3145
rect 9716 3111 9750 3145
rect 9788 3111 9822 3145
rect 9644 3015 9678 3049
rect 9716 3015 9750 3049
rect 9788 3015 9822 3049
rect 9644 2919 9678 2953
rect 9716 2919 9750 2953
rect 9788 2919 9822 2953
rect 9644 2823 9678 2857
rect 9716 2823 9750 2857
rect 9788 2823 9822 2857
rect 9644 2727 9678 2761
rect 9716 2727 9750 2761
rect 9788 2727 9822 2761
rect 9644 2631 9678 2665
rect 9716 2631 9750 2665
rect 9788 2631 9822 2665
rect 9644 2535 9678 2569
rect 9716 2535 9750 2569
rect 9788 2535 9822 2569
rect 9644 2439 9678 2473
rect 9716 2439 9750 2473
rect 9788 2439 9822 2473
rect 9644 2343 9678 2377
rect 9716 2343 9750 2377
rect 9788 2343 9822 2377
rect 9644 2247 9678 2281
rect 9716 2247 9750 2281
rect 9788 2247 9822 2281
rect 9644 2151 9678 2185
rect 9716 2151 9750 2185
rect 9788 2151 9822 2185
rect 9644 2055 9678 2089
rect 9716 2055 9750 2089
rect 9788 2055 9822 2089
rect 9644 1959 9678 1993
rect 9716 1959 9750 1993
rect 9788 1959 9822 1993
rect 9644 1863 9678 1897
rect 9716 1863 9750 1897
rect 9788 1863 9822 1897
rect 9644 1767 9678 1801
rect 9716 1767 9750 1801
rect 9788 1767 9822 1801
rect 9644 1671 9678 1705
rect 9716 1671 9750 1705
rect 9788 1671 9822 1705
rect 9644 1575 9678 1609
rect 9716 1575 9750 1609
rect 9788 1575 9822 1609
rect 9644 1479 9678 1513
rect 9716 1479 9750 1513
rect 9788 1479 9822 1513
rect 9644 1383 9678 1417
rect 9716 1383 9750 1417
rect 9788 1383 9822 1417
rect 9644 1287 9678 1321
rect 9716 1287 9750 1321
rect 9788 1287 9822 1321
rect 9644 1191 9678 1225
rect 9716 1191 9750 1225
rect 9788 1191 9822 1225
rect 9644 1095 9678 1129
rect 9716 1095 9750 1129
rect 9788 1095 9822 1129
rect 9644 999 9678 1033
rect 9716 999 9750 1033
rect 9788 999 9822 1033
rect 9644 903 9678 937
rect 9716 903 9750 937
rect 9788 903 9822 937
rect 9644 807 9678 841
rect 9716 807 9750 841
rect 9788 807 9822 841
rect 9644 711 9678 745
rect 9716 711 9750 745
rect 9788 711 9822 745
rect 9644 615 9678 649
rect 9716 615 9750 649
rect 9788 615 9822 649
rect 10056 3303 10090 3337
rect 10128 3303 10162 3337
rect 10200 3303 10234 3337
rect 10056 3207 10090 3241
rect 10128 3207 10162 3241
rect 10200 3207 10234 3241
rect 10056 3111 10090 3145
rect 10128 3111 10162 3145
rect 10200 3111 10234 3145
rect 10056 3015 10090 3049
rect 10128 3015 10162 3049
rect 10200 3015 10234 3049
rect 10056 2919 10090 2953
rect 10128 2919 10162 2953
rect 10200 2919 10234 2953
rect 10056 2823 10090 2857
rect 10128 2823 10162 2857
rect 10200 2823 10234 2857
rect 10056 2727 10090 2761
rect 10128 2727 10162 2761
rect 10200 2727 10234 2761
rect 10056 2631 10090 2665
rect 10128 2631 10162 2665
rect 10200 2631 10234 2665
rect 10056 2535 10090 2569
rect 10128 2535 10162 2569
rect 10200 2535 10234 2569
rect 10056 2439 10090 2473
rect 10128 2439 10162 2473
rect 10200 2439 10234 2473
rect 10056 2343 10090 2377
rect 10128 2343 10162 2377
rect 10200 2343 10234 2377
rect 10056 2247 10090 2281
rect 10128 2247 10162 2281
rect 10200 2247 10234 2281
rect 10056 2151 10090 2185
rect 10128 2151 10162 2185
rect 10200 2151 10234 2185
rect 10056 2055 10090 2089
rect 10128 2055 10162 2089
rect 10200 2055 10234 2089
rect 10056 1959 10090 1993
rect 10128 1959 10162 1993
rect 10200 1959 10234 1993
rect 10056 1863 10090 1897
rect 10128 1863 10162 1897
rect 10200 1863 10234 1897
rect 10056 1767 10090 1801
rect 10128 1767 10162 1801
rect 10200 1767 10234 1801
rect 10056 1671 10090 1705
rect 10128 1671 10162 1705
rect 10200 1671 10234 1705
rect 10056 1575 10090 1609
rect 10128 1575 10162 1609
rect 10200 1575 10234 1609
rect 10056 1479 10090 1513
rect 10128 1479 10162 1513
rect 10200 1479 10234 1513
rect 10056 1383 10090 1417
rect 10128 1383 10162 1417
rect 10200 1383 10234 1417
rect 10056 1287 10090 1321
rect 10128 1287 10162 1321
rect 10200 1287 10234 1321
rect 10056 1191 10090 1225
rect 10128 1191 10162 1225
rect 10200 1191 10234 1225
rect 10056 1095 10090 1129
rect 10128 1095 10162 1129
rect 10200 1095 10234 1129
rect 10056 999 10090 1033
rect 10128 999 10162 1033
rect 10200 999 10234 1033
rect 10056 903 10090 937
rect 10128 903 10162 937
rect 10200 903 10234 937
rect 10056 807 10090 841
rect 10128 807 10162 841
rect 10200 807 10234 841
rect 10056 711 10090 745
rect 10128 711 10162 745
rect 10200 711 10234 745
rect 10056 615 10090 649
rect 10128 615 10162 649
rect 10200 615 10234 649
rect 10468 3303 10502 3337
rect 10540 3303 10574 3337
rect 10612 3303 10646 3337
rect 10468 3207 10502 3241
rect 10540 3207 10574 3241
rect 10612 3207 10646 3241
rect 10468 3111 10502 3145
rect 10540 3111 10574 3145
rect 10612 3111 10646 3145
rect 10468 3015 10502 3049
rect 10540 3015 10574 3049
rect 10612 3015 10646 3049
rect 10468 2919 10502 2953
rect 10540 2919 10574 2953
rect 10612 2919 10646 2953
rect 10468 2823 10502 2857
rect 10540 2823 10574 2857
rect 10612 2823 10646 2857
rect 10468 2727 10502 2761
rect 10540 2727 10574 2761
rect 10612 2727 10646 2761
rect 10468 2631 10502 2665
rect 10540 2631 10574 2665
rect 10612 2631 10646 2665
rect 10468 2535 10502 2569
rect 10540 2535 10574 2569
rect 10612 2535 10646 2569
rect 10468 2439 10502 2473
rect 10540 2439 10574 2473
rect 10612 2439 10646 2473
rect 10468 2343 10502 2377
rect 10540 2343 10574 2377
rect 10612 2343 10646 2377
rect 10468 2247 10502 2281
rect 10540 2247 10574 2281
rect 10612 2247 10646 2281
rect 10468 2151 10502 2185
rect 10540 2151 10574 2185
rect 10612 2151 10646 2185
rect 10468 2055 10502 2089
rect 10540 2055 10574 2089
rect 10612 2055 10646 2089
rect 10468 1959 10502 1993
rect 10540 1959 10574 1993
rect 10612 1959 10646 1993
rect 10468 1863 10502 1897
rect 10540 1863 10574 1897
rect 10612 1863 10646 1897
rect 10468 1767 10502 1801
rect 10540 1767 10574 1801
rect 10612 1767 10646 1801
rect 10468 1671 10502 1705
rect 10540 1671 10574 1705
rect 10612 1671 10646 1705
rect 10468 1575 10502 1609
rect 10540 1575 10574 1609
rect 10612 1575 10646 1609
rect 10468 1479 10502 1513
rect 10540 1479 10574 1513
rect 10612 1479 10646 1513
rect 10468 1383 10502 1417
rect 10540 1383 10574 1417
rect 10612 1383 10646 1417
rect 10468 1287 10502 1321
rect 10540 1287 10574 1321
rect 10612 1287 10646 1321
rect 10468 1191 10502 1225
rect 10540 1191 10574 1225
rect 10612 1191 10646 1225
rect 10468 1095 10502 1129
rect 10540 1095 10574 1129
rect 10612 1095 10646 1129
rect 10468 999 10502 1033
rect 10540 999 10574 1033
rect 10612 999 10646 1033
rect 10468 903 10502 937
rect 10540 903 10574 937
rect 10612 903 10646 937
rect 10468 807 10502 841
rect 10540 807 10574 841
rect 10612 807 10646 841
rect 10468 711 10502 745
rect 10540 711 10574 745
rect 10612 711 10646 745
rect 10468 615 10502 649
rect 10540 615 10574 649
rect 10612 615 10646 649
rect 10880 3303 10914 3337
rect 10952 3303 10986 3337
rect 11024 3303 11058 3337
rect 10880 3207 10914 3241
rect 10952 3207 10986 3241
rect 11024 3207 11058 3241
rect 10880 3111 10914 3145
rect 10952 3111 10986 3145
rect 11024 3111 11058 3145
rect 10880 3015 10914 3049
rect 10952 3015 10986 3049
rect 11024 3015 11058 3049
rect 10880 2919 10914 2953
rect 10952 2919 10986 2953
rect 11024 2919 11058 2953
rect 10880 2823 10914 2857
rect 10952 2823 10986 2857
rect 11024 2823 11058 2857
rect 10880 2727 10914 2761
rect 10952 2727 10986 2761
rect 11024 2727 11058 2761
rect 10880 2631 10914 2665
rect 10952 2631 10986 2665
rect 11024 2631 11058 2665
rect 10880 2535 10914 2569
rect 10952 2535 10986 2569
rect 11024 2535 11058 2569
rect 10880 2439 10914 2473
rect 10952 2439 10986 2473
rect 11024 2439 11058 2473
rect 10880 2343 10914 2377
rect 10952 2343 10986 2377
rect 11024 2343 11058 2377
rect 10880 2247 10914 2281
rect 10952 2247 10986 2281
rect 11024 2247 11058 2281
rect 10880 2151 10914 2185
rect 10952 2151 10986 2185
rect 11024 2151 11058 2185
rect 10880 2055 10914 2089
rect 10952 2055 10986 2089
rect 11024 2055 11058 2089
rect 10880 1959 10914 1993
rect 10952 1959 10986 1993
rect 11024 1959 11058 1993
rect 10880 1863 10914 1897
rect 10952 1863 10986 1897
rect 11024 1863 11058 1897
rect 10880 1767 10914 1801
rect 10952 1767 10986 1801
rect 11024 1767 11058 1801
rect 10880 1671 10914 1705
rect 10952 1671 10986 1705
rect 11024 1671 11058 1705
rect 10880 1575 10914 1609
rect 10952 1575 10986 1609
rect 11024 1575 11058 1609
rect 10880 1479 10914 1513
rect 10952 1479 10986 1513
rect 11024 1479 11058 1513
rect 10880 1383 10914 1417
rect 10952 1383 10986 1417
rect 11024 1383 11058 1417
rect 10880 1287 10914 1321
rect 10952 1287 10986 1321
rect 11024 1287 11058 1321
rect 10880 1191 10914 1225
rect 10952 1191 10986 1225
rect 11024 1191 11058 1225
rect 10880 1095 10914 1129
rect 10952 1095 10986 1129
rect 11024 1095 11058 1129
rect 10880 999 10914 1033
rect 10952 999 10986 1033
rect 11024 999 11058 1033
rect 10880 903 10914 937
rect 10952 903 10986 937
rect 11024 903 11058 937
rect 10880 807 10914 841
rect 10952 807 10986 841
rect 11024 807 11058 841
rect 10880 711 10914 745
rect 10952 711 10986 745
rect 11024 711 11058 745
rect 10880 615 10914 649
rect 10952 615 10986 649
rect 11024 615 11058 649
rect 11252 3455 11255 3464
rect 11255 3455 11286 3464
rect 11252 3430 11286 3455
rect 11252 3387 11255 3392
rect 11255 3387 11286 3392
rect 11252 3358 11286 3387
rect 11252 3319 11255 3320
rect 11255 3319 11286 3320
rect 11252 3286 11286 3319
rect 11252 3217 11286 3248
rect 11252 3214 11255 3217
rect 11255 3214 11286 3217
rect 11252 3149 11286 3176
rect 11252 3142 11255 3149
rect 11255 3142 11286 3149
rect 11252 3081 11286 3104
rect 11252 3070 11255 3081
rect 11255 3070 11286 3081
rect 11252 3013 11286 3032
rect 11252 2998 11255 3013
rect 11255 2998 11286 3013
rect 11252 2945 11286 2960
rect 11252 2926 11255 2945
rect 11255 2926 11286 2945
rect 11252 2877 11286 2888
rect 11252 2854 11255 2877
rect 11255 2854 11286 2877
rect 11252 2809 11286 2816
rect 11252 2782 11255 2809
rect 11255 2782 11286 2809
rect 11252 2741 11286 2744
rect 11252 2710 11255 2741
rect 11255 2710 11286 2741
rect 11252 2639 11255 2672
rect 11255 2639 11286 2672
rect 11252 2638 11286 2639
rect 11252 2571 11255 2600
rect 11255 2571 11286 2600
rect 11252 2566 11286 2571
rect 11252 2503 11255 2528
rect 11255 2503 11286 2528
rect 11252 2494 11286 2503
rect 11252 2435 11255 2456
rect 11255 2435 11286 2456
rect 11252 2422 11286 2435
rect 11252 2367 11255 2384
rect 11255 2367 11286 2384
rect 11252 2350 11286 2367
rect 11252 2299 11255 2312
rect 11255 2299 11286 2312
rect 11252 2278 11286 2299
rect 11252 2231 11255 2240
rect 11255 2231 11286 2240
rect 11252 2206 11286 2231
rect 11252 2163 11255 2168
rect 11255 2163 11286 2168
rect 11252 2134 11286 2163
rect 11252 2095 11255 2096
rect 11255 2095 11286 2096
rect 11252 2062 11286 2095
rect 11252 1993 11286 2024
rect 11252 1990 11255 1993
rect 11255 1990 11286 1993
rect 11252 1925 11286 1952
rect 11252 1918 11255 1925
rect 11255 1918 11286 1925
rect 11252 1857 11286 1880
rect 11252 1846 11255 1857
rect 11255 1846 11286 1857
rect 11252 1789 11286 1808
rect 11252 1774 11255 1789
rect 11255 1774 11286 1789
rect 11252 1721 11286 1736
rect 11252 1702 11255 1721
rect 11255 1702 11286 1721
rect 11252 1653 11286 1664
rect 11252 1630 11255 1653
rect 11255 1630 11286 1653
rect 11252 1585 11286 1592
rect 11252 1558 11255 1585
rect 11255 1558 11286 1585
rect 11252 1517 11286 1520
rect 11252 1486 11255 1517
rect 11255 1486 11286 1517
rect 11252 1415 11255 1448
rect 11255 1415 11286 1448
rect 11252 1414 11286 1415
rect 11252 1347 11255 1376
rect 11255 1347 11286 1376
rect 11252 1342 11286 1347
rect 11252 1279 11255 1304
rect 11255 1279 11286 1304
rect 11252 1270 11286 1279
rect 11252 1211 11255 1232
rect 11255 1211 11286 1232
rect 11252 1198 11286 1211
rect 11252 1143 11255 1160
rect 11255 1143 11286 1160
rect 11252 1126 11286 1143
rect 11252 1075 11255 1088
rect 11255 1075 11286 1088
rect 11252 1054 11286 1075
rect 11252 1007 11255 1016
rect 11255 1007 11286 1016
rect 11252 982 11286 1007
rect 11252 939 11255 944
rect 11255 939 11286 944
rect 11252 910 11286 939
rect 11252 871 11255 872
rect 11255 871 11286 872
rect 11252 838 11286 871
rect 11252 769 11286 800
rect 11252 766 11255 769
rect 11255 766 11286 769
rect 11252 701 11286 728
rect 11252 694 11255 701
rect 11255 694 11286 701
rect 11252 633 11286 656
rect 11252 622 11255 633
rect 11255 622 11286 633
<< metal1 >>
rect 7233 3666 11313 3670
rect 7233 3614 7290 3666
rect 7342 3614 7355 3666
rect 7407 3614 7419 3666
rect 7471 3614 7483 3666
rect 7535 3614 7547 3666
rect 7599 3664 7611 3666
rect 7663 3664 7675 3666
rect 7727 3664 7739 3666
rect 7791 3664 7803 3666
rect 7855 3664 7867 3666
rect 7608 3630 7611 3664
rect 7855 3630 7862 3664
rect 7599 3614 7611 3630
rect 7663 3614 7675 3630
rect 7727 3614 7739 3630
rect 7791 3614 7803 3630
rect 7855 3614 7867 3630
rect 7919 3614 7931 3666
rect 7983 3614 7995 3666
rect 8047 3614 8059 3666
rect 8111 3664 8123 3666
rect 8175 3664 8187 3666
rect 8239 3664 8251 3666
rect 8303 3664 8315 3666
rect 8367 3664 8379 3666
rect 8431 3664 8443 3666
rect 8112 3630 8123 3664
rect 8184 3630 8187 3664
rect 8431 3630 8438 3664
rect 8111 3614 8123 3630
rect 8175 3614 8187 3630
rect 8239 3614 8251 3630
rect 8303 3614 8315 3630
rect 8367 3614 8379 3630
rect 8431 3614 8443 3630
rect 8495 3614 8507 3666
rect 8559 3614 8571 3666
rect 8623 3614 8635 3666
rect 8687 3664 8699 3666
rect 8751 3664 8763 3666
rect 8815 3664 8827 3666
rect 8879 3664 8891 3666
rect 8943 3664 8955 3666
rect 9007 3664 9019 3666
rect 8688 3630 8699 3664
rect 8760 3630 8763 3664
rect 9007 3630 9014 3664
rect 8687 3614 8699 3630
rect 8751 3614 8763 3630
rect 8815 3614 8827 3630
rect 8879 3614 8891 3630
rect 8943 3614 8955 3630
rect 9007 3614 9019 3630
rect 9071 3614 9083 3666
rect 9135 3614 9147 3666
rect 9199 3614 9211 3666
rect 9263 3664 9275 3666
rect 9327 3664 9339 3666
rect 9391 3664 9403 3666
rect 9455 3664 9467 3666
rect 9519 3664 9531 3666
rect 9583 3664 9595 3666
rect 9264 3630 9275 3664
rect 9336 3630 9339 3664
rect 9583 3630 9590 3664
rect 9263 3614 9275 3630
rect 9327 3614 9339 3630
rect 9391 3614 9403 3630
rect 9455 3614 9467 3630
rect 9519 3614 9531 3630
rect 9583 3614 9595 3630
rect 9647 3614 9659 3666
rect 9711 3614 9723 3666
rect 9775 3614 9787 3666
rect 9839 3664 9851 3666
rect 9903 3664 9915 3666
rect 9967 3664 9979 3666
rect 10031 3664 10043 3666
rect 10095 3664 10107 3666
rect 10159 3664 10171 3666
rect 9840 3630 9851 3664
rect 9912 3630 9915 3664
rect 10159 3630 10166 3664
rect 9839 3614 9851 3630
rect 9903 3614 9915 3630
rect 9967 3614 9979 3630
rect 10031 3614 10043 3630
rect 10095 3614 10107 3630
rect 10159 3614 10171 3630
rect 10223 3614 10235 3666
rect 10287 3614 10299 3666
rect 10351 3614 10363 3666
rect 10415 3664 10427 3666
rect 10479 3664 10491 3666
rect 10543 3664 10555 3666
rect 10607 3664 10619 3666
rect 10671 3664 10683 3666
rect 10735 3664 10747 3666
rect 10416 3630 10427 3664
rect 10488 3630 10491 3664
rect 10735 3630 10742 3664
rect 10415 3614 10427 3630
rect 10479 3614 10491 3630
rect 10543 3614 10555 3630
rect 10607 3614 10619 3630
rect 10671 3614 10683 3630
rect 10735 3614 10747 3630
rect 10799 3614 10811 3666
rect 10863 3664 11313 3666
rect 10863 3630 10886 3664
rect 10920 3630 10958 3664
rect 10992 3630 11030 3664
rect 11064 3630 11102 3664
rect 11136 3630 11174 3664
rect 11208 3630 11313 3664
rect 10863 3614 11313 3630
rect 7233 3578 11313 3614
rect 7233 3526 7290 3578
rect 7342 3536 7355 3578
rect 7342 3526 7350 3536
rect 7407 3526 7419 3578
rect 7471 3526 7483 3578
rect 7535 3526 7547 3578
rect 7599 3526 7611 3578
rect 7663 3526 7675 3578
rect 7727 3526 7739 3578
rect 7791 3526 7803 3578
rect 7855 3526 7867 3578
rect 7919 3526 7931 3578
rect 7983 3526 7995 3578
rect 8047 3526 8059 3578
rect 8111 3526 8123 3578
rect 8175 3526 8187 3578
rect 8239 3526 8251 3578
rect 8303 3526 8315 3578
rect 8367 3526 8379 3578
rect 8431 3526 8443 3578
rect 8495 3526 8507 3578
rect 8559 3526 8571 3578
rect 8623 3526 8635 3578
rect 8687 3526 8699 3578
rect 8751 3526 8763 3578
rect 8815 3526 8827 3578
rect 8879 3526 8891 3578
rect 8943 3526 8955 3578
rect 9007 3526 9019 3578
rect 9071 3526 9083 3578
rect 9135 3526 9147 3578
rect 9199 3526 9211 3578
rect 9263 3526 9275 3578
rect 9327 3526 9339 3578
rect 9391 3526 9403 3578
rect 9455 3526 9467 3578
rect 9519 3526 9531 3578
rect 9583 3526 9595 3578
rect 9647 3526 9659 3578
rect 9711 3526 9723 3578
rect 9775 3526 9787 3578
rect 9839 3526 9851 3578
rect 9903 3526 9915 3578
rect 9967 3526 9979 3578
rect 10031 3526 10043 3578
rect 10095 3526 10107 3578
rect 10159 3526 10171 3578
rect 10223 3526 10235 3578
rect 10287 3526 10299 3578
rect 10351 3526 10363 3578
rect 10415 3526 10427 3578
rect 10479 3526 10491 3578
rect 10543 3526 10555 3578
rect 10607 3526 10619 3578
rect 10671 3526 10683 3578
rect 10735 3526 10747 3578
rect 10799 3526 10811 3578
rect 10863 3536 11313 3578
rect 10863 3526 11252 3536
rect 7233 3502 7350 3526
rect 7384 3516 11252 3526
rect 7384 3502 7445 3516
tri 7445 3502 7459 3516 nw
tri 11197 3502 11211 3516 ne
rect 11211 3502 11252 3516
rect 11286 3502 11313 3536
rect 7233 3464 7411 3502
tri 7411 3468 7445 3502 nw
tri 11211 3482 11231 3502 ne
tri 7575 3468 7583 3476 se
rect 7583 3468 7763 3476
tri 7571 3464 7575 3468 se
rect 7575 3464 7763 3468
tri 7763 3464 7775 3476 sw
tri 7983 3464 7995 3476 se
rect 7995 3464 8175 3476
tri 8175 3464 8187 3476 sw
tri 8395 3464 8407 3476 se
rect 8407 3464 8587 3476
tri 8587 3464 8599 3476 sw
tri 8807 3464 8819 3476 se
rect 8819 3464 8999 3476
tri 8999 3464 9011 3476 sw
tri 9219 3464 9231 3476 se
rect 9231 3464 9411 3476
tri 9411 3464 9423 3476 sw
tri 9631 3464 9643 3476 se
rect 9643 3464 9823 3476
tri 9823 3464 9835 3476 sw
tri 10043 3464 10055 3476 se
rect 10055 3464 10235 3476
tri 10235 3464 10247 3476 sw
tri 10455 3464 10467 3476 se
rect 10467 3464 10647 3476
tri 10647 3464 10659 3476 sw
tri 10867 3464 10879 3476 se
rect 10879 3464 11059 3476
tri 11059 3464 11071 3476 sw
rect 11231 3464 11313 3502
rect 7233 3430 7350 3464
rect 7384 3430 7411 3464
tri 7537 3430 7571 3464 se
rect 7571 3430 7775 3464
tri 7775 3430 7809 3464 sw
tri 7949 3430 7983 3464 se
rect 7983 3430 8187 3464
tri 8187 3430 8221 3464 sw
tri 8361 3430 8395 3464 se
rect 8395 3430 8599 3464
tri 8599 3430 8633 3464 sw
tri 8773 3430 8807 3464 se
rect 8807 3430 9011 3464
tri 9011 3430 9045 3464 sw
tri 9185 3430 9219 3464 se
rect 9219 3430 9423 3464
tri 9423 3430 9457 3464 sw
tri 9597 3430 9631 3464 se
rect 9631 3430 9835 3464
tri 9835 3430 9869 3464 sw
tri 10009 3430 10043 3464 se
rect 10043 3430 10247 3464
tri 10247 3430 10281 3464 sw
tri 10421 3430 10455 3464 se
rect 10455 3430 10659 3464
tri 10659 3430 10693 3464 sw
tri 10833 3430 10867 3464 se
rect 10867 3430 11071 3464
tri 11071 3430 11105 3464 sw
rect 11231 3430 11252 3464
rect 11286 3430 11313 3464
rect 7233 3392 7411 3430
rect 7233 3358 7350 3392
rect 7384 3358 7411 3392
rect 7233 3320 7411 3358
rect 7233 3286 7350 3320
rect 7384 3286 7411 3320
rect 7233 3248 7411 3286
rect 7233 3214 7350 3248
rect 7384 3214 7411 3248
rect 7233 3176 7411 3214
rect 7233 3142 7350 3176
rect 7384 3142 7411 3176
rect 7233 3104 7411 3142
rect 7233 3070 7350 3104
rect 7384 3070 7411 3104
rect 7233 3032 7411 3070
rect 7233 2998 7350 3032
rect 7384 2998 7411 3032
rect 7233 2960 7411 2998
rect 7233 2926 7350 2960
rect 7384 2926 7411 2960
rect 7233 2888 7411 2926
rect 7233 2854 7350 2888
rect 7384 2854 7411 2888
rect 7233 2816 7411 2854
rect 7233 2782 7350 2816
rect 7384 2782 7411 2816
rect 7233 2744 7411 2782
rect 7233 2710 7350 2744
rect 7384 2710 7411 2744
rect 7233 2672 7411 2710
rect 7233 2638 7350 2672
rect 7384 2638 7411 2672
rect 7233 2600 7411 2638
rect 7233 2566 7350 2600
rect 7384 2566 7411 2600
rect 7233 2528 7411 2566
rect 7233 2494 7350 2528
rect 7384 2494 7411 2528
rect 7233 2456 7411 2494
rect 7233 2422 7350 2456
rect 7384 2422 7411 2456
rect 7233 2384 7411 2422
rect 7233 2350 7350 2384
rect 7384 2350 7411 2384
rect 7233 2312 7411 2350
rect 7233 2278 7350 2312
rect 7384 2278 7411 2312
rect 7233 2240 7411 2278
rect 7233 2206 7350 2240
rect 7384 2206 7411 2240
rect 7233 2168 7411 2206
rect 7233 2134 7350 2168
rect 7384 2134 7411 2168
rect 7233 2096 7411 2134
rect 7233 2062 7350 2096
rect 7384 2062 7411 2096
rect 7233 2024 7411 2062
rect 7233 1990 7350 2024
rect 7384 1990 7411 2024
rect 7233 1952 7411 1990
rect 7233 1918 7350 1952
rect 7384 1918 7411 1952
rect 7233 1880 7411 1918
rect 7233 1846 7350 1880
rect 7384 1846 7411 1880
rect 7233 1808 7411 1846
rect 7233 1774 7350 1808
rect 7384 1774 7411 1808
rect 7233 1736 7411 1774
rect 7233 1702 7350 1736
rect 7384 1702 7411 1736
rect 7233 1664 7411 1702
rect 7233 1630 7350 1664
rect 7384 1630 7411 1664
rect 7233 1592 7411 1630
rect 7233 1558 7350 1592
rect 7384 1558 7411 1592
rect 7233 1520 7411 1558
rect 7233 1486 7350 1520
rect 7384 1486 7411 1520
rect 7233 1448 7411 1486
rect 7233 1414 7350 1448
rect 7384 1414 7411 1448
rect 7233 1376 7411 1414
rect 7233 1342 7350 1376
rect 7384 1342 7411 1376
rect 7233 1304 7411 1342
rect 7233 1270 7350 1304
rect 7384 1270 7411 1304
rect 7233 1232 7411 1270
rect 7233 1198 7350 1232
rect 7384 1198 7411 1232
rect 7233 1160 7411 1198
rect 7233 1126 7350 1160
rect 7384 1126 7411 1160
rect 7233 1088 7411 1126
rect 7233 1054 7350 1088
rect 7384 1054 7411 1088
rect 7233 1016 7411 1054
rect 7233 982 7350 1016
rect 7384 982 7411 1016
rect 7233 944 7411 982
rect 7233 910 7350 944
rect 7384 910 7411 944
rect 7233 872 7411 910
rect 7233 838 7350 872
rect 7384 838 7411 872
rect 7233 800 7411 838
rect 7233 766 7350 800
rect 7384 766 7411 800
rect 7233 728 7411 766
rect 7233 694 7350 728
rect 7384 694 7411 728
rect 7233 656 7411 694
rect 7233 622 7350 656
rect 7384 622 7411 656
rect 7233 609 7411 622
tri 7523 3416 7537 3430 se
rect 7537 3416 7809 3430
tri 7809 3416 7823 3430 sw
rect 7523 3410 7823 3416
rect 7523 3358 7524 3410
rect 7576 3358 7606 3410
rect 7658 3358 7688 3410
rect 7740 3358 7770 3410
rect 7822 3358 7823 3410
rect 7523 3344 7823 3358
rect 7523 3292 7524 3344
rect 7576 3337 7606 3344
rect 7658 3337 7688 3344
rect 7740 3337 7770 3344
rect 7576 3303 7584 3337
rect 7762 3303 7770 3337
rect 7576 3292 7606 3303
rect 7658 3292 7688 3303
rect 7740 3292 7770 3303
rect 7822 3292 7823 3344
rect 7523 3278 7823 3292
rect 7523 3226 7524 3278
rect 7576 3241 7606 3278
rect 7658 3241 7688 3278
rect 7740 3241 7770 3278
rect 7576 3226 7584 3241
rect 7762 3226 7770 3241
rect 7822 3226 7823 3278
rect 7523 3212 7584 3226
rect 7618 3212 7656 3226
rect 7690 3212 7728 3226
rect 7762 3212 7823 3226
rect 7523 3160 7524 3212
rect 7576 3207 7584 3212
rect 7762 3207 7770 3212
rect 7576 3160 7606 3207
rect 7658 3160 7688 3207
rect 7740 3160 7770 3207
rect 7822 3160 7823 3212
rect 7523 3146 7823 3160
rect 7523 3094 7524 3146
rect 7576 3145 7606 3146
rect 7658 3145 7688 3146
rect 7740 3145 7770 3146
rect 7576 3111 7584 3145
rect 7762 3111 7770 3145
rect 7576 3094 7606 3111
rect 7658 3094 7688 3111
rect 7740 3094 7770 3111
rect 7822 3094 7823 3146
rect 7523 3079 7823 3094
rect 7523 3027 7524 3079
rect 7576 3049 7606 3079
rect 7658 3049 7688 3079
rect 7740 3049 7770 3079
rect 7576 3027 7584 3049
rect 7762 3027 7770 3049
rect 7822 3027 7823 3079
rect 7523 3015 7584 3027
rect 7618 3015 7656 3027
rect 7690 3015 7728 3027
rect 7762 3015 7823 3027
rect 7523 3012 7823 3015
rect 7523 2960 7524 3012
rect 7576 2960 7606 3012
rect 7658 2960 7688 3012
rect 7740 2960 7770 3012
rect 7822 2960 7823 3012
rect 7523 2953 7823 2960
rect 7523 2945 7584 2953
rect 7618 2945 7656 2953
rect 7690 2945 7728 2953
rect 7762 2945 7823 2953
rect 7523 2893 7524 2945
rect 7576 2919 7584 2945
rect 7762 2919 7770 2945
rect 7576 2893 7606 2919
rect 7658 2893 7688 2919
rect 7740 2893 7770 2919
rect 7822 2893 7823 2945
rect 7523 2878 7823 2893
rect 7523 2826 7524 2878
rect 7576 2857 7606 2878
rect 7658 2857 7688 2878
rect 7740 2857 7770 2878
rect 7576 2826 7584 2857
rect 7762 2826 7770 2857
rect 7822 2826 7823 2878
rect 7523 2823 7584 2826
rect 7618 2823 7656 2826
rect 7690 2823 7728 2826
rect 7762 2823 7823 2826
rect 7523 2811 7823 2823
rect 7523 2759 7524 2811
rect 7576 2761 7606 2811
rect 7658 2761 7688 2811
rect 7740 2761 7770 2811
rect 7576 2759 7584 2761
rect 7762 2759 7770 2761
rect 7822 2759 7823 2811
rect 7523 2744 7584 2759
rect 7618 2744 7656 2759
rect 7690 2744 7728 2759
rect 7762 2744 7823 2759
rect 7523 2692 7524 2744
rect 7576 2727 7584 2744
rect 7762 2727 7770 2744
rect 7576 2692 7606 2727
rect 7658 2692 7688 2727
rect 7740 2692 7770 2727
rect 7822 2692 7823 2744
rect 7523 2677 7823 2692
rect 7523 2625 7524 2677
rect 7576 2665 7606 2677
rect 7658 2665 7688 2677
rect 7740 2665 7770 2677
rect 7576 2631 7584 2665
rect 7762 2631 7770 2665
rect 7576 2625 7606 2631
rect 7658 2625 7688 2631
rect 7740 2625 7770 2631
rect 7822 2625 7823 2677
rect 7523 2610 7823 2625
rect 7523 2558 7524 2610
rect 7576 2569 7606 2610
rect 7658 2569 7688 2610
rect 7740 2569 7770 2610
rect 7576 2558 7584 2569
rect 7762 2558 7770 2569
rect 7822 2558 7823 2610
rect 7523 2543 7584 2558
rect 7618 2543 7656 2558
rect 7690 2543 7728 2558
rect 7762 2543 7823 2558
rect 7523 2491 7524 2543
rect 7576 2535 7584 2543
rect 7762 2535 7770 2543
rect 7576 2491 7606 2535
rect 7658 2491 7688 2535
rect 7740 2491 7770 2535
rect 7822 2491 7823 2543
rect 7523 2476 7823 2491
rect 7523 2424 7524 2476
rect 7576 2473 7606 2476
rect 7658 2473 7688 2476
rect 7740 2473 7770 2476
rect 7576 2439 7584 2473
rect 7762 2439 7770 2473
rect 7576 2424 7606 2439
rect 7658 2424 7688 2439
rect 7740 2424 7770 2439
rect 7822 2424 7823 2476
rect 7523 2409 7823 2424
rect 7523 2357 7524 2409
rect 7576 2377 7606 2409
rect 7658 2377 7688 2409
rect 7740 2377 7770 2409
rect 7576 2357 7584 2377
rect 7762 2357 7770 2377
rect 7822 2357 7823 2409
rect 7523 2343 7584 2357
rect 7618 2343 7656 2357
rect 7690 2343 7728 2357
rect 7762 2343 7823 2357
rect 7523 2342 7823 2343
rect 7523 2290 7524 2342
rect 7576 2290 7606 2342
rect 7658 2290 7688 2342
rect 7740 2290 7770 2342
rect 7822 2290 7823 2342
rect 7523 2281 7823 2290
rect 7523 2275 7584 2281
rect 7618 2275 7656 2281
rect 7690 2275 7728 2281
rect 7762 2275 7823 2281
rect 7523 2223 7524 2275
rect 7576 2247 7584 2275
rect 7762 2247 7770 2275
rect 7576 2223 7606 2247
rect 7658 2223 7688 2247
rect 7740 2223 7770 2247
rect 7822 2223 7823 2275
rect 7523 2208 7823 2223
rect 7523 2156 7524 2208
rect 7576 2185 7606 2208
rect 7658 2185 7688 2208
rect 7740 2185 7770 2208
rect 7576 2156 7584 2185
rect 7762 2156 7770 2185
rect 7822 2156 7823 2208
rect 7523 2151 7584 2156
rect 7618 2151 7656 2156
rect 7690 2151 7728 2156
rect 7762 2151 7823 2156
rect 7523 2141 7823 2151
rect 7523 2089 7524 2141
rect 7576 2089 7606 2141
rect 7658 2089 7688 2141
rect 7740 2089 7770 2141
rect 7822 2089 7823 2141
rect 7523 2074 7584 2089
rect 7618 2074 7656 2089
rect 7690 2074 7728 2089
rect 7762 2074 7823 2089
rect 7523 2022 7524 2074
rect 7576 2055 7584 2074
rect 7762 2055 7770 2074
rect 7576 2022 7606 2055
rect 7658 2022 7688 2055
rect 7740 2022 7770 2055
rect 7822 2022 7823 2074
rect 7523 1993 7823 2022
rect 7523 1959 7584 1993
rect 7618 1959 7656 1993
rect 7690 1959 7728 1993
rect 7762 1959 7823 1993
rect 7523 1897 7823 1959
rect 7523 1863 7584 1897
rect 7618 1863 7656 1897
rect 7690 1863 7728 1897
rect 7762 1863 7823 1897
rect 7523 1801 7823 1863
rect 7523 1767 7584 1801
rect 7618 1767 7656 1801
rect 7690 1767 7728 1801
rect 7762 1767 7823 1801
rect 7523 1705 7823 1767
rect 7523 1671 7584 1705
rect 7618 1671 7656 1705
rect 7690 1671 7728 1705
rect 7762 1671 7823 1705
rect 7523 1609 7823 1671
rect 7523 1575 7584 1609
rect 7618 1575 7656 1609
rect 7690 1575 7728 1609
rect 7762 1575 7823 1609
rect 7523 1513 7823 1575
rect 7523 1479 7584 1513
rect 7618 1479 7656 1513
rect 7690 1479 7728 1513
rect 7762 1479 7823 1513
rect 7523 1417 7823 1479
rect 7523 1383 7584 1417
rect 7618 1383 7656 1417
rect 7690 1383 7728 1417
rect 7762 1383 7823 1417
rect 7523 1321 7823 1383
rect 7523 1287 7584 1321
rect 7618 1287 7656 1321
rect 7690 1287 7728 1321
rect 7762 1287 7823 1321
rect 7523 1225 7823 1287
rect 7523 1191 7584 1225
rect 7618 1191 7656 1225
rect 7690 1191 7728 1225
rect 7762 1191 7823 1225
rect 7523 1129 7823 1191
rect 7523 1095 7584 1129
rect 7618 1095 7656 1129
rect 7690 1095 7728 1129
rect 7762 1095 7823 1129
rect 7523 1033 7823 1095
rect 7523 999 7584 1033
rect 7618 999 7656 1033
rect 7690 999 7728 1033
rect 7762 999 7823 1033
rect 7523 937 7823 999
rect 7523 903 7584 937
rect 7618 903 7656 937
rect 7690 903 7728 937
rect 7762 903 7823 937
rect 7523 841 7823 903
rect 7523 807 7584 841
rect 7618 807 7656 841
rect 7690 807 7728 841
rect 7762 807 7823 841
rect 7523 745 7823 807
rect 7523 711 7584 745
rect 7618 711 7656 745
rect 7690 711 7728 745
rect 7762 711 7823 745
rect 7523 649 7823 711
rect 7523 615 7584 649
rect 7618 615 7656 649
rect 7690 615 7728 649
rect 7762 615 7823 649
rect 7523 536 7823 615
tri 7523 476 7583 536 ne
rect 7583 476 7763 536
tri 7763 476 7823 536 nw
tri 7935 3416 7949 3430 se
rect 7949 3416 8221 3430
tri 8221 3416 8235 3430 sw
rect 7935 3337 8235 3416
rect 7935 3303 7996 3337
rect 8030 3303 8068 3337
rect 8102 3303 8140 3337
rect 8174 3303 8235 3337
rect 7935 3241 8235 3303
rect 7935 3207 7996 3241
rect 8030 3207 8068 3241
rect 8102 3207 8140 3241
rect 8174 3207 8235 3241
rect 7935 3145 8235 3207
rect 7935 3111 7996 3145
rect 8030 3111 8068 3145
rect 8102 3111 8140 3145
rect 8174 3111 8235 3145
rect 7935 3049 8235 3111
rect 7935 3015 7996 3049
rect 8030 3015 8068 3049
rect 8102 3015 8140 3049
rect 8174 3015 8235 3049
rect 7935 2953 8235 3015
rect 7935 2919 7996 2953
rect 8030 2919 8068 2953
rect 8102 2919 8140 2953
rect 8174 2919 8235 2953
rect 7935 2857 8235 2919
rect 7935 2823 7996 2857
rect 8030 2823 8068 2857
rect 8102 2823 8140 2857
rect 8174 2823 8235 2857
rect 7935 2761 8235 2823
rect 7935 2727 7996 2761
rect 8030 2727 8068 2761
rect 8102 2727 8140 2761
rect 8174 2727 8235 2761
rect 7935 2665 8235 2727
rect 7935 2631 7996 2665
rect 8030 2631 8068 2665
rect 8102 2631 8140 2665
rect 8174 2631 8235 2665
rect 7935 2569 8235 2631
rect 7935 2535 7996 2569
rect 8030 2535 8068 2569
rect 8102 2535 8140 2569
rect 8174 2535 8235 2569
rect 7935 2473 8235 2535
rect 7935 2439 7996 2473
rect 8030 2439 8068 2473
rect 8102 2439 8140 2473
rect 8174 2439 8235 2473
rect 7935 2377 8235 2439
rect 7935 2343 7996 2377
rect 8030 2343 8068 2377
rect 8102 2343 8140 2377
rect 8174 2343 8235 2377
rect 7935 2281 8235 2343
rect 7935 2247 7996 2281
rect 8030 2247 8068 2281
rect 8102 2247 8140 2281
rect 8174 2247 8235 2281
rect 7935 2185 8235 2247
rect 7935 2151 7996 2185
rect 8030 2151 8068 2185
rect 8102 2151 8140 2185
rect 8174 2151 8235 2185
rect 7935 2089 8235 2151
rect 7935 2055 7996 2089
rect 8030 2055 8068 2089
rect 8102 2055 8140 2089
rect 8174 2055 8235 2089
rect 7935 1993 8235 2055
rect 7935 1959 7996 1993
rect 8030 1959 8068 1993
rect 8102 1959 8140 1993
rect 8174 1959 8235 1993
rect 7935 1902 8235 1959
rect 7935 1850 7936 1902
rect 7988 1897 8018 1902
rect 8070 1897 8100 1902
rect 8152 1897 8182 1902
rect 7988 1863 7996 1897
rect 8174 1863 8182 1897
rect 7988 1850 8018 1863
rect 8070 1850 8100 1863
rect 8152 1850 8182 1863
rect 8234 1850 8235 1902
rect 7935 1838 8235 1850
rect 7935 1786 7936 1838
rect 7988 1801 8018 1838
rect 8070 1801 8100 1838
rect 8152 1801 8182 1838
rect 7988 1786 7996 1801
rect 8174 1786 8182 1801
rect 8234 1786 8235 1838
rect 7935 1774 7996 1786
rect 8030 1774 8068 1786
rect 8102 1774 8140 1786
rect 8174 1774 8235 1786
rect 7935 1722 7936 1774
rect 7988 1767 7996 1774
rect 8174 1767 8182 1774
rect 7988 1722 8018 1767
rect 8070 1722 8100 1767
rect 8152 1722 8182 1767
rect 8234 1722 8235 1774
rect 7935 1710 8235 1722
rect 7935 1658 7936 1710
rect 7988 1705 8018 1710
rect 8070 1705 8100 1710
rect 8152 1705 8182 1710
rect 7988 1671 7996 1705
rect 8174 1671 8182 1705
rect 7988 1658 8018 1671
rect 8070 1658 8100 1671
rect 8152 1658 8182 1671
rect 8234 1658 8235 1710
rect 7935 1646 8235 1658
rect 7935 1594 7936 1646
rect 7988 1609 8018 1646
rect 8070 1609 8100 1646
rect 8152 1609 8182 1646
rect 7988 1594 7996 1609
rect 8174 1594 8182 1609
rect 8234 1594 8235 1646
rect 7935 1582 7996 1594
rect 8030 1582 8068 1594
rect 8102 1582 8140 1594
rect 8174 1582 8235 1594
rect 7935 1530 7936 1582
rect 7988 1575 7996 1582
rect 8174 1575 8182 1582
rect 7988 1530 8018 1575
rect 8070 1530 8100 1575
rect 8152 1530 8182 1575
rect 8234 1530 8235 1582
rect 7935 1518 8235 1530
rect 7935 1466 7936 1518
rect 7988 1513 8018 1518
rect 8070 1513 8100 1518
rect 8152 1513 8182 1518
rect 7988 1479 7996 1513
rect 8174 1479 8182 1513
rect 7988 1466 8018 1479
rect 8070 1466 8100 1479
rect 8152 1466 8182 1479
rect 8234 1466 8235 1518
rect 7935 1454 8235 1466
rect 7935 1402 7936 1454
rect 7988 1417 8018 1454
rect 8070 1417 8100 1454
rect 8152 1417 8182 1454
rect 7988 1402 7996 1417
rect 8174 1402 8182 1417
rect 8234 1402 8235 1454
rect 7935 1390 7996 1402
rect 8030 1390 8068 1402
rect 8102 1390 8140 1402
rect 8174 1390 8235 1402
rect 7935 1338 7936 1390
rect 7988 1383 7996 1390
rect 8174 1383 8182 1390
rect 7988 1338 8018 1383
rect 8070 1338 8100 1383
rect 8152 1338 8182 1383
rect 8234 1338 8235 1390
rect 7935 1326 8235 1338
rect 7935 1274 7936 1326
rect 7988 1321 8018 1326
rect 8070 1321 8100 1326
rect 8152 1321 8182 1326
rect 7988 1287 7996 1321
rect 8174 1287 8182 1321
rect 7988 1274 8018 1287
rect 8070 1274 8100 1287
rect 8152 1274 8182 1287
rect 8234 1274 8235 1326
rect 7935 1262 8235 1274
rect 7935 1210 7936 1262
rect 7988 1225 8018 1262
rect 8070 1225 8100 1262
rect 8152 1225 8182 1262
rect 7988 1210 7996 1225
rect 8174 1210 8182 1225
rect 8234 1210 8235 1262
rect 7935 1198 7996 1210
rect 8030 1198 8068 1210
rect 8102 1198 8140 1210
rect 8174 1198 8235 1210
rect 7935 1146 7936 1198
rect 7988 1191 7996 1198
rect 8174 1191 8182 1198
rect 7988 1146 8018 1191
rect 8070 1146 8100 1191
rect 8152 1146 8182 1191
rect 8234 1146 8235 1198
rect 7935 1134 8235 1146
rect 7935 1082 7936 1134
rect 7988 1129 8018 1134
rect 8070 1129 8100 1134
rect 8152 1129 8182 1134
rect 7988 1095 7996 1129
rect 8174 1095 8182 1129
rect 7988 1082 8018 1095
rect 8070 1082 8100 1095
rect 8152 1082 8182 1095
rect 8234 1082 8235 1134
rect 7935 1070 8235 1082
rect 7935 1018 7936 1070
rect 7988 1033 8018 1070
rect 8070 1033 8100 1070
rect 8152 1033 8182 1070
rect 7988 1018 7996 1033
rect 8174 1018 8182 1033
rect 8234 1018 8235 1070
rect 7935 1006 7996 1018
rect 8030 1006 8068 1018
rect 8102 1006 8140 1018
rect 8174 1006 8235 1018
rect 7935 954 7936 1006
rect 7988 999 7996 1006
rect 8174 999 8182 1006
rect 7988 954 8018 999
rect 8070 954 8100 999
rect 8152 954 8182 999
rect 8234 954 8235 1006
rect 7935 942 8235 954
rect 7935 890 7936 942
rect 7988 937 8018 942
rect 8070 937 8100 942
rect 8152 937 8182 942
rect 7988 903 7996 937
rect 8174 903 8182 937
rect 7988 890 8018 903
rect 8070 890 8100 903
rect 8152 890 8182 903
rect 8234 890 8235 942
rect 7935 878 8235 890
rect 7935 826 7936 878
rect 7988 841 8018 878
rect 8070 841 8100 878
rect 8152 841 8182 878
rect 7988 826 7996 841
rect 8174 826 8182 841
rect 8234 826 8235 878
rect 7935 814 7996 826
rect 8030 814 8068 826
rect 8102 814 8140 826
rect 8174 814 8235 826
rect 7935 762 7936 814
rect 7988 807 7996 814
rect 8174 807 8182 814
rect 7988 762 8018 807
rect 8070 762 8100 807
rect 8152 762 8182 807
rect 8234 762 8235 814
rect 7935 750 8235 762
rect 7935 698 7936 750
rect 7988 745 8018 750
rect 8070 745 8100 750
rect 8152 745 8182 750
rect 7988 711 7996 745
rect 8174 711 8182 745
rect 7988 698 8018 711
rect 8070 698 8100 711
rect 8152 698 8182 711
rect 8234 698 8235 750
rect 7935 685 8235 698
rect 7935 633 7936 685
rect 7988 649 8018 685
rect 8070 649 8100 685
rect 8152 649 8182 685
rect 7988 633 7996 649
rect 8174 633 8182 649
rect 8234 633 8235 685
rect 7935 620 7996 633
rect 8030 620 8068 633
rect 8102 620 8140 633
rect 8174 620 8235 633
rect 7935 568 7936 620
rect 7988 615 7996 620
rect 8174 615 8182 620
rect 7988 568 8018 615
rect 8070 568 8100 615
rect 8152 568 8182 615
rect 8234 568 8235 620
rect 7935 555 8235 568
tri 7905 476 7935 506 se
rect 7935 503 7936 555
rect 7988 503 8018 555
rect 8070 503 8100 555
rect 8152 503 8182 555
rect 8234 503 8235 555
tri 8347 3416 8361 3430 se
rect 8361 3416 8633 3430
tri 8633 3416 8647 3430 sw
rect 8347 3410 8647 3416
rect 8347 3358 8348 3410
rect 8400 3358 8430 3410
rect 8482 3358 8512 3410
rect 8564 3358 8594 3410
rect 8646 3358 8647 3410
rect 8347 3344 8647 3358
rect 8347 3292 8348 3344
rect 8400 3337 8430 3344
rect 8482 3337 8512 3344
rect 8564 3337 8594 3344
rect 8400 3303 8408 3337
rect 8586 3303 8594 3337
rect 8400 3292 8430 3303
rect 8482 3292 8512 3303
rect 8564 3292 8594 3303
rect 8646 3292 8647 3344
rect 8347 3278 8647 3292
rect 8347 3226 8348 3278
rect 8400 3241 8430 3278
rect 8482 3241 8512 3278
rect 8564 3241 8594 3278
rect 8400 3226 8408 3241
rect 8586 3226 8594 3241
rect 8646 3226 8647 3278
rect 8347 3212 8408 3226
rect 8442 3212 8480 3226
rect 8514 3212 8552 3226
rect 8586 3212 8647 3226
rect 8347 3160 8348 3212
rect 8400 3207 8408 3212
rect 8586 3207 8594 3212
rect 8400 3160 8430 3207
rect 8482 3160 8512 3207
rect 8564 3160 8594 3207
rect 8646 3160 8647 3212
rect 8347 3146 8647 3160
rect 8347 3094 8348 3146
rect 8400 3145 8430 3146
rect 8482 3145 8512 3146
rect 8564 3145 8594 3146
rect 8400 3111 8408 3145
rect 8586 3111 8594 3145
rect 8400 3094 8430 3111
rect 8482 3094 8512 3111
rect 8564 3094 8594 3111
rect 8646 3094 8647 3146
rect 8347 3079 8647 3094
rect 8347 3027 8348 3079
rect 8400 3049 8430 3079
rect 8482 3049 8512 3079
rect 8564 3049 8594 3079
rect 8400 3027 8408 3049
rect 8586 3027 8594 3049
rect 8646 3027 8647 3079
rect 8347 3015 8408 3027
rect 8442 3015 8480 3027
rect 8514 3015 8552 3027
rect 8586 3015 8647 3027
rect 8347 3012 8647 3015
rect 8347 2960 8348 3012
rect 8400 2960 8430 3012
rect 8482 2960 8512 3012
rect 8564 2960 8594 3012
rect 8646 2960 8647 3012
rect 8347 2953 8647 2960
rect 8347 2945 8408 2953
rect 8442 2945 8480 2953
rect 8514 2945 8552 2953
rect 8586 2945 8647 2953
rect 8347 2893 8348 2945
rect 8400 2919 8408 2945
rect 8586 2919 8594 2945
rect 8400 2893 8430 2919
rect 8482 2893 8512 2919
rect 8564 2893 8594 2919
rect 8646 2893 8647 2945
rect 8347 2878 8647 2893
rect 8347 2826 8348 2878
rect 8400 2857 8430 2878
rect 8482 2857 8512 2878
rect 8564 2857 8594 2878
rect 8400 2826 8408 2857
rect 8586 2826 8594 2857
rect 8646 2826 8647 2878
rect 8347 2823 8408 2826
rect 8442 2823 8480 2826
rect 8514 2823 8552 2826
rect 8586 2823 8647 2826
rect 8347 2811 8647 2823
rect 8347 2759 8348 2811
rect 8400 2761 8430 2811
rect 8482 2761 8512 2811
rect 8564 2761 8594 2811
rect 8400 2759 8408 2761
rect 8586 2759 8594 2761
rect 8646 2759 8647 2811
rect 8347 2744 8408 2759
rect 8442 2744 8480 2759
rect 8514 2744 8552 2759
rect 8586 2744 8647 2759
rect 8347 2692 8348 2744
rect 8400 2727 8408 2744
rect 8586 2727 8594 2744
rect 8400 2692 8430 2727
rect 8482 2692 8512 2727
rect 8564 2692 8594 2727
rect 8646 2692 8647 2744
rect 8347 2677 8647 2692
rect 8347 2625 8348 2677
rect 8400 2665 8430 2677
rect 8482 2665 8512 2677
rect 8564 2665 8594 2677
rect 8400 2631 8408 2665
rect 8586 2631 8594 2665
rect 8400 2625 8430 2631
rect 8482 2625 8512 2631
rect 8564 2625 8594 2631
rect 8646 2625 8647 2677
rect 8347 2610 8647 2625
rect 8347 2558 8348 2610
rect 8400 2569 8430 2610
rect 8482 2569 8512 2610
rect 8564 2569 8594 2610
rect 8400 2558 8408 2569
rect 8586 2558 8594 2569
rect 8646 2558 8647 2610
rect 8347 2543 8408 2558
rect 8442 2543 8480 2558
rect 8514 2543 8552 2558
rect 8586 2543 8647 2558
rect 8347 2491 8348 2543
rect 8400 2535 8408 2543
rect 8586 2535 8594 2543
rect 8400 2491 8430 2535
rect 8482 2491 8512 2535
rect 8564 2491 8594 2535
rect 8646 2491 8647 2543
rect 8347 2476 8647 2491
rect 8347 2424 8348 2476
rect 8400 2473 8430 2476
rect 8482 2473 8512 2476
rect 8564 2473 8594 2476
rect 8400 2439 8408 2473
rect 8586 2439 8594 2473
rect 8400 2424 8430 2439
rect 8482 2424 8512 2439
rect 8564 2424 8594 2439
rect 8646 2424 8647 2476
rect 8347 2409 8647 2424
rect 8347 2357 8348 2409
rect 8400 2377 8430 2409
rect 8482 2377 8512 2409
rect 8564 2377 8594 2409
rect 8400 2357 8408 2377
rect 8586 2357 8594 2377
rect 8646 2357 8647 2409
rect 8347 2343 8408 2357
rect 8442 2343 8480 2357
rect 8514 2343 8552 2357
rect 8586 2343 8647 2357
rect 8347 2342 8647 2343
rect 8347 2290 8348 2342
rect 8400 2290 8430 2342
rect 8482 2290 8512 2342
rect 8564 2290 8594 2342
rect 8646 2290 8647 2342
rect 8347 2281 8647 2290
rect 8347 2275 8408 2281
rect 8442 2275 8480 2281
rect 8514 2275 8552 2281
rect 8586 2275 8647 2281
rect 8347 2223 8348 2275
rect 8400 2247 8408 2275
rect 8586 2247 8594 2275
rect 8400 2223 8430 2247
rect 8482 2223 8512 2247
rect 8564 2223 8594 2247
rect 8646 2223 8647 2275
rect 8347 2208 8647 2223
rect 8347 2156 8348 2208
rect 8400 2185 8430 2208
rect 8482 2185 8512 2208
rect 8564 2185 8594 2208
rect 8400 2156 8408 2185
rect 8586 2156 8594 2185
rect 8646 2156 8647 2208
rect 8347 2151 8408 2156
rect 8442 2151 8480 2156
rect 8514 2151 8552 2156
rect 8586 2151 8647 2156
rect 8347 2141 8647 2151
rect 8347 2089 8348 2141
rect 8400 2089 8430 2141
rect 8482 2089 8512 2141
rect 8564 2089 8594 2141
rect 8646 2089 8647 2141
rect 8347 2074 8408 2089
rect 8442 2074 8480 2089
rect 8514 2074 8552 2089
rect 8586 2074 8647 2089
rect 8347 2022 8348 2074
rect 8400 2055 8408 2074
rect 8586 2055 8594 2074
rect 8400 2022 8430 2055
rect 8482 2022 8512 2055
rect 8564 2022 8594 2055
rect 8646 2022 8647 2074
rect 8347 1993 8647 2022
rect 8347 1959 8408 1993
rect 8442 1959 8480 1993
rect 8514 1959 8552 1993
rect 8586 1959 8647 1993
rect 8347 1897 8647 1959
rect 8347 1863 8408 1897
rect 8442 1863 8480 1897
rect 8514 1863 8552 1897
rect 8586 1863 8647 1897
rect 8347 1801 8647 1863
rect 8347 1767 8408 1801
rect 8442 1767 8480 1801
rect 8514 1767 8552 1801
rect 8586 1767 8647 1801
rect 8347 1705 8647 1767
rect 8347 1671 8408 1705
rect 8442 1671 8480 1705
rect 8514 1671 8552 1705
rect 8586 1671 8647 1705
rect 8347 1609 8647 1671
rect 8347 1575 8408 1609
rect 8442 1575 8480 1609
rect 8514 1575 8552 1609
rect 8586 1575 8647 1609
rect 8347 1513 8647 1575
rect 8347 1479 8408 1513
rect 8442 1479 8480 1513
rect 8514 1479 8552 1513
rect 8586 1479 8647 1513
rect 8347 1417 8647 1479
rect 8347 1383 8408 1417
rect 8442 1383 8480 1417
rect 8514 1383 8552 1417
rect 8586 1383 8647 1417
rect 8347 1321 8647 1383
rect 8347 1287 8408 1321
rect 8442 1287 8480 1321
rect 8514 1287 8552 1321
rect 8586 1287 8647 1321
rect 8347 1225 8647 1287
rect 8347 1191 8408 1225
rect 8442 1191 8480 1225
rect 8514 1191 8552 1225
rect 8586 1191 8647 1225
rect 8347 1129 8647 1191
rect 8347 1095 8408 1129
rect 8442 1095 8480 1129
rect 8514 1095 8552 1129
rect 8586 1095 8647 1129
rect 8347 1033 8647 1095
rect 8347 999 8408 1033
rect 8442 999 8480 1033
rect 8514 999 8552 1033
rect 8586 999 8647 1033
rect 8347 937 8647 999
rect 8347 903 8408 937
rect 8442 903 8480 937
rect 8514 903 8552 937
rect 8586 903 8647 937
rect 8347 841 8647 903
rect 8347 807 8408 841
rect 8442 807 8480 841
rect 8514 807 8552 841
rect 8586 807 8647 841
rect 8347 745 8647 807
rect 8347 711 8408 745
rect 8442 711 8480 745
rect 8514 711 8552 745
rect 8586 711 8647 745
rect 8347 649 8647 711
rect 8347 615 8408 649
rect 8442 615 8480 649
rect 8514 615 8552 649
rect 8586 615 8647 649
rect 8347 536 8647 615
tri 8347 506 8377 536 ne
rect 8377 506 8587 536
rect 7935 490 8235 503
rect 7935 476 7936 490
tri 7824 395 7905 476 se
rect 7905 438 7936 476
rect 7988 438 8018 490
rect 8070 438 8100 490
rect 8152 438 8182 490
rect 8234 438 8235 490
rect 7905 425 8235 438
rect 7905 395 7936 425
tri 7793 364 7824 395 se
rect 7824 373 7936 395
rect 7988 373 8018 425
rect 8070 373 8100 425
rect 8152 373 8182 425
rect 8234 395 8235 425
tri 8235 395 8346 506 sw
tri 8377 476 8407 506 ne
rect 8407 476 8587 506
tri 8587 476 8647 536 nw
tri 8759 3416 8773 3430 se
rect 8773 3416 9045 3430
tri 9045 3416 9059 3430 sw
rect 8759 3337 9059 3416
rect 8759 3303 8820 3337
rect 8854 3303 8892 3337
rect 8926 3303 8964 3337
rect 8998 3303 9059 3337
rect 8759 3241 9059 3303
rect 8759 3207 8820 3241
rect 8854 3207 8892 3241
rect 8926 3207 8964 3241
rect 8998 3207 9059 3241
rect 8759 3145 9059 3207
rect 8759 3111 8820 3145
rect 8854 3111 8892 3145
rect 8926 3111 8964 3145
rect 8998 3111 9059 3145
rect 8759 3049 9059 3111
rect 8759 3015 8820 3049
rect 8854 3015 8892 3049
rect 8926 3015 8964 3049
rect 8998 3015 9059 3049
rect 8759 2953 9059 3015
rect 8759 2919 8820 2953
rect 8854 2919 8892 2953
rect 8926 2919 8964 2953
rect 8998 2919 9059 2953
rect 8759 2857 9059 2919
rect 8759 2823 8820 2857
rect 8854 2823 8892 2857
rect 8926 2823 8964 2857
rect 8998 2823 9059 2857
rect 8759 2761 9059 2823
rect 8759 2727 8820 2761
rect 8854 2727 8892 2761
rect 8926 2727 8964 2761
rect 8998 2727 9059 2761
rect 8759 2665 9059 2727
rect 8759 2631 8820 2665
rect 8854 2631 8892 2665
rect 8926 2631 8964 2665
rect 8998 2631 9059 2665
rect 8759 2569 9059 2631
rect 8759 2535 8820 2569
rect 8854 2535 8892 2569
rect 8926 2535 8964 2569
rect 8998 2535 9059 2569
rect 8759 2473 9059 2535
rect 8759 2439 8820 2473
rect 8854 2439 8892 2473
rect 8926 2439 8964 2473
rect 8998 2439 9059 2473
rect 8759 2377 9059 2439
rect 8759 2343 8820 2377
rect 8854 2343 8892 2377
rect 8926 2343 8964 2377
rect 8998 2343 9059 2377
rect 8759 2281 9059 2343
rect 8759 2247 8820 2281
rect 8854 2247 8892 2281
rect 8926 2247 8964 2281
rect 8998 2247 9059 2281
rect 8759 2185 9059 2247
rect 8759 2151 8820 2185
rect 8854 2151 8892 2185
rect 8926 2151 8964 2185
rect 8998 2151 9059 2185
rect 8759 2089 9059 2151
rect 8759 2055 8820 2089
rect 8854 2055 8892 2089
rect 8926 2055 8964 2089
rect 8998 2055 9059 2089
rect 8759 1993 9059 2055
rect 8759 1959 8820 1993
rect 8854 1959 8892 1993
rect 8926 1959 8964 1993
rect 8998 1959 9059 1993
rect 8759 1902 9059 1959
rect 8759 1850 8760 1902
rect 8812 1897 8842 1902
rect 8894 1897 8924 1902
rect 8976 1897 9006 1902
rect 8812 1863 8820 1897
rect 8998 1863 9006 1897
rect 8812 1850 8842 1863
rect 8894 1850 8924 1863
rect 8976 1850 9006 1863
rect 9058 1850 9059 1902
rect 8759 1838 9059 1850
rect 8759 1786 8760 1838
rect 8812 1801 8842 1838
rect 8894 1801 8924 1838
rect 8976 1801 9006 1838
rect 8812 1786 8820 1801
rect 8998 1786 9006 1801
rect 9058 1786 9059 1838
rect 8759 1774 8820 1786
rect 8854 1774 8892 1786
rect 8926 1774 8964 1786
rect 8998 1774 9059 1786
rect 8759 1722 8760 1774
rect 8812 1767 8820 1774
rect 8998 1767 9006 1774
rect 8812 1722 8842 1767
rect 8894 1722 8924 1767
rect 8976 1722 9006 1767
rect 9058 1722 9059 1774
rect 8759 1710 9059 1722
rect 8759 1658 8760 1710
rect 8812 1705 8842 1710
rect 8894 1705 8924 1710
rect 8976 1705 9006 1710
rect 8812 1671 8820 1705
rect 8998 1671 9006 1705
rect 8812 1658 8842 1671
rect 8894 1658 8924 1671
rect 8976 1658 9006 1671
rect 9058 1658 9059 1710
rect 8759 1646 9059 1658
rect 8759 1594 8760 1646
rect 8812 1609 8842 1646
rect 8894 1609 8924 1646
rect 8976 1609 9006 1646
rect 8812 1594 8820 1609
rect 8998 1594 9006 1609
rect 9058 1594 9059 1646
rect 8759 1582 8820 1594
rect 8854 1582 8892 1594
rect 8926 1582 8964 1594
rect 8998 1582 9059 1594
rect 8759 1530 8760 1582
rect 8812 1575 8820 1582
rect 8998 1575 9006 1582
rect 8812 1530 8842 1575
rect 8894 1530 8924 1575
rect 8976 1530 9006 1575
rect 9058 1530 9059 1582
rect 8759 1518 9059 1530
rect 8759 1466 8760 1518
rect 8812 1513 8842 1518
rect 8894 1513 8924 1518
rect 8976 1513 9006 1518
rect 8812 1479 8820 1513
rect 8998 1479 9006 1513
rect 8812 1466 8842 1479
rect 8894 1466 8924 1479
rect 8976 1466 9006 1479
rect 9058 1466 9059 1518
rect 8759 1454 9059 1466
rect 8759 1402 8760 1454
rect 8812 1417 8842 1454
rect 8894 1417 8924 1454
rect 8976 1417 9006 1454
rect 8812 1402 8820 1417
rect 8998 1402 9006 1417
rect 9058 1402 9059 1454
rect 8759 1390 8820 1402
rect 8854 1390 8892 1402
rect 8926 1390 8964 1402
rect 8998 1390 9059 1402
rect 8759 1338 8760 1390
rect 8812 1383 8820 1390
rect 8998 1383 9006 1390
rect 8812 1338 8842 1383
rect 8894 1338 8924 1383
rect 8976 1338 9006 1383
rect 9058 1338 9059 1390
rect 8759 1326 9059 1338
rect 8759 1274 8760 1326
rect 8812 1321 8842 1326
rect 8894 1321 8924 1326
rect 8976 1321 9006 1326
rect 8812 1287 8820 1321
rect 8998 1287 9006 1321
rect 8812 1274 8842 1287
rect 8894 1274 8924 1287
rect 8976 1274 9006 1287
rect 9058 1274 9059 1326
rect 8759 1262 9059 1274
rect 8759 1210 8760 1262
rect 8812 1225 8842 1262
rect 8894 1225 8924 1262
rect 8976 1225 9006 1262
rect 8812 1210 8820 1225
rect 8998 1210 9006 1225
rect 9058 1210 9059 1262
rect 8759 1198 8820 1210
rect 8854 1198 8892 1210
rect 8926 1198 8964 1210
rect 8998 1198 9059 1210
rect 8759 1146 8760 1198
rect 8812 1191 8820 1198
rect 8998 1191 9006 1198
rect 8812 1146 8842 1191
rect 8894 1146 8924 1191
rect 8976 1146 9006 1191
rect 9058 1146 9059 1198
rect 8759 1134 9059 1146
rect 8759 1082 8760 1134
rect 8812 1129 8842 1134
rect 8894 1129 8924 1134
rect 8976 1129 9006 1134
rect 8812 1095 8820 1129
rect 8998 1095 9006 1129
rect 8812 1082 8842 1095
rect 8894 1082 8924 1095
rect 8976 1082 9006 1095
rect 9058 1082 9059 1134
rect 8759 1070 9059 1082
rect 8759 1018 8760 1070
rect 8812 1033 8842 1070
rect 8894 1033 8924 1070
rect 8976 1033 9006 1070
rect 8812 1018 8820 1033
rect 8998 1018 9006 1033
rect 9058 1018 9059 1070
rect 8759 1006 8820 1018
rect 8854 1006 8892 1018
rect 8926 1006 8964 1018
rect 8998 1006 9059 1018
rect 8759 954 8760 1006
rect 8812 999 8820 1006
rect 8998 999 9006 1006
rect 8812 954 8842 999
rect 8894 954 8924 999
rect 8976 954 9006 999
rect 9058 954 9059 1006
rect 8759 942 9059 954
rect 8759 890 8760 942
rect 8812 937 8842 942
rect 8894 937 8924 942
rect 8976 937 9006 942
rect 8812 903 8820 937
rect 8998 903 9006 937
rect 8812 890 8842 903
rect 8894 890 8924 903
rect 8976 890 9006 903
rect 9058 890 9059 942
rect 8759 878 9059 890
rect 8759 826 8760 878
rect 8812 841 8842 878
rect 8894 841 8924 878
rect 8976 841 9006 878
rect 8812 826 8820 841
rect 8998 826 9006 841
rect 9058 826 9059 878
rect 8759 814 8820 826
rect 8854 814 8892 826
rect 8926 814 8964 826
rect 8998 814 9059 826
rect 8759 762 8760 814
rect 8812 807 8820 814
rect 8998 807 9006 814
rect 8812 762 8842 807
rect 8894 762 8924 807
rect 8976 762 9006 807
rect 9058 762 9059 814
rect 8759 750 9059 762
rect 8759 698 8760 750
rect 8812 745 8842 750
rect 8894 745 8924 750
rect 8976 745 9006 750
rect 8812 711 8820 745
rect 8998 711 9006 745
rect 8812 698 8842 711
rect 8894 698 8924 711
rect 8976 698 9006 711
rect 9058 698 9059 750
rect 8759 685 9059 698
rect 8759 633 8760 685
rect 8812 649 8842 685
rect 8894 649 8924 685
rect 8976 649 9006 685
rect 8812 633 8820 649
rect 8998 633 9006 649
rect 9058 633 9059 685
rect 8759 620 8820 633
rect 8854 620 8892 633
rect 8926 620 8964 633
rect 8998 620 9059 633
rect 8759 568 8760 620
rect 8812 615 8820 620
rect 8998 615 9006 620
rect 8812 568 8842 615
rect 8894 568 8924 615
rect 8976 568 9006 615
rect 9058 568 9059 620
rect 8759 555 9059 568
tri 8729 476 8759 506 se
rect 8759 503 8760 555
rect 8812 503 8842 555
rect 8894 503 8924 555
rect 8976 503 9006 555
rect 9058 503 9059 555
tri 9171 3416 9185 3430 se
rect 9185 3416 9457 3430
tri 9457 3416 9471 3430 sw
rect 9171 3410 9471 3416
rect 9171 3358 9172 3410
rect 9224 3358 9254 3410
rect 9306 3358 9336 3410
rect 9388 3358 9418 3410
rect 9470 3358 9471 3410
rect 9171 3344 9471 3358
rect 9171 3292 9172 3344
rect 9224 3337 9254 3344
rect 9306 3337 9336 3344
rect 9388 3337 9418 3344
rect 9224 3303 9232 3337
rect 9410 3303 9418 3337
rect 9224 3292 9254 3303
rect 9306 3292 9336 3303
rect 9388 3292 9418 3303
rect 9470 3292 9471 3344
rect 9171 3278 9471 3292
rect 9171 3226 9172 3278
rect 9224 3241 9254 3278
rect 9306 3241 9336 3278
rect 9388 3241 9418 3278
rect 9224 3226 9232 3241
rect 9410 3226 9418 3241
rect 9470 3226 9471 3278
rect 9171 3212 9232 3226
rect 9266 3212 9304 3226
rect 9338 3212 9376 3226
rect 9410 3212 9471 3226
rect 9171 3160 9172 3212
rect 9224 3207 9232 3212
rect 9410 3207 9418 3212
rect 9224 3160 9254 3207
rect 9306 3160 9336 3207
rect 9388 3160 9418 3207
rect 9470 3160 9471 3212
rect 9171 3146 9471 3160
rect 9171 3094 9172 3146
rect 9224 3145 9254 3146
rect 9306 3145 9336 3146
rect 9388 3145 9418 3146
rect 9224 3111 9232 3145
rect 9410 3111 9418 3145
rect 9224 3094 9254 3111
rect 9306 3094 9336 3111
rect 9388 3094 9418 3111
rect 9470 3094 9471 3146
rect 9171 3079 9471 3094
rect 9171 3027 9172 3079
rect 9224 3049 9254 3079
rect 9306 3049 9336 3079
rect 9388 3049 9418 3079
rect 9224 3027 9232 3049
rect 9410 3027 9418 3049
rect 9470 3027 9471 3079
rect 9171 3015 9232 3027
rect 9266 3015 9304 3027
rect 9338 3015 9376 3027
rect 9410 3015 9471 3027
rect 9171 3012 9471 3015
rect 9171 2960 9172 3012
rect 9224 2960 9254 3012
rect 9306 2960 9336 3012
rect 9388 2960 9418 3012
rect 9470 2960 9471 3012
rect 9171 2953 9471 2960
rect 9171 2945 9232 2953
rect 9266 2945 9304 2953
rect 9338 2945 9376 2953
rect 9410 2945 9471 2953
rect 9171 2893 9172 2945
rect 9224 2919 9232 2945
rect 9410 2919 9418 2945
rect 9224 2893 9254 2919
rect 9306 2893 9336 2919
rect 9388 2893 9418 2919
rect 9470 2893 9471 2945
rect 9171 2878 9471 2893
rect 9171 2826 9172 2878
rect 9224 2857 9254 2878
rect 9306 2857 9336 2878
rect 9388 2857 9418 2878
rect 9224 2826 9232 2857
rect 9410 2826 9418 2857
rect 9470 2826 9471 2878
rect 9171 2823 9232 2826
rect 9266 2823 9304 2826
rect 9338 2823 9376 2826
rect 9410 2823 9471 2826
rect 9171 2811 9471 2823
rect 9171 2759 9172 2811
rect 9224 2761 9254 2811
rect 9306 2761 9336 2811
rect 9388 2761 9418 2811
rect 9224 2759 9232 2761
rect 9410 2759 9418 2761
rect 9470 2759 9471 2811
rect 9171 2744 9232 2759
rect 9266 2744 9304 2759
rect 9338 2744 9376 2759
rect 9410 2744 9471 2759
rect 9171 2692 9172 2744
rect 9224 2727 9232 2744
rect 9410 2727 9418 2744
rect 9224 2692 9254 2727
rect 9306 2692 9336 2727
rect 9388 2692 9418 2727
rect 9470 2692 9471 2744
rect 9171 2677 9471 2692
rect 9171 2625 9172 2677
rect 9224 2665 9254 2677
rect 9306 2665 9336 2677
rect 9388 2665 9418 2677
rect 9224 2631 9232 2665
rect 9410 2631 9418 2665
rect 9224 2625 9254 2631
rect 9306 2625 9336 2631
rect 9388 2625 9418 2631
rect 9470 2625 9471 2677
rect 9171 2610 9471 2625
rect 9171 2558 9172 2610
rect 9224 2569 9254 2610
rect 9306 2569 9336 2610
rect 9388 2569 9418 2610
rect 9224 2558 9232 2569
rect 9410 2558 9418 2569
rect 9470 2558 9471 2610
rect 9171 2543 9232 2558
rect 9266 2543 9304 2558
rect 9338 2543 9376 2558
rect 9410 2543 9471 2558
rect 9171 2491 9172 2543
rect 9224 2535 9232 2543
rect 9410 2535 9418 2543
rect 9224 2491 9254 2535
rect 9306 2491 9336 2535
rect 9388 2491 9418 2535
rect 9470 2491 9471 2543
rect 9171 2476 9471 2491
rect 9171 2424 9172 2476
rect 9224 2473 9254 2476
rect 9306 2473 9336 2476
rect 9388 2473 9418 2476
rect 9224 2439 9232 2473
rect 9410 2439 9418 2473
rect 9224 2424 9254 2439
rect 9306 2424 9336 2439
rect 9388 2424 9418 2439
rect 9470 2424 9471 2476
rect 9171 2409 9471 2424
rect 9171 2357 9172 2409
rect 9224 2377 9254 2409
rect 9306 2377 9336 2409
rect 9388 2377 9418 2409
rect 9224 2357 9232 2377
rect 9410 2357 9418 2377
rect 9470 2357 9471 2409
rect 9171 2343 9232 2357
rect 9266 2343 9304 2357
rect 9338 2343 9376 2357
rect 9410 2343 9471 2357
rect 9171 2342 9471 2343
rect 9171 2290 9172 2342
rect 9224 2290 9254 2342
rect 9306 2290 9336 2342
rect 9388 2290 9418 2342
rect 9470 2290 9471 2342
rect 9171 2281 9471 2290
rect 9171 2275 9232 2281
rect 9266 2275 9304 2281
rect 9338 2275 9376 2281
rect 9410 2275 9471 2281
rect 9171 2223 9172 2275
rect 9224 2247 9232 2275
rect 9410 2247 9418 2275
rect 9224 2223 9254 2247
rect 9306 2223 9336 2247
rect 9388 2223 9418 2247
rect 9470 2223 9471 2275
rect 9171 2208 9471 2223
rect 9171 2156 9172 2208
rect 9224 2185 9254 2208
rect 9306 2185 9336 2208
rect 9388 2185 9418 2208
rect 9224 2156 9232 2185
rect 9410 2156 9418 2185
rect 9470 2156 9471 2208
rect 9171 2151 9232 2156
rect 9266 2151 9304 2156
rect 9338 2151 9376 2156
rect 9410 2151 9471 2156
rect 9171 2141 9471 2151
rect 9171 2089 9172 2141
rect 9224 2089 9254 2141
rect 9306 2089 9336 2141
rect 9388 2089 9418 2141
rect 9470 2089 9471 2141
rect 9171 2074 9232 2089
rect 9266 2074 9304 2089
rect 9338 2074 9376 2089
rect 9410 2074 9471 2089
rect 9171 2022 9172 2074
rect 9224 2055 9232 2074
rect 9410 2055 9418 2074
rect 9224 2022 9254 2055
rect 9306 2022 9336 2055
rect 9388 2022 9418 2055
rect 9470 2022 9471 2074
rect 9171 1993 9471 2022
rect 9171 1959 9232 1993
rect 9266 1959 9304 1993
rect 9338 1959 9376 1993
rect 9410 1959 9471 1993
rect 9171 1897 9471 1959
rect 9171 1863 9232 1897
rect 9266 1863 9304 1897
rect 9338 1863 9376 1897
rect 9410 1863 9471 1897
rect 9171 1801 9471 1863
rect 9171 1767 9232 1801
rect 9266 1767 9304 1801
rect 9338 1767 9376 1801
rect 9410 1767 9471 1801
rect 9171 1705 9471 1767
rect 9171 1671 9232 1705
rect 9266 1671 9304 1705
rect 9338 1671 9376 1705
rect 9410 1671 9471 1705
rect 9171 1609 9471 1671
rect 9171 1575 9232 1609
rect 9266 1575 9304 1609
rect 9338 1575 9376 1609
rect 9410 1575 9471 1609
rect 9171 1513 9471 1575
rect 9171 1479 9232 1513
rect 9266 1479 9304 1513
rect 9338 1479 9376 1513
rect 9410 1479 9471 1513
rect 9171 1417 9471 1479
rect 9171 1383 9232 1417
rect 9266 1383 9304 1417
rect 9338 1383 9376 1417
rect 9410 1383 9471 1417
rect 9171 1321 9471 1383
rect 9171 1287 9232 1321
rect 9266 1287 9304 1321
rect 9338 1287 9376 1321
rect 9410 1287 9471 1321
rect 9171 1225 9471 1287
rect 9171 1191 9232 1225
rect 9266 1191 9304 1225
rect 9338 1191 9376 1225
rect 9410 1191 9471 1225
rect 9171 1129 9471 1191
rect 9171 1095 9232 1129
rect 9266 1095 9304 1129
rect 9338 1095 9376 1129
rect 9410 1095 9471 1129
rect 9171 1033 9471 1095
rect 9171 999 9232 1033
rect 9266 999 9304 1033
rect 9338 999 9376 1033
rect 9410 999 9471 1033
rect 9171 937 9471 999
rect 9171 903 9232 937
rect 9266 903 9304 937
rect 9338 903 9376 937
rect 9410 903 9471 937
rect 9171 841 9471 903
rect 9171 807 9232 841
rect 9266 807 9304 841
rect 9338 807 9376 841
rect 9410 807 9471 841
rect 9171 745 9471 807
rect 9171 711 9232 745
rect 9266 711 9304 745
rect 9338 711 9376 745
rect 9410 711 9471 745
rect 9171 649 9471 711
rect 9171 615 9232 649
rect 9266 615 9304 649
rect 9338 615 9376 649
rect 9410 615 9471 649
rect 9171 536 9471 615
tri 9171 506 9201 536 ne
rect 9201 506 9411 536
rect 8759 490 9059 503
rect 8759 476 8760 490
tri 8648 395 8729 476 se
rect 8729 438 8760 476
rect 8812 438 8842 490
rect 8894 438 8924 490
rect 8976 438 9006 490
rect 9058 438 9059 490
rect 8729 425 9059 438
rect 8729 395 8760 425
rect 8234 373 8346 395
rect 7824 364 8346 373
tri 8346 364 8377 395 sw
tri 8617 364 8648 395 se
rect 8648 373 8760 395
rect 8812 373 8842 425
rect 8894 373 8924 425
rect 8976 373 9006 425
rect 9058 395 9059 425
tri 9059 395 9170 506 sw
tri 9201 476 9231 506 ne
rect 9231 476 9411 506
tri 9411 476 9471 536 nw
tri 9583 3416 9597 3430 se
rect 9597 3416 9869 3430
tri 9869 3416 9883 3430 sw
rect 9583 3337 9883 3416
rect 9583 3303 9644 3337
rect 9678 3303 9716 3337
rect 9750 3303 9788 3337
rect 9822 3303 9883 3337
rect 9583 3241 9883 3303
rect 9583 3207 9644 3241
rect 9678 3207 9716 3241
rect 9750 3207 9788 3241
rect 9822 3207 9883 3241
rect 9583 3145 9883 3207
rect 9583 3111 9644 3145
rect 9678 3111 9716 3145
rect 9750 3111 9788 3145
rect 9822 3111 9883 3145
rect 9583 3049 9883 3111
rect 9583 3015 9644 3049
rect 9678 3015 9716 3049
rect 9750 3015 9788 3049
rect 9822 3015 9883 3049
rect 9583 2953 9883 3015
rect 9583 2919 9644 2953
rect 9678 2919 9716 2953
rect 9750 2919 9788 2953
rect 9822 2919 9883 2953
rect 9583 2857 9883 2919
rect 9583 2823 9644 2857
rect 9678 2823 9716 2857
rect 9750 2823 9788 2857
rect 9822 2823 9883 2857
rect 9583 2761 9883 2823
rect 9583 2727 9644 2761
rect 9678 2727 9716 2761
rect 9750 2727 9788 2761
rect 9822 2727 9883 2761
rect 9583 2665 9883 2727
rect 9583 2631 9644 2665
rect 9678 2631 9716 2665
rect 9750 2631 9788 2665
rect 9822 2631 9883 2665
rect 9583 2569 9883 2631
rect 9583 2535 9644 2569
rect 9678 2535 9716 2569
rect 9750 2535 9788 2569
rect 9822 2535 9883 2569
rect 9583 2473 9883 2535
rect 9583 2439 9644 2473
rect 9678 2439 9716 2473
rect 9750 2439 9788 2473
rect 9822 2439 9883 2473
rect 9583 2377 9883 2439
rect 9583 2343 9644 2377
rect 9678 2343 9716 2377
rect 9750 2343 9788 2377
rect 9822 2343 9883 2377
rect 9583 2281 9883 2343
rect 9583 2247 9644 2281
rect 9678 2247 9716 2281
rect 9750 2247 9788 2281
rect 9822 2247 9883 2281
rect 9583 2185 9883 2247
rect 9583 2151 9644 2185
rect 9678 2151 9716 2185
rect 9750 2151 9788 2185
rect 9822 2151 9883 2185
rect 9583 2089 9883 2151
rect 9583 2055 9644 2089
rect 9678 2055 9716 2089
rect 9750 2055 9788 2089
rect 9822 2055 9883 2089
rect 9583 1993 9883 2055
rect 9583 1959 9644 1993
rect 9678 1959 9716 1993
rect 9750 1959 9788 1993
rect 9822 1959 9883 1993
rect 9583 1902 9883 1959
rect 9583 1850 9584 1902
rect 9636 1897 9666 1902
rect 9718 1897 9748 1902
rect 9800 1897 9830 1902
rect 9636 1863 9644 1897
rect 9822 1863 9830 1897
rect 9636 1850 9666 1863
rect 9718 1850 9748 1863
rect 9800 1850 9830 1863
rect 9882 1850 9883 1902
rect 9583 1838 9883 1850
rect 9583 1786 9584 1838
rect 9636 1801 9666 1838
rect 9718 1801 9748 1838
rect 9800 1801 9830 1838
rect 9636 1786 9644 1801
rect 9822 1786 9830 1801
rect 9882 1786 9883 1838
rect 9583 1774 9644 1786
rect 9678 1774 9716 1786
rect 9750 1774 9788 1786
rect 9822 1774 9883 1786
rect 9583 1722 9584 1774
rect 9636 1767 9644 1774
rect 9822 1767 9830 1774
rect 9636 1722 9666 1767
rect 9718 1722 9748 1767
rect 9800 1722 9830 1767
rect 9882 1722 9883 1774
rect 9583 1710 9883 1722
rect 9583 1658 9584 1710
rect 9636 1705 9666 1710
rect 9718 1705 9748 1710
rect 9800 1705 9830 1710
rect 9636 1671 9644 1705
rect 9822 1671 9830 1705
rect 9636 1658 9666 1671
rect 9718 1658 9748 1671
rect 9800 1658 9830 1671
rect 9882 1658 9883 1710
rect 9583 1646 9883 1658
rect 9583 1594 9584 1646
rect 9636 1609 9666 1646
rect 9718 1609 9748 1646
rect 9800 1609 9830 1646
rect 9636 1594 9644 1609
rect 9822 1594 9830 1609
rect 9882 1594 9883 1646
rect 9583 1582 9644 1594
rect 9678 1582 9716 1594
rect 9750 1582 9788 1594
rect 9822 1582 9883 1594
rect 9583 1530 9584 1582
rect 9636 1575 9644 1582
rect 9822 1575 9830 1582
rect 9636 1530 9666 1575
rect 9718 1530 9748 1575
rect 9800 1530 9830 1575
rect 9882 1530 9883 1582
rect 9583 1518 9883 1530
rect 9583 1466 9584 1518
rect 9636 1513 9666 1518
rect 9718 1513 9748 1518
rect 9800 1513 9830 1518
rect 9636 1479 9644 1513
rect 9822 1479 9830 1513
rect 9636 1466 9666 1479
rect 9718 1466 9748 1479
rect 9800 1466 9830 1479
rect 9882 1466 9883 1518
rect 9583 1454 9883 1466
rect 9583 1402 9584 1454
rect 9636 1417 9666 1454
rect 9718 1417 9748 1454
rect 9800 1417 9830 1454
rect 9636 1402 9644 1417
rect 9822 1402 9830 1417
rect 9882 1402 9883 1454
rect 9583 1390 9644 1402
rect 9678 1390 9716 1402
rect 9750 1390 9788 1402
rect 9822 1390 9883 1402
rect 9583 1338 9584 1390
rect 9636 1383 9644 1390
rect 9822 1383 9830 1390
rect 9636 1338 9666 1383
rect 9718 1338 9748 1383
rect 9800 1338 9830 1383
rect 9882 1338 9883 1390
rect 9583 1326 9883 1338
rect 9583 1274 9584 1326
rect 9636 1321 9666 1326
rect 9718 1321 9748 1326
rect 9800 1321 9830 1326
rect 9636 1287 9644 1321
rect 9822 1287 9830 1321
rect 9636 1274 9666 1287
rect 9718 1274 9748 1287
rect 9800 1274 9830 1287
rect 9882 1274 9883 1326
rect 9583 1262 9883 1274
rect 9583 1210 9584 1262
rect 9636 1225 9666 1262
rect 9718 1225 9748 1262
rect 9800 1225 9830 1262
rect 9636 1210 9644 1225
rect 9822 1210 9830 1225
rect 9882 1210 9883 1262
rect 9583 1198 9644 1210
rect 9678 1198 9716 1210
rect 9750 1198 9788 1210
rect 9822 1198 9883 1210
rect 9583 1146 9584 1198
rect 9636 1191 9644 1198
rect 9822 1191 9830 1198
rect 9636 1146 9666 1191
rect 9718 1146 9748 1191
rect 9800 1146 9830 1191
rect 9882 1146 9883 1198
rect 9583 1134 9883 1146
rect 9583 1082 9584 1134
rect 9636 1129 9666 1134
rect 9718 1129 9748 1134
rect 9800 1129 9830 1134
rect 9636 1095 9644 1129
rect 9822 1095 9830 1129
rect 9636 1082 9666 1095
rect 9718 1082 9748 1095
rect 9800 1082 9830 1095
rect 9882 1082 9883 1134
rect 9583 1070 9883 1082
rect 9583 1018 9584 1070
rect 9636 1033 9666 1070
rect 9718 1033 9748 1070
rect 9800 1033 9830 1070
rect 9636 1018 9644 1033
rect 9822 1018 9830 1033
rect 9882 1018 9883 1070
rect 9583 1006 9644 1018
rect 9678 1006 9716 1018
rect 9750 1006 9788 1018
rect 9822 1006 9883 1018
rect 9583 954 9584 1006
rect 9636 999 9644 1006
rect 9822 999 9830 1006
rect 9636 954 9666 999
rect 9718 954 9748 999
rect 9800 954 9830 999
rect 9882 954 9883 1006
rect 9583 942 9883 954
rect 9583 890 9584 942
rect 9636 937 9666 942
rect 9718 937 9748 942
rect 9800 937 9830 942
rect 9636 903 9644 937
rect 9822 903 9830 937
rect 9636 890 9666 903
rect 9718 890 9748 903
rect 9800 890 9830 903
rect 9882 890 9883 942
rect 9583 878 9883 890
rect 9583 826 9584 878
rect 9636 841 9666 878
rect 9718 841 9748 878
rect 9800 841 9830 878
rect 9636 826 9644 841
rect 9822 826 9830 841
rect 9882 826 9883 878
rect 9583 814 9644 826
rect 9678 814 9716 826
rect 9750 814 9788 826
rect 9822 814 9883 826
rect 9583 762 9584 814
rect 9636 807 9644 814
rect 9822 807 9830 814
rect 9636 762 9666 807
rect 9718 762 9748 807
rect 9800 762 9830 807
rect 9882 762 9883 814
rect 9583 750 9883 762
rect 9583 698 9584 750
rect 9636 745 9666 750
rect 9718 745 9748 750
rect 9800 745 9830 750
rect 9636 711 9644 745
rect 9822 711 9830 745
rect 9636 698 9666 711
rect 9718 698 9748 711
rect 9800 698 9830 711
rect 9882 698 9883 750
rect 9583 685 9883 698
rect 9583 633 9584 685
rect 9636 649 9666 685
rect 9718 649 9748 685
rect 9800 649 9830 685
rect 9636 633 9644 649
rect 9822 633 9830 649
rect 9882 633 9883 685
rect 9583 620 9644 633
rect 9678 620 9716 633
rect 9750 620 9788 633
rect 9822 620 9883 633
rect 9583 568 9584 620
rect 9636 615 9644 620
rect 9822 615 9830 620
rect 9636 568 9666 615
rect 9718 568 9748 615
rect 9800 568 9830 615
rect 9882 568 9883 620
rect 9583 555 9883 568
tri 9553 476 9583 506 se
rect 9583 503 9584 555
rect 9636 503 9666 555
rect 9718 503 9748 555
rect 9800 503 9830 555
rect 9882 503 9883 555
tri 9995 3416 10009 3430 se
rect 10009 3416 10281 3430
tri 10281 3416 10295 3430 sw
rect 9995 3410 10295 3416
rect 9995 3358 9996 3410
rect 10048 3358 10078 3410
rect 10130 3358 10160 3410
rect 10212 3358 10242 3410
rect 10294 3358 10295 3410
rect 9995 3344 10295 3358
rect 9995 3292 9996 3344
rect 10048 3337 10078 3344
rect 10130 3337 10160 3344
rect 10212 3337 10242 3344
rect 10048 3303 10056 3337
rect 10234 3303 10242 3337
rect 10048 3292 10078 3303
rect 10130 3292 10160 3303
rect 10212 3292 10242 3303
rect 10294 3292 10295 3344
rect 9995 3278 10295 3292
rect 9995 3226 9996 3278
rect 10048 3241 10078 3278
rect 10130 3241 10160 3278
rect 10212 3241 10242 3278
rect 10048 3226 10056 3241
rect 10234 3226 10242 3241
rect 10294 3226 10295 3278
rect 9995 3212 10056 3226
rect 10090 3212 10128 3226
rect 10162 3212 10200 3226
rect 10234 3212 10295 3226
rect 9995 3160 9996 3212
rect 10048 3207 10056 3212
rect 10234 3207 10242 3212
rect 10048 3160 10078 3207
rect 10130 3160 10160 3207
rect 10212 3160 10242 3207
rect 10294 3160 10295 3212
rect 9995 3146 10295 3160
rect 9995 3094 9996 3146
rect 10048 3145 10078 3146
rect 10130 3145 10160 3146
rect 10212 3145 10242 3146
rect 10048 3111 10056 3145
rect 10234 3111 10242 3145
rect 10048 3094 10078 3111
rect 10130 3094 10160 3111
rect 10212 3094 10242 3111
rect 10294 3094 10295 3146
rect 9995 3079 10295 3094
rect 9995 3027 9996 3079
rect 10048 3049 10078 3079
rect 10130 3049 10160 3079
rect 10212 3049 10242 3079
rect 10048 3027 10056 3049
rect 10234 3027 10242 3049
rect 10294 3027 10295 3079
rect 9995 3015 10056 3027
rect 10090 3015 10128 3027
rect 10162 3015 10200 3027
rect 10234 3015 10295 3027
rect 9995 3012 10295 3015
rect 9995 2960 9996 3012
rect 10048 2960 10078 3012
rect 10130 2960 10160 3012
rect 10212 2960 10242 3012
rect 10294 2960 10295 3012
rect 9995 2953 10295 2960
rect 9995 2945 10056 2953
rect 10090 2945 10128 2953
rect 10162 2945 10200 2953
rect 10234 2945 10295 2953
rect 9995 2893 9996 2945
rect 10048 2919 10056 2945
rect 10234 2919 10242 2945
rect 10048 2893 10078 2919
rect 10130 2893 10160 2919
rect 10212 2893 10242 2919
rect 10294 2893 10295 2945
rect 9995 2878 10295 2893
rect 9995 2826 9996 2878
rect 10048 2857 10078 2878
rect 10130 2857 10160 2878
rect 10212 2857 10242 2878
rect 10048 2826 10056 2857
rect 10234 2826 10242 2857
rect 10294 2826 10295 2878
rect 9995 2823 10056 2826
rect 10090 2823 10128 2826
rect 10162 2823 10200 2826
rect 10234 2823 10295 2826
rect 9995 2811 10295 2823
rect 9995 2759 9996 2811
rect 10048 2761 10078 2811
rect 10130 2761 10160 2811
rect 10212 2761 10242 2811
rect 10048 2759 10056 2761
rect 10234 2759 10242 2761
rect 10294 2759 10295 2811
rect 9995 2744 10056 2759
rect 10090 2744 10128 2759
rect 10162 2744 10200 2759
rect 10234 2744 10295 2759
rect 9995 2692 9996 2744
rect 10048 2727 10056 2744
rect 10234 2727 10242 2744
rect 10048 2692 10078 2727
rect 10130 2692 10160 2727
rect 10212 2692 10242 2727
rect 10294 2692 10295 2744
rect 9995 2677 10295 2692
rect 9995 2625 9996 2677
rect 10048 2665 10078 2677
rect 10130 2665 10160 2677
rect 10212 2665 10242 2677
rect 10048 2631 10056 2665
rect 10234 2631 10242 2665
rect 10048 2625 10078 2631
rect 10130 2625 10160 2631
rect 10212 2625 10242 2631
rect 10294 2625 10295 2677
rect 9995 2610 10295 2625
rect 9995 2558 9996 2610
rect 10048 2569 10078 2610
rect 10130 2569 10160 2610
rect 10212 2569 10242 2610
rect 10048 2558 10056 2569
rect 10234 2558 10242 2569
rect 10294 2558 10295 2610
rect 9995 2543 10056 2558
rect 10090 2543 10128 2558
rect 10162 2543 10200 2558
rect 10234 2543 10295 2558
rect 9995 2491 9996 2543
rect 10048 2535 10056 2543
rect 10234 2535 10242 2543
rect 10048 2491 10078 2535
rect 10130 2491 10160 2535
rect 10212 2491 10242 2535
rect 10294 2491 10295 2543
rect 9995 2476 10295 2491
rect 9995 2424 9996 2476
rect 10048 2473 10078 2476
rect 10130 2473 10160 2476
rect 10212 2473 10242 2476
rect 10048 2439 10056 2473
rect 10234 2439 10242 2473
rect 10048 2424 10078 2439
rect 10130 2424 10160 2439
rect 10212 2424 10242 2439
rect 10294 2424 10295 2476
rect 9995 2409 10295 2424
rect 9995 2357 9996 2409
rect 10048 2377 10078 2409
rect 10130 2377 10160 2409
rect 10212 2377 10242 2409
rect 10048 2357 10056 2377
rect 10234 2357 10242 2377
rect 10294 2357 10295 2409
rect 9995 2343 10056 2357
rect 10090 2343 10128 2357
rect 10162 2343 10200 2357
rect 10234 2343 10295 2357
rect 9995 2342 10295 2343
rect 9995 2290 9996 2342
rect 10048 2290 10078 2342
rect 10130 2290 10160 2342
rect 10212 2290 10242 2342
rect 10294 2290 10295 2342
rect 9995 2281 10295 2290
rect 9995 2275 10056 2281
rect 10090 2275 10128 2281
rect 10162 2275 10200 2281
rect 10234 2275 10295 2281
rect 9995 2223 9996 2275
rect 10048 2247 10056 2275
rect 10234 2247 10242 2275
rect 10048 2223 10078 2247
rect 10130 2223 10160 2247
rect 10212 2223 10242 2247
rect 10294 2223 10295 2275
rect 9995 2208 10295 2223
rect 9995 2156 9996 2208
rect 10048 2185 10078 2208
rect 10130 2185 10160 2208
rect 10212 2185 10242 2208
rect 10048 2156 10056 2185
rect 10234 2156 10242 2185
rect 10294 2156 10295 2208
rect 9995 2151 10056 2156
rect 10090 2151 10128 2156
rect 10162 2151 10200 2156
rect 10234 2151 10295 2156
rect 9995 2141 10295 2151
rect 9995 2089 9996 2141
rect 10048 2089 10078 2141
rect 10130 2089 10160 2141
rect 10212 2089 10242 2141
rect 10294 2089 10295 2141
rect 9995 2074 10056 2089
rect 10090 2074 10128 2089
rect 10162 2074 10200 2089
rect 10234 2074 10295 2089
rect 9995 2022 9996 2074
rect 10048 2055 10056 2074
rect 10234 2055 10242 2074
rect 10048 2022 10078 2055
rect 10130 2022 10160 2055
rect 10212 2022 10242 2055
rect 10294 2022 10295 2074
rect 9995 1993 10295 2022
rect 9995 1959 10056 1993
rect 10090 1959 10128 1993
rect 10162 1959 10200 1993
rect 10234 1959 10295 1993
rect 9995 1897 10295 1959
rect 9995 1863 10056 1897
rect 10090 1863 10128 1897
rect 10162 1863 10200 1897
rect 10234 1863 10295 1897
rect 9995 1801 10295 1863
rect 9995 1767 10056 1801
rect 10090 1767 10128 1801
rect 10162 1767 10200 1801
rect 10234 1767 10295 1801
rect 9995 1705 10295 1767
rect 9995 1671 10056 1705
rect 10090 1671 10128 1705
rect 10162 1671 10200 1705
rect 10234 1671 10295 1705
rect 9995 1609 10295 1671
rect 9995 1575 10056 1609
rect 10090 1575 10128 1609
rect 10162 1575 10200 1609
rect 10234 1575 10295 1609
rect 9995 1513 10295 1575
rect 9995 1479 10056 1513
rect 10090 1479 10128 1513
rect 10162 1479 10200 1513
rect 10234 1479 10295 1513
rect 9995 1417 10295 1479
rect 9995 1383 10056 1417
rect 10090 1383 10128 1417
rect 10162 1383 10200 1417
rect 10234 1383 10295 1417
rect 9995 1321 10295 1383
rect 9995 1287 10056 1321
rect 10090 1287 10128 1321
rect 10162 1287 10200 1321
rect 10234 1287 10295 1321
rect 9995 1225 10295 1287
rect 9995 1191 10056 1225
rect 10090 1191 10128 1225
rect 10162 1191 10200 1225
rect 10234 1191 10295 1225
rect 9995 1129 10295 1191
rect 9995 1095 10056 1129
rect 10090 1095 10128 1129
rect 10162 1095 10200 1129
rect 10234 1095 10295 1129
rect 9995 1033 10295 1095
rect 9995 999 10056 1033
rect 10090 999 10128 1033
rect 10162 999 10200 1033
rect 10234 999 10295 1033
rect 9995 937 10295 999
rect 9995 903 10056 937
rect 10090 903 10128 937
rect 10162 903 10200 937
rect 10234 903 10295 937
rect 9995 841 10295 903
rect 9995 807 10056 841
rect 10090 807 10128 841
rect 10162 807 10200 841
rect 10234 807 10295 841
rect 9995 745 10295 807
rect 9995 711 10056 745
rect 10090 711 10128 745
rect 10162 711 10200 745
rect 10234 711 10295 745
rect 9995 649 10295 711
rect 9995 615 10056 649
rect 10090 615 10128 649
rect 10162 615 10200 649
rect 10234 615 10295 649
rect 9995 536 10295 615
tri 9995 506 10025 536 ne
rect 10025 506 10235 536
rect 9583 490 9883 503
rect 9583 476 9584 490
tri 9472 395 9553 476 se
rect 9553 438 9584 476
rect 9636 438 9666 490
rect 9718 438 9748 490
rect 9800 438 9830 490
rect 9882 438 9883 490
rect 9553 425 9883 438
rect 9553 395 9584 425
rect 9058 373 9170 395
rect 8648 364 9170 373
tri 9170 364 9201 395 sw
tri 9441 364 9472 395 se
rect 9472 373 9584 395
rect 9636 373 9666 425
rect 9718 373 9748 425
rect 9800 373 9830 425
rect 9882 395 9883 425
tri 9883 395 9994 506 sw
tri 10025 476 10055 506 ne
rect 10055 476 10235 506
tri 10235 476 10295 536 nw
tri 10407 3416 10421 3430 se
rect 10421 3416 10693 3430
tri 10693 3416 10707 3430 sw
rect 10407 3337 10707 3416
rect 10407 3303 10468 3337
rect 10502 3303 10540 3337
rect 10574 3303 10612 3337
rect 10646 3303 10707 3337
rect 10407 3241 10707 3303
rect 10407 3207 10468 3241
rect 10502 3207 10540 3241
rect 10574 3207 10612 3241
rect 10646 3207 10707 3241
rect 10407 3145 10707 3207
rect 10407 3111 10468 3145
rect 10502 3111 10540 3145
rect 10574 3111 10612 3145
rect 10646 3111 10707 3145
rect 10407 3049 10707 3111
rect 10407 3015 10468 3049
rect 10502 3015 10540 3049
rect 10574 3015 10612 3049
rect 10646 3015 10707 3049
rect 10407 2953 10707 3015
rect 10407 2919 10468 2953
rect 10502 2919 10540 2953
rect 10574 2919 10612 2953
rect 10646 2919 10707 2953
rect 10407 2857 10707 2919
rect 10407 2823 10468 2857
rect 10502 2823 10540 2857
rect 10574 2823 10612 2857
rect 10646 2823 10707 2857
rect 10407 2761 10707 2823
rect 10407 2727 10468 2761
rect 10502 2727 10540 2761
rect 10574 2727 10612 2761
rect 10646 2727 10707 2761
rect 10407 2665 10707 2727
rect 10407 2631 10468 2665
rect 10502 2631 10540 2665
rect 10574 2631 10612 2665
rect 10646 2631 10707 2665
rect 10407 2569 10707 2631
rect 10407 2535 10468 2569
rect 10502 2535 10540 2569
rect 10574 2535 10612 2569
rect 10646 2535 10707 2569
rect 10407 2473 10707 2535
rect 10407 2439 10468 2473
rect 10502 2439 10540 2473
rect 10574 2439 10612 2473
rect 10646 2439 10707 2473
rect 10407 2377 10707 2439
rect 10407 2343 10468 2377
rect 10502 2343 10540 2377
rect 10574 2343 10612 2377
rect 10646 2343 10707 2377
rect 10407 2281 10707 2343
rect 10407 2247 10468 2281
rect 10502 2247 10540 2281
rect 10574 2247 10612 2281
rect 10646 2247 10707 2281
rect 10407 2185 10707 2247
rect 10407 2151 10468 2185
rect 10502 2151 10540 2185
rect 10574 2151 10612 2185
rect 10646 2151 10707 2185
rect 10407 2089 10707 2151
rect 10407 2055 10468 2089
rect 10502 2055 10540 2089
rect 10574 2055 10612 2089
rect 10646 2055 10707 2089
rect 10407 1993 10707 2055
rect 10407 1959 10468 1993
rect 10502 1959 10540 1993
rect 10574 1959 10612 1993
rect 10646 1959 10707 1993
rect 10407 1902 10707 1959
rect 10407 1850 10408 1902
rect 10460 1897 10490 1902
rect 10542 1897 10572 1902
rect 10624 1897 10654 1902
rect 10460 1863 10468 1897
rect 10646 1863 10654 1897
rect 10460 1850 10490 1863
rect 10542 1850 10572 1863
rect 10624 1850 10654 1863
rect 10706 1850 10707 1902
rect 10407 1838 10707 1850
rect 10407 1786 10408 1838
rect 10460 1801 10490 1838
rect 10542 1801 10572 1838
rect 10624 1801 10654 1838
rect 10460 1786 10468 1801
rect 10646 1786 10654 1801
rect 10706 1786 10707 1838
rect 10407 1774 10468 1786
rect 10502 1774 10540 1786
rect 10574 1774 10612 1786
rect 10646 1774 10707 1786
rect 10407 1722 10408 1774
rect 10460 1767 10468 1774
rect 10646 1767 10654 1774
rect 10460 1722 10490 1767
rect 10542 1722 10572 1767
rect 10624 1722 10654 1767
rect 10706 1722 10707 1774
rect 10407 1710 10707 1722
rect 10407 1658 10408 1710
rect 10460 1705 10490 1710
rect 10542 1705 10572 1710
rect 10624 1705 10654 1710
rect 10460 1671 10468 1705
rect 10646 1671 10654 1705
rect 10460 1658 10490 1671
rect 10542 1658 10572 1671
rect 10624 1658 10654 1671
rect 10706 1658 10707 1710
rect 10407 1646 10707 1658
rect 10407 1594 10408 1646
rect 10460 1609 10490 1646
rect 10542 1609 10572 1646
rect 10624 1609 10654 1646
rect 10460 1594 10468 1609
rect 10646 1594 10654 1609
rect 10706 1594 10707 1646
rect 10407 1582 10468 1594
rect 10502 1582 10540 1594
rect 10574 1582 10612 1594
rect 10646 1582 10707 1594
rect 10407 1530 10408 1582
rect 10460 1575 10468 1582
rect 10646 1575 10654 1582
rect 10460 1530 10490 1575
rect 10542 1530 10572 1575
rect 10624 1530 10654 1575
rect 10706 1530 10707 1582
rect 10407 1518 10707 1530
rect 10407 1466 10408 1518
rect 10460 1513 10490 1518
rect 10542 1513 10572 1518
rect 10624 1513 10654 1518
rect 10460 1479 10468 1513
rect 10646 1479 10654 1513
rect 10460 1466 10490 1479
rect 10542 1466 10572 1479
rect 10624 1466 10654 1479
rect 10706 1466 10707 1518
rect 10407 1454 10707 1466
rect 10407 1402 10408 1454
rect 10460 1417 10490 1454
rect 10542 1417 10572 1454
rect 10624 1417 10654 1454
rect 10460 1402 10468 1417
rect 10646 1402 10654 1417
rect 10706 1402 10707 1454
rect 10407 1390 10468 1402
rect 10502 1390 10540 1402
rect 10574 1390 10612 1402
rect 10646 1390 10707 1402
rect 10407 1338 10408 1390
rect 10460 1383 10468 1390
rect 10646 1383 10654 1390
rect 10460 1338 10490 1383
rect 10542 1338 10572 1383
rect 10624 1338 10654 1383
rect 10706 1338 10707 1390
rect 10407 1326 10707 1338
rect 10407 1274 10408 1326
rect 10460 1321 10490 1326
rect 10542 1321 10572 1326
rect 10624 1321 10654 1326
rect 10460 1287 10468 1321
rect 10646 1287 10654 1321
rect 10460 1274 10490 1287
rect 10542 1274 10572 1287
rect 10624 1274 10654 1287
rect 10706 1274 10707 1326
rect 10407 1262 10707 1274
rect 10407 1210 10408 1262
rect 10460 1225 10490 1262
rect 10542 1225 10572 1262
rect 10624 1225 10654 1262
rect 10460 1210 10468 1225
rect 10646 1210 10654 1225
rect 10706 1210 10707 1262
rect 10407 1198 10468 1210
rect 10502 1198 10540 1210
rect 10574 1198 10612 1210
rect 10646 1198 10707 1210
rect 10407 1146 10408 1198
rect 10460 1191 10468 1198
rect 10646 1191 10654 1198
rect 10460 1146 10490 1191
rect 10542 1146 10572 1191
rect 10624 1146 10654 1191
rect 10706 1146 10707 1198
rect 10407 1134 10707 1146
rect 10407 1082 10408 1134
rect 10460 1129 10490 1134
rect 10542 1129 10572 1134
rect 10624 1129 10654 1134
rect 10460 1095 10468 1129
rect 10646 1095 10654 1129
rect 10460 1082 10490 1095
rect 10542 1082 10572 1095
rect 10624 1082 10654 1095
rect 10706 1082 10707 1134
rect 10407 1070 10707 1082
rect 10407 1018 10408 1070
rect 10460 1033 10490 1070
rect 10542 1033 10572 1070
rect 10624 1033 10654 1070
rect 10460 1018 10468 1033
rect 10646 1018 10654 1033
rect 10706 1018 10707 1070
rect 10407 1006 10468 1018
rect 10502 1006 10540 1018
rect 10574 1006 10612 1018
rect 10646 1006 10707 1018
rect 10407 954 10408 1006
rect 10460 999 10468 1006
rect 10646 999 10654 1006
rect 10460 954 10490 999
rect 10542 954 10572 999
rect 10624 954 10654 999
rect 10706 954 10707 1006
rect 10407 942 10707 954
rect 10407 890 10408 942
rect 10460 937 10490 942
rect 10542 937 10572 942
rect 10624 937 10654 942
rect 10460 903 10468 937
rect 10646 903 10654 937
rect 10460 890 10490 903
rect 10542 890 10572 903
rect 10624 890 10654 903
rect 10706 890 10707 942
rect 10407 878 10707 890
rect 10407 826 10408 878
rect 10460 841 10490 878
rect 10542 841 10572 878
rect 10624 841 10654 878
rect 10460 826 10468 841
rect 10646 826 10654 841
rect 10706 826 10707 878
rect 10407 814 10468 826
rect 10502 814 10540 826
rect 10574 814 10612 826
rect 10646 814 10707 826
rect 10407 762 10408 814
rect 10460 807 10468 814
rect 10646 807 10654 814
rect 10460 762 10490 807
rect 10542 762 10572 807
rect 10624 762 10654 807
rect 10706 762 10707 814
rect 10407 750 10707 762
rect 10407 698 10408 750
rect 10460 745 10490 750
rect 10542 745 10572 750
rect 10624 745 10654 750
rect 10460 711 10468 745
rect 10646 711 10654 745
rect 10460 698 10490 711
rect 10542 698 10572 711
rect 10624 698 10654 711
rect 10706 698 10707 750
rect 10407 685 10707 698
rect 10407 633 10408 685
rect 10460 649 10490 685
rect 10542 649 10572 685
rect 10624 649 10654 685
rect 10460 633 10468 649
rect 10646 633 10654 649
rect 10706 633 10707 685
rect 10407 620 10468 633
rect 10502 620 10540 633
rect 10574 620 10612 633
rect 10646 620 10707 633
rect 10407 568 10408 620
rect 10460 615 10468 620
rect 10646 615 10654 620
rect 10460 568 10490 615
rect 10542 568 10572 615
rect 10624 568 10654 615
rect 10706 568 10707 620
rect 10407 555 10707 568
tri 10377 476 10407 506 se
rect 10407 503 10408 555
rect 10460 503 10490 555
rect 10542 503 10572 555
rect 10624 503 10654 555
rect 10706 503 10707 555
tri 10819 3416 10833 3430 se
rect 10833 3416 11105 3430
tri 11105 3416 11119 3430 sw
rect 10819 3410 11119 3416
rect 10819 3358 10820 3410
rect 10872 3358 10902 3410
rect 10954 3358 10984 3410
rect 11036 3358 11066 3410
rect 11118 3358 11119 3410
rect 10819 3344 11119 3358
rect 10819 3292 10820 3344
rect 10872 3337 10902 3344
rect 10954 3337 10984 3344
rect 11036 3337 11066 3344
rect 10872 3303 10880 3337
rect 11058 3303 11066 3337
rect 10872 3292 10902 3303
rect 10954 3292 10984 3303
rect 11036 3292 11066 3303
rect 11118 3292 11119 3344
rect 10819 3278 11119 3292
rect 10819 3226 10820 3278
rect 10872 3241 10902 3278
rect 10954 3241 10984 3278
rect 11036 3241 11066 3278
rect 10872 3226 10880 3241
rect 11058 3226 11066 3241
rect 11118 3226 11119 3278
rect 10819 3212 10880 3226
rect 10914 3212 10952 3226
rect 10986 3212 11024 3226
rect 11058 3212 11119 3226
rect 10819 3160 10820 3212
rect 10872 3207 10880 3212
rect 11058 3207 11066 3212
rect 10872 3160 10902 3207
rect 10954 3160 10984 3207
rect 11036 3160 11066 3207
rect 11118 3160 11119 3212
rect 10819 3146 11119 3160
rect 10819 3094 10820 3146
rect 10872 3145 10902 3146
rect 10954 3145 10984 3146
rect 11036 3145 11066 3146
rect 10872 3111 10880 3145
rect 11058 3111 11066 3145
rect 10872 3094 10902 3111
rect 10954 3094 10984 3111
rect 11036 3094 11066 3111
rect 11118 3094 11119 3146
rect 10819 3079 11119 3094
rect 10819 3027 10820 3079
rect 10872 3049 10902 3079
rect 10954 3049 10984 3079
rect 11036 3049 11066 3079
rect 10872 3027 10880 3049
rect 11058 3027 11066 3049
rect 11118 3027 11119 3079
rect 10819 3015 10880 3027
rect 10914 3015 10952 3027
rect 10986 3015 11024 3027
rect 11058 3015 11119 3027
rect 10819 3012 11119 3015
rect 10819 2960 10820 3012
rect 10872 2960 10902 3012
rect 10954 2960 10984 3012
rect 11036 2960 11066 3012
rect 11118 2960 11119 3012
rect 10819 2953 11119 2960
rect 10819 2945 10880 2953
rect 10914 2945 10952 2953
rect 10986 2945 11024 2953
rect 11058 2945 11119 2953
rect 10819 2893 10820 2945
rect 10872 2919 10880 2945
rect 11058 2919 11066 2945
rect 10872 2893 10902 2919
rect 10954 2893 10984 2919
rect 11036 2893 11066 2919
rect 11118 2893 11119 2945
rect 10819 2878 11119 2893
rect 10819 2826 10820 2878
rect 10872 2857 10902 2878
rect 10954 2857 10984 2878
rect 11036 2857 11066 2878
rect 10872 2826 10880 2857
rect 11058 2826 11066 2857
rect 11118 2826 11119 2878
rect 10819 2823 10880 2826
rect 10914 2823 10952 2826
rect 10986 2823 11024 2826
rect 11058 2823 11119 2826
rect 10819 2811 11119 2823
rect 10819 2759 10820 2811
rect 10872 2761 10902 2811
rect 10954 2761 10984 2811
rect 11036 2761 11066 2811
rect 10872 2759 10880 2761
rect 11058 2759 11066 2761
rect 11118 2759 11119 2811
rect 10819 2744 10880 2759
rect 10914 2744 10952 2759
rect 10986 2744 11024 2759
rect 11058 2744 11119 2759
rect 10819 2692 10820 2744
rect 10872 2727 10880 2744
rect 11058 2727 11066 2744
rect 10872 2692 10902 2727
rect 10954 2692 10984 2727
rect 11036 2692 11066 2727
rect 11118 2692 11119 2744
rect 10819 2677 11119 2692
rect 10819 2625 10820 2677
rect 10872 2665 10902 2677
rect 10954 2665 10984 2677
rect 11036 2665 11066 2677
rect 10872 2631 10880 2665
rect 11058 2631 11066 2665
rect 10872 2625 10902 2631
rect 10954 2625 10984 2631
rect 11036 2625 11066 2631
rect 11118 2625 11119 2677
rect 10819 2610 11119 2625
rect 10819 2558 10820 2610
rect 10872 2569 10902 2610
rect 10954 2569 10984 2610
rect 11036 2569 11066 2610
rect 10872 2558 10880 2569
rect 11058 2558 11066 2569
rect 11118 2558 11119 2610
rect 10819 2543 10880 2558
rect 10914 2543 10952 2558
rect 10986 2543 11024 2558
rect 11058 2543 11119 2558
rect 10819 2491 10820 2543
rect 10872 2535 10880 2543
rect 11058 2535 11066 2543
rect 10872 2491 10902 2535
rect 10954 2491 10984 2535
rect 11036 2491 11066 2535
rect 11118 2491 11119 2543
rect 10819 2476 11119 2491
rect 10819 2424 10820 2476
rect 10872 2473 10902 2476
rect 10954 2473 10984 2476
rect 11036 2473 11066 2476
rect 10872 2439 10880 2473
rect 11058 2439 11066 2473
rect 10872 2424 10902 2439
rect 10954 2424 10984 2439
rect 11036 2424 11066 2439
rect 11118 2424 11119 2476
rect 10819 2409 11119 2424
rect 10819 2357 10820 2409
rect 10872 2377 10902 2409
rect 10954 2377 10984 2409
rect 11036 2377 11066 2409
rect 10872 2357 10880 2377
rect 11058 2357 11066 2377
rect 11118 2357 11119 2409
rect 10819 2343 10880 2357
rect 10914 2343 10952 2357
rect 10986 2343 11024 2357
rect 11058 2343 11119 2357
rect 10819 2342 11119 2343
rect 10819 2290 10820 2342
rect 10872 2290 10902 2342
rect 10954 2290 10984 2342
rect 11036 2290 11066 2342
rect 11118 2290 11119 2342
rect 10819 2281 11119 2290
rect 10819 2275 10880 2281
rect 10914 2275 10952 2281
rect 10986 2275 11024 2281
rect 11058 2275 11119 2281
rect 10819 2223 10820 2275
rect 10872 2247 10880 2275
rect 11058 2247 11066 2275
rect 10872 2223 10902 2247
rect 10954 2223 10984 2247
rect 11036 2223 11066 2247
rect 11118 2223 11119 2275
rect 10819 2208 11119 2223
rect 10819 2156 10820 2208
rect 10872 2185 10902 2208
rect 10954 2185 10984 2208
rect 11036 2185 11066 2208
rect 10872 2156 10880 2185
rect 11058 2156 11066 2185
rect 11118 2156 11119 2208
rect 10819 2151 10880 2156
rect 10914 2151 10952 2156
rect 10986 2151 11024 2156
rect 11058 2151 11119 2156
rect 10819 2141 11119 2151
rect 10819 2089 10820 2141
rect 10872 2089 10902 2141
rect 10954 2089 10984 2141
rect 11036 2089 11066 2141
rect 11118 2089 11119 2141
rect 10819 2074 10880 2089
rect 10914 2074 10952 2089
rect 10986 2074 11024 2089
rect 11058 2074 11119 2089
rect 10819 2022 10820 2074
rect 10872 2055 10880 2074
rect 11058 2055 11066 2074
rect 10872 2022 10902 2055
rect 10954 2022 10984 2055
rect 11036 2022 11066 2055
rect 11118 2022 11119 2074
rect 10819 1993 11119 2022
rect 10819 1959 10880 1993
rect 10914 1959 10952 1993
rect 10986 1959 11024 1993
rect 11058 1959 11119 1993
rect 10819 1897 11119 1959
rect 10819 1863 10880 1897
rect 10914 1863 10952 1897
rect 10986 1863 11024 1897
rect 11058 1863 11119 1897
rect 10819 1801 11119 1863
rect 10819 1767 10880 1801
rect 10914 1767 10952 1801
rect 10986 1767 11024 1801
rect 11058 1767 11119 1801
rect 10819 1705 11119 1767
rect 10819 1671 10880 1705
rect 10914 1671 10952 1705
rect 10986 1671 11024 1705
rect 11058 1671 11119 1705
rect 10819 1609 11119 1671
rect 10819 1575 10880 1609
rect 10914 1575 10952 1609
rect 10986 1575 11024 1609
rect 11058 1575 11119 1609
rect 10819 1513 11119 1575
rect 10819 1479 10880 1513
rect 10914 1479 10952 1513
rect 10986 1479 11024 1513
rect 11058 1479 11119 1513
rect 10819 1417 11119 1479
rect 10819 1383 10880 1417
rect 10914 1383 10952 1417
rect 10986 1383 11024 1417
rect 11058 1383 11119 1417
rect 10819 1321 11119 1383
rect 10819 1287 10880 1321
rect 10914 1287 10952 1321
rect 10986 1287 11024 1321
rect 11058 1287 11119 1321
rect 10819 1225 11119 1287
rect 10819 1191 10880 1225
rect 10914 1191 10952 1225
rect 10986 1191 11024 1225
rect 11058 1191 11119 1225
rect 10819 1129 11119 1191
rect 10819 1095 10880 1129
rect 10914 1095 10952 1129
rect 10986 1095 11024 1129
rect 11058 1095 11119 1129
rect 10819 1033 11119 1095
rect 10819 999 10880 1033
rect 10914 999 10952 1033
rect 10986 999 11024 1033
rect 11058 999 11119 1033
rect 10819 937 11119 999
rect 10819 903 10880 937
rect 10914 903 10952 937
rect 10986 903 11024 937
rect 11058 903 11119 937
rect 10819 841 11119 903
rect 10819 807 10880 841
rect 10914 807 10952 841
rect 10986 807 11024 841
rect 11058 807 11119 841
rect 10819 745 11119 807
rect 10819 711 10880 745
rect 10914 711 10952 745
rect 10986 711 11024 745
rect 11058 711 11119 745
rect 10819 649 11119 711
rect 10819 615 10880 649
rect 10914 615 10952 649
rect 10986 615 11024 649
rect 11058 615 11119 649
rect 10819 536 11119 615
rect 11231 3392 11313 3430
rect 11231 3358 11252 3392
rect 11286 3358 11313 3392
rect 11231 3320 11313 3358
rect 11231 3286 11252 3320
rect 11286 3286 11313 3320
rect 11231 3248 11313 3286
rect 11231 3214 11252 3248
rect 11286 3214 11313 3248
rect 11231 3176 11313 3214
rect 11231 3142 11252 3176
rect 11286 3142 11313 3176
rect 11231 3104 11313 3142
rect 11231 3070 11252 3104
rect 11286 3070 11313 3104
rect 11231 3032 11313 3070
rect 11231 2998 11252 3032
rect 11286 2998 11313 3032
rect 11231 2960 11313 2998
rect 11231 2926 11252 2960
rect 11286 2926 11313 2960
rect 11231 2888 11313 2926
rect 11231 2854 11252 2888
rect 11286 2854 11313 2888
rect 11231 2816 11313 2854
rect 11231 2782 11252 2816
rect 11286 2782 11313 2816
rect 11231 2744 11313 2782
rect 11231 2710 11252 2744
rect 11286 2710 11313 2744
rect 11231 2672 11313 2710
rect 11231 2638 11252 2672
rect 11286 2638 11313 2672
rect 11231 2600 11313 2638
rect 11231 2566 11252 2600
rect 11286 2566 11313 2600
rect 11231 2528 11313 2566
rect 11231 2494 11252 2528
rect 11286 2494 11313 2528
rect 11231 2456 11313 2494
rect 11231 2422 11252 2456
rect 11286 2422 11313 2456
rect 11231 2384 11313 2422
rect 11231 2350 11252 2384
rect 11286 2350 11313 2384
rect 11231 2312 11313 2350
rect 11231 2278 11252 2312
rect 11286 2278 11313 2312
rect 11231 2240 11313 2278
rect 11231 2206 11252 2240
rect 11286 2206 11313 2240
rect 11231 2168 11313 2206
rect 11231 2134 11252 2168
rect 11286 2134 11313 2168
rect 11231 2096 11313 2134
rect 11231 2062 11252 2096
rect 11286 2062 11313 2096
rect 11231 2024 11313 2062
rect 11231 1990 11252 2024
rect 11286 1990 11313 2024
rect 11231 1952 11313 1990
rect 11231 1918 11252 1952
rect 11286 1918 11313 1952
rect 11231 1880 11313 1918
rect 11231 1846 11252 1880
rect 11286 1846 11313 1880
rect 11231 1808 11313 1846
rect 11231 1774 11252 1808
rect 11286 1774 11313 1808
rect 11231 1736 11313 1774
rect 11231 1702 11252 1736
rect 11286 1702 11313 1736
rect 11231 1664 11313 1702
rect 11231 1630 11252 1664
rect 11286 1630 11313 1664
rect 11231 1592 11313 1630
rect 11231 1558 11252 1592
rect 11286 1558 11313 1592
rect 11231 1520 11313 1558
rect 11231 1486 11252 1520
rect 11286 1486 11313 1520
rect 11231 1448 11313 1486
rect 11231 1414 11252 1448
rect 11286 1414 11313 1448
rect 11231 1376 11313 1414
rect 11231 1342 11252 1376
rect 11286 1342 11313 1376
rect 11231 1304 11313 1342
rect 11231 1270 11252 1304
rect 11286 1270 11313 1304
rect 11231 1232 11313 1270
rect 11231 1198 11252 1232
rect 11286 1198 11313 1232
rect 11231 1160 11313 1198
rect 11231 1126 11252 1160
rect 11286 1126 11313 1160
rect 11231 1088 11313 1126
rect 11231 1054 11252 1088
rect 11286 1054 11313 1088
rect 11231 1016 11313 1054
rect 11231 982 11252 1016
rect 11286 982 11313 1016
rect 11231 944 11313 982
rect 11231 910 11252 944
rect 11286 910 11313 944
rect 11231 872 11313 910
rect 11231 838 11252 872
rect 11286 838 11313 872
rect 11231 800 11313 838
rect 11231 766 11252 800
rect 11286 766 11313 800
rect 11231 728 11313 766
rect 11231 694 11252 728
rect 11286 694 11313 728
rect 11231 656 11313 694
rect 11231 622 11252 656
rect 11286 622 11313 656
rect 11231 609 11313 622
tri 10819 506 10849 536 ne
rect 10849 506 11059 536
rect 10407 490 10707 503
rect 10407 476 10408 490
tri 10296 395 10377 476 se
rect 10377 438 10408 476
rect 10460 438 10490 490
rect 10542 438 10572 490
rect 10624 438 10654 490
rect 10706 438 10707 490
rect 10377 425 10707 438
rect 10377 395 10408 425
rect 9882 373 9994 395
rect 9472 364 9994 373
tri 9994 364 10025 395 sw
tri 10265 364 10296 395 se
rect 10296 373 10408 395
rect 10460 373 10490 425
rect 10542 373 10572 425
rect 10624 373 10654 425
rect 10706 395 10707 425
tri 10707 395 10818 506 sw
tri 10849 476 10879 506 ne
rect 10879 476 11059 506
tri 11059 476 11119 536 nw
tri 11201 476 11231 506 se
rect 11231 476 11313 506
tri 11120 395 11201 476 se
rect 11201 395 11313 476
rect 10706 373 10818 395
rect 10296 364 10818 373
tri 10818 364 10849 395 sw
tri 11089 364 11120 395 se
rect 11120 364 11313 395
rect 7233 356 11313 364
rect 7233 304 7284 356
rect 7336 304 7349 356
rect 7401 304 7414 356
rect 7466 304 7479 356
rect 7531 304 7544 356
rect 7596 304 7609 356
rect 7661 304 7674 356
rect 7726 304 7739 356
rect 7791 304 7804 356
rect 7856 304 7869 356
rect 7921 304 7934 356
rect 7986 304 7999 356
rect 8051 304 8064 356
rect 8116 304 8129 356
rect 8181 304 8194 356
rect 8246 304 8259 356
rect 8311 304 8324 356
rect 8376 304 8389 356
rect 8441 304 8454 356
rect 8506 304 8519 356
rect 8571 304 8584 356
rect 8636 304 8649 356
rect 8701 304 8714 356
rect 8766 304 8779 356
rect 8831 304 8844 356
rect 8896 304 8909 356
rect 8961 304 8974 356
rect 9026 304 9039 356
rect 9091 304 9104 356
rect 9156 304 9169 356
rect 9221 304 9234 356
rect 9286 304 9299 356
rect 9351 304 9364 356
rect 9416 304 9429 356
rect 9481 304 9494 356
rect 9546 304 9559 356
rect 9611 304 9624 356
rect 9676 304 9689 356
rect 9741 304 9753 356
rect 9805 304 9817 356
rect 9869 304 9881 356
rect 9933 304 9945 356
rect 9997 304 10009 356
rect 10061 304 10073 356
rect 10125 304 10137 356
rect 10189 304 10201 356
rect 10253 304 10265 356
rect 10317 304 10329 356
rect 10381 304 10393 356
rect 10445 304 10457 356
rect 10509 304 10521 356
rect 10573 304 10585 356
rect 10637 304 10649 356
rect 10701 304 11313 356
rect 7233 282 11313 304
rect 7233 230 7284 282
rect 7336 230 7349 282
rect 7401 230 7414 282
rect 7466 230 7479 282
rect 7531 230 7544 282
rect 7596 230 7609 282
rect 7661 230 7674 282
rect 7726 230 7739 282
rect 7791 230 7804 282
rect 7856 230 7869 282
rect 7921 230 7934 282
rect 7986 230 7999 282
rect 8051 230 8064 282
rect 8116 230 8129 282
rect 8181 230 8194 282
rect 8246 230 8259 282
rect 8311 230 8324 282
rect 8376 230 8389 282
rect 8441 230 8454 282
rect 8506 230 8519 282
rect 8571 230 8584 282
rect 8636 230 8649 282
rect 8701 230 8714 282
rect 8766 230 8779 282
rect 8831 230 8844 282
rect 8896 230 8909 282
rect 8961 230 8974 282
rect 9026 230 9039 282
rect 9091 230 9104 282
rect 9156 230 9169 282
rect 9221 230 9234 282
rect 9286 230 9299 282
rect 9351 230 9364 282
rect 9416 230 9429 282
rect 9481 230 9494 282
rect 9546 230 9559 282
rect 9611 230 9624 282
rect 9676 230 9689 282
rect 9741 230 9753 282
rect 9805 230 9817 282
rect 9869 230 9881 282
rect 9933 230 9945 282
rect 9997 230 10009 282
rect 10061 230 10073 282
rect 10125 230 10137 282
rect 10189 230 10201 282
rect 10253 230 10265 282
rect 10317 230 10329 282
rect 10381 230 10393 282
rect 10445 230 10457 282
rect 10509 230 10521 282
rect 10573 230 10585 282
rect 10637 230 10649 282
rect 10701 230 11313 282
rect 7233 208 11313 230
rect 7233 156 7284 208
rect 7336 156 7349 208
rect 7401 156 7414 208
rect 7466 156 7479 208
rect 7531 156 7544 208
rect 7596 156 7609 208
rect 7661 156 7674 208
rect 7726 156 7739 208
rect 7791 156 7804 208
rect 7856 156 7869 208
rect 7921 156 7934 208
rect 7986 156 7999 208
rect 8051 156 8064 208
rect 8116 156 8129 208
rect 8181 156 8194 208
rect 8246 156 8259 208
rect 8311 156 8324 208
rect 8376 156 8389 208
rect 8441 156 8454 208
rect 8506 156 8519 208
rect 8571 156 8584 208
rect 8636 156 8649 208
rect 8701 156 8714 208
rect 8766 156 8779 208
rect 8831 156 8844 208
rect 8896 156 8909 208
rect 8961 156 8974 208
rect 9026 156 9039 208
rect 9091 156 9104 208
rect 9156 156 9169 208
rect 9221 156 9234 208
rect 9286 156 9299 208
rect 9351 156 9364 208
rect 9416 156 9429 208
rect 9481 156 9494 208
rect 9546 156 9559 208
rect 9611 156 9624 208
rect 9676 156 9689 208
rect 9741 156 9753 208
rect 9805 156 9817 208
rect 9869 156 9881 208
rect 9933 156 9945 208
rect 9997 156 10009 208
rect 10061 156 10073 208
rect 10125 156 10137 208
rect 10189 156 10201 208
rect 10253 156 10265 208
rect 10317 156 10329 208
rect 10381 156 10393 208
rect 10445 156 10457 208
rect 10509 156 10521 208
rect 10573 156 10585 208
rect 10637 156 10649 208
rect 10701 156 11313 208
rect 7233 134 11313 156
rect 7233 82 7284 134
rect 7336 82 7349 134
rect 7401 82 7414 134
rect 7466 82 7479 134
rect 7531 82 7544 134
rect 7596 82 7609 134
rect 7661 82 7674 134
rect 7726 82 7739 134
rect 7791 82 7804 134
rect 7856 82 7869 134
rect 7921 82 7934 134
rect 7986 82 7999 134
rect 8051 82 8064 134
rect 8116 82 8129 134
rect 8181 82 8194 134
rect 8246 82 8259 134
rect 8311 82 8324 134
rect 8376 82 8389 134
rect 8441 82 8454 134
rect 8506 82 8519 134
rect 8571 82 8584 134
rect 8636 82 8649 134
rect 8701 82 8714 134
rect 8766 82 8779 134
rect 8831 82 8844 134
rect 8896 82 8909 134
rect 8961 82 8974 134
rect 9026 82 9039 134
rect 9091 82 9104 134
rect 9156 82 9169 134
rect 9221 82 9234 134
rect 9286 82 9299 134
rect 9351 82 9364 134
rect 9416 82 9429 134
rect 9481 82 9494 134
rect 9546 82 9559 134
rect 9611 82 9624 134
rect 9676 82 9689 134
rect 9741 82 9753 134
rect 9805 82 9817 134
rect 9869 82 9881 134
rect 9933 82 9945 134
rect 9997 82 10009 134
rect 10061 82 10073 134
rect 10125 82 10137 134
rect 10189 82 10201 134
rect 10253 82 10265 134
rect 10317 82 10329 134
rect 10381 82 10393 134
rect 10445 82 10457 134
rect 10509 82 10521 134
rect 10573 82 10585 134
rect 10637 82 10649 134
rect 10701 82 11313 134
rect 7233 60 11313 82
rect 7233 8 7284 60
rect 7336 8 7349 60
rect 7401 8 7414 60
rect 7466 8 7479 60
rect 7531 8 7544 60
rect 7596 8 7609 60
rect 7661 8 7674 60
rect 7726 8 7739 60
rect 7791 8 7804 60
rect 7856 8 7869 60
rect 7921 8 7934 60
rect 7986 8 7999 60
rect 8051 8 8064 60
rect 8116 8 8129 60
rect 8181 8 8194 60
rect 8246 8 8259 60
rect 8311 8 8324 60
rect 8376 8 8389 60
rect 8441 8 8454 60
rect 8506 8 8519 60
rect 8571 8 8584 60
rect 8636 8 8649 60
rect 8701 8 8714 60
rect 8766 8 8779 60
rect 8831 8 8844 60
rect 8896 8 8909 60
rect 8961 8 8974 60
rect 9026 8 9039 60
rect 9091 8 9104 60
rect 9156 8 9169 60
rect 9221 8 9234 60
rect 9286 8 9299 60
rect 9351 8 9364 60
rect 9416 8 9429 60
rect 9481 8 9494 60
rect 9546 8 9559 60
rect 9611 8 9624 60
rect 9676 8 9689 60
rect 9741 8 9753 60
rect 9805 8 9817 60
rect 9869 8 9881 60
rect 9933 8 9945 60
rect 9997 8 10009 60
rect 10061 8 10073 60
rect 10125 8 10137 60
rect 10189 8 10201 60
rect 10253 8 10265 60
rect 10317 8 10329 60
rect 10381 8 10393 60
rect 10445 8 10457 60
rect 10509 8 10521 60
rect 10573 8 10585 60
rect 10637 8 10649 60
rect 10701 8 11313 60
rect 7233 0 11313 8
<< via1 >>
rect 7290 3614 7342 3666
rect 7355 3614 7407 3666
rect 7419 3664 7471 3666
rect 7419 3630 7428 3664
rect 7428 3630 7462 3664
rect 7462 3630 7471 3664
rect 7419 3614 7471 3630
rect 7483 3664 7535 3666
rect 7483 3630 7501 3664
rect 7501 3630 7535 3664
rect 7483 3614 7535 3630
rect 7547 3664 7599 3666
rect 7611 3664 7663 3666
rect 7675 3664 7727 3666
rect 7739 3664 7791 3666
rect 7803 3664 7855 3666
rect 7867 3664 7919 3666
rect 7547 3630 7574 3664
rect 7574 3630 7599 3664
rect 7611 3630 7646 3664
rect 7646 3630 7663 3664
rect 7675 3630 7680 3664
rect 7680 3630 7718 3664
rect 7718 3630 7727 3664
rect 7739 3630 7752 3664
rect 7752 3630 7790 3664
rect 7790 3630 7791 3664
rect 7803 3630 7824 3664
rect 7824 3630 7855 3664
rect 7867 3630 7896 3664
rect 7896 3630 7919 3664
rect 7547 3614 7599 3630
rect 7611 3614 7663 3630
rect 7675 3614 7727 3630
rect 7739 3614 7791 3630
rect 7803 3614 7855 3630
rect 7867 3614 7919 3630
rect 7931 3664 7983 3666
rect 7931 3630 7934 3664
rect 7934 3630 7968 3664
rect 7968 3630 7983 3664
rect 7931 3614 7983 3630
rect 7995 3664 8047 3666
rect 7995 3630 8006 3664
rect 8006 3630 8040 3664
rect 8040 3630 8047 3664
rect 7995 3614 8047 3630
rect 8059 3664 8111 3666
rect 8123 3664 8175 3666
rect 8187 3664 8239 3666
rect 8251 3664 8303 3666
rect 8315 3664 8367 3666
rect 8379 3664 8431 3666
rect 8443 3664 8495 3666
rect 8059 3630 8078 3664
rect 8078 3630 8111 3664
rect 8123 3630 8150 3664
rect 8150 3630 8175 3664
rect 8187 3630 8222 3664
rect 8222 3630 8239 3664
rect 8251 3630 8256 3664
rect 8256 3630 8294 3664
rect 8294 3630 8303 3664
rect 8315 3630 8328 3664
rect 8328 3630 8366 3664
rect 8366 3630 8367 3664
rect 8379 3630 8400 3664
rect 8400 3630 8431 3664
rect 8443 3630 8472 3664
rect 8472 3630 8495 3664
rect 8059 3614 8111 3630
rect 8123 3614 8175 3630
rect 8187 3614 8239 3630
rect 8251 3614 8303 3630
rect 8315 3614 8367 3630
rect 8379 3614 8431 3630
rect 8443 3614 8495 3630
rect 8507 3664 8559 3666
rect 8507 3630 8510 3664
rect 8510 3630 8544 3664
rect 8544 3630 8559 3664
rect 8507 3614 8559 3630
rect 8571 3664 8623 3666
rect 8571 3630 8582 3664
rect 8582 3630 8616 3664
rect 8616 3630 8623 3664
rect 8571 3614 8623 3630
rect 8635 3664 8687 3666
rect 8699 3664 8751 3666
rect 8763 3664 8815 3666
rect 8827 3664 8879 3666
rect 8891 3664 8943 3666
rect 8955 3664 9007 3666
rect 9019 3664 9071 3666
rect 8635 3630 8654 3664
rect 8654 3630 8687 3664
rect 8699 3630 8726 3664
rect 8726 3630 8751 3664
rect 8763 3630 8798 3664
rect 8798 3630 8815 3664
rect 8827 3630 8832 3664
rect 8832 3630 8870 3664
rect 8870 3630 8879 3664
rect 8891 3630 8904 3664
rect 8904 3630 8942 3664
rect 8942 3630 8943 3664
rect 8955 3630 8976 3664
rect 8976 3630 9007 3664
rect 9019 3630 9048 3664
rect 9048 3630 9071 3664
rect 8635 3614 8687 3630
rect 8699 3614 8751 3630
rect 8763 3614 8815 3630
rect 8827 3614 8879 3630
rect 8891 3614 8943 3630
rect 8955 3614 9007 3630
rect 9019 3614 9071 3630
rect 9083 3664 9135 3666
rect 9083 3630 9086 3664
rect 9086 3630 9120 3664
rect 9120 3630 9135 3664
rect 9083 3614 9135 3630
rect 9147 3664 9199 3666
rect 9147 3630 9158 3664
rect 9158 3630 9192 3664
rect 9192 3630 9199 3664
rect 9147 3614 9199 3630
rect 9211 3664 9263 3666
rect 9275 3664 9327 3666
rect 9339 3664 9391 3666
rect 9403 3664 9455 3666
rect 9467 3664 9519 3666
rect 9531 3664 9583 3666
rect 9595 3664 9647 3666
rect 9211 3630 9230 3664
rect 9230 3630 9263 3664
rect 9275 3630 9302 3664
rect 9302 3630 9327 3664
rect 9339 3630 9374 3664
rect 9374 3630 9391 3664
rect 9403 3630 9408 3664
rect 9408 3630 9446 3664
rect 9446 3630 9455 3664
rect 9467 3630 9480 3664
rect 9480 3630 9518 3664
rect 9518 3630 9519 3664
rect 9531 3630 9552 3664
rect 9552 3630 9583 3664
rect 9595 3630 9624 3664
rect 9624 3630 9647 3664
rect 9211 3614 9263 3630
rect 9275 3614 9327 3630
rect 9339 3614 9391 3630
rect 9403 3614 9455 3630
rect 9467 3614 9519 3630
rect 9531 3614 9583 3630
rect 9595 3614 9647 3630
rect 9659 3664 9711 3666
rect 9659 3630 9662 3664
rect 9662 3630 9696 3664
rect 9696 3630 9711 3664
rect 9659 3614 9711 3630
rect 9723 3664 9775 3666
rect 9723 3630 9734 3664
rect 9734 3630 9768 3664
rect 9768 3630 9775 3664
rect 9723 3614 9775 3630
rect 9787 3664 9839 3666
rect 9851 3664 9903 3666
rect 9915 3664 9967 3666
rect 9979 3664 10031 3666
rect 10043 3664 10095 3666
rect 10107 3664 10159 3666
rect 10171 3664 10223 3666
rect 9787 3630 9806 3664
rect 9806 3630 9839 3664
rect 9851 3630 9878 3664
rect 9878 3630 9903 3664
rect 9915 3630 9950 3664
rect 9950 3630 9967 3664
rect 9979 3630 9984 3664
rect 9984 3630 10022 3664
rect 10022 3630 10031 3664
rect 10043 3630 10056 3664
rect 10056 3630 10094 3664
rect 10094 3630 10095 3664
rect 10107 3630 10128 3664
rect 10128 3630 10159 3664
rect 10171 3630 10200 3664
rect 10200 3630 10223 3664
rect 9787 3614 9839 3630
rect 9851 3614 9903 3630
rect 9915 3614 9967 3630
rect 9979 3614 10031 3630
rect 10043 3614 10095 3630
rect 10107 3614 10159 3630
rect 10171 3614 10223 3630
rect 10235 3664 10287 3666
rect 10235 3630 10238 3664
rect 10238 3630 10272 3664
rect 10272 3630 10287 3664
rect 10235 3614 10287 3630
rect 10299 3664 10351 3666
rect 10299 3630 10310 3664
rect 10310 3630 10344 3664
rect 10344 3630 10351 3664
rect 10299 3614 10351 3630
rect 10363 3664 10415 3666
rect 10427 3664 10479 3666
rect 10491 3664 10543 3666
rect 10555 3664 10607 3666
rect 10619 3664 10671 3666
rect 10683 3664 10735 3666
rect 10747 3664 10799 3666
rect 10363 3630 10382 3664
rect 10382 3630 10415 3664
rect 10427 3630 10454 3664
rect 10454 3630 10479 3664
rect 10491 3630 10526 3664
rect 10526 3630 10543 3664
rect 10555 3630 10560 3664
rect 10560 3630 10598 3664
rect 10598 3630 10607 3664
rect 10619 3630 10632 3664
rect 10632 3630 10670 3664
rect 10670 3630 10671 3664
rect 10683 3630 10704 3664
rect 10704 3630 10735 3664
rect 10747 3630 10776 3664
rect 10776 3630 10799 3664
rect 10363 3614 10415 3630
rect 10427 3614 10479 3630
rect 10491 3614 10543 3630
rect 10555 3614 10607 3630
rect 10619 3614 10671 3630
rect 10683 3614 10735 3630
rect 10747 3614 10799 3630
rect 10811 3664 10863 3666
rect 10811 3630 10814 3664
rect 10814 3630 10848 3664
rect 10848 3630 10863 3664
rect 10811 3614 10863 3630
rect 7290 3526 7342 3578
rect 7355 3536 7407 3578
rect 7355 3526 7384 3536
rect 7384 3526 7407 3536
rect 7419 3526 7471 3578
rect 7483 3526 7535 3578
rect 7547 3526 7599 3578
rect 7611 3526 7663 3578
rect 7675 3526 7727 3578
rect 7739 3526 7791 3578
rect 7803 3526 7855 3578
rect 7867 3526 7919 3578
rect 7931 3526 7983 3578
rect 7995 3526 8047 3578
rect 8059 3526 8111 3578
rect 8123 3526 8175 3578
rect 8187 3526 8239 3578
rect 8251 3526 8303 3578
rect 8315 3526 8367 3578
rect 8379 3526 8431 3578
rect 8443 3526 8495 3578
rect 8507 3526 8559 3578
rect 8571 3526 8623 3578
rect 8635 3526 8687 3578
rect 8699 3526 8751 3578
rect 8763 3526 8815 3578
rect 8827 3526 8879 3578
rect 8891 3526 8943 3578
rect 8955 3526 9007 3578
rect 9019 3526 9071 3578
rect 9083 3526 9135 3578
rect 9147 3526 9199 3578
rect 9211 3526 9263 3578
rect 9275 3526 9327 3578
rect 9339 3526 9391 3578
rect 9403 3526 9455 3578
rect 9467 3526 9519 3578
rect 9531 3526 9583 3578
rect 9595 3526 9647 3578
rect 9659 3526 9711 3578
rect 9723 3526 9775 3578
rect 9787 3526 9839 3578
rect 9851 3526 9903 3578
rect 9915 3526 9967 3578
rect 9979 3526 10031 3578
rect 10043 3526 10095 3578
rect 10107 3526 10159 3578
rect 10171 3526 10223 3578
rect 10235 3526 10287 3578
rect 10299 3526 10351 3578
rect 10363 3526 10415 3578
rect 10427 3526 10479 3578
rect 10491 3526 10543 3578
rect 10555 3526 10607 3578
rect 10619 3526 10671 3578
rect 10683 3526 10735 3578
rect 10747 3526 10799 3578
rect 10811 3526 10863 3578
rect 7524 3358 7576 3410
rect 7606 3358 7658 3410
rect 7688 3358 7740 3410
rect 7770 3358 7822 3410
rect 7524 3292 7576 3344
rect 7606 3337 7658 3344
rect 7688 3337 7740 3344
rect 7606 3303 7618 3337
rect 7618 3303 7656 3337
rect 7656 3303 7658 3337
rect 7688 3303 7690 3337
rect 7690 3303 7728 3337
rect 7728 3303 7740 3337
rect 7606 3292 7658 3303
rect 7688 3292 7740 3303
rect 7770 3292 7822 3344
rect 7524 3226 7576 3278
rect 7606 3241 7658 3278
rect 7688 3241 7740 3278
rect 7606 3226 7618 3241
rect 7618 3226 7656 3241
rect 7656 3226 7658 3241
rect 7688 3226 7690 3241
rect 7690 3226 7728 3241
rect 7728 3226 7740 3241
rect 7770 3226 7822 3278
rect 7524 3160 7576 3212
rect 7606 3207 7618 3212
rect 7618 3207 7656 3212
rect 7656 3207 7658 3212
rect 7688 3207 7690 3212
rect 7690 3207 7728 3212
rect 7728 3207 7740 3212
rect 7606 3160 7658 3207
rect 7688 3160 7740 3207
rect 7770 3160 7822 3212
rect 7524 3094 7576 3146
rect 7606 3145 7658 3146
rect 7688 3145 7740 3146
rect 7606 3111 7618 3145
rect 7618 3111 7656 3145
rect 7656 3111 7658 3145
rect 7688 3111 7690 3145
rect 7690 3111 7728 3145
rect 7728 3111 7740 3145
rect 7606 3094 7658 3111
rect 7688 3094 7740 3111
rect 7770 3094 7822 3146
rect 7524 3027 7576 3079
rect 7606 3049 7658 3079
rect 7688 3049 7740 3079
rect 7606 3027 7618 3049
rect 7618 3027 7656 3049
rect 7656 3027 7658 3049
rect 7688 3027 7690 3049
rect 7690 3027 7728 3049
rect 7728 3027 7740 3049
rect 7770 3027 7822 3079
rect 7524 2960 7576 3012
rect 7606 2960 7658 3012
rect 7688 2960 7740 3012
rect 7770 2960 7822 3012
rect 7524 2893 7576 2945
rect 7606 2919 7618 2945
rect 7618 2919 7656 2945
rect 7656 2919 7658 2945
rect 7688 2919 7690 2945
rect 7690 2919 7728 2945
rect 7728 2919 7740 2945
rect 7606 2893 7658 2919
rect 7688 2893 7740 2919
rect 7770 2893 7822 2945
rect 7524 2826 7576 2878
rect 7606 2857 7658 2878
rect 7688 2857 7740 2878
rect 7606 2826 7618 2857
rect 7618 2826 7656 2857
rect 7656 2826 7658 2857
rect 7688 2826 7690 2857
rect 7690 2826 7728 2857
rect 7728 2826 7740 2857
rect 7770 2826 7822 2878
rect 7524 2759 7576 2811
rect 7606 2761 7658 2811
rect 7688 2761 7740 2811
rect 7606 2759 7618 2761
rect 7618 2759 7656 2761
rect 7656 2759 7658 2761
rect 7688 2759 7690 2761
rect 7690 2759 7728 2761
rect 7728 2759 7740 2761
rect 7770 2759 7822 2811
rect 7524 2692 7576 2744
rect 7606 2727 7618 2744
rect 7618 2727 7656 2744
rect 7656 2727 7658 2744
rect 7688 2727 7690 2744
rect 7690 2727 7728 2744
rect 7728 2727 7740 2744
rect 7606 2692 7658 2727
rect 7688 2692 7740 2727
rect 7770 2692 7822 2744
rect 7524 2625 7576 2677
rect 7606 2665 7658 2677
rect 7688 2665 7740 2677
rect 7606 2631 7618 2665
rect 7618 2631 7656 2665
rect 7656 2631 7658 2665
rect 7688 2631 7690 2665
rect 7690 2631 7728 2665
rect 7728 2631 7740 2665
rect 7606 2625 7658 2631
rect 7688 2625 7740 2631
rect 7770 2625 7822 2677
rect 7524 2558 7576 2610
rect 7606 2569 7658 2610
rect 7688 2569 7740 2610
rect 7606 2558 7618 2569
rect 7618 2558 7656 2569
rect 7656 2558 7658 2569
rect 7688 2558 7690 2569
rect 7690 2558 7728 2569
rect 7728 2558 7740 2569
rect 7770 2558 7822 2610
rect 7524 2491 7576 2543
rect 7606 2535 7618 2543
rect 7618 2535 7656 2543
rect 7656 2535 7658 2543
rect 7688 2535 7690 2543
rect 7690 2535 7728 2543
rect 7728 2535 7740 2543
rect 7606 2491 7658 2535
rect 7688 2491 7740 2535
rect 7770 2491 7822 2543
rect 7524 2424 7576 2476
rect 7606 2473 7658 2476
rect 7688 2473 7740 2476
rect 7606 2439 7618 2473
rect 7618 2439 7656 2473
rect 7656 2439 7658 2473
rect 7688 2439 7690 2473
rect 7690 2439 7728 2473
rect 7728 2439 7740 2473
rect 7606 2424 7658 2439
rect 7688 2424 7740 2439
rect 7770 2424 7822 2476
rect 7524 2357 7576 2409
rect 7606 2377 7658 2409
rect 7688 2377 7740 2409
rect 7606 2357 7618 2377
rect 7618 2357 7656 2377
rect 7656 2357 7658 2377
rect 7688 2357 7690 2377
rect 7690 2357 7728 2377
rect 7728 2357 7740 2377
rect 7770 2357 7822 2409
rect 7524 2290 7576 2342
rect 7606 2290 7658 2342
rect 7688 2290 7740 2342
rect 7770 2290 7822 2342
rect 7524 2223 7576 2275
rect 7606 2247 7618 2275
rect 7618 2247 7656 2275
rect 7656 2247 7658 2275
rect 7688 2247 7690 2275
rect 7690 2247 7728 2275
rect 7728 2247 7740 2275
rect 7606 2223 7658 2247
rect 7688 2223 7740 2247
rect 7770 2223 7822 2275
rect 7524 2156 7576 2208
rect 7606 2185 7658 2208
rect 7688 2185 7740 2208
rect 7606 2156 7618 2185
rect 7618 2156 7656 2185
rect 7656 2156 7658 2185
rect 7688 2156 7690 2185
rect 7690 2156 7728 2185
rect 7728 2156 7740 2185
rect 7770 2156 7822 2208
rect 7524 2089 7576 2141
rect 7606 2089 7658 2141
rect 7688 2089 7740 2141
rect 7770 2089 7822 2141
rect 7524 2022 7576 2074
rect 7606 2055 7618 2074
rect 7618 2055 7656 2074
rect 7656 2055 7658 2074
rect 7688 2055 7690 2074
rect 7690 2055 7728 2074
rect 7728 2055 7740 2074
rect 7606 2022 7658 2055
rect 7688 2022 7740 2055
rect 7770 2022 7822 2074
rect 7936 1850 7988 1902
rect 8018 1897 8070 1902
rect 8100 1897 8152 1902
rect 8018 1863 8030 1897
rect 8030 1863 8068 1897
rect 8068 1863 8070 1897
rect 8100 1863 8102 1897
rect 8102 1863 8140 1897
rect 8140 1863 8152 1897
rect 8018 1850 8070 1863
rect 8100 1850 8152 1863
rect 8182 1850 8234 1902
rect 7936 1786 7988 1838
rect 8018 1801 8070 1838
rect 8100 1801 8152 1838
rect 8018 1786 8030 1801
rect 8030 1786 8068 1801
rect 8068 1786 8070 1801
rect 8100 1786 8102 1801
rect 8102 1786 8140 1801
rect 8140 1786 8152 1801
rect 8182 1786 8234 1838
rect 7936 1722 7988 1774
rect 8018 1767 8030 1774
rect 8030 1767 8068 1774
rect 8068 1767 8070 1774
rect 8100 1767 8102 1774
rect 8102 1767 8140 1774
rect 8140 1767 8152 1774
rect 8018 1722 8070 1767
rect 8100 1722 8152 1767
rect 8182 1722 8234 1774
rect 7936 1658 7988 1710
rect 8018 1705 8070 1710
rect 8100 1705 8152 1710
rect 8018 1671 8030 1705
rect 8030 1671 8068 1705
rect 8068 1671 8070 1705
rect 8100 1671 8102 1705
rect 8102 1671 8140 1705
rect 8140 1671 8152 1705
rect 8018 1658 8070 1671
rect 8100 1658 8152 1671
rect 8182 1658 8234 1710
rect 7936 1594 7988 1646
rect 8018 1609 8070 1646
rect 8100 1609 8152 1646
rect 8018 1594 8030 1609
rect 8030 1594 8068 1609
rect 8068 1594 8070 1609
rect 8100 1594 8102 1609
rect 8102 1594 8140 1609
rect 8140 1594 8152 1609
rect 8182 1594 8234 1646
rect 7936 1530 7988 1582
rect 8018 1575 8030 1582
rect 8030 1575 8068 1582
rect 8068 1575 8070 1582
rect 8100 1575 8102 1582
rect 8102 1575 8140 1582
rect 8140 1575 8152 1582
rect 8018 1530 8070 1575
rect 8100 1530 8152 1575
rect 8182 1530 8234 1582
rect 7936 1466 7988 1518
rect 8018 1513 8070 1518
rect 8100 1513 8152 1518
rect 8018 1479 8030 1513
rect 8030 1479 8068 1513
rect 8068 1479 8070 1513
rect 8100 1479 8102 1513
rect 8102 1479 8140 1513
rect 8140 1479 8152 1513
rect 8018 1466 8070 1479
rect 8100 1466 8152 1479
rect 8182 1466 8234 1518
rect 7936 1402 7988 1454
rect 8018 1417 8070 1454
rect 8100 1417 8152 1454
rect 8018 1402 8030 1417
rect 8030 1402 8068 1417
rect 8068 1402 8070 1417
rect 8100 1402 8102 1417
rect 8102 1402 8140 1417
rect 8140 1402 8152 1417
rect 8182 1402 8234 1454
rect 7936 1338 7988 1390
rect 8018 1383 8030 1390
rect 8030 1383 8068 1390
rect 8068 1383 8070 1390
rect 8100 1383 8102 1390
rect 8102 1383 8140 1390
rect 8140 1383 8152 1390
rect 8018 1338 8070 1383
rect 8100 1338 8152 1383
rect 8182 1338 8234 1390
rect 7936 1274 7988 1326
rect 8018 1321 8070 1326
rect 8100 1321 8152 1326
rect 8018 1287 8030 1321
rect 8030 1287 8068 1321
rect 8068 1287 8070 1321
rect 8100 1287 8102 1321
rect 8102 1287 8140 1321
rect 8140 1287 8152 1321
rect 8018 1274 8070 1287
rect 8100 1274 8152 1287
rect 8182 1274 8234 1326
rect 7936 1210 7988 1262
rect 8018 1225 8070 1262
rect 8100 1225 8152 1262
rect 8018 1210 8030 1225
rect 8030 1210 8068 1225
rect 8068 1210 8070 1225
rect 8100 1210 8102 1225
rect 8102 1210 8140 1225
rect 8140 1210 8152 1225
rect 8182 1210 8234 1262
rect 7936 1146 7988 1198
rect 8018 1191 8030 1198
rect 8030 1191 8068 1198
rect 8068 1191 8070 1198
rect 8100 1191 8102 1198
rect 8102 1191 8140 1198
rect 8140 1191 8152 1198
rect 8018 1146 8070 1191
rect 8100 1146 8152 1191
rect 8182 1146 8234 1198
rect 7936 1082 7988 1134
rect 8018 1129 8070 1134
rect 8100 1129 8152 1134
rect 8018 1095 8030 1129
rect 8030 1095 8068 1129
rect 8068 1095 8070 1129
rect 8100 1095 8102 1129
rect 8102 1095 8140 1129
rect 8140 1095 8152 1129
rect 8018 1082 8070 1095
rect 8100 1082 8152 1095
rect 8182 1082 8234 1134
rect 7936 1018 7988 1070
rect 8018 1033 8070 1070
rect 8100 1033 8152 1070
rect 8018 1018 8030 1033
rect 8030 1018 8068 1033
rect 8068 1018 8070 1033
rect 8100 1018 8102 1033
rect 8102 1018 8140 1033
rect 8140 1018 8152 1033
rect 8182 1018 8234 1070
rect 7936 954 7988 1006
rect 8018 999 8030 1006
rect 8030 999 8068 1006
rect 8068 999 8070 1006
rect 8100 999 8102 1006
rect 8102 999 8140 1006
rect 8140 999 8152 1006
rect 8018 954 8070 999
rect 8100 954 8152 999
rect 8182 954 8234 1006
rect 7936 890 7988 942
rect 8018 937 8070 942
rect 8100 937 8152 942
rect 8018 903 8030 937
rect 8030 903 8068 937
rect 8068 903 8070 937
rect 8100 903 8102 937
rect 8102 903 8140 937
rect 8140 903 8152 937
rect 8018 890 8070 903
rect 8100 890 8152 903
rect 8182 890 8234 942
rect 7936 826 7988 878
rect 8018 841 8070 878
rect 8100 841 8152 878
rect 8018 826 8030 841
rect 8030 826 8068 841
rect 8068 826 8070 841
rect 8100 826 8102 841
rect 8102 826 8140 841
rect 8140 826 8152 841
rect 8182 826 8234 878
rect 7936 762 7988 814
rect 8018 807 8030 814
rect 8030 807 8068 814
rect 8068 807 8070 814
rect 8100 807 8102 814
rect 8102 807 8140 814
rect 8140 807 8152 814
rect 8018 762 8070 807
rect 8100 762 8152 807
rect 8182 762 8234 814
rect 7936 698 7988 750
rect 8018 745 8070 750
rect 8100 745 8152 750
rect 8018 711 8030 745
rect 8030 711 8068 745
rect 8068 711 8070 745
rect 8100 711 8102 745
rect 8102 711 8140 745
rect 8140 711 8152 745
rect 8018 698 8070 711
rect 8100 698 8152 711
rect 8182 698 8234 750
rect 7936 633 7988 685
rect 8018 649 8070 685
rect 8100 649 8152 685
rect 8018 633 8030 649
rect 8030 633 8068 649
rect 8068 633 8070 649
rect 8100 633 8102 649
rect 8102 633 8140 649
rect 8140 633 8152 649
rect 8182 633 8234 685
rect 7936 568 7988 620
rect 8018 615 8030 620
rect 8030 615 8068 620
rect 8068 615 8070 620
rect 8100 615 8102 620
rect 8102 615 8140 620
rect 8140 615 8152 620
rect 8018 568 8070 615
rect 8100 568 8152 615
rect 8182 568 8234 620
rect 7936 503 7988 555
rect 8018 503 8070 555
rect 8100 503 8152 555
rect 8182 503 8234 555
rect 8348 3358 8400 3410
rect 8430 3358 8482 3410
rect 8512 3358 8564 3410
rect 8594 3358 8646 3410
rect 8348 3292 8400 3344
rect 8430 3337 8482 3344
rect 8512 3337 8564 3344
rect 8430 3303 8442 3337
rect 8442 3303 8480 3337
rect 8480 3303 8482 3337
rect 8512 3303 8514 3337
rect 8514 3303 8552 3337
rect 8552 3303 8564 3337
rect 8430 3292 8482 3303
rect 8512 3292 8564 3303
rect 8594 3292 8646 3344
rect 8348 3226 8400 3278
rect 8430 3241 8482 3278
rect 8512 3241 8564 3278
rect 8430 3226 8442 3241
rect 8442 3226 8480 3241
rect 8480 3226 8482 3241
rect 8512 3226 8514 3241
rect 8514 3226 8552 3241
rect 8552 3226 8564 3241
rect 8594 3226 8646 3278
rect 8348 3160 8400 3212
rect 8430 3207 8442 3212
rect 8442 3207 8480 3212
rect 8480 3207 8482 3212
rect 8512 3207 8514 3212
rect 8514 3207 8552 3212
rect 8552 3207 8564 3212
rect 8430 3160 8482 3207
rect 8512 3160 8564 3207
rect 8594 3160 8646 3212
rect 8348 3094 8400 3146
rect 8430 3145 8482 3146
rect 8512 3145 8564 3146
rect 8430 3111 8442 3145
rect 8442 3111 8480 3145
rect 8480 3111 8482 3145
rect 8512 3111 8514 3145
rect 8514 3111 8552 3145
rect 8552 3111 8564 3145
rect 8430 3094 8482 3111
rect 8512 3094 8564 3111
rect 8594 3094 8646 3146
rect 8348 3027 8400 3079
rect 8430 3049 8482 3079
rect 8512 3049 8564 3079
rect 8430 3027 8442 3049
rect 8442 3027 8480 3049
rect 8480 3027 8482 3049
rect 8512 3027 8514 3049
rect 8514 3027 8552 3049
rect 8552 3027 8564 3049
rect 8594 3027 8646 3079
rect 8348 2960 8400 3012
rect 8430 2960 8482 3012
rect 8512 2960 8564 3012
rect 8594 2960 8646 3012
rect 8348 2893 8400 2945
rect 8430 2919 8442 2945
rect 8442 2919 8480 2945
rect 8480 2919 8482 2945
rect 8512 2919 8514 2945
rect 8514 2919 8552 2945
rect 8552 2919 8564 2945
rect 8430 2893 8482 2919
rect 8512 2893 8564 2919
rect 8594 2893 8646 2945
rect 8348 2826 8400 2878
rect 8430 2857 8482 2878
rect 8512 2857 8564 2878
rect 8430 2826 8442 2857
rect 8442 2826 8480 2857
rect 8480 2826 8482 2857
rect 8512 2826 8514 2857
rect 8514 2826 8552 2857
rect 8552 2826 8564 2857
rect 8594 2826 8646 2878
rect 8348 2759 8400 2811
rect 8430 2761 8482 2811
rect 8512 2761 8564 2811
rect 8430 2759 8442 2761
rect 8442 2759 8480 2761
rect 8480 2759 8482 2761
rect 8512 2759 8514 2761
rect 8514 2759 8552 2761
rect 8552 2759 8564 2761
rect 8594 2759 8646 2811
rect 8348 2692 8400 2744
rect 8430 2727 8442 2744
rect 8442 2727 8480 2744
rect 8480 2727 8482 2744
rect 8512 2727 8514 2744
rect 8514 2727 8552 2744
rect 8552 2727 8564 2744
rect 8430 2692 8482 2727
rect 8512 2692 8564 2727
rect 8594 2692 8646 2744
rect 8348 2625 8400 2677
rect 8430 2665 8482 2677
rect 8512 2665 8564 2677
rect 8430 2631 8442 2665
rect 8442 2631 8480 2665
rect 8480 2631 8482 2665
rect 8512 2631 8514 2665
rect 8514 2631 8552 2665
rect 8552 2631 8564 2665
rect 8430 2625 8482 2631
rect 8512 2625 8564 2631
rect 8594 2625 8646 2677
rect 8348 2558 8400 2610
rect 8430 2569 8482 2610
rect 8512 2569 8564 2610
rect 8430 2558 8442 2569
rect 8442 2558 8480 2569
rect 8480 2558 8482 2569
rect 8512 2558 8514 2569
rect 8514 2558 8552 2569
rect 8552 2558 8564 2569
rect 8594 2558 8646 2610
rect 8348 2491 8400 2543
rect 8430 2535 8442 2543
rect 8442 2535 8480 2543
rect 8480 2535 8482 2543
rect 8512 2535 8514 2543
rect 8514 2535 8552 2543
rect 8552 2535 8564 2543
rect 8430 2491 8482 2535
rect 8512 2491 8564 2535
rect 8594 2491 8646 2543
rect 8348 2424 8400 2476
rect 8430 2473 8482 2476
rect 8512 2473 8564 2476
rect 8430 2439 8442 2473
rect 8442 2439 8480 2473
rect 8480 2439 8482 2473
rect 8512 2439 8514 2473
rect 8514 2439 8552 2473
rect 8552 2439 8564 2473
rect 8430 2424 8482 2439
rect 8512 2424 8564 2439
rect 8594 2424 8646 2476
rect 8348 2357 8400 2409
rect 8430 2377 8482 2409
rect 8512 2377 8564 2409
rect 8430 2357 8442 2377
rect 8442 2357 8480 2377
rect 8480 2357 8482 2377
rect 8512 2357 8514 2377
rect 8514 2357 8552 2377
rect 8552 2357 8564 2377
rect 8594 2357 8646 2409
rect 8348 2290 8400 2342
rect 8430 2290 8482 2342
rect 8512 2290 8564 2342
rect 8594 2290 8646 2342
rect 8348 2223 8400 2275
rect 8430 2247 8442 2275
rect 8442 2247 8480 2275
rect 8480 2247 8482 2275
rect 8512 2247 8514 2275
rect 8514 2247 8552 2275
rect 8552 2247 8564 2275
rect 8430 2223 8482 2247
rect 8512 2223 8564 2247
rect 8594 2223 8646 2275
rect 8348 2156 8400 2208
rect 8430 2185 8482 2208
rect 8512 2185 8564 2208
rect 8430 2156 8442 2185
rect 8442 2156 8480 2185
rect 8480 2156 8482 2185
rect 8512 2156 8514 2185
rect 8514 2156 8552 2185
rect 8552 2156 8564 2185
rect 8594 2156 8646 2208
rect 8348 2089 8400 2141
rect 8430 2089 8482 2141
rect 8512 2089 8564 2141
rect 8594 2089 8646 2141
rect 8348 2022 8400 2074
rect 8430 2055 8442 2074
rect 8442 2055 8480 2074
rect 8480 2055 8482 2074
rect 8512 2055 8514 2074
rect 8514 2055 8552 2074
rect 8552 2055 8564 2074
rect 8430 2022 8482 2055
rect 8512 2022 8564 2055
rect 8594 2022 8646 2074
rect 7936 438 7988 490
rect 8018 438 8070 490
rect 8100 438 8152 490
rect 8182 438 8234 490
rect 7936 373 7988 425
rect 8018 373 8070 425
rect 8100 373 8152 425
rect 8182 373 8234 425
rect 8760 1850 8812 1902
rect 8842 1897 8894 1902
rect 8924 1897 8976 1902
rect 8842 1863 8854 1897
rect 8854 1863 8892 1897
rect 8892 1863 8894 1897
rect 8924 1863 8926 1897
rect 8926 1863 8964 1897
rect 8964 1863 8976 1897
rect 8842 1850 8894 1863
rect 8924 1850 8976 1863
rect 9006 1850 9058 1902
rect 8760 1786 8812 1838
rect 8842 1801 8894 1838
rect 8924 1801 8976 1838
rect 8842 1786 8854 1801
rect 8854 1786 8892 1801
rect 8892 1786 8894 1801
rect 8924 1786 8926 1801
rect 8926 1786 8964 1801
rect 8964 1786 8976 1801
rect 9006 1786 9058 1838
rect 8760 1722 8812 1774
rect 8842 1767 8854 1774
rect 8854 1767 8892 1774
rect 8892 1767 8894 1774
rect 8924 1767 8926 1774
rect 8926 1767 8964 1774
rect 8964 1767 8976 1774
rect 8842 1722 8894 1767
rect 8924 1722 8976 1767
rect 9006 1722 9058 1774
rect 8760 1658 8812 1710
rect 8842 1705 8894 1710
rect 8924 1705 8976 1710
rect 8842 1671 8854 1705
rect 8854 1671 8892 1705
rect 8892 1671 8894 1705
rect 8924 1671 8926 1705
rect 8926 1671 8964 1705
rect 8964 1671 8976 1705
rect 8842 1658 8894 1671
rect 8924 1658 8976 1671
rect 9006 1658 9058 1710
rect 8760 1594 8812 1646
rect 8842 1609 8894 1646
rect 8924 1609 8976 1646
rect 8842 1594 8854 1609
rect 8854 1594 8892 1609
rect 8892 1594 8894 1609
rect 8924 1594 8926 1609
rect 8926 1594 8964 1609
rect 8964 1594 8976 1609
rect 9006 1594 9058 1646
rect 8760 1530 8812 1582
rect 8842 1575 8854 1582
rect 8854 1575 8892 1582
rect 8892 1575 8894 1582
rect 8924 1575 8926 1582
rect 8926 1575 8964 1582
rect 8964 1575 8976 1582
rect 8842 1530 8894 1575
rect 8924 1530 8976 1575
rect 9006 1530 9058 1582
rect 8760 1466 8812 1518
rect 8842 1513 8894 1518
rect 8924 1513 8976 1518
rect 8842 1479 8854 1513
rect 8854 1479 8892 1513
rect 8892 1479 8894 1513
rect 8924 1479 8926 1513
rect 8926 1479 8964 1513
rect 8964 1479 8976 1513
rect 8842 1466 8894 1479
rect 8924 1466 8976 1479
rect 9006 1466 9058 1518
rect 8760 1402 8812 1454
rect 8842 1417 8894 1454
rect 8924 1417 8976 1454
rect 8842 1402 8854 1417
rect 8854 1402 8892 1417
rect 8892 1402 8894 1417
rect 8924 1402 8926 1417
rect 8926 1402 8964 1417
rect 8964 1402 8976 1417
rect 9006 1402 9058 1454
rect 8760 1338 8812 1390
rect 8842 1383 8854 1390
rect 8854 1383 8892 1390
rect 8892 1383 8894 1390
rect 8924 1383 8926 1390
rect 8926 1383 8964 1390
rect 8964 1383 8976 1390
rect 8842 1338 8894 1383
rect 8924 1338 8976 1383
rect 9006 1338 9058 1390
rect 8760 1274 8812 1326
rect 8842 1321 8894 1326
rect 8924 1321 8976 1326
rect 8842 1287 8854 1321
rect 8854 1287 8892 1321
rect 8892 1287 8894 1321
rect 8924 1287 8926 1321
rect 8926 1287 8964 1321
rect 8964 1287 8976 1321
rect 8842 1274 8894 1287
rect 8924 1274 8976 1287
rect 9006 1274 9058 1326
rect 8760 1210 8812 1262
rect 8842 1225 8894 1262
rect 8924 1225 8976 1262
rect 8842 1210 8854 1225
rect 8854 1210 8892 1225
rect 8892 1210 8894 1225
rect 8924 1210 8926 1225
rect 8926 1210 8964 1225
rect 8964 1210 8976 1225
rect 9006 1210 9058 1262
rect 8760 1146 8812 1198
rect 8842 1191 8854 1198
rect 8854 1191 8892 1198
rect 8892 1191 8894 1198
rect 8924 1191 8926 1198
rect 8926 1191 8964 1198
rect 8964 1191 8976 1198
rect 8842 1146 8894 1191
rect 8924 1146 8976 1191
rect 9006 1146 9058 1198
rect 8760 1082 8812 1134
rect 8842 1129 8894 1134
rect 8924 1129 8976 1134
rect 8842 1095 8854 1129
rect 8854 1095 8892 1129
rect 8892 1095 8894 1129
rect 8924 1095 8926 1129
rect 8926 1095 8964 1129
rect 8964 1095 8976 1129
rect 8842 1082 8894 1095
rect 8924 1082 8976 1095
rect 9006 1082 9058 1134
rect 8760 1018 8812 1070
rect 8842 1033 8894 1070
rect 8924 1033 8976 1070
rect 8842 1018 8854 1033
rect 8854 1018 8892 1033
rect 8892 1018 8894 1033
rect 8924 1018 8926 1033
rect 8926 1018 8964 1033
rect 8964 1018 8976 1033
rect 9006 1018 9058 1070
rect 8760 954 8812 1006
rect 8842 999 8854 1006
rect 8854 999 8892 1006
rect 8892 999 8894 1006
rect 8924 999 8926 1006
rect 8926 999 8964 1006
rect 8964 999 8976 1006
rect 8842 954 8894 999
rect 8924 954 8976 999
rect 9006 954 9058 1006
rect 8760 890 8812 942
rect 8842 937 8894 942
rect 8924 937 8976 942
rect 8842 903 8854 937
rect 8854 903 8892 937
rect 8892 903 8894 937
rect 8924 903 8926 937
rect 8926 903 8964 937
rect 8964 903 8976 937
rect 8842 890 8894 903
rect 8924 890 8976 903
rect 9006 890 9058 942
rect 8760 826 8812 878
rect 8842 841 8894 878
rect 8924 841 8976 878
rect 8842 826 8854 841
rect 8854 826 8892 841
rect 8892 826 8894 841
rect 8924 826 8926 841
rect 8926 826 8964 841
rect 8964 826 8976 841
rect 9006 826 9058 878
rect 8760 762 8812 814
rect 8842 807 8854 814
rect 8854 807 8892 814
rect 8892 807 8894 814
rect 8924 807 8926 814
rect 8926 807 8964 814
rect 8964 807 8976 814
rect 8842 762 8894 807
rect 8924 762 8976 807
rect 9006 762 9058 814
rect 8760 698 8812 750
rect 8842 745 8894 750
rect 8924 745 8976 750
rect 8842 711 8854 745
rect 8854 711 8892 745
rect 8892 711 8894 745
rect 8924 711 8926 745
rect 8926 711 8964 745
rect 8964 711 8976 745
rect 8842 698 8894 711
rect 8924 698 8976 711
rect 9006 698 9058 750
rect 8760 633 8812 685
rect 8842 649 8894 685
rect 8924 649 8976 685
rect 8842 633 8854 649
rect 8854 633 8892 649
rect 8892 633 8894 649
rect 8924 633 8926 649
rect 8926 633 8964 649
rect 8964 633 8976 649
rect 9006 633 9058 685
rect 8760 568 8812 620
rect 8842 615 8854 620
rect 8854 615 8892 620
rect 8892 615 8894 620
rect 8924 615 8926 620
rect 8926 615 8964 620
rect 8964 615 8976 620
rect 8842 568 8894 615
rect 8924 568 8976 615
rect 9006 568 9058 620
rect 8760 503 8812 555
rect 8842 503 8894 555
rect 8924 503 8976 555
rect 9006 503 9058 555
rect 9172 3358 9224 3410
rect 9254 3358 9306 3410
rect 9336 3358 9388 3410
rect 9418 3358 9470 3410
rect 9172 3292 9224 3344
rect 9254 3337 9306 3344
rect 9336 3337 9388 3344
rect 9254 3303 9266 3337
rect 9266 3303 9304 3337
rect 9304 3303 9306 3337
rect 9336 3303 9338 3337
rect 9338 3303 9376 3337
rect 9376 3303 9388 3337
rect 9254 3292 9306 3303
rect 9336 3292 9388 3303
rect 9418 3292 9470 3344
rect 9172 3226 9224 3278
rect 9254 3241 9306 3278
rect 9336 3241 9388 3278
rect 9254 3226 9266 3241
rect 9266 3226 9304 3241
rect 9304 3226 9306 3241
rect 9336 3226 9338 3241
rect 9338 3226 9376 3241
rect 9376 3226 9388 3241
rect 9418 3226 9470 3278
rect 9172 3160 9224 3212
rect 9254 3207 9266 3212
rect 9266 3207 9304 3212
rect 9304 3207 9306 3212
rect 9336 3207 9338 3212
rect 9338 3207 9376 3212
rect 9376 3207 9388 3212
rect 9254 3160 9306 3207
rect 9336 3160 9388 3207
rect 9418 3160 9470 3212
rect 9172 3094 9224 3146
rect 9254 3145 9306 3146
rect 9336 3145 9388 3146
rect 9254 3111 9266 3145
rect 9266 3111 9304 3145
rect 9304 3111 9306 3145
rect 9336 3111 9338 3145
rect 9338 3111 9376 3145
rect 9376 3111 9388 3145
rect 9254 3094 9306 3111
rect 9336 3094 9388 3111
rect 9418 3094 9470 3146
rect 9172 3027 9224 3079
rect 9254 3049 9306 3079
rect 9336 3049 9388 3079
rect 9254 3027 9266 3049
rect 9266 3027 9304 3049
rect 9304 3027 9306 3049
rect 9336 3027 9338 3049
rect 9338 3027 9376 3049
rect 9376 3027 9388 3049
rect 9418 3027 9470 3079
rect 9172 2960 9224 3012
rect 9254 2960 9306 3012
rect 9336 2960 9388 3012
rect 9418 2960 9470 3012
rect 9172 2893 9224 2945
rect 9254 2919 9266 2945
rect 9266 2919 9304 2945
rect 9304 2919 9306 2945
rect 9336 2919 9338 2945
rect 9338 2919 9376 2945
rect 9376 2919 9388 2945
rect 9254 2893 9306 2919
rect 9336 2893 9388 2919
rect 9418 2893 9470 2945
rect 9172 2826 9224 2878
rect 9254 2857 9306 2878
rect 9336 2857 9388 2878
rect 9254 2826 9266 2857
rect 9266 2826 9304 2857
rect 9304 2826 9306 2857
rect 9336 2826 9338 2857
rect 9338 2826 9376 2857
rect 9376 2826 9388 2857
rect 9418 2826 9470 2878
rect 9172 2759 9224 2811
rect 9254 2761 9306 2811
rect 9336 2761 9388 2811
rect 9254 2759 9266 2761
rect 9266 2759 9304 2761
rect 9304 2759 9306 2761
rect 9336 2759 9338 2761
rect 9338 2759 9376 2761
rect 9376 2759 9388 2761
rect 9418 2759 9470 2811
rect 9172 2692 9224 2744
rect 9254 2727 9266 2744
rect 9266 2727 9304 2744
rect 9304 2727 9306 2744
rect 9336 2727 9338 2744
rect 9338 2727 9376 2744
rect 9376 2727 9388 2744
rect 9254 2692 9306 2727
rect 9336 2692 9388 2727
rect 9418 2692 9470 2744
rect 9172 2625 9224 2677
rect 9254 2665 9306 2677
rect 9336 2665 9388 2677
rect 9254 2631 9266 2665
rect 9266 2631 9304 2665
rect 9304 2631 9306 2665
rect 9336 2631 9338 2665
rect 9338 2631 9376 2665
rect 9376 2631 9388 2665
rect 9254 2625 9306 2631
rect 9336 2625 9388 2631
rect 9418 2625 9470 2677
rect 9172 2558 9224 2610
rect 9254 2569 9306 2610
rect 9336 2569 9388 2610
rect 9254 2558 9266 2569
rect 9266 2558 9304 2569
rect 9304 2558 9306 2569
rect 9336 2558 9338 2569
rect 9338 2558 9376 2569
rect 9376 2558 9388 2569
rect 9418 2558 9470 2610
rect 9172 2491 9224 2543
rect 9254 2535 9266 2543
rect 9266 2535 9304 2543
rect 9304 2535 9306 2543
rect 9336 2535 9338 2543
rect 9338 2535 9376 2543
rect 9376 2535 9388 2543
rect 9254 2491 9306 2535
rect 9336 2491 9388 2535
rect 9418 2491 9470 2543
rect 9172 2424 9224 2476
rect 9254 2473 9306 2476
rect 9336 2473 9388 2476
rect 9254 2439 9266 2473
rect 9266 2439 9304 2473
rect 9304 2439 9306 2473
rect 9336 2439 9338 2473
rect 9338 2439 9376 2473
rect 9376 2439 9388 2473
rect 9254 2424 9306 2439
rect 9336 2424 9388 2439
rect 9418 2424 9470 2476
rect 9172 2357 9224 2409
rect 9254 2377 9306 2409
rect 9336 2377 9388 2409
rect 9254 2357 9266 2377
rect 9266 2357 9304 2377
rect 9304 2357 9306 2377
rect 9336 2357 9338 2377
rect 9338 2357 9376 2377
rect 9376 2357 9388 2377
rect 9418 2357 9470 2409
rect 9172 2290 9224 2342
rect 9254 2290 9306 2342
rect 9336 2290 9388 2342
rect 9418 2290 9470 2342
rect 9172 2223 9224 2275
rect 9254 2247 9266 2275
rect 9266 2247 9304 2275
rect 9304 2247 9306 2275
rect 9336 2247 9338 2275
rect 9338 2247 9376 2275
rect 9376 2247 9388 2275
rect 9254 2223 9306 2247
rect 9336 2223 9388 2247
rect 9418 2223 9470 2275
rect 9172 2156 9224 2208
rect 9254 2185 9306 2208
rect 9336 2185 9388 2208
rect 9254 2156 9266 2185
rect 9266 2156 9304 2185
rect 9304 2156 9306 2185
rect 9336 2156 9338 2185
rect 9338 2156 9376 2185
rect 9376 2156 9388 2185
rect 9418 2156 9470 2208
rect 9172 2089 9224 2141
rect 9254 2089 9306 2141
rect 9336 2089 9388 2141
rect 9418 2089 9470 2141
rect 9172 2022 9224 2074
rect 9254 2055 9266 2074
rect 9266 2055 9304 2074
rect 9304 2055 9306 2074
rect 9336 2055 9338 2074
rect 9338 2055 9376 2074
rect 9376 2055 9388 2074
rect 9254 2022 9306 2055
rect 9336 2022 9388 2055
rect 9418 2022 9470 2074
rect 8760 438 8812 490
rect 8842 438 8894 490
rect 8924 438 8976 490
rect 9006 438 9058 490
rect 8760 373 8812 425
rect 8842 373 8894 425
rect 8924 373 8976 425
rect 9006 373 9058 425
rect 9584 1850 9636 1902
rect 9666 1897 9718 1902
rect 9748 1897 9800 1902
rect 9666 1863 9678 1897
rect 9678 1863 9716 1897
rect 9716 1863 9718 1897
rect 9748 1863 9750 1897
rect 9750 1863 9788 1897
rect 9788 1863 9800 1897
rect 9666 1850 9718 1863
rect 9748 1850 9800 1863
rect 9830 1850 9882 1902
rect 9584 1786 9636 1838
rect 9666 1801 9718 1838
rect 9748 1801 9800 1838
rect 9666 1786 9678 1801
rect 9678 1786 9716 1801
rect 9716 1786 9718 1801
rect 9748 1786 9750 1801
rect 9750 1786 9788 1801
rect 9788 1786 9800 1801
rect 9830 1786 9882 1838
rect 9584 1722 9636 1774
rect 9666 1767 9678 1774
rect 9678 1767 9716 1774
rect 9716 1767 9718 1774
rect 9748 1767 9750 1774
rect 9750 1767 9788 1774
rect 9788 1767 9800 1774
rect 9666 1722 9718 1767
rect 9748 1722 9800 1767
rect 9830 1722 9882 1774
rect 9584 1658 9636 1710
rect 9666 1705 9718 1710
rect 9748 1705 9800 1710
rect 9666 1671 9678 1705
rect 9678 1671 9716 1705
rect 9716 1671 9718 1705
rect 9748 1671 9750 1705
rect 9750 1671 9788 1705
rect 9788 1671 9800 1705
rect 9666 1658 9718 1671
rect 9748 1658 9800 1671
rect 9830 1658 9882 1710
rect 9584 1594 9636 1646
rect 9666 1609 9718 1646
rect 9748 1609 9800 1646
rect 9666 1594 9678 1609
rect 9678 1594 9716 1609
rect 9716 1594 9718 1609
rect 9748 1594 9750 1609
rect 9750 1594 9788 1609
rect 9788 1594 9800 1609
rect 9830 1594 9882 1646
rect 9584 1530 9636 1582
rect 9666 1575 9678 1582
rect 9678 1575 9716 1582
rect 9716 1575 9718 1582
rect 9748 1575 9750 1582
rect 9750 1575 9788 1582
rect 9788 1575 9800 1582
rect 9666 1530 9718 1575
rect 9748 1530 9800 1575
rect 9830 1530 9882 1582
rect 9584 1466 9636 1518
rect 9666 1513 9718 1518
rect 9748 1513 9800 1518
rect 9666 1479 9678 1513
rect 9678 1479 9716 1513
rect 9716 1479 9718 1513
rect 9748 1479 9750 1513
rect 9750 1479 9788 1513
rect 9788 1479 9800 1513
rect 9666 1466 9718 1479
rect 9748 1466 9800 1479
rect 9830 1466 9882 1518
rect 9584 1402 9636 1454
rect 9666 1417 9718 1454
rect 9748 1417 9800 1454
rect 9666 1402 9678 1417
rect 9678 1402 9716 1417
rect 9716 1402 9718 1417
rect 9748 1402 9750 1417
rect 9750 1402 9788 1417
rect 9788 1402 9800 1417
rect 9830 1402 9882 1454
rect 9584 1338 9636 1390
rect 9666 1383 9678 1390
rect 9678 1383 9716 1390
rect 9716 1383 9718 1390
rect 9748 1383 9750 1390
rect 9750 1383 9788 1390
rect 9788 1383 9800 1390
rect 9666 1338 9718 1383
rect 9748 1338 9800 1383
rect 9830 1338 9882 1390
rect 9584 1274 9636 1326
rect 9666 1321 9718 1326
rect 9748 1321 9800 1326
rect 9666 1287 9678 1321
rect 9678 1287 9716 1321
rect 9716 1287 9718 1321
rect 9748 1287 9750 1321
rect 9750 1287 9788 1321
rect 9788 1287 9800 1321
rect 9666 1274 9718 1287
rect 9748 1274 9800 1287
rect 9830 1274 9882 1326
rect 9584 1210 9636 1262
rect 9666 1225 9718 1262
rect 9748 1225 9800 1262
rect 9666 1210 9678 1225
rect 9678 1210 9716 1225
rect 9716 1210 9718 1225
rect 9748 1210 9750 1225
rect 9750 1210 9788 1225
rect 9788 1210 9800 1225
rect 9830 1210 9882 1262
rect 9584 1146 9636 1198
rect 9666 1191 9678 1198
rect 9678 1191 9716 1198
rect 9716 1191 9718 1198
rect 9748 1191 9750 1198
rect 9750 1191 9788 1198
rect 9788 1191 9800 1198
rect 9666 1146 9718 1191
rect 9748 1146 9800 1191
rect 9830 1146 9882 1198
rect 9584 1082 9636 1134
rect 9666 1129 9718 1134
rect 9748 1129 9800 1134
rect 9666 1095 9678 1129
rect 9678 1095 9716 1129
rect 9716 1095 9718 1129
rect 9748 1095 9750 1129
rect 9750 1095 9788 1129
rect 9788 1095 9800 1129
rect 9666 1082 9718 1095
rect 9748 1082 9800 1095
rect 9830 1082 9882 1134
rect 9584 1018 9636 1070
rect 9666 1033 9718 1070
rect 9748 1033 9800 1070
rect 9666 1018 9678 1033
rect 9678 1018 9716 1033
rect 9716 1018 9718 1033
rect 9748 1018 9750 1033
rect 9750 1018 9788 1033
rect 9788 1018 9800 1033
rect 9830 1018 9882 1070
rect 9584 954 9636 1006
rect 9666 999 9678 1006
rect 9678 999 9716 1006
rect 9716 999 9718 1006
rect 9748 999 9750 1006
rect 9750 999 9788 1006
rect 9788 999 9800 1006
rect 9666 954 9718 999
rect 9748 954 9800 999
rect 9830 954 9882 1006
rect 9584 890 9636 942
rect 9666 937 9718 942
rect 9748 937 9800 942
rect 9666 903 9678 937
rect 9678 903 9716 937
rect 9716 903 9718 937
rect 9748 903 9750 937
rect 9750 903 9788 937
rect 9788 903 9800 937
rect 9666 890 9718 903
rect 9748 890 9800 903
rect 9830 890 9882 942
rect 9584 826 9636 878
rect 9666 841 9718 878
rect 9748 841 9800 878
rect 9666 826 9678 841
rect 9678 826 9716 841
rect 9716 826 9718 841
rect 9748 826 9750 841
rect 9750 826 9788 841
rect 9788 826 9800 841
rect 9830 826 9882 878
rect 9584 762 9636 814
rect 9666 807 9678 814
rect 9678 807 9716 814
rect 9716 807 9718 814
rect 9748 807 9750 814
rect 9750 807 9788 814
rect 9788 807 9800 814
rect 9666 762 9718 807
rect 9748 762 9800 807
rect 9830 762 9882 814
rect 9584 698 9636 750
rect 9666 745 9718 750
rect 9748 745 9800 750
rect 9666 711 9678 745
rect 9678 711 9716 745
rect 9716 711 9718 745
rect 9748 711 9750 745
rect 9750 711 9788 745
rect 9788 711 9800 745
rect 9666 698 9718 711
rect 9748 698 9800 711
rect 9830 698 9882 750
rect 9584 633 9636 685
rect 9666 649 9718 685
rect 9748 649 9800 685
rect 9666 633 9678 649
rect 9678 633 9716 649
rect 9716 633 9718 649
rect 9748 633 9750 649
rect 9750 633 9788 649
rect 9788 633 9800 649
rect 9830 633 9882 685
rect 9584 568 9636 620
rect 9666 615 9678 620
rect 9678 615 9716 620
rect 9716 615 9718 620
rect 9748 615 9750 620
rect 9750 615 9788 620
rect 9788 615 9800 620
rect 9666 568 9718 615
rect 9748 568 9800 615
rect 9830 568 9882 620
rect 9584 503 9636 555
rect 9666 503 9718 555
rect 9748 503 9800 555
rect 9830 503 9882 555
rect 9996 3358 10048 3410
rect 10078 3358 10130 3410
rect 10160 3358 10212 3410
rect 10242 3358 10294 3410
rect 9996 3292 10048 3344
rect 10078 3337 10130 3344
rect 10160 3337 10212 3344
rect 10078 3303 10090 3337
rect 10090 3303 10128 3337
rect 10128 3303 10130 3337
rect 10160 3303 10162 3337
rect 10162 3303 10200 3337
rect 10200 3303 10212 3337
rect 10078 3292 10130 3303
rect 10160 3292 10212 3303
rect 10242 3292 10294 3344
rect 9996 3226 10048 3278
rect 10078 3241 10130 3278
rect 10160 3241 10212 3278
rect 10078 3226 10090 3241
rect 10090 3226 10128 3241
rect 10128 3226 10130 3241
rect 10160 3226 10162 3241
rect 10162 3226 10200 3241
rect 10200 3226 10212 3241
rect 10242 3226 10294 3278
rect 9996 3160 10048 3212
rect 10078 3207 10090 3212
rect 10090 3207 10128 3212
rect 10128 3207 10130 3212
rect 10160 3207 10162 3212
rect 10162 3207 10200 3212
rect 10200 3207 10212 3212
rect 10078 3160 10130 3207
rect 10160 3160 10212 3207
rect 10242 3160 10294 3212
rect 9996 3094 10048 3146
rect 10078 3145 10130 3146
rect 10160 3145 10212 3146
rect 10078 3111 10090 3145
rect 10090 3111 10128 3145
rect 10128 3111 10130 3145
rect 10160 3111 10162 3145
rect 10162 3111 10200 3145
rect 10200 3111 10212 3145
rect 10078 3094 10130 3111
rect 10160 3094 10212 3111
rect 10242 3094 10294 3146
rect 9996 3027 10048 3079
rect 10078 3049 10130 3079
rect 10160 3049 10212 3079
rect 10078 3027 10090 3049
rect 10090 3027 10128 3049
rect 10128 3027 10130 3049
rect 10160 3027 10162 3049
rect 10162 3027 10200 3049
rect 10200 3027 10212 3049
rect 10242 3027 10294 3079
rect 9996 2960 10048 3012
rect 10078 2960 10130 3012
rect 10160 2960 10212 3012
rect 10242 2960 10294 3012
rect 9996 2893 10048 2945
rect 10078 2919 10090 2945
rect 10090 2919 10128 2945
rect 10128 2919 10130 2945
rect 10160 2919 10162 2945
rect 10162 2919 10200 2945
rect 10200 2919 10212 2945
rect 10078 2893 10130 2919
rect 10160 2893 10212 2919
rect 10242 2893 10294 2945
rect 9996 2826 10048 2878
rect 10078 2857 10130 2878
rect 10160 2857 10212 2878
rect 10078 2826 10090 2857
rect 10090 2826 10128 2857
rect 10128 2826 10130 2857
rect 10160 2826 10162 2857
rect 10162 2826 10200 2857
rect 10200 2826 10212 2857
rect 10242 2826 10294 2878
rect 9996 2759 10048 2811
rect 10078 2761 10130 2811
rect 10160 2761 10212 2811
rect 10078 2759 10090 2761
rect 10090 2759 10128 2761
rect 10128 2759 10130 2761
rect 10160 2759 10162 2761
rect 10162 2759 10200 2761
rect 10200 2759 10212 2761
rect 10242 2759 10294 2811
rect 9996 2692 10048 2744
rect 10078 2727 10090 2744
rect 10090 2727 10128 2744
rect 10128 2727 10130 2744
rect 10160 2727 10162 2744
rect 10162 2727 10200 2744
rect 10200 2727 10212 2744
rect 10078 2692 10130 2727
rect 10160 2692 10212 2727
rect 10242 2692 10294 2744
rect 9996 2625 10048 2677
rect 10078 2665 10130 2677
rect 10160 2665 10212 2677
rect 10078 2631 10090 2665
rect 10090 2631 10128 2665
rect 10128 2631 10130 2665
rect 10160 2631 10162 2665
rect 10162 2631 10200 2665
rect 10200 2631 10212 2665
rect 10078 2625 10130 2631
rect 10160 2625 10212 2631
rect 10242 2625 10294 2677
rect 9996 2558 10048 2610
rect 10078 2569 10130 2610
rect 10160 2569 10212 2610
rect 10078 2558 10090 2569
rect 10090 2558 10128 2569
rect 10128 2558 10130 2569
rect 10160 2558 10162 2569
rect 10162 2558 10200 2569
rect 10200 2558 10212 2569
rect 10242 2558 10294 2610
rect 9996 2491 10048 2543
rect 10078 2535 10090 2543
rect 10090 2535 10128 2543
rect 10128 2535 10130 2543
rect 10160 2535 10162 2543
rect 10162 2535 10200 2543
rect 10200 2535 10212 2543
rect 10078 2491 10130 2535
rect 10160 2491 10212 2535
rect 10242 2491 10294 2543
rect 9996 2424 10048 2476
rect 10078 2473 10130 2476
rect 10160 2473 10212 2476
rect 10078 2439 10090 2473
rect 10090 2439 10128 2473
rect 10128 2439 10130 2473
rect 10160 2439 10162 2473
rect 10162 2439 10200 2473
rect 10200 2439 10212 2473
rect 10078 2424 10130 2439
rect 10160 2424 10212 2439
rect 10242 2424 10294 2476
rect 9996 2357 10048 2409
rect 10078 2377 10130 2409
rect 10160 2377 10212 2409
rect 10078 2357 10090 2377
rect 10090 2357 10128 2377
rect 10128 2357 10130 2377
rect 10160 2357 10162 2377
rect 10162 2357 10200 2377
rect 10200 2357 10212 2377
rect 10242 2357 10294 2409
rect 9996 2290 10048 2342
rect 10078 2290 10130 2342
rect 10160 2290 10212 2342
rect 10242 2290 10294 2342
rect 9996 2223 10048 2275
rect 10078 2247 10090 2275
rect 10090 2247 10128 2275
rect 10128 2247 10130 2275
rect 10160 2247 10162 2275
rect 10162 2247 10200 2275
rect 10200 2247 10212 2275
rect 10078 2223 10130 2247
rect 10160 2223 10212 2247
rect 10242 2223 10294 2275
rect 9996 2156 10048 2208
rect 10078 2185 10130 2208
rect 10160 2185 10212 2208
rect 10078 2156 10090 2185
rect 10090 2156 10128 2185
rect 10128 2156 10130 2185
rect 10160 2156 10162 2185
rect 10162 2156 10200 2185
rect 10200 2156 10212 2185
rect 10242 2156 10294 2208
rect 9996 2089 10048 2141
rect 10078 2089 10130 2141
rect 10160 2089 10212 2141
rect 10242 2089 10294 2141
rect 9996 2022 10048 2074
rect 10078 2055 10090 2074
rect 10090 2055 10128 2074
rect 10128 2055 10130 2074
rect 10160 2055 10162 2074
rect 10162 2055 10200 2074
rect 10200 2055 10212 2074
rect 10078 2022 10130 2055
rect 10160 2022 10212 2055
rect 10242 2022 10294 2074
rect 9584 438 9636 490
rect 9666 438 9718 490
rect 9748 438 9800 490
rect 9830 438 9882 490
rect 9584 373 9636 425
rect 9666 373 9718 425
rect 9748 373 9800 425
rect 9830 373 9882 425
rect 10408 1850 10460 1902
rect 10490 1897 10542 1902
rect 10572 1897 10624 1902
rect 10490 1863 10502 1897
rect 10502 1863 10540 1897
rect 10540 1863 10542 1897
rect 10572 1863 10574 1897
rect 10574 1863 10612 1897
rect 10612 1863 10624 1897
rect 10490 1850 10542 1863
rect 10572 1850 10624 1863
rect 10654 1850 10706 1902
rect 10408 1786 10460 1838
rect 10490 1801 10542 1838
rect 10572 1801 10624 1838
rect 10490 1786 10502 1801
rect 10502 1786 10540 1801
rect 10540 1786 10542 1801
rect 10572 1786 10574 1801
rect 10574 1786 10612 1801
rect 10612 1786 10624 1801
rect 10654 1786 10706 1838
rect 10408 1722 10460 1774
rect 10490 1767 10502 1774
rect 10502 1767 10540 1774
rect 10540 1767 10542 1774
rect 10572 1767 10574 1774
rect 10574 1767 10612 1774
rect 10612 1767 10624 1774
rect 10490 1722 10542 1767
rect 10572 1722 10624 1767
rect 10654 1722 10706 1774
rect 10408 1658 10460 1710
rect 10490 1705 10542 1710
rect 10572 1705 10624 1710
rect 10490 1671 10502 1705
rect 10502 1671 10540 1705
rect 10540 1671 10542 1705
rect 10572 1671 10574 1705
rect 10574 1671 10612 1705
rect 10612 1671 10624 1705
rect 10490 1658 10542 1671
rect 10572 1658 10624 1671
rect 10654 1658 10706 1710
rect 10408 1594 10460 1646
rect 10490 1609 10542 1646
rect 10572 1609 10624 1646
rect 10490 1594 10502 1609
rect 10502 1594 10540 1609
rect 10540 1594 10542 1609
rect 10572 1594 10574 1609
rect 10574 1594 10612 1609
rect 10612 1594 10624 1609
rect 10654 1594 10706 1646
rect 10408 1530 10460 1582
rect 10490 1575 10502 1582
rect 10502 1575 10540 1582
rect 10540 1575 10542 1582
rect 10572 1575 10574 1582
rect 10574 1575 10612 1582
rect 10612 1575 10624 1582
rect 10490 1530 10542 1575
rect 10572 1530 10624 1575
rect 10654 1530 10706 1582
rect 10408 1466 10460 1518
rect 10490 1513 10542 1518
rect 10572 1513 10624 1518
rect 10490 1479 10502 1513
rect 10502 1479 10540 1513
rect 10540 1479 10542 1513
rect 10572 1479 10574 1513
rect 10574 1479 10612 1513
rect 10612 1479 10624 1513
rect 10490 1466 10542 1479
rect 10572 1466 10624 1479
rect 10654 1466 10706 1518
rect 10408 1402 10460 1454
rect 10490 1417 10542 1454
rect 10572 1417 10624 1454
rect 10490 1402 10502 1417
rect 10502 1402 10540 1417
rect 10540 1402 10542 1417
rect 10572 1402 10574 1417
rect 10574 1402 10612 1417
rect 10612 1402 10624 1417
rect 10654 1402 10706 1454
rect 10408 1338 10460 1390
rect 10490 1383 10502 1390
rect 10502 1383 10540 1390
rect 10540 1383 10542 1390
rect 10572 1383 10574 1390
rect 10574 1383 10612 1390
rect 10612 1383 10624 1390
rect 10490 1338 10542 1383
rect 10572 1338 10624 1383
rect 10654 1338 10706 1390
rect 10408 1274 10460 1326
rect 10490 1321 10542 1326
rect 10572 1321 10624 1326
rect 10490 1287 10502 1321
rect 10502 1287 10540 1321
rect 10540 1287 10542 1321
rect 10572 1287 10574 1321
rect 10574 1287 10612 1321
rect 10612 1287 10624 1321
rect 10490 1274 10542 1287
rect 10572 1274 10624 1287
rect 10654 1274 10706 1326
rect 10408 1210 10460 1262
rect 10490 1225 10542 1262
rect 10572 1225 10624 1262
rect 10490 1210 10502 1225
rect 10502 1210 10540 1225
rect 10540 1210 10542 1225
rect 10572 1210 10574 1225
rect 10574 1210 10612 1225
rect 10612 1210 10624 1225
rect 10654 1210 10706 1262
rect 10408 1146 10460 1198
rect 10490 1191 10502 1198
rect 10502 1191 10540 1198
rect 10540 1191 10542 1198
rect 10572 1191 10574 1198
rect 10574 1191 10612 1198
rect 10612 1191 10624 1198
rect 10490 1146 10542 1191
rect 10572 1146 10624 1191
rect 10654 1146 10706 1198
rect 10408 1082 10460 1134
rect 10490 1129 10542 1134
rect 10572 1129 10624 1134
rect 10490 1095 10502 1129
rect 10502 1095 10540 1129
rect 10540 1095 10542 1129
rect 10572 1095 10574 1129
rect 10574 1095 10612 1129
rect 10612 1095 10624 1129
rect 10490 1082 10542 1095
rect 10572 1082 10624 1095
rect 10654 1082 10706 1134
rect 10408 1018 10460 1070
rect 10490 1033 10542 1070
rect 10572 1033 10624 1070
rect 10490 1018 10502 1033
rect 10502 1018 10540 1033
rect 10540 1018 10542 1033
rect 10572 1018 10574 1033
rect 10574 1018 10612 1033
rect 10612 1018 10624 1033
rect 10654 1018 10706 1070
rect 10408 954 10460 1006
rect 10490 999 10502 1006
rect 10502 999 10540 1006
rect 10540 999 10542 1006
rect 10572 999 10574 1006
rect 10574 999 10612 1006
rect 10612 999 10624 1006
rect 10490 954 10542 999
rect 10572 954 10624 999
rect 10654 954 10706 1006
rect 10408 890 10460 942
rect 10490 937 10542 942
rect 10572 937 10624 942
rect 10490 903 10502 937
rect 10502 903 10540 937
rect 10540 903 10542 937
rect 10572 903 10574 937
rect 10574 903 10612 937
rect 10612 903 10624 937
rect 10490 890 10542 903
rect 10572 890 10624 903
rect 10654 890 10706 942
rect 10408 826 10460 878
rect 10490 841 10542 878
rect 10572 841 10624 878
rect 10490 826 10502 841
rect 10502 826 10540 841
rect 10540 826 10542 841
rect 10572 826 10574 841
rect 10574 826 10612 841
rect 10612 826 10624 841
rect 10654 826 10706 878
rect 10408 762 10460 814
rect 10490 807 10502 814
rect 10502 807 10540 814
rect 10540 807 10542 814
rect 10572 807 10574 814
rect 10574 807 10612 814
rect 10612 807 10624 814
rect 10490 762 10542 807
rect 10572 762 10624 807
rect 10654 762 10706 814
rect 10408 698 10460 750
rect 10490 745 10542 750
rect 10572 745 10624 750
rect 10490 711 10502 745
rect 10502 711 10540 745
rect 10540 711 10542 745
rect 10572 711 10574 745
rect 10574 711 10612 745
rect 10612 711 10624 745
rect 10490 698 10542 711
rect 10572 698 10624 711
rect 10654 698 10706 750
rect 10408 633 10460 685
rect 10490 649 10542 685
rect 10572 649 10624 685
rect 10490 633 10502 649
rect 10502 633 10540 649
rect 10540 633 10542 649
rect 10572 633 10574 649
rect 10574 633 10612 649
rect 10612 633 10624 649
rect 10654 633 10706 685
rect 10408 568 10460 620
rect 10490 615 10502 620
rect 10502 615 10540 620
rect 10540 615 10542 620
rect 10572 615 10574 620
rect 10574 615 10612 620
rect 10612 615 10624 620
rect 10490 568 10542 615
rect 10572 568 10624 615
rect 10654 568 10706 620
rect 10408 503 10460 555
rect 10490 503 10542 555
rect 10572 503 10624 555
rect 10654 503 10706 555
rect 10820 3358 10872 3410
rect 10902 3358 10954 3410
rect 10984 3358 11036 3410
rect 11066 3358 11118 3410
rect 10820 3292 10872 3344
rect 10902 3337 10954 3344
rect 10984 3337 11036 3344
rect 10902 3303 10914 3337
rect 10914 3303 10952 3337
rect 10952 3303 10954 3337
rect 10984 3303 10986 3337
rect 10986 3303 11024 3337
rect 11024 3303 11036 3337
rect 10902 3292 10954 3303
rect 10984 3292 11036 3303
rect 11066 3292 11118 3344
rect 10820 3226 10872 3278
rect 10902 3241 10954 3278
rect 10984 3241 11036 3278
rect 10902 3226 10914 3241
rect 10914 3226 10952 3241
rect 10952 3226 10954 3241
rect 10984 3226 10986 3241
rect 10986 3226 11024 3241
rect 11024 3226 11036 3241
rect 11066 3226 11118 3278
rect 10820 3160 10872 3212
rect 10902 3207 10914 3212
rect 10914 3207 10952 3212
rect 10952 3207 10954 3212
rect 10984 3207 10986 3212
rect 10986 3207 11024 3212
rect 11024 3207 11036 3212
rect 10902 3160 10954 3207
rect 10984 3160 11036 3207
rect 11066 3160 11118 3212
rect 10820 3094 10872 3146
rect 10902 3145 10954 3146
rect 10984 3145 11036 3146
rect 10902 3111 10914 3145
rect 10914 3111 10952 3145
rect 10952 3111 10954 3145
rect 10984 3111 10986 3145
rect 10986 3111 11024 3145
rect 11024 3111 11036 3145
rect 10902 3094 10954 3111
rect 10984 3094 11036 3111
rect 11066 3094 11118 3146
rect 10820 3027 10872 3079
rect 10902 3049 10954 3079
rect 10984 3049 11036 3079
rect 10902 3027 10914 3049
rect 10914 3027 10952 3049
rect 10952 3027 10954 3049
rect 10984 3027 10986 3049
rect 10986 3027 11024 3049
rect 11024 3027 11036 3049
rect 11066 3027 11118 3079
rect 10820 2960 10872 3012
rect 10902 2960 10954 3012
rect 10984 2960 11036 3012
rect 11066 2960 11118 3012
rect 10820 2893 10872 2945
rect 10902 2919 10914 2945
rect 10914 2919 10952 2945
rect 10952 2919 10954 2945
rect 10984 2919 10986 2945
rect 10986 2919 11024 2945
rect 11024 2919 11036 2945
rect 10902 2893 10954 2919
rect 10984 2893 11036 2919
rect 11066 2893 11118 2945
rect 10820 2826 10872 2878
rect 10902 2857 10954 2878
rect 10984 2857 11036 2878
rect 10902 2826 10914 2857
rect 10914 2826 10952 2857
rect 10952 2826 10954 2857
rect 10984 2826 10986 2857
rect 10986 2826 11024 2857
rect 11024 2826 11036 2857
rect 11066 2826 11118 2878
rect 10820 2759 10872 2811
rect 10902 2761 10954 2811
rect 10984 2761 11036 2811
rect 10902 2759 10914 2761
rect 10914 2759 10952 2761
rect 10952 2759 10954 2761
rect 10984 2759 10986 2761
rect 10986 2759 11024 2761
rect 11024 2759 11036 2761
rect 11066 2759 11118 2811
rect 10820 2692 10872 2744
rect 10902 2727 10914 2744
rect 10914 2727 10952 2744
rect 10952 2727 10954 2744
rect 10984 2727 10986 2744
rect 10986 2727 11024 2744
rect 11024 2727 11036 2744
rect 10902 2692 10954 2727
rect 10984 2692 11036 2727
rect 11066 2692 11118 2744
rect 10820 2625 10872 2677
rect 10902 2665 10954 2677
rect 10984 2665 11036 2677
rect 10902 2631 10914 2665
rect 10914 2631 10952 2665
rect 10952 2631 10954 2665
rect 10984 2631 10986 2665
rect 10986 2631 11024 2665
rect 11024 2631 11036 2665
rect 10902 2625 10954 2631
rect 10984 2625 11036 2631
rect 11066 2625 11118 2677
rect 10820 2558 10872 2610
rect 10902 2569 10954 2610
rect 10984 2569 11036 2610
rect 10902 2558 10914 2569
rect 10914 2558 10952 2569
rect 10952 2558 10954 2569
rect 10984 2558 10986 2569
rect 10986 2558 11024 2569
rect 11024 2558 11036 2569
rect 11066 2558 11118 2610
rect 10820 2491 10872 2543
rect 10902 2535 10914 2543
rect 10914 2535 10952 2543
rect 10952 2535 10954 2543
rect 10984 2535 10986 2543
rect 10986 2535 11024 2543
rect 11024 2535 11036 2543
rect 10902 2491 10954 2535
rect 10984 2491 11036 2535
rect 11066 2491 11118 2543
rect 10820 2424 10872 2476
rect 10902 2473 10954 2476
rect 10984 2473 11036 2476
rect 10902 2439 10914 2473
rect 10914 2439 10952 2473
rect 10952 2439 10954 2473
rect 10984 2439 10986 2473
rect 10986 2439 11024 2473
rect 11024 2439 11036 2473
rect 10902 2424 10954 2439
rect 10984 2424 11036 2439
rect 11066 2424 11118 2476
rect 10820 2357 10872 2409
rect 10902 2377 10954 2409
rect 10984 2377 11036 2409
rect 10902 2357 10914 2377
rect 10914 2357 10952 2377
rect 10952 2357 10954 2377
rect 10984 2357 10986 2377
rect 10986 2357 11024 2377
rect 11024 2357 11036 2377
rect 11066 2357 11118 2409
rect 10820 2290 10872 2342
rect 10902 2290 10954 2342
rect 10984 2290 11036 2342
rect 11066 2290 11118 2342
rect 10820 2223 10872 2275
rect 10902 2247 10914 2275
rect 10914 2247 10952 2275
rect 10952 2247 10954 2275
rect 10984 2247 10986 2275
rect 10986 2247 11024 2275
rect 11024 2247 11036 2275
rect 10902 2223 10954 2247
rect 10984 2223 11036 2247
rect 11066 2223 11118 2275
rect 10820 2156 10872 2208
rect 10902 2185 10954 2208
rect 10984 2185 11036 2208
rect 10902 2156 10914 2185
rect 10914 2156 10952 2185
rect 10952 2156 10954 2185
rect 10984 2156 10986 2185
rect 10986 2156 11024 2185
rect 11024 2156 11036 2185
rect 11066 2156 11118 2208
rect 10820 2089 10872 2141
rect 10902 2089 10954 2141
rect 10984 2089 11036 2141
rect 11066 2089 11118 2141
rect 10820 2022 10872 2074
rect 10902 2055 10914 2074
rect 10914 2055 10952 2074
rect 10952 2055 10954 2074
rect 10984 2055 10986 2074
rect 10986 2055 11024 2074
rect 11024 2055 11036 2074
rect 10902 2022 10954 2055
rect 10984 2022 11036 2055
rect 11066 2022 11118 2074
rect 10408 438 10460 490
rect 10490 438 10542 490
rect 10572 438 10624 490
rect 10654 438 10706 490
rect 10408 373 10460 425
rect 10490 373 10542 425
rect 10572 373 10624 425
rect 10654 373 10706 425
rect 7284 304 7336 356
rect 7349 304 7401 356
rect 7414 304 7466 356
rect 7479 304 7531 356
rect 7544 304 7596 356
rect 7609 304 7661 356
rect 7674 304 7726 356
rect 7739 304 7791 356
rect 7804 304 7856 356
rect 7869 304 7921 356
rect 7934 304 7986 356
rect 7999 304 8051 356
rect 8064 304 8116 356
rect 8129 304 8181 356
rect 8194 304 8246 356
rect 8259 304 8311 356
rect 8324 304 8376 356
rect 8389 304 8441 356
rect 8454 304 8506 356
rect 8519 304 8571 356
rect 8584 304 8636 356
rect 8649 304 8701 356
rect 8714 304 8766 356
rect 8779 304 8831 356
rect 8844 304 8896 356
rect 8909 304 8961 356
rect 8974 304 9026 356
rect 9039 304 9091 356
rect 9104 304 9156 356
rect 9169 304 9221 356
rect 9234 304 9286 356
rect 9299 304 9351 356
rect 9364 304 9416 356
rect 9429 304 9481 356
rect 9494 304 9546 356
rect 9559 304 9611 356
rect 9624 304 9676 356
rect 9689 304 9741 356
rect 9753 304 9805 356
rect 9817 304 9869 356
rect 9881 304 9933 356
rect 9945 304 9997 356
rect 10009 304 10061 356
rect 10073 304 10125 356
rect 10137 304 10189 356
rect 10201 304 10253 356
rect 10265 304 10317 356
rect 10329 304 10381 356
rect 10393 304 10445 356
rect 10457 304 10509 356
rect 10521 304 10573 356
rect 10585 304 10637 356
rect 10649 304 10701 356
rect 7284 230 7336 282
rect 7349 230 7401 282
rect 7414 230 7466 282
rect 7479 230 7531 282
rect 7544 230 7596 282
rect 7609 230 7661 282
rect 7674 230 7726 282
rect 7739 230 7791 282
rect 7804 230 7856 282
rect 7869 230 7921 282
rect 7934 230 7986 282
rect 7999 230 8051 282
rect 8064 230 8116 282
rect 8129 230 8181 282
rect 8194 230 8246 282
rect 8259 230 8311 282
rect 8324 230 8376 282
rect 8389 230 8441 282
rect 8454 230 8506 282
rect 8519 230 8571 282
rect 8584 230 8636 282
rect 8649 230 8701 282
rect 8714 230 8766 282
rect 8779 230 8831 282
rect 8844 230 8896 282
rect 8909 230 8961 282
rect 8974 230 9026 282
rect 9039 230 9091 282
rect 9104 230 9156 282
rect 9169 230 9221 282
rect 9234 230 9286 282
rect 9299 230 9351 282
rect 9364 230 9416 282
rect 9429 230 9481 282
rect 9494 230 9546 282
rect 9559 230 9611 282
rect 9624 230 9676 282
rect 9689 230 9741 282
rect 9753 230 9805 282
rect 9817 230 9869 282
rect 9881 230 9933 282
rect 9945 230 9997 282
rect 10009 230 10061 282
rect 10073 230 10125 282
rect 10137 230 10189 282
rect 10201 230 10253 282
rect 10265 230 10317 282
rect 10329 230 10381 282
rect 10393 230 10445 282
rect 10457 230 10509 282
rect 10521 230 10573 282
rect 10585 230 10637 282
rect 10649 230 10701 282
rect 7284 156 7336 208
rect 7349 156 7401 208
rect 7414 156 7466 208
rect 7479 156 7531 208
rect 7544 156 7596 208
rect 7609 156 7661 208
rect 7674 156 7726 208
rect 7739 156 7791 208
rect 7804 156 7856 208
rect 7869 156 7921 208
rect 7934 156 7986 208
rect 7999 156 8051 208
rect 8064 156 8116 208
rect 8129 156 8181 208
rect 8194 156 8246 208
rect 8259 156 8311 208
rect 8324 156 8376 208
rect 8389 156 8441 208
rect 8454 156 8506 208
rect 8519 156 8571 208
rect 8584 156 8636 208
rect 8649 156 8701 208
rect 8714 156 8766 208
rect 8779 156 8831 208
rect 8844 156 8896 208
rect 8909 156 8961 208
rect 8974 156 9026 208
rect 9039 156 9091 208
rect 9104 156 9156 208
rect 9169 156 9221 208
rect 9234 156 9286 208
rect 9299 156 9351 208
rect 9364 156 9416 208
rect 9429 156 9481 208
rect 9494 156 9546 208
rect 9559 156 9611 208
rect 9624 156 9676 208
rect 9689 156 9741 208
rect 9753 156 9805 208
rect 9817 156 9869 208
rect 9881 156 9933 208
rect 9945 156 9997 208
rect 10009 156 10061 208
rect 10073 156 10125 208
rect 10137 156 10189 208
rect 10201 156 10253 208
rect 10265 156 10317 208
rect 10329 156 10381 208
rect 10393 156 10445 208
rect 10457 156 10509 208
rect 10521 156 10573 208
rect 10585 156 10637 208
rect 10649 156 10701 208
rect 7284 82 7336 134
rect 7349 82 7401 134
rect 7414 82 7466 134
rect 7479 82 7531 134
rect 7544 82 7596 134
rect 7609 82 7661 134
rect 7674 82 7726 134
rect 7739 82 7791 134
rect 7804 82 7856 134
rect 7869 82 7921 134
rect 7934 82 7986 134
rect 7999 82 8051 134
rect 8064 82 8116 134
rect 8129 82 8181 134
rect 8194 82 8246 134
rect 8259 82 8311 134
rect 8324 82 8376 134
rect 8389 82 8441 134
rect 8454 82 8506 134
rect 8519 82 8571 134
rect 8584 82 8636 134
rect 8649 82 8701 134
rect 8714 82 8766 134
rect 8779 82 8831 134
rect 8844 82 8896 134
rect 8909 82 8961 134
rect 8974 82 9026 134
rect 9039 82 9091 134
rect 9104 82 9156 134
rect 9169 82 9221 134
rect 9234 82 9286 134
rect 9299 82 9351 134
rect 9364 82 9416 134
rect 9429 82 9481 134
rect 9494 82 9546 134
rect 9559 82 9611 134
rect 9624 82 9676 134
rect 9689 82 9741 134
rect 9753 82 9805 134
rect 9817 82 9869 134
rect 9881 82 9933 134
rect 9945 82 9997 134
rect 10009 82 10061 134
rect 10073 82 10125 134
rect 10137 82 10189 134
rect 10201 82 10253 134
rect 10265 82 10317 134
rect 10329 82 10381 134
rect 10393 82 10445 134
rect 10457 82 10509 134
rect 10521 82 10573 134
rect 10585 82 10637 134
rect 10649 82 10701 134
rect 7284 8 7336 60
rect 7349 8 7401 60
rect 7414 8 7466 60
rect 7479 8 7531 60
rect 7544 8 7596 60
rect 7609 8 7661 60
rect 7674 8 7726 60
rect 7739 8 7791 60
rect 7804 8 7856 60
rect 7869 8 7921 60
rect 7934 8 7986 60
rect 7999 8 8051 60
rect 8064 8 8116 60
rect 8129 8 8181 60
rect 8194 8 8246 60
rect 8259 8 8311 60
rect 8324 8 8376 60
rect 8389 8 8441 60
rect 8454 8 8506 60
rect 8519 8 8571 60
rect 8584 8 8636 60
rect 8649 8 8701 60
rect 8714 8 8766 60
rect 8779 8 8831 60
rect 8844 8 8896 60
rect 8909 8 8961 60
rect 8974 8 9026 60
rect 9039 8 9091 60
rect 9104 8 9156 60
rect 9169 8 9221 60
rect 9234 8 9286 60
rect 9299 8 9351 60
rect 9364 8 9416 60
rect 9429 8 9481 60
rect 9494 8 9546 60
rect 9559 8 9611 60
rect 9624 8 9676 60
rect 9689 8 9741 60
rect 9753 8 9805 60
rect 9817 8 9869 60
rect 9881 8 9933 60
rect 9945 8 9997 60
rect 10009 8 10061 60
rect 10073 8 10125 60
rect 10137 8 10189 60
rect 10201 8 10253 60
rect 10265 8 10317 60
rect 10329 8 10381 60
rect 10393 8 10445 60
rect 10457 8 10509 60
rect 10521 8 10573 60
rect 10585 8 10637 60
rect 10649 8 10701 60
<< metal2 >>
rect 7161 3614 7290 3666
rect 7342 3614 7355 3666
rect 7407 3614 7419 3666
rect 7471 3614 7483 3666
rect 7535 3614 7547 3666
rect 7599 3614 7611 3666
rect 7663 3614 7675 3666
rect 7727 3614 7739 3666
rect 7791 3614 7803 3666
rect 7855 3614 7867 3666
rect 7919 3614 7931 3666
rect 7983 3614 7995 3666
rect 8047 3614 8059 3666
rect 8111 3614 8123 3666
rect 8175 3614 8187 3666
rect 8239 3614 8251 3666
rect 8303 3614 8315 3666
rect 8367 3614 8379 3666
rect 8431 3614 8443 3666
rect 8495 3614 8507 3666
rect 8559 3614 8571 3666
rect 8623 3614 8635 3666
rect 8687 3614 8699 3666
rect 8751 3614 8763 3666
rect 8815 3614 8827 3666
rect 8879 3614 8891 3666
rect 8943 3614 8955 3666
rect 9007 3614 9019 3666
rect 9071 3614 9083 3666
rect 9135 3614 9147 3666
rect 9199 3614 9211 3666
rect 9263 3614 9275 3666
rect 9327 3614 9339 3666
rect 9391 3614 9403 3666
rect 9455 3614 9467 3666
rect 9519 3614 9531 3666
rect 9583 3614 9595 3666
rect 9647 3614 9659 3666
rect 9711 3614 9723 3666
rect 9775 3614 9787 3666
rect 9839 3614 9851 3666
rect 9903 3614 9915 3666
rect 9967 3614 9979 3666
rect 10031 3614 10043 3666
rect 10095 3614 10107 3666
rect 10159 3614 10171 3666
rect 10223 3614 10235 3666
rect 10287 3614 10299 3666
rect 10351 3614 10363 3666
rect 10415 3614 10427 3666
rect 10479 3614 10491 3666
rect 10543 3614 10555 3666
rect 10607 3614 10619 3666
rect 10671 3614 10683 3666
rect 10735 3614 10747 3666
rect 10799 3614 10811 3666
rect 10863 3614 10869 3666
rect 7161 3578 10869 3614
rect 7161 3526 7290 3578
rect 7342 3526 7355 3578
rect 7407 3526 7419 3578
rect 7471 3526 7483 3578
rect 7535 3526 7547 3578
rect 7599 3526 7611 3578
rect 7663 3526 7675 3578
rect 7727 3526 7739 3578
rect 7791 3526 7803 3578
rect 7855 3526 7867 3578
rect 7919 3526 7931 3578
rect 7983 3526 7995 3578
rect 8047 3526 8059 3578
rect 8111 3526 8123 3578
rect 8175 3526 8187 3578
rect 8239 3526 8251 3578
rect 8303 3526 8315 3578
rect 8367 3526 8379 3578
rect 8431 3526 8443 3578
rect 8495 3526 8507 3578
rect 8559 3526 8571 3578
rect 8623 3526 8635 3578
rect 8687 3526 8699 3578
rect 8751 3526 8763 3578
rect 8815 3526 8827 3578
rect 8879 3526 8891 3578
rect 8943 3526 8955 3578
rect 9007 3526 9019 3578
rect 9071 3526 9083 3578
rect 9135 3526 9147 3578
rect 9199 3526 9211 3578
rect 9263 3526 9275 3578
rect 9327 3526 9339 3578
rect 9391 3526 9403 3578
rect 9455 3526 9467 3578
rect 9519 3526 9531 3578
rect 9583 3526 9595 3578
rect 9647 3526 9659 3578
rect 9711 3526 9723 3578
rect 9775 3526 9787 3578
rect 9839 3526 9851 3578
rect 9903 3526 9915 3578
rect 9967 3526 9979 3578
rect 10031 3526 10043 3578
rect 10095 3526 10107 3578
rect 10159 3526 10171 3578
rect 10223 3526 10235 3578
rect 10287 3526 10299 3578
rect 10351 3526 10363 3578
rect 10415 3526 10427 3578
rect 10479 3526 10491 3578
rect 10543 3526 10555 3578
rect 10607 3526 10619 3578
rect 10671 3526 10683 3578
rect 10735 3526 10747 3578
rect 10799 3526 10811 3578
rect 10863 3526 10869 3578
rect 7161 3410 11119 3416
rect 7161 3358 7524 3410
rect 7576 3358 7606 3410
rect 7658 3358 7688 3410
rect 7740 3358 7770 3410
rect 7822 3358 8348 3410
rect 8400 3358 8430 3410
rect 8482 3358 8512 3410
rect 8564 3358 8594 3410
rect 8646 3358 9172 3410
rect 9224 3358 9254 3410
rect 9306 3358 9336 3410
rect 9388 3358 9418 3410
rect 9470 3358 9996 3410
rect 10048 3358 10078 3410
rect 10130 3358 10160 3410
rect 10212 3358 10242 3410
rect 10294 3358 10820 3410
rect 10872 3358 10902 3410
rect 10954 3358 10984 3410
rect 11036 3358 11066 3410
rect 11118 3358 11119 3410
rect 7161 3344 11119 3358
rect 7161 3292 7524 3344
rect 7576 3292 7606 3344
rect 7658 3292 7688 3344
rect 7740 3292 7770 3344
rect 7822 3292 8348 3344
rect 8400 3292 8430 3344
rect 8482 3292 8512 3344
rect 8564 3292 8594 3344
rect 8646 3292 9172 3344
rect 9224 3292 9254 3344
rect 9306 3292 9336 3344
rect 9388 3292 9418 3344
rect 9470 3292 9996 3344
rect 10048 3292 10078 3344
rect 10130 3292 10160 3344
rect 10212 3292 10242 3344
rect 10294 3292 10820 3344
rect 10872 3292 10902 3344
rect 10954 3292 10984 3344
rect 11036 3292 11066 3344
rect 11118 3292 11119 3344
rect 7161 3278 11119 3292
rect 7161 3226 7524 3278
rect 7576 3226 7606 3278
rect 7658 3226 7688 3278
rect 7740 3226 7770 3278
rect 7822 3226 8348 3278
rect 8400 3226 8430 3278
rect 8482 3226 8512 3278
rect 8564 3226 8594 3278
rect 8646 3226 9172 3278
rect 9224 3226 9254 3278
rect 9306 3226 9336 3278
rect 9388 3226 9418 3278
rect 9470 3226 9996 3278
rect 10048 3226 10078 3278
rect 10130 3226 10160 3278
rect 10212 3226 10242 3278
rect 10294 3226 10820 3278
rect 10872 3226 10902 3278
rect 10954 3226 10984 3278
rect 11036 3226 11066 3278
rect 11118 3226 11119 3278
rect 7161 3212 11119 3226
rect 7161 3160 7524 3212
rect 7576 3160 7606 3212
rect 7658 3160 7688 3212
rect 7740 3160 7770 3212
rect 7822 3160 8348 3212
rect 8400 3160 8430 3212
rect 8482 3160 8512 3212
rect 8564 3160 8594 3212
rect 8646 3160 9172 3212
rect 9224 3160 9254 3212
rect 9306 3160 9336 3212
rect 9388 3160 9418 3212
rect 9470 3160 9996 3212
rect 10048 3160 10078 3212
rect 10130 3160 10160 3212
rect 10212 3160 10242 3212
rect 10294 3160 10820 3212
rect 10872 3160 10902 3212
rect 10954 3160 10984 3212
rect 11036 3160 11066 3212
rect 11118 3160 11119 3212
rect 7161 3146 11119 3160
rect 7161 3094 7524 3146
rect 7576 3094 7606 3146
rect 7658 3094 7688 3146
rect 7740 3094 7770 3146
rect 7822 3094 8348 3146
rect 8400 3094 8430 3146
rect 8482 3094 8512 3146
rect 8564 3094 8594 3146
rect 8646 3094 9172 3146
rect 9224 3094 9254 3146
rect 9306 3094 9336 3146
rect 9388 3094 9418 3146
rect 9470 3094 9996 3146
rect 10048 3094 10078 3146
rect 10130 3094 10160 3146
rect 10212 3094 10242 3146
rect 10294 3094 10820 3146
rect 10872 3094 10902 3146
rect 10954 3094 10984 3146
rect 11036 3094 11066 3146
rect 11118 3094 11119 3146
rect 7161 3079 11119 3094
rect 7161 3027 7524 3079
rect 7576 3027 7606 3079
rect 7658 3027 7688 3079
rect 7740 3027 7770 3079
rect 7822 3027 8348 3079
rect 8400 3027 8430 3079
rect 8482 3027 8512 3079
rect 8564 3027 8594 3079
rect 8646 3027 9172 3079
rect 9224 3027 9254 3079
rect 9306 3027 9336 3079
rect 9388 3027 9418 3079
rect 9470 3027 9996 3079
rect 10048 3027 10078 3079
rect 10130 3027 10160 3079
rect 10212 3027 10242 3079
rect 10294 3027 10820 3079
rect 10872 3027 10902 3079
rect 10954 3027 10984 3079
rect 11036 3027 11066 3079
rect 11118 3027 11119 3079
rect 7161 3012 11119 3027
rect 7161 2960 7524 3012
rect 7576 2960 7606 3012
rect 7658 2960 7688 3012
rect 7740 2960 7770 3012
rect 7822 2960 8348 3012
rect 8400 2960 8430 3012
rect 8482 2960 8512 3012
rect 8564 2960 8594 3012
rect 8646 2960 9172 3012
rect 9224 2960 9254 3012
rect 9306 2960 9336 3012
rect 9388 2960 9418 3012
rect 9470 2960 9996 3012
rect 10048 2960 10078 3012
rect 10130 2960 10160 3012
rect 10212 2960 10242 3012
rect 10294 2960 10820 3012
rect 10872 2960 10902 3012
rect 10954 2960 10984 3012
rect 11036 2960 11066 3012
rect 11118 2960 11119 3012
rect 7161 2945 11119 2960
rect 7161 2893 7524 2945
rect 7576 2893 7606 2945
rect 7658 2893 7688 2945
rect 7740 2893 7770 2945
rect 7822 2893 8348 2945
rect 8400 2893 8430 2945
rect 8482 2893 8512 2945
rect 8564 2893 8594 2945
rect 8646 2893 9172 2945
rect 9224 2893 9254 2945
rect 9306 2893 9336 2945
rect 9388 2893 9418 2945
rect 9470 2893 9996 2945
rect 10048 2893 10078 2945
rect 10130 2893 10160 2945
rect 10212 2893 10242 2945
rect 10294 2893 10820 2945
rect 10872 2893 10902 2945
rect 10954 2893 10984 2945
rect 11036 2893 11066 2945
rect 11118 2893 11119 2945
rect 7161 2878 11119 2893
rect 7161 2826 7524 2878
rect 7576 2826 7606 2878
rect 7658 2826 7688 2878
rect 7740 2826 7770 2878
rect 7822 2826 8348 2878
rect 8400 2826 8430 2878
rect 8482 2826 8512 2878
rect 8564 2826 8594 2878
rect 8646 2826 9172 2878
rect 9224 2826 9254 2878
rect 9306 2826 9336 2878
rect 9388 2826 9418 2878
rect 9470 2826 9996 2878
rect 10048 2826 10078 2878
rect 10130 2826 10160 2878
rect 10212 2826 10242 2878
rect 10294 2826 10820 2878
rect 10872 2826 10902 2878
rect 10954 2826 10984 2878
rect 11036 2826 11066 2878
rect 11118 2826 11119 2878
rect 7161 2811 11119 2826
rect 7161 2759 7524 2811
rect 7576 2759 7606 2811
rect 7658 2759 7688 2811
rect 7740 2759 7770 2811
rect 7822 2759 8348 2811
rect 8400 2759 8430 2811
rect 8482 2759 8512 2811
rect 8564 2759 8594 2811
rect 8646 2759 9172 2811
rect 9224 2759 9254 2811
rect 9306 2759 9336 2811
rect 9388 2759 9418 2811
rect 9470 2759 9996 2811
rect 10048 2759 10078 2811
rect 10130 2759 10160 2811
rect 10212 2759 10242 2811
rect 10294 2759 10820 2811
rect 10872 2759 10902 2811
rect 10954 2759 10984 2811
rect 11036 2759 11066 2811
rect 11118 2759 11119 2811
rect 7161 2744 11119 2759
rect 7161 2692 7524 2744
rect 7576 2692 7606 2744
rect 7658 2692 7688 2744
rect 7740 2692 7770 2744
rect 7822 2692 8348 2744
rect 8400 2692 8430 2744
rect 8482 2692 8512 2744
rect 8564 2692 8594 2744
rect 8646 2692 9172 2744
rect 9224 2692 9254 2744
rect 9306 2692 9336 2744
rect 9388 2692 9418 2744
rect 9470 2692 9996 2744
rect 10048 2692 10078 2744
rect 10130 2692 10160 2744
rect 10212 2692 10242 2744
rect 10294 2692 10820 2744
rect 10872 2692 10902 2744
rect 10954 2692 10984 2744
rect 11036 2692 11066 2744
rect 11118 2692 11119 2744
rect 7161 2677 11119 2692
rect 7161 2625 7524 2677
rect 7576 2625 7606 2677
rect 7658 2625 7688 2677
rect 7740 2625 7770 2677
rect 7822 2625 8348 2677
rect 8400 2625 8430 2677
rect 8482 2625 8512 2677
rect 8564 2625 8594 2677
rect 8646 2625 9172 2677
rect 9224 2625 9254 2677
rect 9306 2625 9336 2677
rect 9388 2625 9418 2677
rect 9470 2625 9996 2677
rect 10048 2625 10078 2677
rect 10130 2625 10160 2677
rect 10212 2625 10242 2677
rect 10294 2625 10820 2677
rect 10872 2625 10902 2677
rect 10954 2625 10984 2677
rect 11036 2625 11066 2677
rect 11118 2625 11119 2677
rect 7161 2610 11119 2625
rect 7161 2558 7524 2610
rect 7576 2558 7606 2610
rect 7658 2558 7688 2610
rect 7740 2558 7770 2610
rect 7822 2558 8348 2610
rect 8400 2558 8430 2610
rect 8482 2558 8512 2610
rect 8564 2558 8594 2610
rect 8646 2558 9172 2610
rect 9224 2558 9254 2610
rect 9306 2558 9336 2610
rect 9388 2558 9418 2610
rect 9470 2558 9996 2610
rect 10048 2558 10078 2610
rect 10130 2558 10160 2610
rect 10212 2558 10242 2610
rect 10294 2558 10820 2610
rect 10872 2558 10902 2610
rect 10954 2558 10984 2610
rect 11036 2558 11066 2610
rect 11118 2558 11119 2610
rect 7161 2543 11119 2558
rect 7161 2491 7524 2543
rect 7576 2491 7606 2543
rect 7658 2491 7688 2543
rect 7740 2491 7770 2543
rect 7822 2491 8348 2543
rect 8400 2491 8430 2543
rect 8482 2491 8512 2543
rect 8564 2491 8594 2543
rect 8646 2491 9172 2543
rect 9224 2491 9254 2543
rect 9306 2491 9336 2543
rect 9388 2491 9418 2543
rect 9470 2491 9996 2543
rect 10048 2491 10078 2543
rect 10130 2491 10160 2543
rect 10212 2491 10242 2543
rect 10294 2491 10820 2543
rect 10872 2491 10902 2543
rect 10954 2491 10984 2543
rect 11036 2491 11066 2543
rect 11118 2491 11119 2543
rect 7161 2476 11119 2491
rect 7161 2424 7524 2476
rect 7576 2424 7606 2476
rect 7658 2424 7688 2476
rect 7740 2424 7770 2476
rect 7822 2424 8348 2476
rect 8400 2424 8430 2476
rect 8482 2424 8512 2476
rect 8564 2424 8594 2476
rect 8646 2424 9172 2476
rect 9224 2424 9254 2476
rect 9306 2424 9336 2476
rect 9388 2424 9418 2476
rect 9470 2424 9996 2476
rect 10048 2424 10078 2476
rect 10130 2424 10160 2476
rect 10212 2424 10242 2476
rect 10294 2424 10820 2476
rect 10872 2424 10902 2476
rect 10954 2424 10984 2476
rect 11036 2424 11066 2476
rect 11118 2424 11119 2476
rect 7161 2409 11119 2424
rect 7161 2357 7524 2409
rect 7576 2357 7606 2409
rect 7658 2357 7688 2409
rect 7740 2357 7770 2409
rect 7822 2357 8348 2409
rect 8400 2357 8430 2409
rect 8482 2357 8512 2409
rect 8564 2357 8594 2409
rect 8646 2357 9172 2409
rect 9224 2357 9254 2409
rect 9306 2357 9336 2409
rect 9388 2357 9418 2409
rect 9470 2357 9996 2409
rect 10048 2357 10078 2409
rect 10130 2357 10160 2409
rect 10212 2357 10242 2409
rect 10294 2357 10820 2409
rect 10872 2357 10902 2409
rect 10954 2357 10984 2409
rect 11036 2357 11066 2409
rect 11118 2357 11119 2409
rect 7161 2342 11119 2357
rect 7161 2290 7524 2342
rect 7576 2290 7606 2342
rect 7658 2290 7688 2342
rect 7740 2290 7770 2342
rect 7822 2290 8348 2342
rect 8400 2290 8430 2342
rect 8482 2290 8512 2342
rect 8564 2290 8594 2342
rect 8646 2290 9172 2342
rect 9224 2290 9254 2342
rect 9306 2290 9336 2342
rect 9388 2290 9418 2342
rect 9470 2290 9996 2342
rect 10048 2290 10078 2342
rect 10130 2290 10160 2342
rect 10212 2290 10242 2342
rect 10294 2290 10820 2342
rect 10872 2290 10902 2342
rect 10954 2290 10984 2342
rect 11036 2290 11066 2342
rect 11118 2290 11119 2342
rect 7161 2275 11119 2290
rect 7161 2223 7524 2275
rect 7576 2223 7606 2275
rect 7658 2223 7688 2275
rect 7740 2223 7770 2275
rect 7822 2223 8348 2275
rect 8400 2223 8430 2275
rect 8482 2223 8512 2275
rect 8564 2223 8594 2275
rect 8646 2223 9172 2275
rect 9224 2223 9254 2275
rect 9306 2223 9336 2275
rect 9388 2223 9418 2275
rect 9470 2223 9996 2275
rect 10048 2223 10078 2275
rect 10130 2223 10160 2275
rect 10212 2223 10242 2275
rect 10294 2223 10820 2275
rect 10872 2223 10902 2275
rect 10954 2223 10984 2275
rect 11036 2223 11066 2275
rect 11118 2223 11119 2275
rect 7161 2208 11119 2223
rect 7161 2156 7524 2208
rect 7576 2156 7606 2208
rect 7658 2156 7688 2208
rect 7740 2156 7770 2208
rect 7822 2156 8348 2208
rect 8400 2156 8430 2208
rect 8482 2156 8512 2208
rect 8564 2156 8594 2208
rect 8646 2156 9172 2208
rect 9224 2156 9254 2208
rect 9306 2156 9336 2208
rect 9388 2156 9418 2208
rect 9470 2156 9996 2208
rect 10048 2156 10078 2208
rect 10130 2156 10160 2208
rect 10212 2156 10242 2208
rect 10294 2156 10820 2208
rect 10872 2156 10902 2208
rect 10954 2156 10984 2208
rect 11036 2156 11066 2208
rect 11118 2156 11119 2208
rect 7161 2141 11119 2156
rect 7161 2089 7524 2141
rect 7576 2089 7606 2141
rect 7658 2089 7688 2141
rect 7740 2089 7770 2141
rect 7822 2089 8348 2141
rect 8400 2089 8430 2141
rect 8482 2089 8512 2141
rect 8564 2089 8594 2141
rect 8646 2089 9172 2141
rect 9224 2089 9254 2141
rect 9306 2089 9336 2141
rect 9388 2089 9418 2141
rect 9470 2089 9996 2141
rect 10048 2089 10078 2141
rect 10130 2089 10160 2141
rect 10212 2089 10242 2141
rect 10294 2089 10820 2141
rect 10872 2089 10902 2141
rect 10954 2089 10984 2141
rect 11036 2089 11066 2141
rect 11118 2089 11119 2141
rect 7161 2074 11119 2089
rect 7161 2022 7524 2074
rect 7576 2022 7606 2074
rect 7658 2022 7688 2074
rect 7740 2022 7770 2074
rect 7822 2022 8348 2074
rect 8400 2022 8430 2074
rect 8482 2022 8512 2074
rect 8564 2022 8594 2074
rect 8646 2022 9172 2074
rect 9224 2022 9254 2074
rect 9306 2022 9336 2074
rect 9388 2022 9418 2074
rect 9470 2022 9996 2074
rect 10048 2022 10078 2074
rect 10130 2022 10160 2074
rect 10212 2022 10242 2074
rect 10294 2022 10820 2074
rect 10872 2022 10902 2074
rect 10954 2022 10984 2074
rect 11036 2022 11066 2074
rect 11118 2022 11119 2074
rect 7161 2016 11119 2022
rect 7161 1902 11141 1908
rect 7161 1850 7936 1902
rect 7988 1850 8018 1902
rect 8070 1850 8100 1902
rect 8152 1850 8182 1902
rect 8234 1850 8760 1902
rect 8812 1850 8842 1902
rect 8894 1850 8924 1902
rect 8976 1850 9006 1902
rect 9058 1850 9584 1902
rect 9636 1850 9666 1902
rect 9718 1850 9748 1902
rect 9800 1850 9830 1902
rect 9882 1850 10408 1902
rect 10460 1850 10490 1902
rect 10542 1850 10572 1902
rect 10624 1850 10654 1902
rect 10706 1850 11141 1902
rect 7161 1838 11141 1850
rect 7161 1786 7936 1838
rect 7988 1786 8018 1838
rect 8070 1786 8100 1838
rect 8152 1786 8182 1838
rect 8234 1786 8760 1838
rect 8812 1786 8842 1838
rect 8894 1786 8924 1838
rect 8976 1786 9006 1838
rect 9058 1786 9584 1838
rect 9636 1786 9666 1838
rect 9718 1786 9748 1838
rect 9800 1786 9830 1838
rect 9882 1786 10408 1838
rect 10460 1786 10490 1838
rect 10542 1786 10572 1838
rect 10624 1786 10654 1838
rect 10706 1786 11141 1838
rect 7161 1774 11141 1786
rect 7161 1722 7936 1774
rect 7988 1722 8018 1774
rect 8070 1722 8100 1774
rect 8152 1722 8182 1774
rect 8234 1722 8760 1774
rect 8812 1722 8842 1774
rect 8894 1722 8924 1774
rect 8976 1722 9006 1774
rect 9058 1722 9584 1774
rect 9636 1722 9666 1774
rect 9718 1722 9748 1774
rect 9800 1722 9830 1774
rect 9882 1722 10408 1774
rect 10460 1722 10490 1774
rect 10542 1722 10572 1774
rect 10624 1722 10654 1774
rect 10706 1722 11141 1774
rect 7161 1710 11141 1722
rect 7161 1658 7936 1710
rect 7988 1658 8018 1710
rect 8070 1658 8100 1710
rect 8152 1658 8182 1710
rect 8234 1658 8760 1710
rect 8812 1658 8842 1710
rect 8894 1658 8924 1710
rect 8976 1658 9006 1710
rect 9058 1658 9584 1710
rect 9636 1658 9666 1710
rect 9718 1658 9748 1710
rect 9800 1658 9830 1710
rect 9882 1658 10408 1710
rect 10460 1658 10490 1710
rect 10542 1658 10572 1710
rect 10624 1658 10654 1710
rect 10706 1658 11141 1710
rect 7161 1646 11141 1658
rect 7161 1594 7936 1646
rect 7988 1594 8018 1646
rect 8070 1594 8100 1646
rect 8152 1594 8182 1646
rect 8234 1594 8760 1646
rect 8812 1594 8842 1646
rect 8894 1594 8924 1646
rect 8976 1594 9006 1646
rect 9058 1594 9584 1646
rect 9636 1594 9666 1646
rect 9718 1594 9748 1646
rect 9800 1594 9830 1646
rect 9882 1594 10408 1646
rect 10460 1594 10490 1646
rect 10542 1594 10572 1646
rect 10624 1594 10654 1646
rect 10706 1594 11141 1646
rect 7161 1582 11141 1594
rect 7161 1530 7936 1582
rect 7988 1530 8018 1582
rect 8070 1530 8100 1582
rect 8152 1530 8182 1582
rect 8234 1530 8760 1582
rect 8812 1530 8842 1582
rect 8894 1530 8924 1582
rect 8976 1530 9006 1582
rect 9058 1530 9584 1582
rect 9636 1530 9666 1582
rect 9718 1530 9748 1582
rect 9800 1530 9830 1582
rect 9882 1530 10408 1582
rect 10460 1530 10490 1582
rect 10542 1530 10572 1582
rect 10624 1530 10654 1582
rect 10706 1530 11141 1582
rect 7161 1518 11141 1530
rect 7161 1466 7936 1518
rect 7988 1466 8018 1518
rect 8070 1466 8100 1518
rect 8152 1466 8182 1518
rect 8234 1466 8760 1518
rect 8812 1466 8842 1518
rect 8894 1466 8924 1518
rect 8976 1466 9006 1518
rect 9058 1466 9584 1518
rect 9636 1466 9666 1518
rect 9718 1466 9748 1518
rect 9800 1466 9830 1518
rect 9882 1466 10408 1518
rect 10460 1466 10490 1518
rect 10542 1466 10572 1518
rect 10624 1466 10654 1518
rect 10706 1466 11141 1518
rect 7161 1454 11141 1466
rect 7161 1402 7936 1454
rect 7988 1402 8018 1454
rect 8070 1402 8100 1454
rect 8152 1402 8182 1454
rect 8234 1402 8760 1454
rect 8812 1402 8842 1454
rect 8894 1402 8924 1454
rect 8976 1402 9006 1454
rect 9058 1402 9584 1454
rect 9636 1402 9666 1454
rect 9718 1402 9748 1454
rect 9800 1402 9830 1454
rect 9882 1402 10408 1454
rect 10460 1402 10490 1454
rect 10542 1402 10572 1454
rect 10624 1402 10654 1454
rect 10706 1402 11141 1454
rect 7161 1390 11141 1402
rect 7161 1338 7936 1390
rect 7988 1338 8018 1390
rect 8070 1338 8100 1390
rect 8152 1338 8182 1390
rect 8234 1338 8760 1390
rect 8812 1338 8842 1390
rect 8894 1338 8924 1390
rect 8976 1338 9006 1390
rect 9058 1338 9584 1390
rect 9636 1338 9666 1390
rect 9718 1338 9748 1390
rect 9800 1338 9830 1390
rect 9882 1338 10408 1390
rect 10460 1338 10490 1390
rect 10542 1338 10572 1390
rect 10624 1338 10654 1390
rect 10706 1338 11141 1390
rect 7161 1326 11141 1338
rect 7161 1274 7936 1326
rect 7988 1274 8018 1326
rect 8070 1274 8100 1326
rect 8152 1274 8182 1326
rect 8234 1274 8760 1326
rect 8812 1274 8842 1326
rect 8894 1274 8924 1326
rect 8976 1274 9006 1326
rect 9058 1274 9584 1326
rect 9636 1274 9666 1326
rect 9718 1274 9748 1326
rect 9800 1274 9830 1326
rect 9882 1274 10408 1326
rect 10460 1274 10490 1326
rect 10542 1274 10572 1326
rect 10624 1274 10654 1326
rect 10706 1274 11141 1326
rect 7161 1262 11141 1274
rect 7161 1210 7936 1262
rect 7988 1210 8018 1262
rect 8070 1210 8100 1262
rect 8152 1210 8182 1262
rect 8234 1210 8760 1262
rect 8812 1210 8842 1262
rect 8894 1210 8924 1262
rect 8976 1210 9006 1262
rect 9058 1210 9584 1262
rect 9636 1210 9666 1262
rect 9718 1210 9748 1262
rect 9800 1210 9830 1262
rect 9882 1210 10408 1262
rect 10460 1210 10490 1262
rect 10542 1210 10572 1262
rect 10624 1210 10654 1262
rect 10706 1210 11141 1262
rect 7161 1198 11141 1210
rect 7161 1146 7936 1198
rect 7988 1146 8018 1198
rect 8070 1146 8100 1198
rect 8152 1146 8182 1198
rect 8234 1146 8760 1198
rect 8812 1146 8842 1198
rect 8894 1146 8924 1198
rect 8976 1146 9006 1198
rect 9058 1146 9584 1198
rect 9636 1146 9666 1198
rect 9718 1146 9748 1198
rect 9800 1146 9830 1198
rect 9882 1146 10408 1198
rect 10460 1146 10490 1198
rect 10542 1146 10572 1198
rect 10624 1146 10654 1198
rect 10706 1146 11141 1198
rect 7161 1134 11141 1146
rect 7161 1082 7936 1134
rect 7988 1082 8018 1134
rect 8070 1082 8100 1134
rect 8152 1082 8182 1134
rect 8234 1082 8760 1134
rect 8812 1082 8842 1134
rect 8894 1082 8924 1134
rect 8976 1082 9006 1134
rect 9058 1082 9584 1134
rect 9636 1082 9666 1134
rect 9718 1082 9748 1134
rect 9800 1082 9830 1134
rect 9882 1082 10408 1134
rect 10460 1082 10490 1134
rect 10542 1082 10572 1134
rect 10624 1082 10654 1134
rect 10706 1082 11141 1134
rect 7161 1070 11141 1082
rect 7161 1018 7936 1070
rect 7988 1018 8018 1070
rect 8070 1018 8100 1070
rect 8152 1018 8182 1070
rect 8234 1018 8760 1070
rect 8812 1018 8842 1070
rect 8894 1018 8924 1070
rect 8976 1018 9006 1070
rect 9058 1018 9584 1070
rect 9636 1018 9666 1070
rect 9718 1018 9748 1070
rect 9800 1018 9830 1070
rect 9882 1018 10408 1070
rect 10460 1018 10490 1070
rect 10542 1018 10572 1070
rect 10624 1018 10654 1070
rect 10706 1018 11141 1070
rect 7161 1006 11141 1018
rect 7161 954 7936 1006
rect 7988 954 8018 1006
rect 8070 954 8100 1006
rect 8152 954 8182 1006
rect 8234 954 8760 1006
rect 8812 954 8842 1006
rect 8894 954 8924 1006
rect 8976 954 9006 1006
rect 9058 954 9584 1006
rect 9636 954 9666 1006
rect 9718 954 9748 1006
rect 9800 954 9830 1006
rect 9882 954 10408 1006
rect 10460 954 10490 1006
rect 10542 954 10572 1006
rect 10624 954 10654 1006
rect 10706 954 11141 1006
rect 7161 942 11141 954
rect 7161 890 7936 942
rect 7988 890 8018 942
rect 8070 890 8100 942
rect 8152 890 8182 942
rect 8234 890 8760 942
rect 8812 890 8842 942
rect 8894 890 8924 942
rect 8976 890 9006 942
rect 9058 890 9584 942
rect 9636 890 9666 942
rect 9718 890 9748 942
rect 9800 890 9830 942
rect 9882 890 10408 942
rect 10460 890 10490 942
rect 10542 890 10572 942
rect 10624 890 10654 942
rect 10706 890 11141 942
rect 7161 878 11141 890
rect 7161 826 7936 878
rect 7988 826 8018 878
rect 8070 826 8100 878
rect 8152 826 8182 878
rect 8234 826 8760 878
rect 8812 826 8842 878
rect 8894 826 8924 878
rect 8976 826 9006 878
rect 9058 826 9584 878
rect 9636 826 9666 878
rect 9718 826 9748 878
rect 9800 826 9830 878
rect 9882 826 10408 878
rect 10460 826 10490 878
rect 10542 826 10572 878
rect 10624 826 10654 878
rect 10706 826 11141 878
rect 7161 814 11141 826
rect 7161 762 7936 814
rect 7988 762 8018 814
rect 8070 762 8100 814
rect 8152 762 8182 814
rect 8234 762 8760 814
rect 8812 762 8842 814
rect 8894 762 8924 814
rect 8976 762 9006 814
rect 9058 762 9584 814
rect 9636 762 9666 814
rect 9718 762 9748 814
rect 9800 762 9830 814
rect 9882 762 10408 814
rect 10460 762 10490 814
rect 10542 762 10572 814
rect 10624 762 10654 814
rect 10706 762 11141 814
rect 7161 750 11141 762
rect 7161 698 7936 750
rect 7988 698 8018 750
rect 8070 698 8100 750
rect 8152 698 8182 750
rect 8234 698 8760 750
rect 8812 698 8842 750
rect 8894 698 8924 750
rect 8976 698 9006 750
rect 9058 698 9584 750
rect 9636 698 9666 750
rect 9718 698 9748 750
rect 9800 698 9830 750
rect 9882 698 10408 750
rect 10460 698 10490 750
rect 10542 698 10572 750
rect 10624 698 10654 750
rect 10706 698 11141 750
rect 7161 685 11141 698
rect 7161 633 7936 685
rect 7988 633 8018 685
rect 8070 633 8100 685
rect 8152 633 8182 685
rect 8234 633 8760 685
rect 8812 633 8842 685
rect 8894 633 8924 685
rect 8976 633 9006 685
rect 9058 633 9584 685
rect 9636 633 9666 685
rect 9718 633 9748 685
rect 9800 633 9830 685
rect 9882 633 10408 685
rect 10460 633 10490 685
rect 10542 633 10572 685
rect 10624 633 10654 685
rect 10706 633 11141 685
rect 7161 620 11141 633
rect 7161 568 7936 620
rect 7988 568 8018 620
rect 8070 568 8100 620
rect 8152 568 8182 620
rect 8234 568 8760 620
rect 8812 568 8842 620
rect 8894 568 8924 620
rect 8976 568 9006 620
rect 9058 568 9584 620
rect 9636 568 9666 620
rect 9718 568 9748 620
rect 9800 568 9830 620
rect 9882 568 10408 620
rect 10460 568 10490 620
rect 10542 568 10572 620
rect 10624 568 10654 620
rect 10706 568 11141 620
rect 7161 555 11141 568
rect 7161 503 7936 555
rect 7988 503 8018 555
rect 8070 503 8100 555
rect 8152 503 8182 555
rect 8234 503 8760 555
rect 8812 503 8842 555
rect 8894 503 8924 555
rect 8976 503 9006 555
rect 9058 503 9584 555
rect 9636 503 9666 555
rect 9718 503 9748 555
rect 9800 503 9830 555
rect 9882 503 10408 555
rect 10460 503 10490 555
rect 10542 503 10572 555
rect 10624 503 10654 555
rect 10706 503 11141 555
rect 7161 490 11141 503
rect 7161 438 7936 490
rect 7988 438 8018 490
rect 8070 438 8100 490
rect 8152 438 8182 490
rect 8234 438 8760 490
rect 8812 438 8842 490
rect 8894 438 8924 490
rect 8976 438 9006 490
rect 9058 438 9584 490
rect 9636 438 9666 490
rect 9718 438 9748 490
rect 9800 438 9830 490
rect 9882 438 10408 490
rect 10460 438 10490 490
rect 10542 438 10572 490
rect 10624 438 10654 490
rect 10706 438 11141 490
rect 7161 425 11141 438
rect 7161 373 7936 425
rect 7988 373 8018 425
rect 8070 373 8100 425
rect 8152 373 8182 425
rect 8234 373 8760 425
rect 8812 373 8842 425
rect 8894 373 8924 425
rect 8976 373 9006 425
rect 9058 373 9584 425
rect 9636 373 9666 425
rect 9718 373 9748 425
rect 9800 373 9830 425
rect 9882 373 10408 425
rect 10460 373 10490 425
rect 10542 373 10572 425
rect 10624 373 10654 425
rect 10706 373 11141 425
rect 7161 356 11141 373
rect 7161 304 7284 356
rect 7336 304 7349 356
rect 7401 304 7414 356
rect 7466 304 7479 356
rect 7531 304 7544 356
rect 7596 304 7609 356
rect 7661 304 7674 356
rect 7726 304 7739 356
rect 7791 304 7804 356
rect 7856 304 7869 356
rect 7921 304 7934 356
rect 7986 304 7999 356
rect 8051 304 8064 356
rect 8116 304 8129 356
rect 8181 304 8194 356
rect 8246 304 8259 356
rect 8311 304 8324 356
rect 8376 304 8389 356
rect 8441 304 8454 356
rect 8506 304 8519 356
rect 8571 304 8584 356
rect 8636 304 8649 356
rect 8701 304 8714 356
rect 8766 304 8779 356
rect 8831 304 8844 356
rect 8896 304 8909 356
rect 8961 304 8974 356
rect 9026 304 9039 356
rect 9091 304 9104 356
rect 9156 304 9169 356
rect 9221 304 9234 356
rect 9286 304 9299 356
rect 9351 304 9364 356
rect 9416 304 9429 356
rect 9481 304 9494 356
rect 9546 304 9559 356
rect 9611 304 9624 356
rect 9676 304 9689 356
rect 9741 304 9753 356
rect 9805 304 9817 356
rect 9869 304 9881 356
rect 9933 304 9945 356
rect 9997 304 10009 356
rect 10061 304 10073 356
rect 10125 304 10137 356
rect 10189 304 10201 356
rect 10253 304 10265 356
rect 10317 304 10329 356
rect 10381 304 10393 356
rect 10445 304 10457 356
rect 10509 304 10521 356
rect 10573 304 10585 356
rect 10637 304 10649 356
rect 10701 304 11141 356
rect 7161 282 11141 304
rect 7161 230 7284 282
rect 7336 230 7349 282
rect 7401 230 7414 282
rect 7466 230 7479 282
rect 7531 230 7544 282
rect 7596 230 7609 282
rect 7661 230 7674 282
rect 7726 230 7739 282
rect 7791 230 7804 282
rect 7856 230 7869 282
rect 7921 230 7934 282
rect 7986 230 7999 282
rect 8051 230 8064 282
rect 8116 230 8129 282
rect 8181 230 8194 282
rect 8246 230 8259 282
rect 8311 230 8324 282
rect 8376 230 8389 282
rect 8441 230 8454 282
rect 8506 230 8519 282
rect 8571 230 8584 282
rect 8636 230 8649 282
rect 8701 230 8714 282
rect 8766 230 8779 282
rect 8831 230 8844 282
rect 8896 230 8909 282
rect 8961 230 8974 282
rect 9026 230 9039 282
rect 9091 230 9104 282
rect 9156 230 9169 282
rect 9221 230 9234 282
rect 9286 230 9299 282
rect 9351 230 9364 282
rect 9416 230 9429 282
rect 9481 230 9494 282
rect 9546 230 9559 282
rect 9611 230 9624 282
rect 9676 230 9689 282
rect 9741 230 9753 282
rect 9805 230 9817 282
rect 9869 230 9881 282
rect 9933 230 9945 282
rect 9997 230 10009 282
rect 10061 230 10073 282
rect 10125 230 10137 282
rect 10189 230 10201 282
rect 10253 230 10265 282
rect 10317 230 10329 282
rect 10381 230 10393 282
rect 10445 230 10457 282
rect 10509 230 10521 282
rect 10573 230 10585 282
rect 10637 230 10649 282
rect 10701 230 11141 282
rect 7161 208 11141 230
rect 7161 156 7284 208
rect 7336 156 7349 208
rect 7401 156 7414 208
rect 7466 156 7479 208
rect 7531 156 7544 208
rect 7596 156 7609 208
rect 7661 156 7674 208
rect 7726 156 7739 208
rect 7791 156 7804 208
rect 7856 156 7869 208
rect 7921 156 7934 208
rect 7986 156 7999 208
rect 8051 156 8064 208
rect 8116 156 8129 208
rect 8181 156 8194 208
rect 8246 156 8259 208
rect 8311 156 8324 208
rect 8376 156 8389 208
rect 8441 156 8454 208
rect 8506 156 8519 208
rect 8571 156 8584 208
rect 8636 156 8649 208
rect 8701 156 8714 208
rect 8766 156 8779 208
rect 8831 156 8844 208
rect 8896 156 8909 208
rect 8961 156 8974 208
rect 9026 156 9039 208
rect 9091 156 9104 208
rect 9156 156 9169 208
rect 9221 156 9234 208
rect 9286 156 9299 208
rect 9351 156 9364 208
rect 9416 156 9429 208
rect 9481 156 9494 208
rect 9546 156 9559 208
rect 9611 156 9624 208
rect 9676 156 9689 208
rect 9741 156 9753 208
rect 9805 156 9817 208
rect 9869 156 9881 208
rect 9933 156 9945 208
rect 9997 156 10009 208
rect 10061 156 10073 208
rect 10125 156 10137 208
rect 10189 156 10201 208
rect 10253 156 10265 208
rect 10317 156 10329 208
rect 10381 156 10393 208
rect 10445 156 10457 208
rect 10509 156 10521 208
rect 10573 156 10585 208
rect 10637 156 10649 208
rect 10701 156 11141 208
rect 7161 134 11141 156
rect 7161 82 7284 134
rect 7336 82 7349 134
rect 7401 82 7414 134
rect 7466 82 7479 134
rect 7531 82 7544 134
rect 7596 82 7609 134
rect 7661 82 7674 134
rect 7726 82 7739 134
rect 7791 82 7804 134
rect 7856 82 7869 134
rect 7921 82 7934 134
rect 7986 82 7999 134
rect 8051 82 8064 134
rect 8116 82 8129 134
rect 8181 82 8194 134
rect 8246 82 8259 134
rect 8311 82 8324 134
rect 8376 82 8389 134
rect 8441 82 8454 134
rect 8506 82 8519 134
rect 8571 82 8584 134
rect 8636 82 8649 134
rect 8701 82 8714 134
rect 8766 82 8779 134
rect 8831 82 8844 134
rect 8896 82 8909 134
rect 8961 82 8974 134
rect 9026 82 9039 134
rect 9091 82 9104 134
rect 9156 82 9169 134
rect 9221 82 9234 134
rect 9286 82 9299 134
rect 9351 82 9364 134
rect 9416 82 9429 134
rect 9481 82 9494 134
rect 9546 82 9559 134
rect 9611 82 9624 134
rect 9676 82 9689 134
rect 9741 82 9753 134
rect 9805 82 9817 134
rect 9869 82 9881 134
rect 9933 82 9945 134
rect 9997 82 10009 134
rect 10061 82 10073 134
rect 10125 82 10137 134
rect 10189 82 10201 134
rect 10253 82 10265 134
rect 10317 82 10329 134
rect 10381 82 10393 134
rect 10445 82 10457 134
rect 10509 82 10521 134
rect 10573 82 10585 134
rect 10637 82 10649 134
rect 10701 82 11141 134
rect 7161 60 11141 82
rect 7161 8 7284 60
rect 7336 8 7349 60
rect 7401 8 7414 60
rect 7466 8 7479 60
rect 7531 8 7544 60
rect 7596 8 7609 60
rect 7661 8 7674 60
rect 7726 8 7739 60
rect 7791 8 7804 60
rect 7856 8 7869 60
rect 7921 8 7934 60
rect 7986 8 7999 60
rect 8051 8 8064 60
rect 8116 8 8129 60
rect 8181 8 8194 60
rect 8246 8 8259 60
rect 8311 8 8324 60
rect 8376 8 8389 60
rect 8441 8 8454 60
rect 8506 8 8519 60
rect 8571 8 8584 60
rect 8636 8 8649 60
rect 8701 8 8714 60
rect 8766 8 8779 60
rect 8831 8 8844 60
rect 8896 8 8909 60
rect 8961 8 8974 60
rect 9026 8 9039 60
rect 9091 8 9104 60
rect 9156 8 9169 60
rect 9221 8 9234 60
rect 9286 8 9299 60
rect 9351 8 9364 60
rect 9416 8 9429 60
rect 9481 8 9494 60
rect 9546 8 9559 60
rect 9611 8 9624 60
rect 9676 8 9689 60
rect 9741 8 9753 60
rect 9805 8 9817 60
rect 9869 8 9881 60
rect 9933 8 9945 60
rect 9997 8 10009 60
rect 10061 8 10073 60
rect 10125 8 10137 60
rect 10189 8 10201 60
rect 10253 8 10265 60
rect 10317 8 10329 60
rect 10381 8 10393 60
rect 10445 8 10457 60
rect 10509 8 10521 60
rect 10573 8 10585 60
rect 10637 8 10649 60
rect 10701 8 11141 60
rect 7161 0 11141 8
<< properties >>
string GDS_END 5229174
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 4969970
<< end >>
