magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 0 0 856 806
<< pmoslvt >>
rect 204 102 274 704
rect 330 102 400 704
rect 456 102 526 704
rect 582 102 652 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 274 692 330 704
rect 274 658 285 692
rect 319 658 330 692
rect 274 624 330 658
rect 274 590 285 624
rect 319 590 330 624
rect 274 556 330 590
rect 274 522 285 556
rect 319 522 330 556
rect 274 488 330 522
rect 274 454 285 488
rect 319 454 330 488
rect 274 420 330 454
rect 274 386 285 420
rect 319 386 330 420
rect 274 352 330 386
rect 274 318 285 352
rect 319 318 330 352
rect 274 284 330 318
rect 274 250 285 284
rect 319 250 330 284
rect 274 216 330 250
rect 274 182 285 216
rect 319 182 330 216
rect 274 148 330 182
rect 274 114 285 148
rect 319 114 330 148
rect 274 102 330 114
rect 400 692 456 704
rect 400 658 411 692
rect 445 658 456 692
rect 400 624 456 658
rect 400 590 411 624
rect 445 590 456 624
rect 400 556 456 590
rect 400 522 411 556
rect 445 522 456 556
rect 400 488 456 522
rect 400 454 411 488
rect 445 454 456 488
rect 400 420 456 454
rect 400 386 411 420
rect 445 386 456 420
rect 400 352 456 386
rect 400 318 411 352
rect 445 318 456 352
rect 400 284 456 318
rect 400 250 411 284
rect 445 250 456 284
rect 400 216 456 250
rect 400 182 411 216
rect 445 182 456 216
rect 400 148 456 182
rect 400 114 411 148
rect 445 114 456 148
rect 400 102 456 114
rect 526 692 582 704
rect 526 658 537 692
rect 571 658 582 692
rect 526 624 582 658
rect 526 590 537 624
rect 571 590 582 624
rect 526 556 582 590
rect 526 522 537 556
rect 571 522 582 556
rect 526 488 582 522
rect 526 454 537 488
rect 571 454 582 488
rect 526 420 582 454
rect 526 386 537 420
rect 571 386 582 420
rect 526 352 582 386
rect 526 318 537 352
rect 571 318 582 352
rect 526 284 582 318
rect 526 250 537 284
rect 571 250 582 284
rect 526 216 582 250
rect 526 182 537 216
rect 571 182 582 216
rect 526 148 582 182
rect 526 114 537 148
rect 571 114 582 148
rect 526 102 582 114
rect 652 692 708 704
rect 652 658 663 692
rect 697 658 708 692
rect 652 624 708 658
rect 652 590 663 624
rect 697 590 708 624
rect 652 556 708 590
rect 652 522 663 556
rect 697 522 708 556
rect 652 488 708 522
rect 652 454 663 488
rect 697 454 708 488
rect 652 420 708 454
rect 652 386 663 420
rect 697 386 708 420
rect 652 352 708 386
rect 652 318 663 352
rect 697 318 708 352
rect 652 284 708 318
rect 652 250 663 284
rect 697 250 708 284
rect 652 216 708 250
rect 652 182 663 216
rect 697 182 708 216
rect 652 148 708 182
rect 652 114 663 148
rect 697 114 708 148
rect 652 102 708 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 285 658 319 692
rect 285 590 319 624
rect 285 522 319 556
rect 285 454 319 488
rect 285 386 319 420
rect 285 318 319 352
rect 285 250 319 284
rect 285 182 319 216
rect 285 114 319 148
rect 411 658 445 692
rect 411 590 445 624
rect 411 522 445 556
rect 411 454 445 488
rect 411 386 445 420
rect 411 318 445 352
rect 411 250 445 284
rect 411 182 445 216
rect 411 114 445 148
rect 537 658 571 692
rect 537 590 571 624
rect 537 522 571 556
rect 537 454 571 488
rect 537 386 571 420
rect 537 318 571 352
rect 537 250 571 284
rect 537 182 571 216
rect 537 114 571 148
rect 663 658 697 692
rect 663 590 697 624
rect 663 522 697 556
rect 663 454 697 488
rect 663 386 697 420
rect 663 318 697 352
rect 663 250 697 284
rect 663 182 697 216
rect 663 114 697 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 762 658 820 704
rect 762 624 774 658
rect 808 624 820 658
rect 762 590 820 624
rect 762 556 774 590
rect 808 556 820 590
rect 762 522 820 556
rect 762 488 774 522
rect 808 488 820 522
rect 762 454 820 488
rect 762 420 774 454
rect 808 420 820 454
rect 762 386 820 420
rect 762 352 774 386
rect 808 352 820 386
rect 762 318 820 352
rect 762 284 774 318
rect 808 284 820 318
rect 762 250 820 284
rect 762 216 774 250
rect 808 216 820 250
rect 762 182 820 216
rect 762 148 774 182
rect 808 148 820 182
rect 762 102 820 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 774 624 808 658
rect 774 556 808 590
rect 774 488 808 522
rect 774 420 808 454
rect 774 352 808 386
rect 774 284 808 318
rect 774 216 808 250
rect 774 148 808 182
<< poly >>
rect 191 786 665 806
rect 191 752 207 786
rect 241 752 275 786
rect 309 752 343 786
rect 377 752 411 786
rect 445 752 479 786
rect 513 752 547 786
rect 581 752 615 786
rect 649 752 665 786
rect 191 736 665 752
rect 204 704 274 736
rect 330 704 400 736
rect 456 704 526 736
rect 582 704 652 736
rect 204 70 274 102
rect 330 70 400 102
rect 456 70 526 102
rect 582 70 652 102
rect 191 54 665 70
rect 191 20 207 54
rect 241 20 275 54
rect 309 20 343 54
rect 377 20 411 54
rect 445 20 479 54
rect 513 20 547 54
rect 581 20 615 54
rect 649 20 665 54
rect 191 0 665 20
<< polycont >>
rect 207 752 241 786
rect 275 752 309 786
rect 343 752 377 786
rect 411 752 445 786
rect 479 752 513 786
rect 547 752 581 786
rect 615 752 649 786
rect 207 20 241 54
rect 275 20 309 54
rect 343 20 377 54
rect 411 20 445 54
rect 479 20 513 54
rect 547 20 581 54
rect 615 20 649 54
<< locali >>
rect 191 752 195 786
rect 241 752 267 786
rect 309 752 339 786
rect 377 752 411 786
rect 445 752 479 786
rect 517 752 547 786
rect 589 752 615 786
rect 661 752 665 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 285 692 319 708
rect 285 624 319 638
rect 285 556 319 566
rect 285 488 319 494
rect 285 420 319 422
rect 285 384 319 386
rect 285 312 319 318
rect 285 240 319 250
rect 285 168 319 182
rect 285 98 319 114
rect 411 692 445 708
rect 411 624 445 638
rect 411 556 445 566
rect 411 488 445 494
rect 411 420 445 422
rect 411 384 445 386
rect 411 312 445 318
rect 411 240 445 250
rect 411 168 445 182
rect 411 98 445 114
rect 537 692 571 708
rect 537 624 571 638
rect 537 556 571 566
rect 537 488 571 494
rect 537 420 571 422
rect 537 384 571 386
rect 537 312 571 318
rect 537 240 571 250
rect 537 168 571 182
rect 537 98 571 114
rect 663 692 697 708
rect 663 624 697 638
rect 663 556 697 566
rect 663 488 697 494
rect 663 420 697 422
rect 663 384 697 386
rect 663 312 697 318
rect 663 240 697 250
rect 663 168 697 182
rect 774 672 808 674
rect 774 600 808 624
rect 774 528 808 556
rect 774 456 808 488
rect 774 386 808 420
rect 774 318 808 350
rect 774 250 808 278
rect 774 182 808 206
rect 774 132 808 134
rect 663 98 697 114
rect 191 20 195 54
rect 241 20 267 54
rect 309 20 339 54
rect 377 20 411 54
rect 445 20 479 54
rect 517 20 547 54
rect 589 20 615 54
rect 661 20 665 54
<< viali >>
rect 195 752 207 786
rect 207 752 229 786
rect 267 752 275 786
rect 275 752 301 786
rect 339 752 343 786
rect 343 752 373 786
rect 411 752 445 786
rect 483 752 513 786
rect 513 752 517 786
rect 555 752 581 786
rect 581 752 589 786
rect 627 752 649 786
rect 649 752 661 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 285 658 319 672
rect 285 638 319 658
rect 285 590 319 600
rect 285 566 319 590
rect 285 522 319 528
rect 285 494 319 522
rect 285 454 319 456
rect 285 422 319 454
rect 285 352 319 384
rect 285 350 319 352
rect 285 284 319 312
rect 285 278 319 284
rect 285 216 319 240
rect 285 206 319 216
rect 285 148 319 168
rect 285 134 319 148
rect 411 658 445 672
rect 411 638 445 658
rect 411 590 445 600
rect 411 566 445 590
rect 411 522 445 528
rect 411 494 445 522
rect 411 454 445 456
rect 411 422 445 454
rect 411 352 445 384
rect 411 350 445 352
rect 411 284 445 312
rect 411 278 445 284
rect 411 216 445 240
rect 411 206 445 216
rect 411 148 445 168
rect 411 134 445 148
rect 537 658 571 672
rect 537 638 571 658
rect 537 590 571 600
rect 537 566 571 590
rect 537 522 571 528
rect 537 494 571 522
rect 537 454 571 456
rect 537 422 571 454
rect 537 352 571 384
rect 537 350 571 352
rect 537 284 571 312
rect 537 278 571 284
rect 537 216 571 240
rect 537 206 571 216
rect 537 148 571 168
rect 537 134 571 148
rect 663 658 697 672
rect 663 638 697 658
rect 663 590 697 600
rect 663 566 697 590
rect 663 522 697 528
rect 663 494 697 522
rect 663 454 697 456
rect 663 422 697 454
rect 663 352 697 384
rect 663 350 697 352
rect 663 284 697 312
rect 663 278 697 284
rect 663 216 697 240
rect 663 206 697 216
rect 663 148 697 168
rect 663 134 697 148
rect 774 658 808 672
rect 774 638 808 658
rect 774 590 808 600
rect 774 566 808 590
rect 774 522 808 528
rect 774 494 808 522
rect 774 454 808 456
rect 774 422 808 454
rect 774 352 808 384
rect 774 350 808 352
rect 774 284 808 312
rect 774 278 808 284
rect 774 216 808 240
rect 774 206 808 216
rect 774 148 808 168
rect 774 134 808 148
rect 195 20 207 54
rect 207 20 229 54
rect 267 20 275 54
rect 275 20 301 54
rect 339 20 343 54
rect 343 20 373 54
rect 411 20 445 54
rect 483 20 513 54
rect 513 20 517 54
rect 555 20 581 54
rect 581 20 589 54
rect 627 20 649 54
rect 649 20 661 54
<< metal1 >>
rect 183 786 673 806
rect 183 752 195 786
rect 229 752 267 786
rect 301 752 339 786
rect 373 752 411 786
rect 445 752 483 786
rect 517 752 555 786
rect 589 752 627 786
rect 661 752 673 786
rect 183 740 673 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 276 678 328 684
rect 276 614 328 626
rect 276 550 328 562
rect 276 494 285 498
rect 319 494 328 498
rect 276 486 328 494
rect 276 422 285 434
rect 319 422 328 434
rect 276 384 328 422
rect 276 350 285 384
rect 319 350 328 384
rect 276 312 328 350
rect 276 278 285 312
rect 319 278 328 312
rect 276 240 328 278
rect 276 206 285 240
rect 319 206 328 240
rect 276 168 328 206
rect 276 134 285 168
rect 319 134 328 168
rect 276 122 328 134
rect 402 672 454 684
rect 402 638 411 672
rect 445 638 454 672
rect 402 600 454 638
rect 402 566 411 600
rect 445 566 454 600
rect 402 528 454 566
rect 402 494 411 528
rect 445 494 454 528
rect 402 456 454 494
rect 402 422 411 456
rect 445 422 454 456
rect 402 384 454 422
rect 402 372 411 384
rect 445 372 454 384
rect 402 312 454 320
rect 402 308 411 312
rect 445 308 454 312
rect 402 244 454 256
rect 402 180 454 192
rect 402 122 454 128
rect 528 678 580 684
rect 528 614 580 626
rect 528 550 580 562
rect 528 494 537 498
rect 571 494 580 498
rect 528 486 580 494
rect 528 422 537 434
rect 571 422 580 434
rect 528 384 580 422
rect 528 350 537 384
rect 571 350 580 384
rect 528 312 580 350
rect 528 278 537 312
rect 571 278 580 312
rect 528 240 580 278
rect 528 206 537 240
rect 571 206 580 240
rect 528 168 580 206
rect 528 134 537 168
rect 571 134 580 168
rect 528 122 580 134
rect 654 672 706 684
rect 654 638 663 672
rect 697 638 706 672
rect 654 600 706 638
rect 654 566 663 600
rect 697 566 706 600
rect 654 528 706 566
rect 654 494 663 528
rect 697 494 706 528
rect 654 456 706 494
rect 654 422 663 456
rect 697 422 706 456
rect 654 384 706 422
rect 654 372 663 384
rect 697 372 706 384
rect 654 312 706 320
rect 654 308 663 312
rect 697 308 706 312
rect 654 244 706 256
rect 654 180 706 192
rect 654 122 706 128
rect 762 672 820 684
rect 762 638 774 672
rect 808 638 820 672
rect 762 600 820 638
rect 762 566 774 600
rect 808 566 820 600
rect 762 528 820 566
rect 762 494 774 528
rect 808 494 820 528
rect 762 456 820 494
rect 762 422 774 456
rect 808 422 820 456
rect 762 384 820 422
rect 762 350 774 384
rect 808 350 820 384
rect 762 312 820 350
rect 762 278 774 312
rect 808 278 820 312
rect 762 240 820 278
rect 762 206 774 240
rect 808 206 820 240
rect 762 168 820 206
rect 762 134 774 168
rect 808 134 820 168
rect 762 122 820 134
rect 183 54 673 66
rect 183 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 673 54
rect 183 0 673 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 276 672 328 678
rect 276 638 285 672
rect 285 638 319 672
rect 319 638 328 672
rect 276 626 328 638
rect 276 600 328 614
rect 276 566 285 600
rect 285 566 319 600
rect 319 566 328 600
rect 276 562 328 566
rect 276 528 328 550
rect 276 498 285 528
rect 285 498 319 528
rect 319 498 328 528
rect 276 456 328 486
rect 276 434 285 456
rect 285 434 319 456
rect 319 434 328 456
rect 402 350 411 372
rect 411 350 445 372
rect 445 350 454 372
rect 402 320 454 350
rect 402 278 411 308
rect 411 278 445 308
rect 445 278 454 308
rect 402 256 454 278
rect 402 240 454 244
rect 402 206 411 240
rect 411 206 445 240
rect 445 206 454 240
rect 402 192 454 206
rect 402 168 454 180
rect 402 134 411 168
rect 411 134 445 168
rect 445 134 454 168
rect 402 128 454 134
rect 528 672 580 678
rect 528 638 537 672
rect 537 638 571 672
rect 571 638 580 672
rect 528 626 580 638
rect 528 600 580 614
rect 528 566 537 600
rect 537 566 571 600
rect 571 566 580 600
rect 528 562 580 566
rect 528 528 580 550
rect 528 498 537 528
rect 537 498 571 528
rect 571 498 580 528
rect 528 456 580 486
rect 528 434 537 456
rect 537 434 571 456
rect 571 434 580 456
rect 654 350 663 372
rect 663 350 697 372
rect 697 350 706 372
rect 654 320 706 350
rect 654 278 663 308
rect 663 278 697 308
rect 697 278 706 308
rect 654 256 706 278
rect 654 240 706 244
rect 654 206 663 240
rect 663 206 697 240
rect 697 206 706 240
rect 654 192 706 206
rect 654 168 706 180
rect 654 134 663 168
rect 663 134 697 168
rect 697 134 706 168
rect 654 128 706 134
<< metal2 >>
rect 10 678 846 684
rect 10 626 276 678
rect 328 626 528 678
rect 580 626 846 678
rect 10 614 846 626
rect 10 562 276 614
rect 328 562 528 614
rect 580 562 846 614
rect 10 550 846 562
rect 10 498 276 550
rect 328 498 528 550
rect 580 498 846 550
rect 10 486 846 498
rect 10 434 276 486
rect 328 434 528 486
rect 580 434 846 486
rect 10 428 846 434
rect 10 372 846 378
rect 10 320 150 372
rect 202 320 402 372
rect 454 320 654 372
rect 706 320 846 372
rect 10 308 846 320
rect 10 256 150 308
rect 202 256 402 308
rect 454 256 654 308
rect 706 256 846 308
rect 10 244 846 256
rect 10 192 150 244
rect 202 192 402 244
rect 454 192 654 244
rect 706 192 846 244
rect 10 180 846 192
rect 10 128 150 180
rect 202 128 402 180
rect 454 128 654 180
rect 706 128 846 180
rect 10 122 846 128
<< labels >>
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
port 2 nsew
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
port 3 nsew
flabel metal1 s 762 122 820 138 3 FreeSans 300 90 0 0 BULK
port 4 nsew
flabel metal1 s 183 0 673 66 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 183 740 673 806 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9931810
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9916306
<< end >>
