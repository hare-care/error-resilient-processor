magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 37 41 311 203
rect 37 17 63 41
rect 29 -17 63 17
<< scnmos >>
rect 120 67 150 177
rect 198 67 228 177
<< scpmoshvt >>
rect 106 297 156 497
rect 212 297 262 497
<< ndiff >>
rect 63 133 120 177
rect 63 99 75 133
rect 109 99 120 133
rect 63 67 120 99
rect 150 67 198 177
rect 228 133 285 177
rect 228 99 239 133
rect 273 99 285 133
rect 228 67 285 99
<< pdiff >>
rect 53 485 106 497
rect 53 451 61 485
rect 95 451 106 485
rect 53 417 106 451
rect 53 383 61 417
rect 95 383 106 417
rect 53 297 106 383
rect 156 471 212 497
rect 156 437 167 471
rect 201 437 212 471
rect 156 351 212 437
rect 156 317 167 351
rect 201 317 212 351
rect 156 297 212 317
rect 262 485 340 497
rect 262 451 298 485
rect 332 451 340 485
rect 262 414 340 451
rect 262 380 298 414
rect 332 380 340 414
rect 262 343 340 380
rect 262 309 298 343
rect 332 309 340 343
rect 262 297 340 309
<< ndiffc >>
rect 75 99 109 133
rect 239 99 273 133
<< pdiffc >>
rect 61 451 95 485
rect 61 383 95 417
rect 167 437 201 471
rect 167 317 201 351
rect 298 451 332 485
rect 298 380 332 414
rect 298 309 332 343
<< poly >>
rect 106 497 156 523
rect 212 497 262 523
rect 106 263 156 297
rect 29 249 156 263
rect 29 215 86 249
rect 120 234 156 249
rect 212 234 262 297
rect 120 215 262 234
rect 29 199 262 215
rect 120 177 150 199
rect 198 198 262 199
rect 198 177 228 198
rect 120 41 150 67
rect 198 41 228 67
<< polycont >>
rect 86 215 120 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 45 525 348 527
rect 45 485 111 525
rect 45 451 61 485
rect 95 451 111 485
rect 45 417 111 451
rect 45 383 61 417
rect 95 383 111 417
rect 45 367 111 383
rect 162 471 247 491
rect 162 437 167 471
rect 201 437 247 471
rect 162 351 247 437
rect 29 249 120 333
rect 29 215 86 249
rect 29 199 120 215
rect 162 317 167 351
rect 201 317 247 351
rect 162 150 247 317
rect 288 485 348 525
rect 288 451 298 485
rect 332 451 348 485
rect 288 414 348 451
rect 288 380 298 414
rect 332 380 348 414
rect 288 343 348 380
rect 288 309 298 343
rect 332 309 348 343
rect 288 291 348 309
rect 59 133 125 149
rect 59 99 75 133
rect 109 99 125 133
rect 59 17 125 99
rect 162 133 289 150
rect 162 99 239 133
rect 273 99 289 133
rect 162 63 289 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 213 85 247 119 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 clkinvlp_2
rlabel metal1 s 0 -48 368 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 3336944
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3333354
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
