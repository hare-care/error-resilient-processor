magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -36 679 1160 1471
<< pwell >>
rect 988 25 1090 159
<< psubdiff >>
rect 1014 109 1064 133
rect 1014 75 1022 109
rect 1056 75 1064 109
rect 1014 51 1064 75
<< nsubdiff >>
rect 1014 1339 1064 1363
rect 1014 1305 1022 1339
rect 1056 1305 1064 1339
rect 1014 1281 1064 1305
<< psubdiffcont >>
rect 1022 75 1056 109
<< nsubdiffcont >>
rect 1022 1305 1056 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1124 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 918 1130 952 1397
rect 1022 1339 1056 1397
rect 1022 1289 1056 1305
rect 64 724 98 740
rect 64 674 98 690
rect 490 724 524 1096
rect 490 690 541 724
rect 490 318 524 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 918 17 952 218
rect 1022 109 1056 125
rect 1022 17 1056 75
rect 0 -17 1124 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1694700623
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1694700623
transform 1 0 1014 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1694700623
transform 1 0 1014 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m8_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m8_w2_000_sli_dli_da_p_0
timestamp 1694700623
transform 1 0 54 0 1 51
box -26 -26 932 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m8_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m8_w2_000_sli_dli_da_p_0
timestamp 1694700623
transform 1 0 54 0 1 963
box -59 -56 965 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 524 707 524 707 4 Z
rlabel locali s 562 0 562 0 4 gnd
rlabel locali s 562 1414 562 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1124 1414
string GDS_END 375618
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 373236
<< end >>
