magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 30 -17 64 21
<< locali >>
rect 106 357 309 493
rect 18 199 72 265
rect 18 137 69 199
rect 106 165 140 357
rect 174 199 248 323
rect 282 199 340 323
rect 386 199 445 493
rect 515 199 627 265
rect 103 131 169 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 299 72 527
rect 539 299 627 527
rect 203 131 505 165
rect 203 97 269 131
rect 18 51 269 97
rect 303 17 437 97
rect 471 75 505 131
rect 539 17 627 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 515 199 627 265 6 A1
port 1 nsew signal input
rlabel locali s 386 199 445 493 6 A2
port 2 nsew signal input
rlabel locali s 282 199 340 323 6 A3
port 3 nsew signal input
rlabel locali s 18 137 69 199 6 B1
port 4 nsew signal input
rlabel locali s 18 199 72 265 6 B1
port 4 nsew signal input
rlabel locali s 174 199 248 323 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 131 169 165 6 Y
port 10 nsew signal output
rlabel locali s 106 165 140 357 6 Y
port 10 nsew signal output
rlabel locali s 106 357 309 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1487606
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1480930
<< end >>
