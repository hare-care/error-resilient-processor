magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< obsm2 >>
rect -7432 31006 -987 33506
tri -987 31006 1513 33506 sw
tri -2023 28004 979 31006 ne
rect 979 30504 1513 31006
tri 1513 30504 2015 31006 sw
rect 979 28004 7787 30504
rect -7432 25002 -987 27502
tri -987 25002 1513 27502 sw
tri -2023 22000 979 25002 ne
rect 979 24500 1513 25002
tri 1513 24500 2015 25002 sw
rect 979 22000 7787 24500
rect 19408 -1250 37508 1250
tri -2023 -28004 979 -25002 se
rect 979 -27502 7675 -25002
rect 979 -28004 1513 -27502
tri 1513 -28004 2015 -27502 nw
rect -7544 -30504 -987 -28004
tri -987 -30504 1513 -28004 nw
tri -2023 -34008 979 -31006 se
rect 979 -33506 7675 -31006
rect 979 -34008 1513 -33506
tri 1513 -34008 2015 -33506 nw
rect -7544 -36508 -987 -34008
tri -987 -36508 1513 -34008 nw
<< obsm3 >>
tri -17624 34008 -15124 36508 se
rect -15124 34008 15124 36508
tri -20049 31583 -17624 34008 se
rect -17624 33506 -14590 34008
tri -14590 33506 -14088 34008 nw
tri 14088 33506 14590 34008 ne
rect 14590 33506 15124 34008
tri 15124 33506 18126 36508 sw
rect -17624 32804 -15292 33506
tri -15292 32804 -14590 33506 nw
tri -14583 32804 -13881 33506 se
rect -13881 33286 -2268 33506
tri -2268 33286 -2048 33506 sw
rect -13881 32804 -2048 33286
rect -17624 32095 -16001 32804
tri -16001 32095 -15292 32804 nw
tri -15292 32095 -14583 32804 se
rect -14583 32095 -2048 32804
rect -17624 31583 -16513 32095
tri -16513 31583 -16001 32095 nw
tri -15804 31583 -15292 32095 se
rect -15292 31583 -2048 32095
tri -23307 28325 -20049 31583 se
rect -20049 31327 -16769 31583
tri -16769 31327 -16513 31583 nw
tri -16060 31327 -15804 31583 se
rect -15804 31327 -2048 31583
rect -20049 30679 -17417 31327
tri -17417 30679 -16769 31327 nw
tri -16708 30679 -16060 31327 se
rect -16060 31226 -2048 31327
rect -16060 31006 -2268 31226
tri -2268 31006 -2048 31226 nw
rect -16060 30679 -13172 31006
tri -13172 30679 -12845 31006 nw
rect -20049 29970 -18126 30679
tri -18126 29970 -17417 30679 nw
tri -17417 29970 -16708 30679 se
rect -16708 29970 -13881 30679
tri -13881 29970 -13172 30679 nw
tri -2015 30504 987 33506 se
rect 987 32804 13881 33506
tri 13881 32804 14583 33506 sw
tri 14590 32804 15292 33506 ne
rect 15292 32804 18126 33506
tri 18126 32804 18828 33506 sw
rect 987 32270 14583 32804
tri 14583 32270 15117 32804 sw
tri 15292 32270 15826 32804 ne
rect 15826 32270 18828 32804
tri 18828 32270 19362 32804 sw
rect 987 31561 15117 32270
tri 15117 31561 15826 32270 sw
tri 15826 31561 16535 32270 ne
rect 16535 31561 19362 32270
rect 987 31006 15826 31561
rect 987 30504 1521 31006
tri 1521 30504 2023 31006 nw
tri -13171 29970 -12637 30504 se
rect -12637 30317 1334 30504
tri 1334 30317 1521 30504 nw
rect -12637 29970 706 30317
rect -20049 29268 -18828 29970
tri -18828 29268 -18126 29970 nw
tri -18119 29268 -17417 29970 se
rect -17417 29268 -14583 29970
tri -14583 29268 -13881 29970 nw
tri -13873 29268 -13171 29970 se
rect -13171 29689 706 29970
tri 706 29689 1334 30317 nw
tri 2403 30284 2623 30504 se
rect 2623 30317 12637 30504
tri 12637 30317 12824 30504 sw
tri 12845 30317 13534 31006 ne
rect 13534 30852 15826 31006
tri 15826 30852 16535 31561 sw
tri 16535 30852 17244 31561 ne
rect 17244 30852 19362 31561
rect 13534 30317 16535 30852
rect 2623 30284 12824 30317
rect 2403 29689 12824 30284
tri 12824 29689 13452 30317 sw
tri 13534 29689 14162 30317 ne
rect 14162 30143 16535 30317
tri 16535 30143 17244 30852 sw
tri 17244 30143 17953 30852 ne
rect 17953 30143 19362 30852
rect 14162 29689 17244 30143
rect -13171 29268 -979 29689
rect -20049 28581 -19515 29268
tri -19515 28581 -18828 29268 nw
tri -18806 28581 -18119 29268 se
rect -18119 28581 -15292 29268
rect -20049 28325 -19771 28581
tri -19771 28325 -19515 28581 nw
tri -19062 28325 -18806 28581 se
rect -18806 28559 -15292 28581
tri -15292 28559 -14583 29268 nw
tri -14582 28559 -13873 29268 se
rect -13873 28559 -979 29268
rect -18806 28325 -15999 28559
tri -26309 25323 -23307 28325 se
rect -23307 27852 -20244 28325
tri -20244 27852 -19771 28325 nw
tri -19535 27852 -19062 28325 se
rect -19062 27852 -15999 28325
tri -15999 27852 -15292 28559 nw
tri -15289 27852 -14582 28559 se
rect -14582 28004 -979 28559
tri -979 28004 706 29689 nw
rect 2403 29075 13452 29689
tri 13452 29075 14066 29689 sw
tri 14162 29075 14776 29689 ne
rect 14776 29436 17244 29689
tri 17244 29436 17951 30143 sw
tri 17953 29436 18660 30143 ne
rect 18660 29436 19362 30143
rect 14776 29075 17951 29436
rect 2403 28558 14066 29075
tri 14066 28558 14583 29075 sw
tri 14776 28558 15293 29075 ne
rect 15293 28734 17951 29075
tri 17951 28734 18653 29436 sw
tri 18660 28734 19362 29436 ne
tri 19362 28734 22898 32270 sw
rect 15293 28558 18653 28734
rect 2403 28224 14583 28558
tri 2403 28025 2602 28224 ne
rect 2602 28025 14583 28224
tri 2602 28004 2623 28025 ne
rect 2623 28004 14583 28025
tri 14583 28004 15137 28558 sw
tri 15293 28224 15627 28558 ne
rect 15627 28224 18653 28558
tri 15627 28004 15847 28224 ne
rect 15847 28025 18653 28224
tri 18653 28025 19362 28734 sw
tri 19362 28025 20071 28734 ne
rect 20071 28025 22898 28734
rect 15847 28004 19362 28025
rect -14582 27852 -12103 28004
rect -23307 27143 -20953 27852
tri -20953 27143 -20244 27852 nw
tri -20244 27143 -19535 27852 se
rect -19535 27143 -16708 27852
tri -16708 27143 -15999 27852 nw
tri -15998 27143 -15289 27852 se
rect -15289 27502 -12103 27852
tri -12103 27502 -11601 28004 nw
tri 11601 27502 12103 28004 ne
rect 12103 27502 15137 28004
tri 15137 27502 15639 28004 sw
tri 15847 27502 16349 28004 ne
rect 16349 27502 19362 28004
rect -15289 27143 -12637 27502
rect -23307 26434 -21662 27143
tri -21662 26434 -20953 27143 nw
tri -20953 26434 -20244 27143 se
rect -20244 26434 -17417 27143
tri -17417 26434 -16708 27143 nw
tri -16707 26434 -15998 27143 se
rect -15998 26968 -12637 27143
tri -12637 26968 -12103 27502 nw
tri -11928 26968 -11394 27502 se
rect -11394 27282 -2268 27502
tri -2268 27282 -2048 27502 sw
rect -11394 26968 -2048 27282
rect -15998 26434 -13174 26968
rect -23307 25732 -22364 26434
tri -22364 25732 -21662 26434 nw
tri -21655 25732 -20953 26434 se
rect -20953 25732 -18119 26434
tri -18119 25732 -17417 26434 nw
tri -17409 25732 -16707 26434 se
rect -16707 26431 -13174 26434
tri -13174 26431 -12637 26968 nw
tri -12465 26431 -11928 26968 se
rect -11928 26431 -2048 26968
rect -16707 25732 -13873 26431
tri -13873 25732 -13174 26431 nw
tri -13164 25732 -12465 26431 se
rect -12465 25732 -2048 26431
rect -23307 25323 -23073 25732
tri -29436 22196 -26309 25323 se
rect -26309 25023 -23073 25323
tri -23073 25023 -22364 25732 nw
tri -22364 25023 -21655 25732 se
rect -21655 25023 -18828 25732
tri -18828 25023 -18119 25732 nw
tri -18118 25023 -17409 25732 se
rect -17409 25323 -14282 25732
tri -14282 25323 -13873 25732 nw
tri -13573 25323 -13164 25732 se
rect -13164 25323 -2048 25732
rect -17409 25023 -14583 25323
rect -26309 24316 -23780 25023
tri -23780 24316 -23073 25023 nw
tri -23071 24316 -22364 25023 se
rect -22364 24316 -19535 25023
tri -19535 24316 -18828 25023 nw
tri -18825 24316 -18118 25023 se
rect -18118 25022 -14583 25023
tri -14583 25022 -14282 25323 nw
tri -13874 25022 -13573 25323 se
rect -13573 25222 -2048 25323
rect -13573 25022 -2268 25222
rect -18118 24489 -15116 25022
tri -15116 24489 -14583 25022 nw
tri -14407 24489 -13874 25022 se
rect -13874 25002 -2268 25022
tri -2268 25002 -2048 25222 nw
rect -13874 24489 -10871 25002
tri -10871 24489 -10358 25002 nw
tri -2015 24500 987 27502 se
rect 987 26793 11394 27502
tri 11394 26793 12103 27502 sw
tri 12103 26793 12812 27502 ne
rect 12812 26793 15639 27502
tri 15639 26793 16348 27502 sw
tri 16349 26793 17058 27502 ne
rect 17058 27316 19362 27502
tri 19362 27316 20071 28025 sw
tri 20071 27491 20605 28025 ne
rect 20605 27491 22898 28025
tri 20605 27316 20780 27491 ne
rect 20780 27316 22898 27491
rect 17058 26793 20071 27316
rect 987 26247 12103 26793
tri 12103 26247 12649 26793 sw
tri 12812 26247 13358 26793 ne
rect 13358 26247 16348 26793
tri 16348 26247 16894 26793 sw
tri 17058 26247 17604 26793 ne
rect 17604 26607 20071 26793
tri 20071 26607 20780 27316 sw
tri 20780 26607 21489 27316 ne
rect 21489 26607 22898 27316
rect 17604 26247 20780 26607
rect 987 25538 12649 26247
tri 12649 25538 13358 26247 sw
tri 13358 25538 14067 26247 ne
rect 14067 25538 16894 26247
tri 16894 25538 17603 26247 sw
tri 17604 25538 18313 26247 ne
rect 18313 25900 20780 26247
tri 20780 25900 21487 26607 sw
tri 21489 25900 22196 26607 ne
rect 22196 25900 22898 26607
rect 18313 25538 21487 25900
rect 987 25002 13358 25538
rect 987 24500 1521 25002
tri 1521 24500 2023 25002 nw
tri -10161 24489 -10150 24500 se
rect -10150 24489 1315 24500
rect -18118 24316 -15682 24489
rect -26309 23607 -24489 24316
tri -24489 23607 -23780 24316 nw
tri -23780 23607 -23071 24316 se
rect -23071 24179 -19672 24316
tri -19672 24179 -19535 24316 nw
tri -18962 24179 -18825 24316 se
rect -18825 24179 -15682 24316
rect -23071 23607 -20244 24179
tri -20244 23607 -19672 24179 nw
tri -19534 23607 -18962 24179 se
rect -18962 23923 -15682 24179
tri -15682 23923 -15116 24489 nw
tri -14973 23923 -14407 24489 se
rect -14407 23923 -11437 24489
tri -11437 23923 -10871 24489 nw
tri -10727 23923 -10161 24489 se
rect -10161 24294 1315 24489
tri 1315 24294 1521 24500 nw
rect -10161 23923 706 24294
rect -18962 23607 -16360 23923
rect -26309 22898 -25198 23607
tri -25198 22898 -24489 23607 nw
tri -24489 22898 -23780 23607 se
rect -23780 22898 -20953 23607
tri -20953 22898 -20244 23607 nw
tri -20243 22898 -19534 23607 se
rect -19534 23245 -16360 23607
tri -16360 23245 -15682 23923 nw
tri -15651 23245 -14973 23923 se
rect -14973 23245 -12115 23923
tri -12115 23245 -11437 23923 nw
tri -11405 23245 -10727 23923 se
rect -10727 23685 706 23923
tri 706 23685 1315 24294 nw
tri 2403 24280 2623 24500 se
rect 2623 24294 10150 24500
tri 10150 24294 10356 24500 sw
tri 10358 24294 11066 25002 ne
rect 11066 24829 13358 25002
tri 13358 24829 14067 25538 sw
tri 14067 24829 14776 25538 ne
rect 14776 24829 17603 25538
tri 17603 24829 18312 25538 sw
tri 18313 24829 19022 25538 ne
rect 19022 25198 21487 25538
tri 21487 25198 22189 25900 sw
tri 22196 25198 22898 25900 ne
tri 22898 25198 26434 28734 sw
rect 19022 24829 22189 25198
rect 11066 24294 14067 24829
tri 14067 24294 14602 24829 sw
tri 14776 24294 15311 24829 ne
rect 15311 24489 18312 24829
tri 18312 24489 18652 24829 sw
tri 19022 24489 19362 24829 ne
rect 19362 24489 22189 24829
tri 22189 24489 22898 25198 sw
tri 22898 24489 23607 25198 ne
rect 23607 24489 26434 25198
rect 15311 24294 18652 24489
rect 2623 24280 10356 24294
rect 2403 23685 10356 24280
tri 10356 23685 10965 24294 sw
tri 11066 23685 11675 24294 ne
rect 11675 23966 14602 24294
tri 14602 23966 14930 24294 sw
tri 15311 23966 15639 24294 ne
rect 15639 23966 18652 24294
rect 11675 23685 14930 23966
rect -10727 23245 92 23685
rect -19534 22898 -17028 23245
rect -26309 22196 -25900 22898
tri -25900 22196 -25198 22898 nw
tri -25191 22196 -24489 22898 se
rect -24489 22196 -21655 22898
tri -21655 22196 -20953 22898 nw
tri -20945 22196 -20243 22898 se
rect -20243 22577 -17028 22898
tri -17028 22577 -16360 23245 nw
tri -16319 22577 -15651 23245 se
rect -15651 22577 -12783 23245
tri -12783 22577 -12115 23245 nw
tri -12073 22577 -11405 23245 se
rect -11405 23071 92 23245
tri 92 23071 706 23685 nw
rect 2403 23071 10965 23685
tri 10965 23071 11579 23685 sw
tri 11675 23432 11928 23685 ne
rect 11928 23432 14930 23685
tri 14930 23432 15464 23966 sw
tri 15639 23432 16173 23966 ne
rect 16173 23780 18652 23966
tri 18652 23780 19361 24489 sw
tri 19362 23780 20071 24489 ne
rect 20071 23780 22898 24489
tri 22898 23780 23607 24489 sw
tri 23607 23955 24141 24489 ne
rect 24141 23955 26434 24489
tri 24141 23780 24316 23955 ne
rect 24316 23780 26434 23955
rect 16173 23432 19361 23780
tri 11928 23071 12289 23432 ne
rect 12289 23071 15464 23432
rect -11405 22577 -979 23071
rect -20243 22196 -17603 22577
tri -32972 18660 -29436 22196 se
rect -29436 21487 -26609 22196
tri -26609 21487 -25900 22196 nw
tri -25900 21487 -25191 22196 se
rect -25191 21487 -22364 22196
tri -22364 21487 -21655 22196 nw
tri -21654 21487 -20945 22196 se
rect -20945 22002 -17603 22196
tri -17603 22002 -17028 22577 nw
tri -16894 22002 -16319 22577 se
rect -16319 22002 -13358 22577
tri -13358 22002 -12783 22577 nw
rect -20945 21487 -18119 22002
rect -29436 20780 -27316 21487
tri -27316 20780 -26609 21487 nw
tri -26607 20780 -25900 21487 se
rect -25900 20780 -23071 21487
tri -23071 20780 -22364 21487 nw
tri -22361 20780 -21654 21487 se
rect -21654 21486 -18119 21487
tri -18119 21486 -17603 22002 nw
tri -17410 21486 -16894 22002 se
rect -16894 21487 -13873 22002
tri -13873 21487 -13358 22002 nw
tri -12650 22000 -12073 22577 se
rect -12073 22000 -979 22577
tri -979 22000 92 23071 nw
rect 2403 22364 11579 23071
tri 11579 22364 12286 23071 sw
tri 12289 22898 12462 23071 ne
rect 12462 22898 15464 23071
tri 15464 22898 15998 23432 sw
tri 16173 22898 16707 23432 ne
rect 16707 23245 19361 23432
tri 19361 23245 19896 23780 sw
tri 20071 23245 20606 23780 ne
rect 20606 23245 23607 23780
rect 16707 22898 19896 23245
rect 2403 22220 12286 22364
tri 12286 22220 12430 22364 sw
tri 12462 22220 13140 22898 ne
rect 13140 22220 15998 22898
tri 2403 22000 2623 22220 ne
rect 2623 22000 12430 22220
tri 12430 22000 12650 22220 sw
tri 13140 22196 13164 22220 ne
rect 13164 22196 15998 22220
tri 15998 22196 16700 22898 sw
tri 16707 22196 17409 22898 ne
rect 17409 22535 19896 22898
tri 19896 22535 20606 23245 sw
tri 20606 22711 21140 23245 ne
rect 21140 23071 23607 23245
tri 23607 23071 24316 23780 sw
tri 24316 23071 25025 23780 ne
rect 25025 23071 26434 23780
rect 21140 22711 24316 23071
rect 17409 22196 20606 22535
tri 13164 22000 13360 22196 ne
rect 13360 22002 16700 22196
tri 16700 22002 16894 22196 sw
tri 17409 22002 17603 22196 ne
rect 17603 22002 20606 22196
tri 20606 22002 21139 22535 sw
tri 21140 22002 21849 22711 ne
rect 21849 22364 24316 22711
tri 24316 22364 25023 23071 sw
tri 25025 22364 25732 23071 ne
rect 25732 22364 26434 23071
rect 21849 22002 25023 22364
rect 13360 22000 16894 22002
tri -13163 21487 -12650 22000 se
rect -12650 21487 -12454 22000
rect -16894 21486 -14221 21487
rect -21654 20953 -18652 21486
tri -18652 20953 -18119 21486 nw
tri -17943 20953 -17410 21486 se
rect -17410 21139 -14221 21486
tri -14221 21139 -13873 21487 nw
tri -13511 21139 -13163 21487 se
rect -13163 21139 -12454 21487
rect -17410 20953 -14930 21139
rect -21654 20780 -19175 20953
rect -29436 20071 -28025 20780
tri -28025 20071 -27316 20780 nw
tri -27316 20071 -26607 20780 se
rect -26607 20071 -23780 20780
tri -23780 20071 -23071 20780 nw
tri -23070 20071 -22361 20780 se
rect -22361 20430 -19175 20780
tri -19175 20430 -18652 20953 nw
tri -18466 20430 -17943 20953 se
rect -17943 20430 -14930 20953
tri -14930 20430 -14221 21139 nw
tri -14220 20430 -13511 21139 se
rect -13511 20430 -12454 21139
rect -22361 20071 -19709 20430
rect -29436 19362 -28734 20071
tri -28734 19362 -28025 20071 nw
tri -28025 19362 -27316 20071 se
rect -27316 19362 -24489 20071
tri -24489 19362 -23780 20071 nw
tri -23779 19362 -23070 20071 se
rect -23070 19896 -19709 20071
tri -19709 19896 -19175 20430 nw
tri -19000 19896 -18466 20430 se
rect -18466 19896 -15464 20430
tri -15464 19896 -14930 20430 nw
tri -14754 19896 -14220 20430 se
rect -14220 19896 -12454 20430
rect -23070 19362 -20243 19896
tri -20243 19362 -19709 19896 nw
tri -19534 19362 -19000 19896 se
rect -19000 19362 -15998 19896
tri -15998 19362 -15464 19896 nw
tri -15288 19362 -14754 19896 se
rect -14754 19362 -12454 19896
tri -29436 18660 -28734 19362 nw
tri -28727 18660 -28025 19362 se
rect -28025 18660 -25191 19362
tri -25191 18660 -24489 19362 nw
tri -24481 18660 -23779 19362 se
rect -23779 18660 -20945 19362
tri -20945 18660 -20243 19362 nw
tri -20236 18660 -19534 19362 se
rect -19534 18660 -16700 19362
tri -16700 18660 -15998 19362 nw
tri -15990 18660 -15288 19362 se
rect -15288 18660 -12454 19362
tri -12454 18660 -9114 22000 nw
tri -36508 15124 -32972 18660 se
rect -32972 17951 -30145 18660
tri -30145 17951 -29436 18660 nw
tri -29436 17951 -28727 18660 se
rect -28727 17951 -25900 18660
tri -25900 17951 -25191 18660 nw
tri -25190 17951 -24481 18660 se
rect -24481 17951 -21654 18660
tri -21654 17951 -20945 18660 nw
tri -20945 17951 -20236 18660 se
rect -20236 17951 -17409 18660
tri -17409 17951 -16700 18660 nw
tri -16699 17951 -15990 18660 se
rect -15990 17951 -15288 18660
rect -32972 17244 -30852 17951
tri -30852 17244 -30145 17951 nw
tri -30143 17244 -29436 17951 se
rect -29436 17244 -26607 17951
tri -26607 17244 -25900 17951 nw
tri -25897 17244 -25190 17951 se
rect -25190 17417 -22188 17951
tri -22188 17417 -21654 17951 nw
tri -21479 17417 -20945 17951 se
rect -20945 17603 -17757 17951
tri -17757 17603 -17409 17951 nw
tri -17047 17603 -16699 17951 se
rect -16699 17603 -15288 17951
rect -20945 17417 -18466 17603
rect -25190 17244 -22711 17417
rect -32972 16535 -31561 17244
tri -31561 16535 -30852 17244 nw
tri -30852 16535 -30143 17244 se
rect -30143 16535 -27316 17244
tri -27316 16535 -26607 17244 nw
tri -26606 16535 -25897 17244 se
rect -25897 16894 -22711 17244
tri -22711 16894 -22188 17417 nw
tri -22002 16894 -21479 17417 se
rect -21479 16894 -18466 17417
tri -18466 16894 -17757 17603 nw
tri -17756 16894 -17047 17603 se
rect -17047 16894 -15288 17603
rect -25897 16535 -23245 16894
rect -32972 15826 -32270 16535
tri -32270 15826 -31561 16535 nw
tri -31561 15826 -30852 16535 se
rect -30852 15826 -28025 16535
tri -28025 15826 -27316 16535 nw
tri -27315 15826 -26606 16535 se
rect -26606 16360 -23245 16535
tri -23245 16360 -22711 16894 nw
tri -22536 16360 -22002 16894 se
rect -22002 16360 -19000 16894
tri -19000 16360 -18466 16894 nw
tri -18290 16360 -17756 16894 se
rect -17756 16360 -15288 16894
rect -26606 15826 -23779 16360
tri -23779 15826 -23245 16360 nw
tri -23070 15826 -22536 16360 se
rect -22536 15826 -19534 16360
tri -19534 15826 -19000 16360 nw
tri -18824 15826 -18290 16360 se
rect -18290 15826 -15288 16360
tri -15288 15826 -12454 18660 nw
tri 9114 18466 12648 22000 ne
rect 12648 21468 12650 22000
tri 12650 21468 13182 22000 sw
tri 13360 21468 13892 22000 ne
rect 13892 21468 16894 22000
rect 12648 20758 13182 21468
tri 13182 20758 13892 21468 sw
tri 13892 20758 14602 21468 ne
rect 14602 21293 16894 21468
tri 16894 21293 17603 22002 sw
tri 17603 21293 18312 22002 ne
rect 18312 21293 21139 22002
tri 21139 21293 21848 22002 sw
tri 21849 21293 22558 22002 ne
rect 22558 21662 25023 22002
tri 25023 21662 25725 22364 sw
tri 25732 21662 26434 22364 ne
tri 26434 21662 29970 25198 sw
rect 22558 21293 25725 21662
rect 14602 20758 17603 21293
tri 17603 20758 18138 21293 sw
tri 18312 20758 18847 21293 ne
rect 18847 20953 21848 21293
tri 21848 20953 22188 21293 sw
tri 22558 20953 22898 21293 ne
rect 22898 20953 25725 21293
tri 25725 20953 26434 21662 sw
tri 26434 20953 27143 21662 ne
rect 27143 20953 29970 21662
rect 18847 20758 22188 20953
rect 12648 20048 13892 20758
tri 13892 20048 14602 20758 sw
tri 14602 20048 15312 20758 ne
rect 15312 20244 18138 20758
tri 18138 20244 18652 20758 sw
tri 18847 20244 19361 20758 ne
rect 19361 20244 22188 20758
tri 22188 20244 22897 20953 sw
tri 22898 20244 23607 20953 ne
rect 23607 20244 26434 20953
tri 26434 20244 27143 20953 sw
tri 27143 20419 27677 20953 ne
rect 27677 20419 29970 20953
tri 27677 20244 27852 20419 ne
rect 27852 20244 29970 20419
rect 15312 20048 18652 20244
rect 12648 19362 14602 20048
tri 14602 19362 15288 20048 sw
tri 15312 19362 15998 20048 ne
rect 15998 19709 18652 20048
tri 18652 19709 19187 20244 sw
tri 19361 19709 19896 20244 ne
rect 19896 19709 22897 20244
tri 22897 19709 23432 20244 sw
tri 23607 19709 24142 20244 ne
rect 24142 19709 27143 20244
rect 15998 19362 19187 19709
rect 12648 18660 15288 19362
tri 15288 18660 15990 19362 sw
tri 15998 18660 16700 19362 ne
rect 16700 19175 19187 19362
tri 19187 19175 19721 19709 sw
tri 19896 19175 20430 19709 ne
rect 20430 19175 23432 19709
rect 16700 18660 19721 19175
rect 12648 18466 15990 18660
tri 15990 18466 16184 18660 sw
tri 16700 18466 16894 18660 ne
rect 16894 18466 19721 18660
tri 19721 18466 20430 19175 sw
tri 20430 18660 20945 19175 ne
rect 20945 18999 23432 19175
tri 23432 18999 24142 19709 sw
tri 24142 19175 24676 19709 ne
rect 24676 19535 27143 19709
tri 27143 19535 27852 20244 sw
tri 27852 19535 28561 20244 ne
rect 28561 19535 29970 20244
rect 24676 19175 27852 19535
rect 20945 18660 24142 18999
tri 20945 18466 21139 18660 ne
rect 21139 18466 24142 18660
tri 24142 18466 24675 18999 sw
tri 24676 18466 25385 19175 ne
rect 25385 18828 27852 19175
tri 27852 18828 28559 19535 sw
tri 28561 18828 29268 19535 ne
rect 29268 18828 29970 19535
rect 25385 18466 28559 18828
tri -32972 15124 -32270 15826 nw
tri -32263 15124 -31561 15826 se
rect -31561 15124 -28727 15826
tri -28727 15124 -28025 15826 nw
tri -28017 15124 -27315 15826 se
rect -27315 15124 -24481 15826
tri -24481 15124 -23779 15826 nw
tri -23772 15124 -23070 15826 se
rect -23070 15124 -20236 15826
tri -20236 15124 -19534 15826 nw
tri -19526 15124 -18824 15826 se
rect -18824 15124 -18477 15826
rect -36508 14590 -33506 15124
tri -33506 14590 -32972 15124 nw
tri -32797 14590 -32263 15124 se
rect -32263 14590 -29261 15124
tri -29261 14590 -28727 15124 nw
tri -28551 14590 -28017 15124 se
rect -28017 14590 -25190 15124
rect -36508 -14590 -34008 14590
tri -34008 14088 -33506 14590 nw
tri -33506 13881 -32797 14590 se
rect -32797 14088 -29763 14590
tri -29763 14088 -29261 14590 nw
tri -29053 14088 -28551 14590 se
rect -28551 14415 -25190 14590
tri -25190 14415 -24481 15124 nw
tri -24481 14415 -23772 15124 se
rect -23772 14415 -20945 15124
tri -20945 14415 -20236 15124 nw
tri -20235 14415 -19526 15124 se
rect -19526 14415 -18477 15124
rect -28551 14088 -25517 14415
tri -25517 14088 -25190 14415 nw
tri -24808 14088 -24481 14415 se
rect -24481 14088 -21293 14415
rect -32797 13881 -30317 14088
rect -33506 13534 -30317 13881
tri -30317 13534 -29763 14088 nw
tri -29607 13534 -29053 14088 se
rect -29053 13534 -26071 14088
tri -26071 13534 -25517 14088 nw
tri -25362 13534 -24808 14088 se
rect -24808 14067 -21293 14088
tri -21293 14067 -20945 14415 nw
tri -20583 14067 -20235 14415 se
rect -20235 14067 -18477 14415
rect -24808 13534 -22002 14067
rect -33506 -13347 -31006 13534
tri -31006 12845 -30317 13534 nw
tri -30296 12845 -29607 13534 se
rect -29607 12845 -26760 13534
tri -26760 12845 -26071 13534 nw
tri -26051 12845 -25362 13534 se
rect -25362 13358 -22002 13534
tri -22002 13358 -21293 14067 nw
tri -21292 13358 -20583 14067 se
rect -20583 13358 -18477 14067
rect -25362 12845 -22536 13358
tri -30504 12637 -30296 12845 se
rect -30296 12637 -26968 12845
tri -26968 12637 -26760 12845 nw
tri -26259 12637 -26051 12845 se
rect -26051 12824 -22536 12845
tri -22536 12824 -22002 13358 nw
tri -21826 12824 -21292 13358 se
rect -21292 12824 -18477 13358
rect -26051 12637 -22723 12824
tri -22723 12637 -22536 12824 nw
tri -22013 12637 -21826 12824 se
rect -21826 12637 -18477 12824
tri -18477 12637 -15288 15826 nw
tri 12648 14930 16184 18466 ne
tri 16184 17932 16718 18466 sw
tri 16894 17932 17428 18466 ne
rect 17428 17932 20430 18466
rect 16184 17222 16718 17932
tri 16718 17222 17428 17932 sw
tri 17428 17222 18138 17932 ne
rect 18138 17757 20430 17932
tri 20430 17757 21139 18466 sw
tri 21139 17757 21848 18466 ne
rect 21848 17757 24675 18466
tri 24675 17757 25384 18466 sw
tri 25385 17757 26094 18466 ne
rect 26094 18126 28559 18466
tri 28559 18126 29261 18828 sw
tri 29268 18126 29970 18828 ne
tri 29970 18126 33506 21662 sw
rect 26094 17757 29261 18126
rect 18138 17222 21139 17757
tri 21139 17222 21674 17757 sw
tri 21848 17222 22383 17757 ne
rect 22383 17417 25384 17757
tri 25384 17417 25724 17757 sw
tri 26094 17417 26434 17757 ne
rect 26434 17417 29261 17757
tri 29261 17417 29970 18126 sw
tri 29970 17417 30679 18126 ne
rect 30679 17417 33506 18126
rect 22383 17222 25724 17417
rect 16184 16512 17428 17222
tri 17428 16512 18138 17222 sw
tri 18138 16512 18848 17222 ne
rect 18848 16708 21674 17222
tri 21674 16708 22188 17222 sw
tri 22383 16708 22897 17222 ne
rect 22897 16708 25724 17222
tri 25724 16708 26433 17417 sw
tri 26434 16708 27143 17417 ne
rect 27143 16708 29970 17417
tri 29970 16708 30679 17417 sw
tri 30679 16883 31213 17417 ne
rect 31213 16883 33506 17417
tri 31213 16708 31388 16883 ne
rect 31388 16708 33506 16883
rect 18848 16512 22188 16708
rect 16184 15826 18138 16512
tri 18138 15826 18824 16512 sw
tri 18848 15826 19534 16512 ne
rect 19534 16173 22188 16512
tri 22188 16173 22723 16708 sw
tri 22897 16173 23432 16708 ne
rect 23432 16173 26433 16708
tri 26433 16173 26968 16708 sw
tri 27143 16173 27678 16708 ne
rect 27678 16173 30679 16708
rect 19534 15826 22723 16173
rect 16184 15124 18824 15826
tri 18824 15124 19526 15826 sw
tri 19534 15124 20236 15826 ne
rect 20236 15639 22723 15826
tri 22723 15639 23257 16173 sw
tri 23432 15639 23966 16173 ne
rect 23966 15639 26968 16173
rect 20236 15124 23257 15639
rect 16184 14930 19526 15124
tri 19526 14930 19720 15124 sw
tri 20236 14930 20430 15124 ne
rect 20430 14930 23257 15124
tri 23257 14930 23966 15639 sw
tri 23966 15124 24481 15639 ne
rect 24481 15463 26968 15639
tri 26968 15463 27678 16173 sw
tri 27678 15639 28212 16173 ne
rect 28212 15999 30679 16173
tri 30679 15999 31388 16708 sw
tri 31388 15999 32097 16708 ne
rect 32097 15999 33506 16708
rect 28212 15639 31388 15999
rect 24481 15124 27678 15463
tri 24481 14930 24675 15124 ne
rect 24675 14930 27678 15124
tri 27678 14930 28211 15463 sw
tri 28212 14930 28921 15639 ne
rect 28921 15292 31388 15639
tri 31388 15292 32095 15999 sw
tri 32097 15292 32804 15999 ne
rect 32804 15292 33506 15999
rect 28921 14930 32095 15292
rect -30504 12103 -27502 12637
tri -27502 12103 -26968 12637 nw
tri -26793 12103 -26259 12637 se
rect -26259 12103 -23257 12637
tri -23257 12103 -22723 12637 nw
tri -22547 12103 -22013 12637 se
rect -22013 12103 -19187 12637
rect -30504 -12103 -28004 12103
tri -28004 11601 -27502 12103 nw
tri -27502 11394 -26793 12103 se
rect -26793 11601 -23759 12103
tri -23759 11601 -23257 12103 nw
tri -23049 11601 -22547 12103 se
rect -22547 11927 -19187 12103
tri -19187 11927 -18477 12637 nw
rect -22547 11601 -22000 11927
rect -26793 11394 -24294 11601
rect -27502 11066 -24294 11394
tri -24294 11066 -23759 11601 nw
tri -23584 11066 -23049 11601 se
rect -23049 11066 -22000 11601
rect -27502 -10860 -25002 11066
tri -25002 10358 -24294 11066 nw
tri -24292 10358 -23584 11066 se
rect -23584 10358 -22000 11066
tri -24500 10150 -24292 10358 se
rect -24292 10150 -22000 10358
rect -24500 1250 -22000 10150
tri -22000 9114 -19187 11927 nw
tri 16184 11394 19720 14930 ne
tri 19720 14396 20254 14930 sw
tri 20430 14396 20964 14930 ne
rect 20964 14396 23966 14930
rect 19720 13686 20254 14396
tri 20254 13686 20964 14396 sw
tri 20964 13686 21674 14396 ne
rect 21674 14221 23966 14396
tri 23966 14221 24675 14930 sw
tri 24675 14221 25384 14930 ne
rect 25384 14221 28211 14930
tri 28211 14221 28920 14930 sw
tri 28921 14221 29630 14930 ne
rect 29630 14590 32095 14930
tri 32095 14590 32797 15292 sw
tri 32804 14590 33506 15292 ne
tri 33506 15124 36508 18126 sw
rect 33506 14590 36508 15124
rect 29630 14221 32797 14590
rect 21674 13686 24675 14221
tri 24675 13686 25210 14221 sw
tri 25384 13686 25919 14221 ne
rect 25919 13881 28920 14221
tri 28920 13881 29260 14221 sw
tri 29630 13881 29970 14221 ne
rect 29970 13881 32797 14221
tri 32797 13881 33506 14590 sw
tri 33506 14088 34008 14590 ne
rect 25919 13686 29260 13881
rect 19720 12976 20964 13686
tri 20964 12976 21674 13686 sw
tri 21674 12976 22384 13686 ne
rect 22384 13172 25210 13686
tri 25210 13172 25724 13686 sw
tri 25919 13172 26433 13686 ne
rect 26433 13172 29260 13686
tri 29260 13172 29969 13881 sw
tri 29970 13172 30679 13881 ne
rect 30679 13172 33506 13881
rect 22384 12976 25724 13172
rect 19720 12637 21674 12976
tri 21674 12637 22013 12976 sw
tri 22384 12637 22723 12976 ne
rect 22723 12637 25724 12976
tri 25724 12637 26259 13172 sw
tri 26433 12637 26968 13172 ne
rect 26968 12637 29969 13172
tri 29969 12637 30504 13172 sw
tri 30679 12845 31006 13172 ne
rect 19720 11927 22013 12637
tri 22013 11927 22723 12637 sw
tri 22723 11927 23433 12637 ne
rect 23433 12103 26259 12637
tri 26259 12103 26793 12637 sw
tri 26968 12103 27502 12637 ne
rect 27502 12103 30504 12637
rect 23433 11927 26793 12103
rect 19720 11394 22723 11927
tri 22723 11394 23256 11927 sw
tri 23433 11601 23759 11927 ne
rect 23759 11601 26793 11927
tri 23759 11394 23966 11601 ne
rect 23966 11394 26793 11601
tri 26793 11394 27502 12103 sw
tri 27502 11601 28004 12103 ne
tri 19720 9114 22000 11394 ne
rect 22000 10860 23256 11394
tri 23256 10860 23790 11394 sw
tri 23966 10860 24500 11394 ne
rect 24500 10860 27502 11394
rect 22000 10150 23790 10860
tri 23790 10150 24500 10860 sw
tri 24500 10358 25002 10860 ne
rect -24500 -1250 21000 1250
rect -24500 -10150 -22000 -1250
tri -25002 -10860 -24500 -10358 sw
tri -24500 -10860 -23790 -10150 ne
rect -23790 -10860 -22000 -10150
rect -27502 -11394 -24500 -10860
tri -24500 -11394 -23966 -10860 sw
tri -23790 -11394 -23256 -10860 ne
rect -23256 -11394 -22000 -10860
tri -28004 -12103 -27502 -11601 sw
tri -27502 -12103 -26793 -11394 ne
rect -26793 -12103 -23966 -11394
tri -23966 -12103 -23257 -11394 sw
tri -23256 -12103 -22547 -11394 ne
rect -22547 -12103 -22000 -11394
rect -30504 -12637 -27502 -12103
tri -27502 -12637 -26968 -12103 sw
tri -26793 -12637 -26259 -12103 ne
rect -26259 -12637 -23257 -12103
tri -23257 -12637 -22723 -12103 sw
tri -22547 -12637 -22013 -12103 ne
rect -22013 -12637 -22000 -12103
tri -22000 -12637 -18477 -9114 sw
tri 18477 -12637 22000 -9114 se
rect 22000 -10150 24500 10150
rect 22000 -10358 24292 -10150
tri 24292 -10358 24500 -10150 nw
rect 22000 -11066 23584 -10358
tri 23584 -11066 24292 -10358 nw
tri 24294 -11066 25002 -10358 se
rect 25002 -11066 27502 10860
rect 22000 -11601 23049 -11066
tri 23049 -11601 23584 -11066 nw
tri 23759 -11601 24294 -11066 se
rect 24294 -11394 27502 -11066
rect 24294 -11601 26793 -11394
rect 22000 -11927 22723 -11601
tri 22723 -11927 23049 -11601 nw
tri 23433 -11927 23759 -11601 se
rect 23759 -11927 26793 -11601
rect 22000 -12637 22013 -11927
tri 22013 -12637 22723 -11927 nw
tri 22723 -12637 23433 -11927 se
rect 23433 -12103 26793 -11927
tri 26793 -12103 27502 -11394 nw
tri 27502 -12103 28004 -11601 se
rect 28004 -12103 30504 12103
rect 23433 -12637 26259 -12103
tri 26259 -12637 26793 -12103 nw
tri 26968 -12637 27502 -12103 se
rect 27502 -12637 30504 -12103
tri -31006 -13347 -30504 -12845 sw
tri -30504 -13347 -29794 -12637 ne
rect -29794 -13172 -26968 -12637
tri -26968 -13172 -26433 -12637 sw
tri -26259 -13172 -25724 -12637 ne
rect -25724 -13172 -22723 -12637
tri -22723 -13172 -22188 -12637 sw
tri -22013 -13172 -21478 -12637 ne
rect -21478 -13172 -18477 -12637
rect -29794 -13347 -26433 -13172
rect -33506 -13881 -30504 -13347
tri -30504 -13881 -29970 -13347 sw
tri -29794 -13881 -29260 -13347 ne
rect -29260 -13881 -26433 -13347
tri -26433 -13881 -25724 -13172 sw
tri -25724 -13881 -25015 -13172 ne
rect -25015 -13881 -22188 -13172
tri -22188 -13881 -21479 -13172 sw
tri -21478 -13881 -20769 -13172 ne
rect -20769 -13881 -18477 -13172
tri -34008 -14590 -33506 -14088 sw
tri -33506 -14590 -32797 -13881 ne
rect -32797 -14590 -29970 -13881
tri -29970 -14590 -29261 -13881 sw
tri -29260 -14590 -28551 -13881 ne
rect -28551 -14414 -25724 -13881
tri -25724 -14414 -25191 -13881 sw
tri -25015 -14414 -24482 -13881 ne
rect -24482 -14396 -21479 -13881
tri -21479 -14396 -20964 -13881 sw
tri -20769 -14396 -20254 -13881 ne
rect -20254 -14396 -18477 -13881
rect -24482 -14414 -20964 -14396
rect -28551 -14590 -25191 -14414
rect -36508 -15124 -33506 -14590
tri -36508 -17417 -34215 -15124 ne
rect -34215 -15292 -33506 -15124
tri -33506 -15292 -32804 -14590 sw
tri -32797 -15292 -32095 -14590 ne
rect -32095 -15292 -29261 -14590
tri -29261 -15292 -28559 -14590 sw
tri -28551 -15292 -27849 -14590 ne
rect -27849 -14930 -25191 -14590
tri -25191 -14930 -24675 -14414 sw
tri -24482 -14930 -23966 -14414 ne
rect -23966 -14930 -20964 -14414
tri -20964 -14930 -20430 -14396 sw
tri -20254 -14930 -19720 -14396 ne
rect -19720 -14930 -18477 -14396
rect -27849 -15292 -24675 -14930
rect -34215 -16001 -32804 -15292
tri -32804 -16001 -32095 -15292 sw
tri -32095 -16001 -31386 -15292 ne
rect -31386 -16001 -28559 -15292
tri -28559 -16001 -27850 -15292 sw
tri -27849 -16001 -27140 -15292 ne
rect -27140 -15639 -24675 -15292
tri -24675 -15639 -23966 -14930 sw
tri -23966 -15639 -23257 -14930 ne
rect -23257 -15639 -20430 -14930
tri -20430 -15639 -19721 -14930 sw
tri -19720 -15639 -19011 -14930 ne
rect -19011 -15639 -18477 -14930
rect -27140 -16001 -23966 -15639
rect -34215 -16708 -32095 -16001
tri -32095 -16708 -31388 -16001 sw
tri -31386 -16708 -30679 -16001 ne
rect -30679 -16708 -27850 -16001
tri -27850 -16708 -27143 -16001 sw
tri -27140 -16708 -26433 -16001 ne
rect -26433 -16173 -23966 -16001
tri -23966 -16173 -23432 -15639 sw
tri -23257 -16173 -22723 -15639 ne
rect -22723 -16173 -19721 -15639
tri -19721 -16173 -19187 -15639 sw
tri -19011 -16173 -18477 -15639 ne
tri -18477 -16173 -14941 -12637 sw
tri 15288 -15826 18477 -12637 se
rect 18477 -12845 21805 -12637
tri 21805 -12845 22013 -12637 nw
tri 22515 -12845 22723 -12637 se
rect 22723 -12845 26051 -12637
tri 26051 -12845 26259 -12637 nw
tri 26760 -12845 26968 -12637 se
rect 26968 -12845 30296 -12637
tri 30296 -12845 30504 -12637 nw
rect 18477 -13358 21292 -12845
tri 21292 -13358 21805 -12845 nw
tri 22002 -13358 22515 -12845 se
rect 22515 -13358 25538 -12845
tri 25538 -13358 26051 -12845 nw
tri 26247 -13358 26760 -12845 se
rect 26760 -13358 29783 -12845
tri 29783 -13358 30296 -12845 nw
tri 30493 -13358 31006 -12845 se
rect 31006 -13358 33506 13172
rect 34008 5500 36508 14590
rect 34008 3000 37508 5500
rect 18477 -13892 20758 -13358
tri 20758 -13892 21292 -13358 nw
tri 21468 -13892 22002 -13358 se
rect 22002 -13892 25004 -13358
tri 25004 -13892 25538 -13358 nw
tri 25713 -13892 26247 -13358 se
rect 26247 -13892 29074 -13358
rect 18477 -14602 20048 -13892
tri 20048 -14602 20758 -13892 nw
tri 20758 -14602 21468 -13892 se
rect 21468 -14088 24808 -13892
tri 24808 -14088 25004 -13892 nw
tri 25517 -14088 25713 -13892 se
rect 25713 -14067 29074 -13892
tri 29074 -14067 29783 -13358 nw
tri 29784 -14067 30493 -13358 se
rect 30493 -13881 33506 -13358
rect 30493 -14067 32797 -13881
rect 25713 -14088 28726 -14067
rect 21468 -14602 24294 -14088
tri 24294 -14602 24808 -14088 nw
tri 25003 -14602 25517 -14088 se
rect 25517 -14415 28726 -14088
tri 28726 -14415 29074 -14067 nw
tri 29436 -14415 29784 -14067 se
rect 29784 -14415 32797 -14067
rect 25517 -14602 28017 -14415
rect 18477 -15292 19358 -14602
tri 19358 -15292 20048 -14602 nw
tri 20068 -15292 20758 -14602 se
rect 20758 -15292 23604 -14602
tri 23604 -15292 24294 -14602 nw
tri 24313 -15292 25003 -14602 se
rect 25003 -15124 28017 -14602
tri 28017 -15124 28726 -14415 nw
tri 28727 -15124 29436 -14415 se
rect 29436 -14590 32797 -14415
tri 32797 -14590 33506 -13881 nw
rect 34008 -5500 37508 -3000
tri 33506 -14590 34008 -14088 se
rect 34008 -14590 36508 -5500
rect 29436 -15124 32263 -14590
tri 32263 -15124 32797 -14590 nw
tri 32972 -15124 33506 -14590 se
rect 33506 -15124 36508 -14590
rect 25003 -15292 27315 -15124
rect 18477 -15826 18824 -15292
tri 18824 -15826 19358 -15292 nw
tri 19534 -15826 20068 -15292 se
rect 20068 -15826 23070 -15292
tri 23070 -15826 23604 -15292 nw
tri 23779 -15826 24313 -15292 se
rect 24313 -15826 27315 -15292
tri 27315 -15826 28017 -15124 nw
tri 28025 -15826 28727 -15124 se
rect 28727 -15826 31561 -15124
tri 31561 -15826 32263 -15124 nw
tri 32270 -15826 32972 -15124 se
rect 32972 -15826 33513 -15124
rect -26433 -16708 -23432 -16173
tri -23432 -16708 -22897 -16173 sw
tri -22723 -16708 -22188 -16173 ne
rect -22188 -16708 -19187 -16173
tri -19187 -16708 -18652 -16173 sw
tri -18477 -16708 -17942 -16173 ne
rect -17942 -16708 -14941 -16173
rect -34215 -17417 -31388 -16708
tri -31388 -17417 -30679 -16708 sw
tri -30679 -17417 -29970 -16708 ne
rect -29970 -17417 -27143 -16708
tri -27143 -17417 -26434 -16708 sw
tri -26433 -17417 -25724 -16708 ne
rect -25724 -17417 -22897 -16708
tri -22897 -17417 -22188 -16708 sw
tri -22188 -17417 -21479 -16708 ne
rect -21479 -17417 -18652 -16708
tri -18652 -17417 -17943 -16708 sw
tri -17942 -17417 -17233 -16708 ne
rect -17233 -17417 -14941 -16708
tri -34215 -20953 -30679 -17417 ne
tri -30679 -18126 -29970 -17417 sw
tri -29970 -18126 -29261 -17417 ne
rect -29261 -18126 -26434 -17417
tri -26434 -18126 -25725 -17417 sw
tri -25724 -18126 -25015 -17417 ne
rect -25015 -17950 -22188 -17417
tri -22188 -17950 -21655 -17417 sw
tri -21479 -17950 -20946 -17417 ne
rect -20946 -17932 -17943 -17417
tri -17943 -17932 -17428 -17417 sw
tri -17233 -17932 -16718 -17417 ne
rect -16718 -17932 -14941 -17417
rect -20946 -17950 -17428 -17932
rect -25015 -18126 -21655 -17950
rect -30679 -18828 -29970 -18126
tri -29970 -18828 -29268 -18126 sw
tri -29261 -18828 -28559 -18126 ne
rect -28559 -18828 -25725 -18126
tri -25725 -18828 -25023 -18126 sw
tri -25015 -18828 -24313 -18126 ne
rect -24313 -18466 -21655 -18126
tri -21655 -18466 -21139 -17950 sw
tri -20946 -18466 -20430 -17950 ne
rect -20430 -18466 -17428 -17950
tri -17428 -18466 -16894 -17932 sw
tri -16718 -18466 -16184 -17932 ne
rect -16184 -18466 -14941 -17932
rect -24313 -18828 -21139 -18466
rect -30679 -19537 -29268 -18828
tri -29268 -19537 -28559 -18828 sw
tri -28559 -19537 -27850 -18828 ne
rect -27850 -19537 -25023 -18828
tri -25023 -19537 -24314 -18828 sw
tri -24313 -19537 -23604 -18828 ne
rect -23604 -19175 -21139 -18828
tri -21139 -19175 -20430 -18466 sw
tri -20430 -19175 -19721 -18466 ne
rect -19721 -19175 -16894 -18466
tri -16894 -19175 -16185 -18466 sw
tri -16184 -19175 -15475 -18466 ne
rect -15475 -19175 -14941 -18466
rect -23604 -19537 -20430 -19175
rect -30679 -20244 -28559 -19537
tri -28559 -20244 -27852 -19537 sw
tri -27850 -20244 -27143 -19537 ne
rect -27143 -20244 -24314 -19537
tri -24314 -20244 -23607 -19537 sw
tri -23604 -20244 -22897 -19537 ne
rect -22897 -19709 -20430 -19537
tri -20430 -19709 -19896 -19175 sw
tri -19721 -19709 -19187 -19175 ne
rect -19187 -19709 -16185 -19175
tri -16185 -19709 -15651 -19175 sw
tri -15475 -19709 -14941 -19175 ne
tri -14941 -19709 -11405 -16173 sw
tri 11752 -19362 15288 -15826 se
rect 15288 -16360 18290 -15826
tri 18290 -16360 18824 -15826 nw
tri 19000 -16360 19534 -15826 se
rect 19534 -16360 22536 -15826
tri 22536 -16360 23070 -15826 nw
tri 23245 -16360 23779 -15826 se
rect 23779 -16360 26781 -15826
tri 26781 -16360 27315 -15826 nw
tri 27491 -16360 28025 -15826 se
rect 28025 -16360 30852 -15826
rect 15288 -16894 17756 -16360
tri 17756 -16894 18290 -16360 nw
tri 18466 -16894 19000 -16360 se
rect 19000 -16894 22002 -16360
tri 22002 -16894 22536 -16360 nw
tri 22711 -16894 23245 -16360 se
rect 23245 -16894 26247 -16360
tri 26247 -16894 26781 -16360 nw
tri 26957 -16894 27491 -16360 se
rect 27491 -16535 30852 -16360
tri 30852 -16535 31561 -15826 nw
tri 31736 -16360 32270 -15826 se
rect 32270 -16360 33513 -15826
tri 31561 -16535 31736 -16360 se
rect 31736 -16535 33513 -16360
rect 27491 -16894 30143 -16535
rect 15288 -17428 17222 -16894
tri 17222 -17428 17756 -16894 nw
tri 17932 -17428 18466 -16894 se
rect 18466 -17428 21293 -16894
rect 15288 -18138 16512 -17428
tri 16512 -18138 17222 -17428 nw
tri 17222 -18138 17932 -17428 se
rect 17932 -17603 21293 -17428
tri 21293 -17603 22002 -16894 nw
tri 22002 -17603 22711 -16894 se
rect 22711 -17603 25538 -16894
tri 25538 -17603 26247 -16894 nw
tri 26248 -17603 26957 -16894 se
rect 26957 -17244 30143 -16894
tri 30143 -17244 30852 -16535 nw
tri 30852 -17244 31561 -16535 se
rect 31561 -17244 33513 -16535
rect 26957 -17603 29437 -17244
rect 17932 -18138 20758 -17603
tri 20758 -18138 21293 -17603 nw
tri 21467 -18138 22002 -17603 se
rect 22002 -17951 25190 -17603
tri 25190 -17951 25538 -17603 nw
tri 25900 -17951 26248 -17603 se
rect 26248 -17950 29437 -17603
tri 29437 -17950 30143 -17244 nw
tri 30146 -17950 30852 -17244 se
rect 30852 -17950 33513 -17244
rect 26248 -17951 29268 -17950
rect 22002 -18138 24481 -17951
rect 15288 -18828 15822 -18138
tri 15822 -18828 16512 -18138 nw
tri 16532 -18828 17222 -18138 se
rect 17222 -18828 20068 -18138
tri 20068 -18828 20758 -18138 nw
tri 20777 -18828 21467 -18138 se
rect 21467 -18660 24481 -18138
tri 24481 -18660 25190 -17951 nw
tri 25191 -18660 25900 -17951 se
rect 25900 -18119 29268 -17951
tri 29268 -18119 29437 -17950 nw
tri 29977 -18119 30146 -17950 se
rect 30146 -18119 33513 -17950
tri 33513 -18119 36508 -15124 nw
rect 25900 -18660 28727 -18119
tri 28727 -18660 29268 -18119 nw
tri 29436 -18660 29977 -18119 se
rect 29977 -18660 32804 -18119
rect 21467 -18828 23779 -18660
tri 15288 -19362 15822 -18828 nw
tri 15998 -19362 16532 -18828 se
rect 16532 -19362 19534 -18828
tri 19534 -19362 20068 -18828 nw
tri 20243 -19362 20777 -18828 se
rect 20777 -19362 23779 -18828
tri 23779 -19362 24481 -18660 nw
tri 24489 -19362 25191 -18660 se
rect 25191 -19362 28025 -18660
tri 28025 -19362 28727 -18660 nw
tri 28734 -19362 29436 -18660 se
rect 29436 -18828 32804 -18660
tri 32804 -18828 33513 -18119 nw
rect 29436 -19362 29977 -18828
rect -22897 -20244 -19896 -19709
tri -19896 -20244 -19361 -19709 sw
tri -19187 -20244 -18652 -19709 ne
rect -18652 -20244 -15651 -19709
tri -15651 -20244 -15116 -19709 sw
tri -14941 -20244 -14406 -19709 ne
rect -14406 -20244 -11405 -19709
rect -30679 -20953 -27852 -20244
tri -27852 -20953 -27143 -20244 sw
tri -27143 -20953 -26434 -20244 ne
rect -26434 -20953 -23607 -20244
tri -23607 -20953 -22898 -20244 sw
tri -22897 -20953 -22188 -20244 ne
rect -22188 -20953 -19361 -20244
tri -19361 -20953 -18652 -20244 sw
tri -18652 -20953 -17943 -20244 ne
rect -17943 -20953 -15116 -20244
tri -15116 -20953 -14407 -20244 sw
tri -14406 -20953 -13697 -20244 ne
rect -13697 -20953 -11405 -20244
tri -30679 -24489 -27143 -20953 ne
tri -27143 -21662 -26434 -20953 sw
tri -26434 -21662 -25725 -20953 ne
rect -25725 -21662 -22898 -20953
tri -22898 -21662 -22189 -20953 sw
tri -22188 -21662 -21479 -20953 ne
rect -21479 -21486 -18652 -20953
tri -18652 -21486 -18119 -20953 sw
tri -17943 -21486 -17410 -20953 ne
rect -17410 -21468 -14407 -20953
tri -14407 -21468 -13892 -20953 sw
tri -13697 -21468 -13182 -20953 ne
rect -13182 -21468 -11405 -20953
rect -17410 -21486 -13892 -21468
rect -21479 -21662 -18119 -21486
rect -27143 -22364 -26434 -21662
tri -26434 -22364 -25732 -21662 sw
tri -25725 -22364 -25023 -21662 ne
rect -25023 -22364 -22189 -21662
tri -22189 -22364 -21487 -21662 sw
tri -21479 -22364 -20777 -21662 ne
rect -20777 -22002 -18119 -21662
tri -18119 -22002 -17603 -21486 sw
tri -17410 -22002 -16894 -21486 ne
rect -16894 -22002 -13892 -21486
tri -13892 -22002 -13358 -21468 sw
tri -13182 -22002 -12648 -21468 ne
rect -12648 -22000 -11405 -21468
tri -11405 -22000 -9114 -19709 sw
tri 9114 -22000 11752 -19362 se
rect 11752 -19896 14754 -19362
tri 14754 -19896 15288 -19362 nw
tri 15464 -19896 15998 -19362 se
rect 15998 -19896 19000 -19362
tri 19000 -19896 19534 -19362 nw
tri 19709 -19896 20243 -19362 se
rect 20243 -19896 23245 -19362
tri 23245 -19896 23779 -19362 nw
tri 23955 -19896 24489 -19362 se
rect 24489 -19896 27316 -19362
rect 11752 -20430 14220 -19896
tri 14220 -20430 14754 -19896 nw
tri 14930 -20430 15464 -19896 se
rect 15464 -20430 18466 -19896
tri 18466 -20430 19000 -19896 nw
tri 19175 -20430 19709 -19896 se
rect 19709 -20430 22711 -19896
tri 22711 -20430 23245 -19896 nw
tri 23421 -20430 23955 -19896 se
rect 23955 -20071 27316 -19896
tri 27316 -20071 28025 -19362 nw
tri 28200 -19896 28734 -19362 se
rect 28734 -19896 29977 -19362
tri 28025 -20071 28200 -19896 se
rect 28200 -20071 29977 -19896
rect 23955 -20430 26607 -20071
rect 11752 -20964 13686 -20430
tri 13686 -20964 14220 -20430 nw
tri 14396 -20964 14930 -20430 se
rect 14930 -20964 17757 -20430
rect 11752 -21674 12976 -20964
tri 12976 -21674 13686 -20964 nw
tri 13686 -21674 14396 -20964 se
rect 14396 -21139 17757 -20964
tri 17757 -21139 18466 -20430 nw
tri 18466 -21139 19175 -20430 se
rect 19175 -21139 22002 -20430
tri 22002 -21139 22711 -20430 nw
tri 22712 -21139 23421 -20430 se
rect 23421 -20780 26607 -20430
tri 26607 -20780 27316 -20071 nw
tri 27316 -20780 28025 -20071 se
rect 28025 -20780 29977 -20071
rect 23421 -21139 25901 -20780
rect 14396 -21674 17222 -21139
tri 17222 -21674 17757 -21139 nw
tri 17931 -21674 18466 -21139 se
rect 18466 -21487 21654 -21139
tri 21654 -21487 22002 -21139 nw
tri 22364 -21487 22712 -21139 se
rect 22712 -21486 25901 -21139
tri 25901 -21486 26607 -20780 nw
tri 26610 -21486 27316 -20780 se
rect 27316 -21486 29977 -20780
rect 22712 -21487 25732 -21486
rect 18466 -21674 20945 -21487
rect 11752 -22000 12286 -21674
rect -12648 -22002 12286 -22000
rect -20777 -22364 -17603 -22002
rect -27143 -23073 -25732 -22364
tri -25732 -23073 -25023 -22364 sw
tri -25023 -23073 -24314 -22364 ne
rect -24314 -23073 -21487 -22364
tri -21487 -23073 -20778 -22364 sw
tri -20777 -23073 -20068 -22364 ne
rect -20068 -22711 -17603 -22364
tri -17603 -22711 -16894 -22002 sw
tri -16894 -22711 -16185 -22002 ne
rect -16185 -22711 -13358 -22002
tri -13358 -22711 -12649 -22002 sw
tri -12648 -22711 -11939 -22002 ne
rect -11939 -22364 12286 -22002
tri 12286 -22364 12976 -21674 nw
tri 12996 -22364 13686 -21674 se
rect 13686 -22364 16532 -21674
tri 16532 -22364 17222 -21674 nw
tri 17241 -22364 17931 -21674 se
rect 17931 -22196 20945 -21674
tri 20945 -22196 21654 -21487 nw
tri 21655 -22196 22364 -21487 se
rect 22364 -21655 25732 -21487
tri 25732 -21655 25901 -21486 nw
tri 26441 -21655 26610 -21486 se
rect 26610 -21655 29977 -21486
tri 29977 -21655 32804 -18828 nw
rect 22364 -22196 25191 -21655
tri 25191 -22196 25732 -21655 nw
tri 25900 -22196 26441 -21655 se
rect 26441 -22196 29268 -21655
rect 17931 -22364 20243 -22196
rect -11939 -22711 11752 -22364
rect -20068 -23073 -16894 -22711
rect -27143 -23780 -25023 -23073
tri -25023 -23780 -24316 -23073 sw
tri -24314 -23780 -23607 -23073 ne
rect -23607 -23780 -20778 -23073
tri -20778 -23780 -20071 -23073 sw
tri -20068 -23780 -19361 -23073 ne
rect -19361 -23245 -16894 -23073
tri -16894 -23245 -16360 -22711 sw
tri -16185 -23245 -15651 -22711 ne
rect -15651 -23245 -12649 -22711
tri -12649 -23245 -12115 -22711 sw
tri -11939 -23245 -11405 -22711 ne
rect -11405 -22898 11752 -22711
tri 11752 -22898 12286 -22364 nw
tri 12462 -22898 12996 -22364 se
rect 12996 -22898 15998 -22364
tri 15998 -22898 16532 -22364 nw
tri 16707 -22898 17241 -22364 se
rect 17241 -22898 20243 -22364
tri 20243 -22898 20945 -22196 nw
tri 20953 -22898 21655 -22196 se
rect 21655 -22898 24489 -22196
tri 24489 -22898 25191 -22196 nw
tri 25198 -22898 25900 -22196 se
rect 25900 -22364 29268 -22196
tri 29268 -22364 29977 -21655 nw
rect 25900 -22898 26441 -22364
rect -11405 -23245 11218 -22898
rect -19361 -23780 -16360 -23245
tri -16360 -23780 -15825 -23245 sw
tri -15651 -23780 -15116 -23245 ne
rect -15116 -23780 -12115 -23245
tri -12115 -23780 -11580 -23245 sw
tri -11405 -23780 -10870 -23245 ne
rect -10870 -23432 11218 -23245
tri 11218 -23432 11752 -22898 nw
tri 11928 -23432 12462 -22898 se
rect 12462 -23432 15464 -22898
tri 15464 -23432 15998 -22898 nw
tri 16173 -23432 16707 -22898 se
rect 16707 -23432 19709 -22898
tri 19709 -23432 20243 -22898 nw
tri 20419 -23432 20953 -22898 se
rect 20953 -23432 23780 -22898
rect -10870 -23780 10684 -23432
rect -27143 -24489 -24316 -23780
tri -24316 -24489 -23607 -23780 sw
tri -23607 -24489 -22898 -23780 ne
rect -22898 -24489 -20071 -23780
tri -20071 -24489 -19362 -23780 sw
tri -19361 -24489 -18652 -23780 ne
rect -18652 -24489 -15825 -23780
tri -15825 -24489 -15116 -23780 sw
tri -15116 -24489 -14407 -23780 ne
rect -14407 -24489 -11580 -23780
tri -11580 -24489 -10871 -23780 sw
tri -10870 -24489 -10161 -23780 ne
rect -10161 -23966 10684 -23780
tri 10684 -23966 11218 -23432 nw
tri 11394 -23966 11928 -23432 se
rect 11928 -23966 14930 -23432
tri 14930 -23966 15464 -23432 nw
tri 15639 -23966 16173 -23432 se
rect 16173 -23966 19175 -23432
tri 19175 -23966 19709 -23432 nw
tri 19885 -23966 20419 -23432 se
rect 20419 -23607 23780 -23432
tri 23780 -23607 24489 -22898 nw
tri 24664 -23432 25198 -22898 se
rect 25198 -23432 26441 -22898
tri 24489 -23607 24664 -23432 se
rect 24664 -23607 26441 -23432
rect 20419 -23966 23071 -23607
rect -10161 -24489 10150 -23966
tri -27143 -28025 -23607 -24489 ne
tri -23607 -25198 -22898 -24489 sw
tri -22898 -25198 -22189 -24489 ne
rect -22189 -25198 -19362 -24489
tri -19362 -25198 -18653 -24489 sw
tri -18652 -25198 -17943 -24489 ne
rect -17943 -25022 -15116 -24489
tri -15116 -25022 -14583 -24489 sw
tri -14407 -25022 -13874 -24489 ne
rect -13874 -25002 -10871 -24489
tri -10871 -25002 -10358 -24489 sw
tri -10161 -24500 -10150 -24489 ne
rect -10150 -24500 10150 -24489
tri 10150 -24500 10684 -23966 nw
tri 10860 -24500 11394 -23966 se
rect 11394 -24500 14396 -23966
tri 14396 -24500 14930 -23966 nw
tri 15105 -24500 15639 -23966 se
rect 15639 -24500 18466 -23966
tri 10358 -25002 10860 -24500 se
rect 10860 -25002 13894 -24500
tri 13894 -25002 14396 -24500 nw
tri 14603 -25002 15105 -24500 se
rect 15105 -24675 18466 -24500
tri 18466 -24675 19175 -23966 nw
tri 19176 -24675 19885 -23966 se
rect 19885 -24316 23071 -23966
tri 23071 -24316 23780 -23607 nw
tri 23780 -24316 24489 -23607 se
rect 24489 -24316 26441 -23607
rect 19885 -24675 22365 -24316
rect 15105 -25002 18118 -24675
rect -13874 -25022 -979 -25002
rect -17943 -25198 -14583 -25022
rect -23607 -25900 -22898 -25198
tri -22898 -25900 -22196 -25198 sw
tri -22189 -25900 -21487 -25198 ne
rect -21487 -25900 -18653 -25198
tri -18653 -25900 -17951 -25198 sw
tri -17943 -25900 -17241 -25198 ne
rect -17241 -25580 -14583 -25198
tri -14583 -25580 -14025 -25022 sw
tri -13874 -25580 -13316 -25022 ne
rect -13316 -25580 -979 -25022
rect -17241 -25900 -14025 -25580
rect -23607 -26609 -22196 -25900
tri -22196 -26609 -21487 -25900 sw
tri -21487 -26609 -20778 -25900 ne
rect -20778 -26609 -17951 -25900
tri -17951 -26609 -17242 -25900 sw
tri -17241 -26609 -16532 -25900 ne
rect -16532 -26247 -14025 -25900
tri -14025 -26247 -13358 -25580 sw
tri -13316 -25732 -13164 -25580 ne
rect -13164 -25732 -979 -25580
tri -13164 -26247 -12649 -25732 ne
rect -12649 -26247 -979 -25732
rect -16532 -26609 -13358 -26247
rect -23607 -27316 -21487 -26609
tri -21487 -27316 -20780 -26609 sw
tri -20778 -27316 -20071 -26609 ne
rect -20071 -27316 -17242 -26609
tri -17242 -27316 -16535 -26609 sw
tri -16532 -27316 -15825 -26609 ne
rect -15825 -26926 -13358 -26609
tri -13358 -26926 -12679 -26247 sw
tri -12649 -26926 -11970 -26247 ne
rect -11970 -26926 -979 -26247
rect -15825 -27316 -12679 -26926
rect -23607 -28025 -20780 -27316
tri -20780 -28025 -20071 -27316 sw
tri -20071 -28025 -19362 -27316 ne
rect -19362 -28025 -16535 -27316
tri -16535 -28025 -15826 -27316 sw
tri -15825 -28025 -15116 -27316 ne
rect -15116 -27502 -12679 -27316
tri -12679 -27502 -12103 -26926 sw
tri -11970 -27502 -11394 -26926 ne
rect -11394 -27502 -979 -26926
rect -15116 -28004 -12103 -27502
tri -12103 -28004 -11601 -27502 sw
rect -15116 -28025 -2380 -28004
tri -23607 -31561 -20071 -28025 ne
tri -20071 -28734 -19362 -28025 sw
tri -19362 -28734 -18653 -28025 ne
rect -18653 -28734 -15826 -28025
tri -15826 -28734 -15117 -28025 sw
tri -15116 -28734 -14407 -28025 ne
rect -14407 -28224 -2380 -28025
tri -2380 -28224 -2160 -28004 sw
tri -2015 -28224 -1293 -27502 ne
rect -1293 -28004 -979 -27502
tri -979 -28004 2023 -25002 sw
tri 2291 -25222 2511 -25002 se
rect 2511 -25222 13316 -25002
rect 2291 -25580 13316 -25222
tri 13316 -25580 13894 -25002 nw
tri 14025 -25580 14603 -25002 se
rect 14603 -25023 18118 -25002
tri 18118 -25023 18466 -24675 nw
tri 18828 -25023 19176 -24675 se
rect 19176 -25022 22365 -24675
tri 22365 -25022 23071 -24316 nw
tri 23074 -25022 23780 -24316 se
rect 23780 -25022 26441 -24316
rect 19176 -25023 22196 -25022
rect 14603 -25580 17409 -25023
rect 2291 -26247 12649 -25580
tri 12649 -26247 13316 -25580 nw
tri 13358 -26247 14025 -25580 se
rect 14025 -25732 17409 -25580
tri 17409 -25732 18118 -25023 nw
tri 18119 -25732 18828 -25023 se
rect 18828 -25191 22196 -25023
tri 22196 -25191 22365 -25022 nw
tri 22905 -25191 23074 -25022 se
rect 23074 -25191 26441 -25022
tri 26441 -25191 29268 -22364 nw
rect 18828 -25732 21655 -25191
tri 21655 -25732 22196 -25191 nw
tri 22364 -25732 22905 -25191 se
rect 22905 -25732 25732 -25191
rect 14025 -26247 16707 -25732
rect 2291 -26926 11970 -26247
tri 11970 -26926 12649 -26247 nw
tri 12679 -26926 13358 -26247 se
rect 13358 -26434 16707 -26247
tri 16707 -26434 17409 -25732 nw
tri 17417 -26434 18119 -25732 se
rect 18119 -26434 20953 -25732
tri 20953 -26434 21655 -25732 nw
tri 21662 -26434 22364 -25732 se
rect 22364 -25900 25732 -25732
tri 25732 -25900 26441 -25191 nw
rect 22364 -26434 22905 -25900
rect 13358 -26926 16173 -26434
rect 2291 -27282 11394 -26926
tri 2291 -27502 2511 -27282 ne
rect 2511 -27502 11394 -27282
tri 11394 -27502 11970 -26926 nw
tri 12103 -27502 12679 -26926 se
rect 12679 -26968 16173 -26926
tri 16173 -26968 16707 -26434 nw
tri 16883 -26968 17417 -26434 se
rect 17417 -26968 20244 -26434
rect 12679 -27502 15639 -26968
tri 15639 -27502 16173 -26968 nw
tri 16349 -27502 16883 -26968 se
rect 16883 -27143 20244 -26968
tri 20244 -27143 20953 -26434 nw
tri 21128 -26968 21662 -26434 se
rect 21662 -26968 22905 -26434
tri 20953 -27143 21128 -26968 se
rect 21128 -27143 22905 -26968
rect 16883 -27502 19709 -27143
tri 11601 -28004 12103 -27502 se
rect 12103 -28004 15116 -27502
rect -1293 -28025 15116 -28004
tri 15116 -28025 15639 -27502 nw
tri 15826 -28025 16349 -27502 se
rect 16349 -27678 19709 -27502
tri 19709 -27678 20244 -27143 nw
tri 20418 -27678 20953 -27143 se
rect 20953 -27678 22905 -27143
rect 16349 -28004 19383 -27678
tri 19383 -28004 19709 -27678 nw
tri 20092 -28004 20418 -27678 se
rect 20418 -28004 22905 -27678
rect 16349 -28025 18829 -28004
rect -1293 -28224 14583 -28025
rect -14407 -28734 -2160 -28224
tri -1293 -28581 -936 -28224 ne
rect -936 -28558 14583 -28224
tri 14583 -28558 15116 -28025 nw
tri 15293 -28558 15826 -28025 se
rect 15826 -28558 18829 -28025
tri 18829 -28558 19383 -28004 nw
tri 19538 -28558 20092 -28004 se
rect 20092 -28558 22905 -28004
rect -936 -28581 13873 -28558
rect -20071 -29436 -19362 -28734
tri -19362 -29436 -18660 -28734 sw
tri -18653 -29436 -17951 -28734 ne
rect -17951 -29436 -15117 -28734
tri -15117 -29436 -14415 -28734 sw
tri -14407 -29436 -13705 -28734 ne
rect -13705 -29436 -2160 -28734
tri -936 -29268 -249 -28581 ne
rect -249 -29268 13873 -28581
tri 13873 -29268 14583 -28558 nw
tri 14583 -29268 15293 -28558 se
rect 15293 -28727 18660 -28558
tri 18660 -28727 18829 -28558 nw
tri 19369 -28727 19538 -28558 se
rect 19538 -28727 22905 -28558
tri 22905 -28727 25732 -25900 nw
rect 15293 -29268 18119 -28727
tri 18119 -29268 18660 -28727 nw
tri 18828 -29268 19369 -28727 se
rect 19369 -29268 22196 -28727
rect -20071 -30145 -18660 -29436
tri -18660 -30145 -17951 -29436 sw
tri -17951 -30145 -17242 -29436 ne
rect -17242 -30145 -14415 -29436
tri -14415 -30145 -13706 -29436 sw
tri -13705 -30145 -12996 -29436 ne
rect -12996 -30145 -2160 -29436
tri -249 -29970 453 -29268 ne
rect 453 -29970 13171 -29268
tri 13171 -29970 13873 -29268 nw
tri 13881 -29970 14583 -29268 se
rect 14583 -29970 17417 -29268
tri 17417 -29970 18119 -29268 nw
tri 18126 -29970 18828 -29268 se
rect 18828 -29436 22196 -29268
tri 22196 -29436 22905 -28727 nw
rect 18828 -29970 19369 -29436
rect -20071 -30852 -17951 -30145
tri -17951 -30852 -17244 -30145 sw
tri -17242 -30852 -16535 -30145 ne
rect -16535 -30852 -13706 -30145
tri -13706 -30852 -12999 -30145 sw
tri -12996 -30504 -12637 -30145 ne
rect -12637 -30284 -2160 -30145
tri 453 -30284 767 -29970 ne
rect 767 -30284 12637 -29970
rect -12637 -30504 -2380 -30284
tri -2380 -30504 -2160 -30284 nw
tri 767 -30317 800 -30284 ne
rect 800 -30317 12637 -30284
tri 800 -30504 987 -30317 ne
rect 987 -30504 12637 -30317
tri 12637 -30504 13171 -29970 nw
tri 13347 -30504 13881 -29970 se
rect 13881 -30504 16883 -29970
tri 16883 -30504 17417 -29970 nw
tri 17592 -30504 18126 -29970 se
rect 18126 -30504 19369 -29970
rect -20071 -31561 -17244 -30852
tri -17244 -31561 -16535 -30852 sw
tri -16535 -31561 -15826 -30852 ne
rect -15826 -31006 -12999 -30852
tri -12999 -31006 -12845 -30852 sw
tri 12845 -31006 13347 -30504 se
rect 13347 -31006 16381 -30504
tri 16381 -31006 16883 -30504 nw
tri 17090 -31006 17592 -30504 se
rect 17592 -31006 19369 -30504
rect -15826 -31561 -979 -31006
tri -20071 -35079 -16553 -31561 ne
rect -16553 -32270 -16535 -31561
tri -16535 -32270 -15826 -31561 sw
tri -15826 -32270 -15117 -31561 ne
rect -15117 -32270 -979 -31561
rect -16553 -32972 -15826 -32270
tri -15826 -32972 -15124 -32270 sw
tri -15117 -32972 -14415 -32270 ne
rect -14415 -32972 -979 -32270
rect -16553 -33506 -15124 -32972
tri -15124 -33506 -14590 -32972 sw
tri -14415 -33506 -13881 -32972 ne
rect -13881 -33506 -979 -32972
rect -16553 -34008 -14590 -33506
tri -14590 -34008 -14088 -33506 sw
rect -16553 -34228 -2380 -34008
tri -2380 -34228 -2160 -34008 sw
tri -2015 -34228 -1293 -33506 ne
rect -1293 -34008 -979 -33506
tri -979 -34008 2023 -31006 sw
tri 2291 -31226 2511 -31006 se
rect 2511 -31226 16161 -31006
tri 16161 -31226 16381 -31006 nw
tri 16870 -31226 17090 -31006 se
rect 17090 -31226 19369 -31006
rect 2291 -31561 15826 -31226
tri 15826 -31561 16161 -31226 nw
tri 16535 -31561 16870 -31226 se
rect 16870 -31561 19369 -31226
rect 2291 -32270 15117 -31561
tri 15117 -32270 15826 -31561 nw
tri 15826 -32270 16535 -31561 se
rect 16535 -32263 19369 -31561
tri 19369 -32263 22196 -29436 nw
rect 16535 -32270 18660 -32263
rect 2291 -32972 14415 -32270
tri 14415 -32972 15117 -32270 nw
tri 15124 -32972 15826 -32270 se
rect 15826 -32972 18660 -32270
tri 18660 -32972 19369 -32263 nw
rect 2291 -33286 13881 -32972
tri 2291 -33506 2511 -33286 ne
rect 2511 -33506 13881 -33286
tri 13881 -33506 14415 -32972 nw
tri 14590 -33506 15124 -32972 se
tri 14088 -34008 14590 -33506 se
rect 14590 -34008 15124 -33506
rect -1293 -34228 15124 -34008
rect -16553 -35079 -2160 -34228
tri -1293 -35079 -442 -34228 ne
rect -442 -35079 15124 -34228
tri -16553 -36508 -15124 -35079 ne
rect -15124 -36288 -2160 -35079
tri -442 -36288 767 -35079 ne
rect 767 -36288 15124 -35079
rect -15124 -36508 -2380 -36288
tri -2380 -36508 -2160 -36288 nw
tri 767 -36508 987 -36288 ne
rect 987 -36508 15124 -36288
tri 15124 -36508 18660 -32972 nw
<< properties >>
string FIXED_BBOX -36508 -36508 37508 36508
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil3
string library sky130
string parameter m=1
string GDS_END 10411016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10379748
<< end >>
