magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< metal1 >>
rect 1500 1959 1530 2011
rect 1702 1959 1732 2011
rect 6492 1959 6522 2011
rect 6694 1959 6724 2011
rect 11484 1959 11514 2011
rect 11686 1959 11716 2011
rect 16476 1959 16506 2011
rect 16678 1959 16708 2011
rect 21468 1959 21498 2011
rect 21670 1959 21700 2011
rect 26460 1959 26490 2011
rect 26662 1959 26692 2011
rect 31452 1959 31482 2011
rect 31654 1959 31684 2011
rect 36444 1959 36474 2011
rect 36646 1959 36676 2011
rect 1615 1604 1667 1610
rect 1615 1546 1667 1552
rect 6607 1604 6659 1610
rect 6607 1546 6659 1552
rect 11599 1604 11651 1610
rect 11599 1546 11651 1552
rect 16591 1604 16643 1610
rect 16591 1546 16643 1552
rect 21583 1604 21635 1610
rect 21583 1546 21635 1552
rect 26575 1604 26627 1610
rect 26575 1546 26627 1552
rect 31567 1604 31619 1610
rect 31567 1546 31619 1552
rect 36559 1604 36611 1610
rect 36559 1546 36611 1552
rect 1604 1167 1656 1173
rect 1604 1109 1656 1115
rect 6596 1167 6648 1173
rect 6596 1109 6648 1115
rect 11588 1167 11640 1173
rect 11588 1109 11640 1115
rect 16580 1167 16632 1173
rect 16580 1109 16632 1115
rect 21572 1167 21624 1173
rect 21572 1109 21624 1115
rect 26564 1167 26616 1173
rect 26564 1109 26616 1115
rect 31556 1167 31608 1173
rect 31556 1109 31608 1115
rect 36548 1167 36600 1173
rect 36548 1109 36600 1115
rect 1725 836 1777 842
rect 1725 778 1777 784
rect 6717 836 6769 842
rect 6717 778 6769 784
rect 11709 836 11761 842
rect 11709 778 11761 784
rect 16701 836 16753 842
rect 16701 778 16753 784
rect 21693 836 21745 842
rect 21693 778 21745 784
rect 26685 836 26737 842
rect 26685 778 26737 784
rect 31677 836 31729 842
rect 31677 778 31729 784
rect 36669 836 36721 842
rect 36669 778 36721 784
rect 1610 633 1662 639
rect 1610 575 1662 581
rect 6602 633 6654 639
rect 6602 575 6654 581
rect 11594 633 11646 639
rect 11594 575 11646 581
rect 16586 633 16638 639
rect 16586 575 16638 581
rect 21578 633 21630 639
rect 21578 575 21630 581
rect 26570 633 26622 639
rect 26570 575 26622 581
rect 31562 633 31614 639
rect 31562 575 31614 581
rect 36554 633 36606 639
rect 36554 575 36606 581
rect 1624 217 1676 223
rect 1624 159 1676 165
rect 6616 217 6668 223
rect 6616 159 6668 165
rect 11608 217 11660 223
rect 11608 159 11660 165
rect 16600 217 16652 223
rect 16600 159 16652 165
rect 21592 217 21644 223
rect 21592 159 21644 165
rect 26584 217 26636 223
rect 26584 159 26636 165
rect 31576 217 31628 223
rect 31576 159 31628 165
rect 36568 217 36620 223
rect 36568 159 36620 165
rect 1473 94 40785 128
rect 1629 4 1689 60
rect 6621 4 6681 60
rect 11613 4 11673 60
rect 16605 4 16665 60
rect 21597 4 21657 60
rect 26589 4 26649 60
rect 31581 4 31641 60
rect 36573 4 36633 60
<< via1 >>
rect 1615 1552 1667 1604
rect 6607 1552 6659 1604
rect 11599 1552 11651 1604
rect 16591 1552 16643 1604
rect 21583 1552 21635 1604
rect 26575 1552 26627 1604
rect 31567 1552 31619 1604
rect 36559 1552 36611 1604
rect 1604 1115 1656 1167
rect 6596 1115 6648 1167
rect 11588 1115 11640 1167
rect 16580 1115 16632 1167
rect 21572 1115 21624 1167
rect 26564 1115 26616 1167
rect 31556 1115 31608 1167
rect 36548 1115 36600 1167
rect 1725 784 1777 836
rect 6717 784 6769 836
rect 11709 784 11761 836
rect 16701 784 16753 836
rect 21693 784 21745 836
rect 26685 784 26737 836
rect 31677 784 31729 836
rect 36669 784 36721 836
rect 1610 581 1662 633
rect 6602 581 6654 633
rect 11594 581 11646 633
rect 16586 581 16638 633
rect 21578 581 21630 633
rect 26570 581 26622 633
rect 31562 581 31614 633
rect 36554 581 36606 633
rect 1624 165 1676 217
rect 6616 165 6668 217
rect 11608 165 11660 217
rect 16600 165 16652 217
rect 21592 165 21644 217
rect 26584 165 26636 217
rect 31576 165 31628 217
rect 36568 165 36620 217
<< metal2 >>
rect 1613 1606 1669 1615
rect 1613 1541 1669 1550
rect 6605 1606 6661 1615
rect 6605 1541 6661 1550
rect 11597 1606 11653 1615
rect 11597 1541 11653 1550
rect 16589 1606 16645 1615
rect 16589 1541 16645 1550
rect 21581 1606 21637 1615
rect 21581 1541 21637 1550
rect 26573 1606 26629 1615
rect 26573 1541 26629 1550
rect 31565 1606 31621 1615
rect 31565 1541 31621 1550
rect 36557 1606 36613 1615
rect 36557 1541 36613 1550
rect 1602 1169 1658 1178
rect 1602 1104 1658 1113
rect 6594 1169 6650 1178
rect 6594 1104 6650 1113
rect 11586 1169 11642 1178
rect 11586 1104 11642 1113
rect 16578 1169 16634 1178
rect 16578 1104 16634 1113
rect 21570 1169 21626 1178
rect 21570 1104 21626 1113
rect 26562 1169 26618 1178
rect 26562 1104 26618 1113
rect 31554 1169 31610 1178
rect 31554 1104 31610 1113
rect 36546 1169 36602 1178
rect 36546 1104 36602 1113
rect 1723 837 1779 846
rect 1723 772 1779 781
rect 6715 837 6771 846
rect 6715 772 6771 781
rect 11707 837 11763 846
rect 11707 772 11763 781
rect 16699 837 16755 846
rect 16699 772 16755 781
rect 21691 837 21747 846
rect 21691 772 21747 781
rect 26683 837 26739 846
rect 26683 772 26739 781
rect 31675 837 31731 846
rect 31675 772 31731 781
rect 36667 837 36723 846
rect 36667 772 36723 781
rect 1608 635 1664 644
rect 1608 570 1664 579
rect 6600 635 6656 644
rect 6600 570 6656 579
rect 11592 635 11648 644
rect 11592 570 11648 579
rect 16584 635 16640 644
rect 16584 570 16640 579
rect 21576 635 21632 644
rect 21576 570 21632 579
rect 26568 635 26624 644
rect 26568 570 26624 579
rect 31560 635 31616 644
rect 31560 570 31616 579
rect 36552 635 36608 644
rect 36552 570 36608 579
rect 1622 219 1678 228
rect 1622 154 1678 163
rect 6614 219 6670 228
rect 6614 154 6670 163
rect 11606 219 11662 228
rect 11606 154 11662 163
rect 16598 219 16654 228
rect 16598 154 16654 163
rect 21590 219 21646 228
rect 21590 154 21646 163
rect 26582 219 26638 228
rect 26582 154 26638 163
rect 31574 219 31630 228
rect 31574 154 31630 163
rect 36566 219 36622 228
rect 36566 154 36622 163
<< via2 >>
rect 1613 1604 1669 1606
rect 1613 1552 1615 1604
rect 1615 1552 1667 1604
rect 1667 1552 1669 1604
rect 1613 1550 1669 1552
rect 6605 1604 6661 1606
rect 6605 1552 6607 1604
rect 6607 1552 6659 1604
rect 6659 1552 6661 1604
rect 6605 1550 6661 1552
rect 11597 1604 11653 1606
rect 11597 1552 11599 1604
rect 11599 1552 11651 1604
rect 11651 1552 11653 1604
rect 11597 1550 11653 1552
rect 16589 1604 16645 1606
rect 16589 1552 16591 1604
rect 16591 1552 16643 1604
rect 16643 1552 16645 1604
rect 16589 1550 16645 1552
rect 21581 1604 21637 1606
rect 21581 1552 21583 1604
rect 21583 1552 21635 1604
rect 21635 1552 21637 1604
rect 21581 1550 21637 1552
rect 26573 1604 26629 1606
rect 26573 1552 26575 1604
rect 26575 1552 26627 1604
rect 26627 1552 26629 1604
rect 26573 1550 26629 1552
rect 31565 1604 31621 1606
rect 31565 1552 31567 1604
rect 31567 1552 31619 1604
rect 31619 1552 31621 1604
rect 31565 1550 31621 1552
rect 36557 1604 36613 1606
rect 36557 1552 36559 1604
rect 36559 1552 36611 1604
rect 36611 1552 36613 1604
rect 36557 1550 36613 1552
rect 1602 1167 1658 1169
rect 1602 1115 1604 1167
rect 1604 1115 1656 1167
rect 1656 1115 1658 1167
rect 1602 1113 1658 1115
rect 6594 1167 6650 1169
rect 6594 1115 6596 1167
rect 6596 1115 6648 1167
rect 6648 1115 6650 1167
rect 6594 1113 6650 1115
rect 11586 1167 11642 1169
rect 11586 1115 11588 1167
rect 11588 1115 11640 1167
rect 11640 1115 11642 1167
rect 11586 1113 11642 1115
rect 16578 1167 16634 1169
rect 16578 1115 16580 1167
rect 16580 1115 16632 1167
rect 16632 1115 16634 1167
rect 16578 1113 16634 1115
rect 21570 1167 21626 1169
rect 21570 1115 21572 1167
rect 21572 1115 21624 1167
rect 21624 1115 21626 1167
rect 21570 1113 21626 1115
rect 26562 1167 26618 1169
rect 26562 1115 26564 1167
rect 26564 1115 26616 1167
rect 26616 1115 26618 1167
rect 26562 1113 26618 1115
rect 31554 1167 31610 1169
rect 31554 1115 31556 1167
rect 31556 1115 31608 1167
rect 31608 1115 31610 1167
rect 31554 1113 31610 1115
rect 36546 1167 36602 1169
rect 36546 1115 36548 1167
rect 36548 1115 36600 1167
rect 36600 1115 36602 1167
rect 36546 1113 36602 1115
rect 1723 836 1779 837
rect 1723 784 1725 836
rect 1725 784 1777 836
rect 1777 784 1779 836
rect 1723 781 1779 784
rect 6715 836 6771 837
rect 6715 784 6717 836
rect 6717 784 6769 836
rect 6769 784 6771 836
rect 6715 781 6771 784
rect 11707 836 11763 837
rect 11707 784 11709 836
rect 11709 784 11761 836
rect 11761 784 11763 836
rect 11707 781 11763 784
rect 16699 836 16755 837
rect 16699 784 16701 836
rect 16701 784 16753 836
rect 16753 784 16755 836
rect 16699 781 16755 784
rect 21691 836 21747 837
rect 21691 784 21693 836
rect 21693 784 21745 836
rect 21745 784 21747 836
rect 21691 781 21747 784
rect 26683 836 26739 837
rect 26683 784 26685 836
rect 26685 784 26737 836
rect 26737 784 26739 836
rect 26683 781 26739 784
rect 31675 836 31731 837
rect 31675 784 31677 836
rect 31677 784 31729 836
rect 31729 784 31731 836
rect 31675 781 31731 784
rect 36667 836 36723 837
rect 36667 784 36669 836
rect 36669 784 36721 836
rect 36721 784 36723 836
rect 36667 781 36723 784
rect 1608 633 1664 635
rect 1608 581 1610 633
rect 1610 581 1662 633
rect 1662 581 1664 633
rect 1608 579 1664 581
rect 6600 633 6656 635
rect 6600 581 6602 633
rect 6602 581 6654 633
rect 6654 581 6656 633
rect 6600 579 6656 581
rect 11592 633 11648 635
rect 11592 581 11594 633
rect 11594 581 11646 633
rect 11646 581 11648 633
rect 11592 579 11648 581
rect 16584 633 16640 635
rect 16584 581 16586 633
rect 16586 581 16638 633
rect 16638 581 16640 633
rect 16584 579 16640 581
rect 21576 633 21632 635
rect 21576 581 21578 633
rect 21578 581 21630 633
rect 21630 581 21632 633
rect 21576 579 21632 581
rect 26568 633 26624 635
rect 26568 581 26570 633
rect 26570 581 26622 633
rect 26622 581 26624 633
rect 26568 579 26624 581
rect 31560 633 31616 635
rect 31560 581 31562 633
rect 31562 581 31614 633
rect 31614 581 31616 633
rect 31560 579 31616 581
rect 36552 633 36608 635
rect 36552 581 36554 633
rect 36554 581 36606 633
rect 36606 581 36608 633
rect 36552 579 36608 581
rect 1622 217 1678 219
rect 1622 165 1624 217
rect 1624 165 1676 217
rect 1676 165 1678 217
rect 1622 163 1678 165
rect 6614 217 6670 219
rect 6614 165 6616 217
rect 6616 165 6668 217
rect 6668 165 6670 217
rect 6614 163 6670 165
rect 11606 217 11662 219
rect 11606 165 11608 217
rect 11608 165 11660 217
rect 11660 165 11662 217
rect 11606 163 11662 165
rect 16598 217 16654 219
rect 16598 165 16600 217
rect 16600 165 16652 217
rect 16652 165 16654 217
rect 16598 163 16654 165
rect 21590 217 21646 219
rect 21590 165 21592 217
rect 21592 165 21644 217
rect 21644 165 21646 217
rect 21590 163 21646 165
rect 26582 217 26638 219
rect 26582 165 26584 217
rect 26584 165 26636 217
rect 26636 165 26638 217
rect 26582 163 26638 165
rect 31574 217 31630 219
rect 31574 165 31576 217
rect 31576 165 31628 217
rect 31628 165 31630 217
rect 31574 163 31630 165
rect 36566 217 36622 219
rect 36566 165 36568 217
rect 36568 165 36620 217
rect 36620 165 36622 217
rect 36566 163 36622 165
<< metal3 >>
rect 1592 1606 1690 1627
rect 1592 1550 1613 1606
rect 1669 1550 1690 1606
rect 1592 1529 1690 1550
rect 6584 1606 6682 1627
rect 6584 1550 6605 1606
rect 6661 1550 6682 1606
rect 6584 1529 6682 1550
rect 11576 1606 11674 1627
rect 11576 1550 11597 1606
rect 11653 1550 11674 1606
rect 11576 1529 11674 1550
rect 16568 1606 16666 1627
rect 16568 1550 16589 1606
rect 16645 1550 16666 1606
rect 16568 1529 16666 1550
rect 21560 1606 21658 1627
rect 21560 1550 21581 1606
rect 21637 1550 21658 1606
rect 21560 1529 21658 1550
rect 26552 1606 26650 1627
rect 26552 1550 26573 1606
rect 26629 1550 26650 1606
rect 26552 1529 26650 1550
rect 31544 1606 31642 1627
rect 31544 1550 31565 1606
rect 31621 1550 31642 1606
rect 31544 1529 31642 1550
rect 36536 1606 36634 1627
rect 36536 1550 36557 1606
rect 36613 1550 36634 1606
rect 36536 1529 36634 1550
rect 1581 1169 1679 1190
rect 1581 1113 1602 1169
rect 1658 1113 1679 1169
rect 1581 1092 1679 1113
rect 6573 1169 6671 1190
rect 6573 1113 6594 1169
rect 6650 1113 6671 1169
rect 6573 1092 6671 1113
rect 11565 1169 11663 1190
rect 11565 1113 11586 1169
rect 11642 1113 11663 1169
rect 11565 1092 11663 1113
rect 16557 1169 16655 1190
rect 16557 1113 16578 1169
rect 16634 1113 16655 1169
rect 16557 1092 16655 1113
rect 21549 1169 21647 1190
rect 21549 1113 21570 1169
rect 21626 1113 21647 1169
rect 21549 1092 21647 1113
rect 26541 1169 26639 1190
rect 26541 1113 26562 1169
rect 26618 1113 26639 1169
rect 26541 1092 26639 1113
rect 31533 1169 31631 1190
rect 31533 1113 31554 1169
rect 31610 1113 31631 1169
rect 31533 1092 31631 1113
rect 36525 1169 36623 1190
rect 36525 1113 36546 1169
rect 36602 1113 36623 1169
rect 36525 1092 36623 1113
rect 1702 837 1800 858
rect 1702 781 1723 837
rect 1779 781 1800 837
rect 1702 760 1800 781
rect 6694 837 6792 858
rect 6694 781 6715 837
rect 6771 781 6792 837
rect 6694 760 6792 781
rect 11686 837 11784 858
rect 11686 781 11707 837
rect 11763 781 11784 837
rect 11686 760 11784 781
rect 16678 837 16776 858
rect 16678 781 16699 837
rect 16755 781 16776 837
rect 16678 760 16776 781
rect 21670 837 21768 858
rect 21670 781 21691 837
rect 21747 781 21768 837
rect 21670 760 21768 781
rect 26662 837 26760 858
rect 26662 781 26683 837
rect 26739 781 26760 837
rect 26662 760 26760 781
rect 31654 837 31752 858
rect 31654 781 31675 837
rect 31731 781 31752 837
rect 31654 760 31752 781
rect 36646 837 36744 858
rect 36646 781 36667 837
rect 36723 781 36744 837
rect 36646 760 36744 781
rect 1587 635 1685 656
rect 1587 579 1608 635
rect 1664 579 1685 635
rect 1587 558 1685 579
rect 6579 635 6677 656
rect 6579 579 6600 635
rect 6656 579 6677 635
rect 6579 558 6677 579
rect 11571 635 11669 656
rect 11571 579 11592 635
rect 11648 579 11669 635
rect 11571 558 11669 579
rect 16563 635 16661 656
rect 16563 579 16584 635
rect 16640 579 16661 635
rect 16563 558 16661 579
rect 21555 635 21653 656
rect 21555 579 21576 635
rect 21632 579 21653 635
rect 21555 558 21653 579
rect 26547 635 26645 656
rect 26547 579 26568 635
rect 26624 579 26645 635
rect 26547 558 26645 579
rect 31539 635 31637 656
rect 31539 579 31560 635
rect 31616 579 31637 635
rect 31539 558 31637 579
rect 36531 635 36629 656
rect 36531 579 36552 635
rect 36608 579 36629 635
rect 36531 558 36629 579
rect 1601 219 1699 240
rect 1601 163 1622 219
rect 1678 163 1699 219
rect 1601 142 1699 163
rect 6593 219 6691 240
rect 6593 163 6614 219
rect 6670 163 6691 219
rect 6593 142 6691 163
rect 11585 219 11683 240
rect 11585 163 11606 219
rect 11662 163 11683 219
rect 11585 142 11683 163
rect 16577 219 16675 240
rect 16577 163 16598 219
rect 16654 163 16675 219
rect 16577 142 16675 163
rect 21569 219 21667 240
rect 21569 163 21590 219
rect 21646 163 21667 219
rect 21569 142 21667 163
rect 26561 219 26659 240
rect 26561 163 26582 219
rect 26638 163 26659 219
rect 26561 142 26659 163
rect 31553 219 31651 240
rect 31553 163 31574 219
rect 31630 163 31651 219
rect 31553 142 31651 163
rect 36545 219 36643 240
rect 36545 163 36566 219
rect 36622 163 36643 219
rect 36545 142 36643 163
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_0
timestamp 1694700623
transform 1 0 36318 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_1
timestamp 1694700623
transform 1 0 31326 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_2
timestamp 1694700623
transform 1 0 26334 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_3
timestamp 1694700623
transform 1 0 21342 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_4
timestamp 1694700623
transform 1 0 16350 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_5
timestamp 1694700623
transform 1 0 11358 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_6
timestamp 1694700623
transform 1 0 6366 0 1 0
box -376 4 880 2011
use sky130_fd_bd_sram__openram_write_driver_1  sky130_fd_bd_sram__openram_write_driver_7
timestamp 1694700623
transform 1 0 1374 0 1 0
box -376 4 880 2011
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_0
timestamp 1694700623
transform 1 0 36559 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_1
timestamp 1694700623
transform 1 0 36669 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_2
timestamp 1694700623
transform 1 0 36554 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_3
timestamp 1694700623
transform 1 0 36548 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_4
timestamp 1694700623
transform 1 0 36568 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_5
timestamp 1694700623
transform 1 0 31567 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_6
timestamp 1694700623
transform 1 0 31677 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_7
timestamp 1694700623
transform 1 0 31562 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_8
timestamp 1694700623
transform 1 0 31556 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_9
timestamp 1694700623
transform 1 0 31576 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_10
timestamp 1694700623
transform 1 0 26575 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_11
timestamp 1694700623
transform 1 0 26685 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_12
timestamp 1694700623
transform 1 0 26570 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_13
timestamp 1694700623
transform 1 0 26564 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_14
timestamp 1694700623
transform 1 0 26584 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_15
timestamp 1694700623
transform 1 0 21583 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_16
timestamp 1694700623
transform 1 0 21693 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_17
timestamp 1694700623
transform 1 0 21578 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_18
timestamp 1694700623
transform 1 0 21572 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_19
timestamp 1694700623
transform 1 0 21592 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_20
timestamp 1694700623
transform 1 0 16591 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_21
timestamp 1694700623
transform 1 0 16701 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_22
timestamp 1694700623
transform 1 0 16586 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_23
timestamp 1694700623
transform 1 0 16580 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_24
timestamp 1694700623
transform 1 0 16600 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_25
timestamp 1694700623
transform 1 0 11599 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_26
timestamp 1694700623
transform 1 0 11709 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_27
timestamp 1694700623
transform 1 0 11594 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_28
timestamp 1694700623
transform 1 0 11588 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_29
timestamp 1694700623
transform 1 0 11608 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_30
timestamp 1694700623
transform 1 0 6607 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_31
timestamp 1694700623
transform 1 0 6717 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_32
timestamp 1694700623
transform 1 0 6602 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_33
timestamp 1694700623
transform 1 0 6596 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_34
timestamp 1694700623
transform 1 0 6616 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_35
timestamp 1694700623
transform 1 0 1615 0 1 1546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_36
timestamp 1694700623
transform 1 0 1725 0 1 778
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_37
timestamp 1694700623
transform 1 0 1610 0 1 575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_38
timestamp 1694700623
transform 1 0 1604 0 1 1109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_21_39
timestamp 1694700623
transform 1 0 1624 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_0
timestamp 1694700623
transform 1 0 36552 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_1
timestamp 1694700623
transform 1 0 36662 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_2
timestamp 1694700623
transform 1 0 36547 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_3
timestamp 1694700623
transform 1 0 36541 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_4
timestamp 1694700623
transform 1 0 36561 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_5
timestamp 1694700623
transform 1 0 31560 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_6
timestamp 1694700623
transform 1 0 31670 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_7
timestamp 1694700623
transform 1 0 31555 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_8
timestamp 1694700623
transform 1 0 31549 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_9
timestamp 1694700623
transform 1 0 31569 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_10
timestamp 1694700623
transform 1 0 26568 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_11
timestamp 1694700623
transform 1 0 26678 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_12
timestamp 1694700623
transform 1 0 26563 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_13
timestamp 1694700623
transform 1 0 26557 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_14
timestamp 1694700623
transform 1 0 26577 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_15
timestamp 1694700623
transform 1 0 21576 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_16
timestamp 1694700623
transform 1 0 21686 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_17
timestamp 1694700623
transform 1 0 21571 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_18
timestamp 1694700623
transform 1 0 21565 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_19
timestamp 1694700623
transform 1 0 21585 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_20
timestamp 1694700623
transform 1 0 16584 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_21
timestamp 1694700623
transform 1 0 16694 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_22
timestamp 1694700623
transform 1 0 16579 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_23
timestamp 1694700623
transform 1 0 16573 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_24
timestamp 1694700623
transform 1 0 16593 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_25
timestamp 1694700623
transform 1 0 11592 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_26
timestamp 1694700623
transform 1 0 11702 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_27
timestamp 1694700623
transform 1 0 11587 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_28
timestamp 1694700623
transform 1 0 11581 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_29
timestamp 1694700623
transform 1 0 11601 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_30
timestamp 1694700623
transform 1 0 6600 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_31
timestamp 1694700623
transform 1 0 6710 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_32
timestamp 1694700623
transform 1 0 6595 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_33
timestamp 1694700623
transform 1 0 6589 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_34
timestamp 1694700623
transform 1 0 6609 0 1 154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_35
timestamp 1694700623
transform 1 0 1608 0 1 1541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_36
timestamp 1694700623
transform 1 0 1718 0 1 772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_37
timestamp 1694700623
transform 1 0 1603 0 1 570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_38
timestamp 1694700623
transform 1 0 1597 0 1 1104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_22_39
timestamp 1694700623
transform 1 0 1617 0 1 154
box 0 0 1 1
<< labels >>
rlabel metal3 s 6593 142 6691 240 4 vdd
port 1 nsew
rlabel metal3 s 11585 142 11683 240 4 vdd
port 1 nsew
rlabel metal3 s 16577 142 16675 240 4 vdd
port 1 nsew
rlabel metal3 s 26541 1092 26639 1190 4 vdd
port 1 nsew
rlabel metal3 s 21549 1092 21647 1190 4 vdd
port 1 nsew
rlabel metal3 s 36545 142 36643 240 4 vdd
port 1 nsew
rlabel metal3 s 26561 142 26659 240 4 vdd
port 1 nsew
rlabel metal3 s 6573 1092 6671 1190 4 vdd
port 1 nsew
rlabel metal3 s 36525 1092 36623 1190 4 vdd
port 1 nsew
rlabel metal3 s 31553 142 31651 240 4 vdd
port 1 nsew
rlabel metal3 s 16557 1092 16655 1190 4 vdd
port 1 nsew
rlabel metal3 s 11565 1092 11663 1190 4 vdd
port 1 nsew
rlabel metal3 s 1581 1092 1679 1190 4 vdd
port 1 nsew
rlabel metal3 s 21569 142 21667 240 4 vdd
port 1 nsew
rlabel metal3 s 31533 1092 31631 1190 4 vdd
port 1 nsew
rlabel metal3 s 1601 142 1699 240 4 vdd
port 1 nsew
rlabel metal3 s 11686 760 11784 858 4 gnd
port 2 nsew
rlabel metal3 s 21670 760 21768 858 4 gnd
port 2 nsew
rlabel metal3 s 1587 558 1685 656 4 gnd
port 2 nsew
rlabel metal3 s 21555 558 21653 656 4 gnd
port 2 nsew
rlabel metal3 s 31544 1529 31642 1627 4 gnd
port 2 nsew
rlabel metal3 s 36531 558 36629 656 4 gnd
port 2 nsew
rlabel metal3 s 31539 558 31637 656 4 gnd
port 2 nsew
rlabel metal3 s 26552 1529 26650 1627 4 gnd
port 2 nsew
rlabel metal3 s 1592 1529 1690 1627 4 gnd
port 2 nsew
rlabel metal3 s 6579 558 6677 656 4 gnd
port 2 nsew
rlabel metal3 s 31654 760 31752 858 4 gnd
port 2 nsew
rlabel metal3 s 6694 760 6792 858 4 gnd
port 2 nsew
rlabel metal3 s 16568 1529 16666 1627 4 gnd
port 2 nsew
rlabel metal3 s 26662 760 26760 858 4 gnd
port 2 nsew
rlabel metal3 s 1702 760 1800 858 4 gnd
port 2 nsew
rlabel metal3 s 6584 1529 6682 1627 4 gnd
port 2 nsew
rlabel metal3 s 11571 558 11669 656 4 gnd
port 2 nsew
rlabel metal3 s 16563 558 16661 656 4 gnd
port 2 nsew
rlabel metal3 s 21560 1529 21658 1627 4 gnd
port 2 nsew
rlabel metal3 s 26547 558 26645 656 4 gnd
port 2 nsew
rlabel metal3 s 36536 1529 36634 1627 4 gnd
port 2 nsew
rlabel metal3 s 16678 760 16776 858 4 gnd
port 2 nsew
rlabel metal3 s 11576 1529 11674 1627 4 gnd
port 2 nsew
rlabel metal3 s 36646 760 36744 858 4 gnd
port 2 nsew
rlabel metal1 s 1629 4 1689 60 4 data_0
port 3 nsew
rlabel metal1 s 1500 1959 1530 2011 4 bl_0
port 4 nsew
rlabel metal1 s 1702 1959 1732 2011 4 br_0
port 5 nsew
rlabel metal1 s 6621 4 6681 60 4 data_1
port 6 nsew
rlabel metal1 s 6492 1959 6522 2011 4 bl_1
port 7 nsew
rlabel metal1 s 6694 1959 6724 2011 4 br_1
port 8 nsew
rlabel metal1 s 11613 4 11673 60 4 data_2
port 9 nsew
rlabel metal1 s 11484 1959 11514 2011 4 bl_2
port 10 nsew
rlabel metal1 s 11686 1959 11716 2011 4 br_2
port 11 nsew
rlabel metal1 s 16605 4 16665 60 4 data_3
port 12 nsew
rlabel metal1 s 16476 1959 16506 2011 4 bl_3
port 13 nsew
rlabel metal1 s 16678 1959 16708 2011 4 br_3
port 14 nsew
rlabel metal1 s 21597 4 21657 60 4 data_4
port 15 nsew
rlabel metal1 s 21468 1959 21498 2011 4 bl_4
port 16 nsew
rlabel metal1 s 21670 1959 21700 2011 4 br_4
port 17 nsew
rlabel metal1 s 26589 4 26649 60 4 data_5
port 18 nsew
rlabel metal1 s 26460 1959 26490 2011 4 bl_5
port 19 nsew
rlabel metal1 s 26662 1959 26692 2011 4 br_5
port 20 nsew
rlabel metal1 s 31581 4 31641 60 4 data_6
port 21 nsew
rlabel metal1 s 31452 1959 31482 2011 4 bl_6
port 22 nsew
rlabel metal1 s 31654 1959 31684 2011 4 br_6
port 23 nsew
rlabel metal1 s 36573 4 36633 60 4 data_7
port 24 nsew
rlabel metal1 s 36444 1959 36474 2011 4 bl_7
port 25 nsew
rlabel metal1 s 36646 1959 36676 2011 4 br_7
port 26 nsew
rlabel metal1 s 1473 94 40785 128 4 en_0
port 27 nsew
<< properties >>
string FIXED_BBOX 0 0 36818 2011
string GDS_END 1072706
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 1052208
<< end >>
