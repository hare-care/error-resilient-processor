magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< dnwell >>
rect 11252 4817 20055 4870
rect 11208 3302 20055 4817
rect 2105 1401 9491 2545
rect 23973 1960 26586 2130
rect 2105 -406 18943 1401
rect 23973 751 28048 1960
rect 15534 -1206 18943 -406
rect 15552 -1280 18943 -1206
rect 25211 -2096 28048 751
rect 25161 -3505 28048 -2096
rect 23973 -10735 28048 -3505
<< nwell >>
rect 455 3027 7939 5038
rect 8416 4817 20135 4983
rect 8416 4138 11478 4817
rect 19025 4138 19270 4817
rect 19825 4138 20135 4817
rect 8416 3508 11414 4138
rect 19849 3508 20135 4138
rect 8416 3222 20135 3508
rect 8416 2980 11368 3222
rect 16905 3006 20135 3222
rect 8416 2902 10403 2980
rect 508 -2515 1640 2618
rect 2025 2339 9571 2625
rect 2025 -200 2311 2339
rect 9285 1481 9571 2339
rect 16905 2506 19165 3006
rect 19760 2470 20135 3006
rect 19760 1648 20278 2470
rect 23838 1924 28132 2159
rect 23838 1872 25371 1924
rect 9285 1195 19023 1481
rect 2025 -486 15758 -200
rect 15472 -1074 15758 -486
rect 18737 -1074 19023 1195
rect 15472 -1360 19023 -1074
rect 23838 1152 25277 1872
rect 26227 1754 28132 1924
rect 23838 -8171 24177 1152
rect 27114 1059 28132 1754
rect 26828 8 28132 1059
rect 26683 -1156 28132 8
rect 23838 -8355 24179 -8171
rect 26796 -8344 28132 -1156
rect 23838 -10178 24177 -8355
rect 23838 -10526 24912 -10178
rect 27144 -10480 28132 -8344
rect 26548 -10526 28132 -10480
rect 23838 -11477 28132 -10526
rect 2949 -17766 3443 -17034
rect 2506 -18981 3000 -17849
<< pwell >>
rect 11526 3572 19787 3658
rect 10462 2838 16470 2881
rect 2402 2193 7042 2279
rect 2402 2171 4450 2193
rect 2398 1042 4450 2171
rect 4636 1980 6688 2193
rect 7477 1980 8529 2271
rect 4636 1630 8553 1980
rect 4636 1042 6688 1630
rect 9690 2436 16470 2838
rect 9690 2320 19071 2436
rect 9690 1566 19611 2320
rect 2372 -10 7076 1042
rect 2372 -118 6948 -10
rect 7390 -35 7922 1417
rect 20226 1226 20312 1478
rect 13050 1060 15102 1103
rect 16318 1060 16420 1111
rect 8142 974 8228 992
rect 13050 974 16420 1060
rect 8142 722 16420 974
rect 8142 -78 12738 722
rect 13050 453 16420 722
rect 13050 203 15763 453
rect 16318 203 16420 453
rect 13050 57 16420 203
rect 12652 -121 12738 -78
rect 13092 -97 16420 57
rect 18370 -42 18622 372
rect 15850 -903 16420 -97
rect 15848 -1005 16420 -903
rect 25761 1176 25847 1811
rect 380 -11133 1099 -3205
rect 2590 -10210 3004 -9558
<< pmos >>
rect 916 4709 1716 4819
rect 1772 4709 1972 4819
rect 2028 4709 2228 4819
rect 2284 4709 2484 4819
rect 2540 4709 2740 4819
rect 2796 4709 2996 4819
rect 3052 4709 3252 4819
rect 3308 4709 3508 4819
rect 3564 4709 3764 4819
rect 3820 4709 4020 4819
rect 4076 4709 4276 4819
rect 4332 4709 4532 4819
rect 4588 4709 4788 4819
rect 4844 4709 5044 4819
rect 5100 4709 5300 4819
rect 5356 4709 5556 4819
rect 5612 4709 5812 4819
rect 5868 4709 6068 4819
rect 6124 4709 6324 4819
rect 6380 4709 6580 4819
rect 6636 4709 6836 4819
rect 6892 4709 7692 4819
rect 916 4291 1716 4401
rect 1772 4291 1972 4401
rect 2028 4291 2228 4401
rect 2284 4291 2484 4401
rect 2540 4291 2740 4401
rect 2796 4291 2996 4401
rect 3052 4291 3252 4401
rect 3308 4291 3508 4401
rect 3564 4291 3764 4401
rect 3820 4291 4020 4401
rect 4076 4291 4276 4401
rect 4332 4291 4532 4401
rect 4588 4291 4788 4401
rect 4844 4291 5044 4401
rect 5100 4291 5300 4401
rect 5356 4291 5556 4401
rect 5612 4291 5812 4401
rect 5868 4291 6068 4401
rect 6124 4291 6324 4401
rect 6380 4291 6580 4401
rect 6636 4291 6836 4401
rect 6892 4291 7692 4401
rect 916 3699 1716 3809
rect 1772 3699 1972 3809
rect 2028 3699 2228 3809
rect 2284 3699 2484 3809
rect 2540 3699 2740 3809
rect 2796 3699 2996 3809
rect 3052 3699 3252 3809
rect 3308 3699 3508 3809
rect 3564 3699 3764 3809
rect 3820 3699 4020 3809
rect 4076 3699 4276 3809
rect 4332 3699 4532 3809
rect 4588 3699 4788 3809
rect 4844 3699 5044 3809
rect 5100 3699 5300 3809
rect 5356 3699 5556 3809
rect 5612 3699 5812 3809
rect 5868 3699 6068 3809
rect 6124 3699 6324 3809
rect 6380 3699 6580 3809
rect 6636 3699 6836 3809
rect 6892 3699 7692 3809
rect 916 3281 1716 3391
rect 1772 3281 1972 3391
rect 2028 3281 2228 3391
rect 2284 3281 2484 3391
rect 2540 3281 2740 3391
rect 2796 3281 2996 3391
rect 3052 3281 3252 3391
rect 3308 3281 3508 3391
rect 3564 3281 3764 3391
rect 3820 3281 4020 3391
rect 4076 3281 4276 3391
rect 4332 3281 4532 3391
rect 4588 3281 4788 3391
rect 4844 3281 5044 3391
rect 5100 3281 5300 3391
rect 5356 3281 5556 3391
rect 5612 3281 5812 3391
rect 5868 3281 6068 3391
rect 6124 3281 6324 3391
rect 6380 3281 6580 3391
rect 6636 3281 6836 3391
rect 6892 3281 7692 3391
<< mvnmos >>
rect 7503 2092 8503 2192
rect 6874 1870 8474 1954
rect 6874 1656 8474 1740
rect 2451 16 2551 1016
rect 2607 16 2707 1016
rect 2763 16 2863 1016
rect 2919 16 3019 1016
rect 3075 16 3175 1016
rect 3231 16 3331 1016
rect 3387 16 3487 1016
rect 3543 16 3643 1016
rect 3823 16 3923 1016
rect 3979 16 4079 1016
rect 4135 16 4235 1016
rect 4291 16 4391 1016
rect 4447 16 4547 1016
rect 4603 16 4703 1016
rect 4759 16 4859 1016
rect 4915 16 5015 1016
rect 5071 16 5171 1016
rect 5227 16 5327 1016
rect 5383 16 5483 1016
rect 5713 16 5813 1016
rect 5869 16 5969 1016
rect 6025 16 6125 1016
rect 6181 16 6281 1016
rect 6461 16 6561 1016
rect 6741 16 6841 1016
rect 6897 16 6997 1016
rect 8329 -52 8429 948
rect 8485 -52 8585 948
rect 8641 -52 8741 948
rect 8797 -52 8897 948
rect 8953 -52 9053 948
rect 9109 -52 9209 948
rect 9265 -52 9365 948
rect 9421 -52 9521 948
rect 9577 -52 9677 948
rect 9733 -52 9833 948
rect 9889 -52 9989 948
rect 10045 -52 10145 948
rect 10201 -52 10301 948
rect 10357 -52 10457 948
rect 10782 -52 11182 948
rect 11238 -52 11638 948
rect 11694 -52 12094 948
rect 12150 -52 12550 948
rect 12828 748 12948 948
rect 18396 193 18596 293
rect 15929 -823 16029 177
rect 16085 -823 16185 177
rect 18396 37 18596 137
rect 2669 -10184 2769 -9584
rect 2825 -10184 2925 -9584
<< mvpmos >>
rect 8759 3804 8859 4804
rect 8915 3804 9015 4804
rect 9071 3804 9171 4804
rect 9227 3804 9327 4804
rect 9507 3804 9607 4804
rect 9787 3804 9887 4804
rect 9943 3804 10043 4804
rect 10376 3804 10476 4804
rect 10532 3804 10632 4804
rect 10688 3804 10788 4804
rect 10844 3804 10944 4804
rect 11000 3804 11100 4804
rect 10624 3477 10824 3561
rect 8893 3364 9893 3464
rect 8893 3208 9893 3308
rect 10152 3225 11152 3325
rect 16971 3064 17571 3184
rect 17843 3034 17943 3234
rect 17999 3034 18099 3234
rect 18327 3034 18427 3234
rect 18483 3034 18583 3234
rect 18789 3034 18889 3234
rect 18945 3034 19045 3234
rect 574 2288 1574 2388
rect 574 1696 1574 1796
rect 574 1540 1574 1640
rect 18086 2738 19086 2838
rect 574 1134 1574 1234
rect 574 978 1574 1078
rect 574 822 1574 922
rect 574 666 1574 766
rect 574 510 1574 610
rect 574 354 1574 454
rect 574 198 1574 298
rect 574 42 1574 142
rect 574 -114 1574 -14
rect 574 -270 1574 -170
rect 574 -426 1574 -326
rect 574 -582 1574 -482
rect 574 -738 1574 -638
rect 574 -1179 1574 -1079
rect 574 -1335 1574 -1235
rect 574 -1491 1574 -1391
rect 574 -1647 1574 -1547
rect 574 -1803 1574 -1703
rect 574 -1959 1574 -1859
rect 574 -2115 1574 -2015
rect 574 -2271 1574 -2171
rect 3068 -17700 3168 -17100
rect 3224 -17700 3324 -17100
rect 2625 -18915 2725 -17915
rect 2781 -18915 2881 -17915
<< mvnnmos >>
rect 2424 1912 4424 2092
rect 2424 1676 4424 1856
rect 4662 1912 6662 2092
rect 4662 1676 6662 1856
rect 2424 1440 4424 1620
rect 2424 1204 4424 1384
rect 4662 1204 6662 1384
rect 13076 844 15076 1024
rect 15268 834 15448 1034
rect 15504 834 15684 1034
rect 15740 834 15920 1034
rect 15976 834 16156 1034
rect 13076 608 15076 788
rect 13076 372 15076 552
rect 15268 479 15448 679
rect 15504 479 15684 679
rect 15740 479 15920 679
rect 15976 479 16156 679
rect 13076 136 15076 316
rect 15268 94 15448 294
rect 15504 94 15684 294
<< nmoslvt >>
rect 7469 -9 7499 1391
rect 7555 -9 7585 1391
rect 7641 -9 7671 1391
rect 7727 -9 7757 1391
rect 7813 -9 7843 1391
<< ndiff >>
rect 7416 1329 7469 1391
rect 7416 1295 7424 1329
rect 7458 1295 7469 1329
rect 7416 1261 7469 1295
rect 7416 1227 7424 1261
rect 7458 1227 7469 1261
rect 7416 1193 7469 1227
rect 7416 1159 7424 1193
rect 7458 1159 7469 1193
rect 7416 1125 7469 1159
rect 7416 1091 7424 1125
rect 7458 1091 7469 1125
rect 7416 1057 7469 1091
rect 7416 1023 7424 1057
rect 7458 1023 7469 1057
rect 7416 989 7469 1023
rect 7416 955 7424 989
rect 7458 955 7469 989
rect 7416 921 7469 955
rect 7416 887 7424 921
rect 7458 887 7469 921
rect 7416 853 7469 887
rect 7416 819 7424 853
rect 7458 819 7469 853
rect 7416 785 7469 819
rect 7416 751 7424 785
rect 7458 751 7469 785
rect 7416 717 7469 751
rect 7416 683 7424 717
rect 7458 683 7469 717
rect 7416 649 7469 683
rect 7416 615 7424 649
rect 7458 615 7469 649
rect 7416 581 7469 615
rect 7416 547 7424 581
rect 7458 547 7469 581
rect 7416 513 7469 547
rect 7416 479 7424 513
rect 7458 479 7469 513
rect 7416 445 7469 479
rect 7416 411 7424 445
rect 7458 411 7469 445
rect 7416 377 7469 411
rect 7416 343 7424 377
rect 7458 343 7469 377
rect 7416 309 7469 343
rect 7416 275 7424 309
rect 7458 275 7469 309
rect 7416 241 7469 275
rect 7416 207 7424 241
rect 7458 207 7469 241
rect 7416 173 7469 207
rect 7416 139 7424 173
rect 7458 139 7469 173
rect 7416 105 7469 139
rect 7416 71 7424 105
rect 7458 71 7469 105
rect 7416 37 7469 71
rect 7416 3 7424 37
rect 7458 3 7469 37
rect 7416 -9 7469 3
rect 7499 1329 7555 1391
rect 7499 1295 7510 1329
rect 7544 1295 7555 1329
rect 7499 1261 7555 1295
rect 7499 1227 7510 1261
rect 7544 1227 7555 1261
rect 7499 1193 7555 1227
rect 7499 1159 7510 1193
rect 7544 1159 7555 1193
rect 7499 1125 7555 1159
rect 7499 1091 7510 1125
rect 7544 1091 7555 1125
rect 7499 1057 7555 1091
rect 7499 1023 7510 1057
rect 7544 1023 7555 1057
rect 7499 989 7555 1023
rect 7499 955 7510 989
rect 7544 955 7555 989
rect 7499 921 7555 955
rect 7499 887 7510 921
rect 7544 887 7555 921
rect 7499 853 7555 887
rect 7499 819 7510 853
rect 7544 819 7555 853
rect 7499 785 7555 819
rect 7499 751 7510 785
rect 7544 751 7555 785
rect 7499 717 7555 751
rect 7499 683 7510 717
rect 7544 683 7555 717
rect 7499 649 7555 683
rect 7499 615 7510 649
rect 7544 615 7555 649
rect 7499 581 7555 615
rect 7499 547 7510 581
rect 7544 547 7555 581
rect 7499 513 7555 547
rect 7499 479 7510 513
rect 7544 479 7555 513
rect 7499 445 7555 479
rect 7499 411 7510 445
rect 7544 411 7555 445
rect 7499 377 7555 411
rect 7499 343 7510 377
rect 7544 343 7555 377
rect 7499 309 7555 343
rect 7499 275 7510 309
rect 7544 275 7555 309
rect 7499 241 7555 275
rect 7499 207 7510 241
rect 7544 207 7555 241
rect 7499 173 7555 207
rect 7499 139 7510 173
rect 7544 139 7555 173
rect 7499 105 7555 139
rect 7499 71 7510 105
rect 7544 71 7555 105
rect 7499 37 7555 71
rect 7499 3 7510 37
rect 7544 3 7555 37
rect 7499 -9 7555 3
rect 7585 1329 7641 1391
rect 7585 1295 7596 1329
rect 7630 1295 7641 1329
rect 7585 1261 7641 1295
rect 7585 1227 7596 1261
rect 7630 1227 7641 1261
rect 7585 1193 7641 1227
rect 7585 1159 7596 1193
rect 7630 1159 7641 1193
rect 7585 1125 7641 1159
rect 7585 1091 7596 1125
rect 7630 1091 7641 1125
rect 7585 1057 7641 1091
rect 7585 1023 7596 1057
rect 7630 1023 7641 1057
rect 7585 989 7641 1023
rect 7585 955 7596 989
rect 7630 955 7641 989
rect 7585 921 7641 955
rect 7585 887 7596 921
rect 7630 887 7641 921
rect 7585 853 7641 887
rect 7585 819 7596 853
rect 7630 819 7641 853
rect 7585 785 7641 819
rect 7585 751 7596 785
rect 7630 751 7641 785
rect 7585 717 7641 751
rect 7585 683 7596 717
rect 7630 683 7641 717
rect 7585 649 7641 683
rect 7585 615 7596 649
rect 7630 615 7641 649
rect 7585 581 7641 615
rect 7585 547 7596 581
rect 7630 547 7641 581
rect 7585 513 7641 547
rect 7585 479 7596 513
rect 7630 479 7641 513
rect 7585 445 7641 479
rect 7585 411 7596 445
rect 7630 411 7641 445
rect 7585 377 7641 411
rect 7585 343 7596 377
rect 7630 343 7641 377
rect 7585 309 7641 343
rect 7585 275 7596 309
rect 7630 275 7641 309
rect 7585 241 7641 275
rect 7585 207 7596 241
rect 7630 207 7641 241
rect 7585 173 7641 207
rect 7585 139 7596 173
rect 7630 139 7641 173
rect 7585 105 7641 139
rect 7585 71 7596 105
rect 7630 71 7641 105
rect 7585 37 7641 71
rect 7585 3 7596 37
rect 7630 3 7641 37
rect 7585 -9 7641 3
rect 7671 1329 7727 1391
rect 7671 1295 7682 1329
rect 7716 1295 7727 1329
rect 7671 1261 7727 1295
rect 7671 1227 7682 1261
rect 7716 1227 7727 1261
rect 7671 1193 7727 1227
rect 7671 1159 7682 1193
rect 7716 1159 7727 1193
rect 7671 1125 7727 1159
rect 7671 1091 7682 1125
rect 7716 1091 7727 1125
rect 7671 1057 7727 1091
rect 7671 1023 7682 1057
rect 7716 1023 7727 1057
rect 7671 989 7727 1023
rect 7671 955 7682 989
rect 7716 955 7727 989
rect 7671 921 7727 955
rect 7671 887 7682 921
rect 7716 887 7727 921
rect 7671 853 7727 887
rect 7671 819 7682 853
rect 7716 819 7727 853
rect 7671 785 7727 819
rect 7671 751 7682 785
rect 7716 751 7727 785
rect 7671 717 7727 751
rect 7671 683 7682 717
rect 7716 683 7727 717
rect 7671 649 7727 683
rect 7671 615 7682 649
rect 7716 615 7727 649
rect 7671 581 7727 615
rect 7671 547 7682 581
rect 7716 547 7727 581
rect 7671 513 7727 547
rect 7671 479 7682 513
rect 7716 479 7727 513
rect 7671 445 7727 479
rect 7671 411 7682 445
rect 7716 411 7727 445
rect 7671 377 7727 411
rect 7671 343 7682 377
rect 7716 343 7727 377
rect 7671 309 7727 343
rect 7671 275 7682 309
rect 7716 275 7727 309
rect 7671 241 7727 275
rect 7671 207 7682 241
rect 7716 207 7727 241
rect 7671 173 7727 207
rect 7671 139 7682 173
rect 7716 139 7727 173
rect 7671 105 7727 139
rect 7671 71 7682 105
rect 7716 71 7727 105
rect 7671 37 7727 71
rect 7671 3 7682 37
rect 7716 3 7727 37
rect 7671 -9 7727 3
rect 7757 1329 7813 1391
rect 7757 1295 7768 1329
rect 7802 1295 7813 1329
rect 7757 1261 7813 1295
rect 7757 1227 7768 1261
rect 7802 1227 7813 1261
rect 7757 1193 7813 1227
rect 7757 1159 7768 1193
rect 7802 1159 7813 1193
rect 7757 1125 7813 1159
rect 7757 1091 7768 1125
rect 7802 1091 7813 1125
rect 7757 1057 7813 1091
rect 7757 1023 7768 1057
rect 7802 1023 7813 1057
rect 7757 989 7813 1023
rect 7757 955 7768 989
rect 7802 955 7813 989
rect 7757 921 7813 955
rect 7757 887 7768 921
rect 7802 887 7813 921
rect 7757 853 7813 887
rect 7757 819 7768 853
rect 7802 819 7813 853
rect 7757 785 7813 819
rect 7757 751 7768 785
rect 7802 751 7813 785
rect 7757 717 7813 751
rect 7757 683 7768 717
rect 7802 683 7813 717
rect 7757 649 7813 683
rect 7757 615 7768 649
rect 7802 615 7813 649
rect 7757 581 7813 615
rect 7757 547 7768 581
rect 7802 547 7813 581
rect 7757 513 7813 547
rect 7757 479 7768 513
rect 7802 479 7813 513
rect 7757 445 7813 479
rect 7757 411 7768 445
rect 7802 411 7813 445
rect 7757 377 7813 411
rect 7757 343 7768 377
rect 7802 343 7813 377
rect 7757 309 7813 343
rect 7757 275 7768 309
rect 7802 275 7813 309
rect 7757 241 7813 275
rect 7757 207 7768 241
rect 7802 207 7813 241
rect 7757 173 7813 207
rect 7757 139 7768 173
rect 7802 139 7813 173
rect 7757 105 7813 139
rect 7757 71 7768 105
rect 7802 71 7813 105
rect 7757 37 7813 71
rect 7757 3 7768 37
rect 7802 3 7813 37
rect 7757 -9 7813 3
rect 7843 1329 7896 1391
rect 7843 1295 7854 1329
rect 7888 1295 7896 1329
rect 7843 1261 7896 1295
rect 7843 1227 7854 1261
rect 7888 1227 7896 1261
rect 7843 1193 7896 1227
rect 7843 1159 7854 1193
rect 7888 1159 7896 1193
rect 7843 1125 7896 1159
rect 7843 1091 7854 1125
rect 7888 1091 7896 1125
rect 7843 1057 7896 1091
rect 7843 1023 7854 1057
rect 7888 1023 7896 1057
rect 7843 989 7896 1023
rect 7843 955 7854 989
rect 7888 955 7896 989
rect 7843 921 7896 955
rect 7843 887 7854 921
rect 7888 887 7896 921
rect 7843 853 7896 887
rect 7843 819 7854 853
rect 7888 819 7896 853
rect 7843 785 7896 819
rect 7843 751 7854 785
rect 7888 751 7896 785
rect 7843 717 7896 751
rect 7843 683 7854 717
rect 7888 683 7896 717
rect 7843 649 7896 683
rect 7843 615 7854 649
rect 7888 615 7896 649
rect 7843 581 7896 615
rect 7843 547 7854 581
rect 7888 547 7896 581
rect 7843 513 7896 547
rect 7843 479 7854 513
rect 7888 479 7896 513
rect 7843 445 7896 479
rect 7843 411 7854 445
rect 7888 411 7896 445
rect 7843 377 7896 411
rect 7843 343 7854 377
rect 7888 343 7896 377
rect 7843 309 7896 343
rect 7843 275 7854 309
rect 7888 275 7896 309
rect 7843 241 7896 275
rect 7843 207 7854 241
rect 7888 207 7896 241
rect 7843 173 7896 207
rect 7843 139 7854 173
rect 7888 139 7896 173
rect 7843 105 7896 139
rect 7843 71 7854 105
rect 7888 71 7896 105
rect 7843 37 7896 71
rect 7843 3 7854 37
rect 7888 3 7896 37
rect 7843 -9 7896 3
<< pdiff >>
rect 863 4807 916 4819
rect 863 4773 871 4807
rect 905 4773 916 4807
rect 863 4709 916 4773
rect 1716 4807 1772 4819
rect 1716 4773 1727 4807
rect 1761 4773 1772 4807
rect 1716 4709 1772 4773
rect 1972 4807 2028 4819
rect 1972 4773 1983 4807
rect 2017 4773 2028 4807
rect 1972 4709 2028 4773
rect 2228 4807 2284 4819
rect 2228 4773 2239 4807
rect 2273 4773 2284 4807
rect 2228 4709 2284 4773
rect 2484 4807 2540 4819
rect 2484 4773 2495 4807
rect 2529 4773 2540 4807
rect 2484 4709 2540 4773
rect 2740 4807 2796 4819
rect 2740 4773 2751 4807
rect 2785 4773 2796 4807
rect 2740 4709 2796 4773
rect 2996 4807 3052 4819
rect 2996 4773 3007 4807
rect 3041 4773 3052 4807
rect 2996 4709 3052 4773
rect 3252 4807 3308 4819
rect 3252 4773 3263 4807
rect 3297 4773 3308 4807
rect 3252 4709 3308 4773
rect 3508 4807 3564 4819
rect 3508 4773 3519 4807
rect 3553 4773 3564 4807
rect 3508 4709 3564 4773
rect 3764 4807 3820 4819
rect 3764 4773 3775 4807
rect 3809 4773 3820 4807
rect 3764 4709 3820 4773
rect 4020 4807 4076 4819
rect 4020 4773 4031 4807
rect 4065 4773 4076 4807
rect 4020 4709 4076 4773
rect 4276 4807 4332 4819
rect 4276 4773 4287 4807
rect 4321 4773 4332 4807
rect 4276 4709 4332 4773
rect 4532 4807 4588 4819
rect 4532 4773 4543 4807
rect 4577 4773 4588 4807
rect 4532 4709 4588 4773
rect 4788 4807 4844 4819
rect 4788 4773 4799 4807
rect 4833 4773 4844 4807
rect 4788 4709 4844 4773
rect 5044 4807 5100 4819
rect 5044 4773 5055 4807
rect 5089 4773 5100 4807
rect 5044 4709 5100 4773
rect 5300 4807 5356 4819
rect 5300 4773 5311 4807
rect 5345 4773 5356 4807
rect 5300 4709 5356 4773
rect 5556 4807 5612 4819
rect 5556 4773 5567 4807
rect 5601 4773 5612 4807
rect 5556 4709 5612 4773
rect 5812 4807 5868 4819
rect 5812 4773 5823 4807
rect 5857 4773 5868 4807
rect 5812 4709 5868 4773
rect 6068 4807 6124 4819
rect 6068 4773 6079 4807
rect 6113 4773 6124 4807
rect 6068 4709 6124 4773
rect 6324 4807 6380 4819
rect 6324 4773 6335 4807
rect 6369 4773 6380 4807
rect 6324 4709 6380 4773
rect 6580 4807 6636 4819
rect 6580 4773 6591 4807
rect 6625 4773 6636 4807
rect 6580 4709 6636 4773
rect 6836 4807 6892 4819
rect 6836 4773 6847 4807
rect 6881 4773 6892 4807
rect 6836 4709 6892 4773
rect 7692 4807 7745 4819
rect 7692 4773 7703 4807
rect 7737 4773 7745 4807
rect 7692 4709 7745 4773
rect 863 4337 916 4401
rect 863 4303 871 4337
rect 905 4303 916 4337
rect 863 4291 916 4303
rect 1716 4337 1772 4401
rect 1716 4303 1727 4337
rect 1761 4303 1772 4337
rect 1716 4291 1772 4303
rect 1972 4337 2028 4401
rect 1972 4303 1983 4337
rect 2017 4303 2028 4337
rect 1972 4291 2028 4303
rect 2228 4337 2284 4401
rect 2228 4303 2239 4337
rect 2273 4303 2284 4337
rect 2228 4291 2284 4303
rect 2484 4337 2540 4401
rect 2484 4303 2495 4337
rect 2529 4303 2540 4337
rect 2484 4291 2540 4303
rect 2740 4337 2796 4401
rect 2740 4303 2751 4337
rect 2785 4303 2796 4337
rect 2740 4291 2796 4303
rect 2996 4337 3052 4401
rect 2996 4303 3007 4337
rect 3041 4303 3052 4337
rect 2996 4291 3052 4303
rect 3252 4337 3308 4401
rect 3252 4303 3263 4337
rect 3297 4303 3308 4337
rect 3252 4291 3308 4303
rect 3508 4337 3564 4401
rect 3508 4303 3519 4337
rect 3553 4303 3564 4337
rect 3508 4291 3564 4303
rect 3764 4337 3820 4401
rect 3764 4303 3775 4337
rect 3809 4303 3820 4337
rect 3764 4291 3820 4303
rect 4020 4337 4076 4401
rect 4020 4303 4031 4337
rect 4065 4303 4076 4337
rect 4020 4291 4076 4303
rect 4276 4337 4332 4401
rect 4276 4303 4287 4337
rect 4321 4303 4332 4337
rect 4276 4291 4332 4303
rect 4532 4337 4588 4401
rect 4532 4303 4543 4337
rect 4577 4303 4588 4337
rect 4532 4291 4588 4303
rect 4788 4337 4844 4401
rect 4788 4303 4799 4337
rect 4833 4303 4844 4337
rect 4788 4291 4844 4303
rect 5044 4337 5100 4401
rect 5044 4303 5055 4337
rect 5089 4303 5100 4337
rect 5044 4291 5100 4303
rect 5300 4337 5356 4401
rect 5300 4303 5311 4337
rect 5345 4303 5356 4337
rect 5300 4291 5356 4303
rect 5556 4337 5612 4401
rect 5556 4303 5567 4337
rect 5601 4303 5612 4337
rect 5556 4291 5612 4303
rect 5812 4337 5868 4401
rect 5812 4303 5823 4337
rect 5857 4303 5868 4337
rect 5812 4291 5868 4303
rect 6068 4337 6124 4401
rect 6068 4303 6079 4337
rect 6113 4303 6124 4337
rect 6068 4291 6124 4303
rect 6324 4337 6380 4401
rect 6324 4303 6335 4337
rect 6369 4303 6380 4337
rect 6324 4291 6380 4303
rect 6580 4337 6636 4401
rect 6580 4303 6591 4337
rect 6625 4303 6636 4337
rect 6580 4291 6636 4303
rect 6836 4337 6892 4401
rect 6836 4303 6847 4337
rect 6881 4303 6892 4337
rect 6836 4291 6892 4303
rect 7692 4337 7745 4401
rect 7692 4303 7703 4337
rect 7737 4303 7745 4337
rect 7692 4291 7745 4303
rect 863 3797 916 3809
rect 863 3763 871 3797
rect 905 3763 916 3797
rect 863 3699 916 3763
rect 1716 3797 1772 3809
rect 1716 3763 1727 3797
rect 1761 3763 1772 3797
rect 1716 3699 1772 3763
rect 1972 3797 2028 3809
rect 1972 3763 1983 3797
rect 2017 3763 2028 3797
rect 1972 3699 2028 3763
rect 2228 3797 2284 3809
rect 2228 3763 2239 3797
rect 2273 3763 2284 3797
rect 2228 3699 2284 3763
rect 2484 3797 2540 3809
rect 2484 3763 2495 3797
rect 2529 3763 2540 3797
rect 2484 3699 2540 3763
rect 2740 3797 2796 3809
rect 2740 3763 2751 3797
rect 2785 3763 2796 3797
rect 2740 3699 2796 3763
rect 2996 3797 3052 3809
rect 2996 3763 3007 3797
rect 3041 3763 3052 3797
rect 2996 3699 3052 3763
rect 3252 3797 3308 3809
rect 3252 3763 3263 3797
rect 3297 3763 3308 3797
rect 3252 3699 3308 3763
rect 3508 3797 3564 3809
rect 3508 3763 3519 3797
rect 3553 3763 3564 3797
rect 3508 3699 3564 3763
rect 3764 3797 3820 3809
rect 3764 3763 3775 3797
rect 3809 3763 3820 3797
rect 3764 3699 3820 3763
rect 4020 3797 4076 3809
rect 4020 3763 4031 3797
rect 4065 3763 4076 3797
rect 4020 3699 4076 3763
rect 4276 3797 4332 3809
rect 4276 3763 4287 3797
rect 4321 3763 4332 3797
rect 4276 3699 4332 3763
rect 4532 3797 4588 3809
rect 4532 3763 4543 3797
rect 4577 3763 4588 3797
rect 4532 3699 4588 3763
rect 4788 3797 4844 3809
rect 4788 3763 4799 3797
rect 4833 3763 4844 3797
rect 4788 3699 4844 3763
rect 5044 3797 5100 3809
rect 5044 3763 5055 3797
rect 5089 3763 5100 3797
rect 5044 3699 5100 3763
rect 5300 3797 5356 3809
rect 5300 3763 5311 3797
rect 5345 3763 5356 3797
rect 5300 3699 5356 3763
rect 5556 3797 5612 3809
rect 5556 3763 5567 3797
rect 5601 3763 5612 3797
rect 5556 3699 5612 3763
rect 5812 3797 5868 3809
rect 5812 3763 5823 3797
rect 5857 3763 5868 3797
rect 5812 3699 5868 3763
rect 6068 3797 6124 3809
rect 6068 3763 6079 3797
rect 6113 3763 6124 3797
rect 6068 3699 6124 3763
rect 6324 3797 6380 3809
rect 6324 3763 6335 3797
rect 6369 3763 6380 3797
rect 6324 3699 6380 3763
rect 6580 3797 6636 3809
rect 6580 3763 6591 3797
rect 6625 3763 6636 3797
rect 6580 3699 6636 3763
rect 6836 3797 6892 3809
rect 6836 3763 6847 3797
rect 6881 3763 6892 3797
rect 6836 3699 6892 3763
rect 7692 3797 7745 3809
rect 7692 3763 7703 3797
rect 7737 3763 7745 3797
rect 7692 3699 7745 3763
rect 863 3327 916 3391
rect 863 3293 871 3327
rect 905 3293 916 3327
rect 863 3281 916 3293
rect 1716 3327 1772 3391
rect 1716 3293 1727 3327
rect 1761 3293 1772 3327
rect 1716 3281 1772 3293
rect 1972 3327 2028 3391
rect 1972 3293 1983 3327
rect 2017 3293 2028 3327
rect 1972 3281 2028 3293
rect 2228 3327 2284 3391
rect 2228 3293 2239 3327
rect 2273 3293 2284 3327
rect 2228 3281 2284 3293
rect 2484 3327 2540 3391
rect 2484 3293 2495 3327
rect 2529 3293 2540 3327
rect 2484 3281 2540 3293
rect 2740 3327 2796 3391
rect 2740 3293 2751 3327
rect 2785 3293 2796 3327
rect 2740 3281 2796 3293
rect 2996 3327 3052 3391
rect 2996 3293 3007 3327
rect 3041 3293 3052 3327
rect 2996 3281 3052 3293
rect 3252 3327 3308 3391
rect 3252 3293 3263 3327
rect 3297 3293 3308 3327
rect 3252 3281 3308 3293
rect 3508 3327 3564 3391
rect 3508 3293 3519 3327
rect 3553 3293 3564 3327
rect 3508 3281 3564 3293
rect 3764 3327 3820 3391
rect 3764 3293 3775 3327
rect 3809 3293 3820 3327
rect 3764 3281 3820 3293
rect 4020 3327 4076 3391
rect 4020 3293 4031 3327
rect 4065 3293 4076 3327
rect 4020 3281 4076 3293
rect 4276 3327 4332 3391
rect 4276 3293 4287 3327
rect 4321 3293 4332 3327
rect 4276 3281 4332 3293
rect 4532 3327 4588 3391
rect 4532 3293 4543 3327
rect 4577 3293 4588 3327
rect 4532 3281 4588 3293
rect 4788 3327 4844 3391
rect 4788 3293 4799 3327
rect 4833 3293 4844 3327
rect 4788 3281 4844 3293
rect 5044 3327 5100 3391
rect 5044 3293 5055 3327
rect 5089 3293 5100 3327
rect 5044 3281 5100 3293
rect 5300 3327 5356 3391
rect 5300 3293 5311 3327
rect 5345 3293 5356 3327
rect 5300 3281 5356 3293
rect 5556 3327 5612 3391
rect 5556 3293 5567 3327
rect 5601 3293 5612 3327
rect 5556 3281 5612 3293
rect 5812 3327 5868 3391
rect 5812 3293 5823 3327
rect 5857 3293 5868 3327
rect 5812 3281 5868 3293
rect 6068 3327 6124 3391
rect 6068 3293 6079 3327
rect 6113 3293 6124 3327
rect 6068 3281 6124 3293
rect 6324 3327 6380 3391
rect 6324 3293 6335 3327
rect 6369 3293 6380 3327
rect 6324 3281 6380 3293
rect 6580 3327 6636 3391
rect 6580 3293 6591 3327
rect 6625 3293 6636 3327
rect 6580 3281 6636 3293
rect 6836 3327 6892 3391
rect 6836 3293 6847 3327
rect 6881 3293 6892 3327
rect 6836 3281 6892 3293
rect 7692 3327 7745 3391
rect 7692 3293 7703 3327
rect 7737 3293 7745 3327
rect 7692 3281 7745 3293
<< mvndiff >>
rect 7503 2237 8503 2245
rect 7503 2203 7515 2237
rect 7549 2203 7583 2237
rect 7617 2203 7651 2237
rect 7685 2203 7719 2237
rect 7753 2203 7787 2237
rect 7821 2203 7855 2237
rect 7889 2203 7923 2237
rect 7957 2203 7991 2237
rect 8025 2203 8059 2237
rect 8093 2203 8127 2237
rect 8161 2203 8195 2237
rect 8229 2203 8263 2237
rect 8297 2203 8331 2237
rect 8365 2203 8399 2237
rect 8433 2203 8503 2237
rect 7503 2192 8503 2203
rect 2424 2137 4424 2145
rect 2424 2103 2436 2137
rect 2470 2103 2504 2137
rect 2538 2103 2572 2137
rect 2606 2103 2640 2137
rect 2674 2103 2708 2137
rect 2742 2103 2776 2137
rect 2810 2103 2844 2137
rect 2878 2103 2912 2137
rect 2946 2103 2980 2137
rect 3014 2103 3048 2137
rect 3082 2103 3116 2137
rect 3150 2103 3184 2137
rect 3218 2103 3252 2137
rect 3286 2103 3320 2137
rect 3354 2103 3388 2137
rect 3422 2103 3456 2137
rect 3490 2103 3524 2137
rect 3558 2103 3592 2137
rect 3626 2103 3660 2137
rect 3694 2103 3728 2137
rect 3762 2103 3796 2137
rect 3830 2103 3864 2137
rect 3898 2103 3932 2137
rect 3966 2103 4000 2137
rect 4034 2103 4068 2137
rect 4102 2103 4136 2137
rect 4170 2103 4204 2137
rect 4238 2103 4272 2137
rect 4306 2103 4340 2137
rect 4374 2103 4424 2137
rect 2424 2092 4424 2103
rect 4662 2137 6662 2145
rect 4662 2103 4712 2137
rect 4746 2103 4780 2137
rect 4814 2103 4848 2137
rect 4882 2103 4916 2137
rect 4950 2103 4984 2137
rect 5018 2103 5052 2137
rect 5086 2103 5120 2137
rect 5154 2103 5188 2137
rect 5222 2103 5256 2137
rect 5290 2103 5324 2137
rect 5358 2103 5392 2137
rect 5426 2103 5460 2137
rect 5494 2103 5528 2137
rect 5562 2103 5596 2137
rect 5630 2103 5664 2137
rect 5698 2103 5732 2137
rect 5766 2103 5800 2137
rect 5834 2103 5868 2137
rect 5902 2103 5936 2137
rect 5970 2103 6004 2137
rect 6038 2103 6072 2137
rect 6106 2103 6140 2137
rect 6174 2103 6208 2137
rect 6242 2103 6276 2137
rect 6310 2103 6344 2137
rect 6378 2103 6412 2137
rect 6446 2103 6480 2137
rect 6514 2103 6548 2137
rect 6582 2103 6616 2137
rect 6650 2103 6662 2137
rect 4662 2092 6662 2103
rect 2424 1901 4424 1912
rect 2424 1867 2436 1901
rect 2470 1867 2504 1901
rect 2538 1867 2572 1901
rect 2606 1867 2640 1901
rect 2674 1867 2708 1901
rect 2742 1867 2776 1901
rect 2810 1867 2844 1901
rect 2878 1867 2912 1901
rect 2946 1867 2980 1901
rect 3014 1867 3048 1901
rect 3082 1867 3116 1901
rect 3150 1867 3184 1901
rect 3218 1867 3252 1901
rect 3286 1867 3320 1901
rect 3354 1867 3388 1901
rect 3422 1867 3456 1901
rect 3490 1867 3524 1901
rect 3558 1867 3592 1901
rect 3626 1867 3660 1901
rect 3694 1867 3728 1901
rect 3762 1867 3796 1901
rect 3830 1867 3864 1901
rect 3898 1867 3932 1901
rect 3966 1867 4000 1901
rect 4034 1867 4068 1901
rect 4102 1867 4136 1901
rect 4170 1867 4204 1901
rect 4238 1867 4272 1901
rect 4306 1867 4340 1901
rect 4374 1867 4424 1901
rect 2424 1856 4424 1867
rect 7503 2081 8503 2092
rect 7503 2047 7515 2081
rect 7549 2047 7583 2081
rect 7617 2047 7651 2081
rect 7685 2047 7719 2081
rect 7753 2047 7787 2081
rect 7821 2047 7855 2081
rect 7889 2047 7923 2081
rect 7957 2047 7991 2081
rect 8025 2047 8059 2081
rect 8093 2047 8127 2081
rect 8161 2047 8195 2081
rect 8229 2047 8263 2081
rect 8297 2047 8331 2081
rect 8365 2047 8399 2081
rect 8433 2047 8503 2081
rect 7503 2039 8503 2047
rect 6821 1942 6874 1954
rect 4662 1901 6662 1912
rect 4662 1867 4712 1901
rect 4746 1867 4780 1901
rect 4814 1867 4848 1901
rect 4882 1867 4916 1901
rect 4950 1867 4984 1901
rect 5018 1867 5052 1901
rect 5086 1867 5120 1901
rect 5154 1867 5188 1901
rect 5222 1867 5256 1901
rect 5290 1867 5324 1901
rect 5358 1867 5392 1901
rect 5426 1867 5460 1901
rect 5494 1867 5528 1901
rect 5562 1867 5596 1901
rect 5630 1867 5664 1901
rect 5698 1867 5732 1901
rect 5766 1867 5800 1901
rect 5834 1867 5868 1901
rect 5902 1867 5936 1901
rect 5970 1867 6004 1901
rect 6038 1867 6072 1901
rect 6106 1867 6140 1901
rect 6174 1867 6208 1901
rect 6242 1867 6276 1901
rect 6310 1867 6344 1901
rect 6378 1867 6412 1901
rect 6446 1867 6480 1901
rect 6514 1867 6548 1901
rect 6582 1867 6616 1901
rect 6650 1867 6662 1901
rect 6821 1908 6829 1942
rect 6863 1908 6874 1942
rect 6821 1870 6874 1908
rect 8474 1942 8527 1954
rect 8474 1908 8485 1942
rect 8519 1908 8527 1942
rect 8474 1870 8527 1908
rect 4662 1856 6662 1867
rect 6821 1702 6874 1740
rect 2424 1665 4424 1676
rect 2424 1631 2436 1665
rect 2470 1631 2504 1665
rect 2538 1631 2572 1665
rect 2606 1631 2640 1665
rect 2674 1631 2708 1665
rect 2742 1631 2776 1665
rect 2810 1631 2844 1665
rect 2878 1631 2912 1665
rect 2946 1631 2980 1665
rect 3014 1631 3048 1665
rect 3082 1631 3116 1665
rect 3150 1631 3184 1665
rect 3218 1631 3252 1665
rect 3286 1631 3320 1665
rect 3354 1631 3388 1665
rect 3422 1631 3456 1665
rect 3490 1631 3524 1665
rect 3558 1631 3592 1665
rect 3626 1631 3660 1665
rect 3694 1631 3728 1665
rect 3762 1631 3796 1665
rect 3830 1631 3864 1665
rect 3898 1631 3932 1665
rect 3966 1631 4000 1665
rect 4034 1631 4068 1665
rect 4102 1631 4136 1665
rect 4170 1631 4204 1665
rect 4238 1631 4272 1665
rect 4306 1631 4340 1665
rect 4374 1631 4424 1665
rect 2424 1620 4424 1631
rect 4662 1665 6662 1676
rect 4662 1631 4712 1665
rect 4746 1631 4780 1665
rect 4814 1631 4848 1665
rect 4882 1631 4916 1665
rect 4950 1631 4984 1665
rect 5018 1631 5052 1665
rect 5086 1631 5120 1665
rect 5154 1631 5188 1665
rect 5222 1631 5256 1665
rect 5290 1631 5324 1665
rect 5358 1631 5392 1665
rect 5426 1631 5460 1665
rect 5494 1631 5528 1665
rect 5562 1631 5596 1665
rect 5630 1631 5664 1665
rect 5698 1631 5732 1665
rect 5766 1631 5800 1665
rect 5834 1631 5868 1665
rect 5902 1631 5936 1665
rect 5970 1631 6004 1665
rect 6038 1631 6072 1665
rect 6106 1631 6140 1665
rect 6174 1631 6208 1665
rect 6242 1631 6276 1665
rect 6310 1631 6344 1665
rect 6378 1631 6412 1665
rect 6446 1631 6480 1665
rect 6514 1631 6548 1665
rect 6582 1631 6616 1665
rect 6650 1631 6662 1665
rect 6821 1668 6829 1702
rect 6863 1668 6874 1702
rect 6821 1656 6874 1668
rect 8474 1702 8527 1740
rect 8474 1668 8485 1702
rect 8519 1668 8527 1702
rect 8474 1656 8527 1668
rect 4662 1623 6662 1631
rect 10626 2710 10671 2743
rect 10626 2676 10637 2710
rect 10626 2643 10671 2676
rect 10626 2188 10668 2221
rect 10626 2154 10634 2188
rect 10626 2121 10668 2154
rect 2424 1429 4424 1440
rect 2424 1395 2436 1429
rect 2470 1395 2504 1429
rect 2538 1395 2572 1429
rect 2606 1395 2640 1429
rect 2674 1395 2708 1429
rect 2742 1395 2776 1429
rect 2810 1395 2844 1429
rect 2878 1395 2912 1429
rect 2946 1395 2980 1429
rect 3014 1395 3048 1429
rect 3082 1395 3116 1429
rect 3150 1395 3184 1429
rect 3218 1395 3252 1429
rect 3286 1395 3320 1429
rect 3354 1395 3388 1429
rect 3422 1395 3456 1429
rect 3490 1395 3524 1429
rect 3558 1395 3592 1429
rect 3626 1395 3660 1429
rect 3694 1395 3728 1429
rect 3762 1395 3796 1429
rect 3830 1395 3864 1429
rect 3898 1395 3932 1429
rect 3966 1395 4000 1429
rect 4034 1395 4068 1429
rect 4102 1395 4136 1429
rect 4170 1395 4204 1429
rect 4238 1395 4272 1429
rect 4306 1395 4340 1429
rect 4374 1395 4424 1429
rect 2424 1384 4424 1395
rect 4662 1429 6662 1437
rect 4662 1395 4712 1429
rect 4746 1395 4780 1429
rect 4814 1395 4848 1429
rect 4882 1395 4916 1429
rect 4950 1395 4984 1429
rect 5018 1395 5052 1429
rect 5086 1395 5120 1429
rect 5154 1395 5188 1429
rect 5222 1395 5256 1429
rect 5290 1395 5324 1429
rect 5358 1395 5392 1429
rect 5426 1395 5460 1429
rect 5494 1395 5528 1429
rect 5562 1395 5596 1429
rect 5630 1395 5664 1429
rect 5698 1395 5732 1429
rect 5766 1395 5800 1429
rect 5834 1395 5868 1429
rect 5902 1395 5936 1429
rect 5970 1395 6004 1429
rect 6038 1395 6072 1429
rect 6106 1395 6140 1429
rect 6174 1395 6208 1429
rect 6242 1395 6276 1429
rect 6310 1395 6344 1429
rect 6378 1395 6412 1429
rect 6446 1395 6480 1429
rect 6514 1395 6548 1429
rect 6582 1395 6616 1429
rect 6650 1395 6662 1429
rect 4662 1384 6662 1395
rect 2424 1193 4424 1204
rect 2424 1159 2436 1193
rect 2470 1159 2504 1193
rect 2538 1159 2572 1193
rect 2606 1159 2640 1193
rect 2674 1159 2708 1193
rect 2742 1159 2776 1193
rect 2810 1159 2844 1193
rect 2878 1159 2912 1193
rect 2946 1159 2980 1193
rect 3014 1159 3048 1193
rect 3082 1159 3116 1193
rect 3150 1159 3184 1193
rect 3218 1159 3252 1193
rect 3286 1159 3320 1193
rect 3354 1159 3388 1193
rect 3422 1159 3456 1193
rect 3490 1159 3524 1193
rect 3558 1159 3592 1193
rect 3626 1159 3660 1193
rect 3694 1159 3728 1193
rect 3762 1159 3796 1193
rect 3830 1159 3864 1193
rect 3898 1159 3932 1193
rect 3966 1159 4000 1193
rect 4034 1159 4068 1193
rect 4102 1159 4136 1193
rect 4170 1159 4204 1193
rect 4238 1159 4272 1193
rect 4306 1159 4340 1193
rect 4374 1159 4424 1193
rect 2424 1151 4424 1159
rect 4662 1193 6662 1204
rect 4662 1159 4712 1193
rect 4746 1159 4780 1193
rect 4814 1159 4848 1193
rect 4882 1159 4916 1193
rect 4950 1159 4984 1193
rect 5018 1159 5052 1193
rect 5086 1159 5120 1193
rect 5154 1159 5188 1193
rect 5222 1159 5256 1193
rect 5290 1159 5324 1193
rect 5358 1159 5392 1193
rect 5426 1159 5460 1193
rect 5494 1159 5528 1193
rect 5562 1159 5596 1193
rect 5630 1159 5664 1193
rect 5698 1159 5732 1193
rect 5766 1159 5800 1193
rect 5834 1159 5868 1193
rect 5902 1159 5936 1193
rect 5970 1159 6004 1193
rect 6038 1159 6072 1193
rect 6106 1159 6140 1193
rect 6174 1159 6208 1193
rect 6242 1159 6276 1193
rect 6310 1159 6344 1193
rect 6378 1159 6412 1193
rect 6446 1159 6480 1193
rect 6514 1159 6548 1193
rect 6582 1159 6616 1193
rect 6650 1159 6662 1193
rect 4662 1151 6662 1159
rect 2398 946 2451 1016
rect 2398 912 2406 946
rect 2440 912 2451 946
rect 2398 878 2451 912
rect 2398 844 2406 878
rect 2440 844 2451 878
rect 2398 810 2451 844
rect 2398 776 2406 810
rect 2440 776 2451 810
rect 2398 742 2451 776
rect 2398 708 2406 742
rect 2440 708 2451 742
rect 2398 674 2451 708
rect 2398 640 2406 674
rect 2440 640 2451 674
rect 2398 606 2451 640
rect 2398 572 2406 606
rect 2440 572 2451 606
rect 2398 538 2451 572
rect 2398 504 2406 538
rect 2440 504 2451 538
rect 2398 470 2451 504
rect 2398 436 2406 470
rect 2440 436 2451 470
rect 2398 402 2451 436
rect 2398 368 2406 402
rect 2440 368 2451 402
rect 2398 334 2451 368
rect 2398 300 2406 334
rect 2440 300 2451 334
rect 2398 266 2451 300
rect 2398 232 2406 266
rect 2440 232 2451 266
rect 2398 198 2451 232
rect 2398 164 2406 198
rect 2440 164 2451 198
rect 2398 130 2451 164
rect 2398 96 2406 130
rect 2440 96 2451 130
rect 2398 62 2451 96
rect 2398 28 2406 62
rect 2440 28 2451 62
rect 2398 16 2451 28
rect 2551 946 2607 1016
rect 2551 912 2562 946
rect 2596 912 2607 946
rect 2551 878 2607 912
rect 2551 844 2562 878
rect 2596 844 2607 878
rect 2551 810 2607 844
rect 2551 776 2562 810
rect 2596 776 2607 810
rect 2551 742 2607 776
rect 2551 708 2562 742
rect 2596 708 2607 742
rect 2551 674 2607 708
rect 2551 640 2562 674
rect 2596 640 2607 674
rect 2551 606 2607 640
rect 2551 572 2562 606
rect 2596 572 2607 606
rect 2551 538 2607 572
rect 2551 504 2562 538
rect 2596 504 2607 538
rect 2551 470 2607 504
rect 2551 436 2562 470
rect 2596 436 2607 470
rect 2551 402 2607 436
rect 2551 368 2562 402
rect 2596 368 2607 402
rect 2551 334 2607 368
rect 2551 300 2562 334
rect 2596 300 2607 334
rect 2551 266 2607 300
rect 2551 232 2562 266
rect 2596 232 2607 266
rect 2551 198 2607 232
rect 2551 164 2562 198
rect 2596 164 2607 198
rect 2551 130 2607 164
rect 2551 96 2562 130
rect 2596 96 2607 130
rect 2551 62 2607 96
rect 2551 28 2562 62
rect 2596 28 2607 62
rect 2551 16 2607 28
rect 2707 946 2763 1016
rect 2707 912 2718 946
rect 2752 912 2763 946
rect 2707 878 2763 912
rect 2707 844 2718 878
rect 2752 844 2763 878
rect 2707 810 2763 844
rect 2707 776 2718 810
rect 2752 776 2763 810
rect 2707 742 2763 776
rect 2707 708 2718 742
rect 2752 708 2763 742
rect 2707 674 2763 708
rect 2707 640 2718 674
rect 2752 640 2763 674
rect 2707 606 2763 640
rect 2707 572 2718 606
rect 2752 572 2763 606
rect 2707 538 2763 572
rect 2707 504 2718 538
rect 2752 504 2763 538
rect 2707 470 2763 504
rect 2707 436 2718 470
rect 2752 436 2763 470
rect 2707 402 2763 436
rect 2707 368 2718 402
rect 2752 368 2763 402
rect 2707 334 2763 368
rect 2707 300 2718 334
rect 2752 300 2763 334
rect 2707 266 2763 300
rect 2707 232 2718 266
rect 2752 232 2763 266
rect 2707 198 2763 232
rect 2707 164 2718 198
rect 2752 164 2763 198
rect 2707 130 2763 164
rect 2707 96 2718 130
rect 2752 96 2763 130
rect 2707 62 2763 96
rect 2707 28 2718 62
rect 2752 28 2763 62
rect 2707 16 2763 28
rect 2863 946 2919 1016
rect 2863 912 2874 946
rect 2908 912 2919 946
rect 2863 878 2919 912
rect 2863 844 2874 878
rect 2908 844 2919 878
rect 2863 810 2919 844
rect 2863 776 2874 810
rect 2908 776 2919 810
rect 2863 742 2919 776
rect 2863 708 2874 742
rect 2908 708 2919 742
rect 2863 674 2919 708
rect 2863 640 2874 674
rect 2908 640 2919 674
rect 2863 606 2919 640
rect 2863 572 2874 606
rect 2908 572 2919 606
rect 2863 538 2919 572
rect 2863 504 2874 538
rect 2908 504 2919 538
rect 2863 470 2919 504
rect 2863 436 2874 470
rect 2908 436 2919 470
rect 2863 402 2919 436
rect 2863 368 2874 402
rect 2908 368 2919 402
rect 2863 334 2919 368
rect 2863 300 2874 334
rect 2908 300 2919 334
rect 2863 266 2919 300
rect 2863 232 2874 266
rect 2908 232 2919 266
rect 2863 198 2919 232
rect 2863 164 2874 198
rect 2908 164 2919 198
rect 2863 130 2919 164
rect 2863 96 2874 130
rect 2908 96 2919 130
rect 2863 62 2919 96
rect 2863 28 2874 62
rect 2908 28 2919 62
rect 2863 16 2919 28
rect 3019 946 3075 1016
rect 3019 912 3030 946
rect 3064 912 3075 946
rect 3019 878 3075 912
rect 3019 844 3030 878
rect 3064 844 3075 878
rect 3019 810 3075 844
rect 3019 776 3030 810
rect 3064 776 3075 810
rect 3019 742 3075 776
rect 3019 708 3030 742
rect 3064 708 3075 742
rect 3019 674 3075 708
rect 3019 640 3030 674
rect 3064 640 3075 674
rect 3019 606 3075 640
rect 3019 572 3030 606
rect 3064 572 3075 606
rect 3019 538 3075 572
rect 3019 504 3030 538
rect 3064 504 3075 538
rect 3019 470 3075 504
rect 3019 436 3030 470
rect 3064 436 3075 470
rect 3019 402 3075 436
rect 3019 368 3030 402
rect 3064 368 3075 402
rect 3019 334 3075 368
rect 3019 300 3030 334
rect 3064 300 3075 334
rect 3019 266 3075 300
rect 3019 232 3030 266
rect 3064 232 3075 266
rect 3019 198 3075 232
rect 3019 164 3030 198
rect 3064 164 3075 198
rect 3019 130 3075 164
rect 3019 96 3030 130
rect 3064 96 3075 130
rect 3019 62 3075 96
rect 3019 28 3030 62
rect 3064 28 3075 62
rect 3019 16 3075 28
rect 3175 946 3231 1016
rect 3175 912 3186 946
rect 3220 912 3231 946
rect 3175 878 3231 912
rect 3175 844 3186 878
rect 3220 844 3231 878
rect 3175 810 3231 844
rect 3175 776 3186 810
rect 3220 776 3231 810
rect 3175 742 3231 776
rect 3175 708 3186 742
rect 3220 708 3231 742
rect 3175 674 3231 708
rect 3175 640 3186 674
rect 3220 640 3231 674
rect 3175 606 3231 640
rect 3175 572 3186 606
rect 3220 572 3231 606
rect 3175 538 3231 572
rect 3175 504 3186 538
rect 3220 504 3231 538
rect 3175 470 3231 504
rect 3175 436 3186 470
rect 3220 436 3231 470
rect 3175 402 3231 436
rect 3175 368 3186 402
rect 3220 368 3231 402
rect 3175 334 3231 368
rect 3175 300 3186 334
rect 3220 300 3231 334
rect 3175 266 3231 300
rect 3175 232 3186 266
rect 3220 232 3231 266
rect 3175 198 3231 232
rect 3175 164 3186 198
rect 3220 164 3231 198
rect 3175 130 3231 164
rect 3175 96 3186 130
rect 3220 96 3231 130
rect 3175 62 3231 96
rect 3175 28 3186 62
rect 3220 28 3231 62
rect 3175 16 3231 28
rect 3331 946 3387 1016
rect 3331 912 3342 946
rect 3376 912 3387 946
rect 3331 878 3387 912
rect 3331 844 3342 878
rect 3376 844 3387 878
rect 3331 810 3387 844
rect 3331 776 3342 810
rect 3376 776 3387 810
rect 3331 742 3387 776
rect 3331 708 3342 742
rect 3376 708 3387 742
rect 3331 674 3387 708
rect 3331 640 3342 674
rect 3376 640 3387 674
rect 3331 606 3387 640
rect 3331 572 3342 606
rect 3376 572 3387 606
rect 3331 538 3387 572
rect 3331 504 3342 538
rect 3376 504 3387 538
rect 3331 470 3387 504
rect 3331 436 3342 470
rect 3376 436 3387 470
rect 3331 402 3387 436
rect 3331 368 3342 402
rect 3376 368 3387 402
rect 3331 334 3387 368
rect 3331 300 3342 334
rect 3376 300 3387 334
rect 3331 266 3387 300
rect 3331 232 3342 266
rect 3376 232 3387 266
rect 3331 198 3387 232
rect 3331 164 3342 198
rect 3376 164 3387 198
rect 3331 130 3387 164
rect 3331 96 3342 130
rect 3376 96 3387 130
rect 3331 62 3387 96
rect 3331 28 3342 62
rect 3376 28 3387 62
rect 3331 16 3387 28
rect 3487 946 3543 1016
rect 3487 912 3498 946
rect 3532 912 3543 946
rect 3487 878 3543 912
rect 3487 844 3498 878
rect 3532 844 3543 878
rect 3487 810 3543 844
rect 3487 776 3498 810
rect 3532 776 3543 810
rect 3487 742 3543 776
rect 3487 708 3498 742
rect 3532 708 3543 742
rect 3487 674 3543 708
rect 3487 640 3498 674
rect 3532 640 3543 674
rect 3487 606 3543 640
rect 3487 572 3498 606
rect 3532 572 3543 606
rect 3487 538 3543 572
rect 3487 504 3498 538
rect 3532 504 3543 538
rect 3487 470 3543 504
rect 3487 436 3498 470
rect 3532 436 3543 470
rect 3487 402 3543 436
rect 3487 368 3498 402
rect 3532 368 3543 402
rect 3487 334 3543 368
rect 3487 300 3498 334
rect 3532 300 3543 334
rect 3487 266 3543 300
rect 3487 232 3498 266
rect 3532 232 3543 266
rect 3487 198 3543 232
rect 3487 164 3498 198
rect 3532 164 3543 198
rect 3487 130 3543 164
rect 3487 96 3498 130
rect 3532 96 3543 130
rect 3487 62 3543 96
rect 3487 28 3498 62
rect 3532 28 3543 62
rect 3487 16 3543 28
rect 3643 946 3696 1016
rect 3643 912 3654 946
rect 3688 912 3696 946
rect 3643 878 3696 912
rect 3643 844 3654 878
rect 3688 844 3696 878
rect 3643 810 3696 844
rect 3643 776 3654 810
rect 3688 776 3696 810
rect 3643 742 3696 776
rect 3643 708 3654 742
rect 3688 708 3696 742
rect 3643 674 3696 708
rect 3643 640 3654 674
rect 3688 640 3696 674
rect 3643 606 3696 640
rect 3643 572 3654 606
rect 3688 572 3696 606
rect 3643 538 3696 572
rect 3643 504 3654 538
rect 3688 504 3696 538
rect 3643 470 3696 504
rect 3643 436 3654 470
rect 3688 436 3696 470
rect 3643 402 3696 436
rect 3643 368 3654 402
rect 3688 368 3696 402
rect 3643 334 3696 368
rect 3643 300 3654 334
rect 3688 300 3696 334
rect 3643 266 3696 300
rect 3643 232 3654 266
rect 3688 232 3696 266
rect 3643 198 3696 232
rect 3643 164 3654 198
rect 3688 164 3696 198
rect 3643 130 3696 164
rect 3643 96 3654 130
rect 3688 96 3696 130
rect 3643 62 3696 96
rect 3643 28 3654 62
rect 3688 28 3696 62
rect 3643 16 3696 28
rect 3770 946 3823 1016
rect 3770 912 3778 946
rect 3812 912 3823 946
rect 3770 878 3823 912
rect 3770 844 3778 878
rect 3812 844 3823 878
rect 3770 810 3823 844
rect 3770 776 3778 810
rect 3812 776 3823 810
rect 3770 742 3823 776
rect 3770 708 3778 742
rect 3812 708 3823 742
rect 3770 674 3823 708
rect 3770 640 3778 674
rect 3812 640 3823 674
rect 3770 606 3823 640
rect 3770 572 3778 606
rect 3812 572 3823 606
rect 3770 538 3823 572
rect 3770 504 3778 538
rect 3812 504 3823 538
rect 3770 470 3823 504
rect 3770 436 3778 470
rect 3812 436 3823 470
rect 3770 402 3823 436
rect 3770 368 3778 402
rect 3812 368 3823 402
rect 3770 334 3823 368
rect 3770 300 3778 334
rect 3812 300 3823 334
rect 3770 266 3823 300
rect 3770 232 3778 266
rect 3812 232 3823 266
rect 3770 198 3823 232
rect 3770 164 3778 198
rect 3812 164 3823 198
rect 3770 130 3823 164
rect 3770 96 3778 130
rect 3812 96 3823 130
rect 3770 62 3823 96
rect 3770 28 3778 62
rect 3812 28 3823 62
rect 3770 16 3823 28
rect 3923 946 3979 1016
rect 3923 912 3934 946
rect 3968 912 3979 946
rect 3923 878 3979 912
rect 3923 844 3934 878
rect 3968 844 3979 878
rect 3923 810 3979 844
rect 3923 776 3934 810
rect 3968 776 3979 810
rect 3923 742 3979 776
rect 3923 708 3934 742
rect 3968 708 3979 742
rect 3923 674 3979 708
rect 3923 640 3934 674
rect 3968 640 3979 674
rect 3923 606 3979 640
rect 3923 572 3934 606
rect 3968 572 3979 606
rect 3923 538 3979 572
rect 3923 504 3934 538
rect 3968 504 3979 538
rect 3923 470 3979 504
rect 3923 436 3934 470
rect 3968 436 3979 470
rect 3923 402 3979 436
rect 3923 368 3934 402
rect 3968 368 3979 402
rect 3923 334 3979 368
rect 3923 300 3934 334
rect 3968 300 3979 334
rect 3923 266 3979 300
rect 3923 232 3934 266
rect 3968 232 3979 266
rect 3923 198 3979 232
rect 3923 164 3934 198
rect 3968 164 3979 198
rect 3923 130 3979 164
rect 3923 96 3934 130
rect 3968 96 3979 130
rect 3923 62 3979 96
rect 3923 28 3934 62
rect 3968 28 3979 62
rect 3923 16 3979 28
rect 4079 946 4135 1016
rect 4079 912 4090 946
rect 4124 912 4135 946
rect 4079 878 4135 912
rect 4079 844 4090 878
rect 4124 844 4135 878
rect 4079 810 4135 844
rect 4079 776 4090 810
rect 4124 776 4135 810
rect 4079 742 4135 776
rect 4079 708 4090 742
rect 4124 708 4135 742
rect 4079 674 4135 708
rect 4079 640 4090 674
rect 4124 640 4135 674
rect 4079 606 4135 640
rect 4079 572 4090 606
rect 4124 572 4135 606
rect 4079 538 4135 572
rect 4079 504 4090 538
rect 4124 504 4135 538
rect 4079 470 4135 504
rect 4079 436 4090 470
rect 4124 436 4135 470
rect 4079 402 4135 436
rect 4079 368 4090 402
rect 4124 368 4135 402
rect 4079 334 4135 368
rect 4079 300 4090 334
rect 4124 300 4135 334
rect 4079 266 4135 300
rect 4079 232 4090 266
rect 4124 232 4135 266
rect 4079 198 4135 232
rect 4079 164 4090 198
rect 4124 164 4135 198
rect 4079 130 4135 164
rect 4079 96 4090 130
rect 4124 96 4135 130
rect 4079 62 4135 96
rect 4079 28 4090 62
rect 4124 28 4135 62
rect 4079 16 4135 28
rect 4235 946 4291 1016
rect 4235 912 4246 946
rect 4280 912 4291 946
rect 4235 878 4291 912
rect 4235 844 4246 878
rect 4280 844 4291 878
rect 4235 810 4291 844
rect 4235 776 4246 810
rect 4280 776 4291 810
rect 4235 742 4291 776
rect 4235 708 4246 742
rect 4280 708 4291 742
rect 4235 674 4291 708
rect 4235 640 4246 674
rect 4280 640 4291 674
rect 4235 606 4291 640
rect 4235 572 4246 606
rect 4280 572 4291 606
rect 4235 538 4291 572
rect 4235 504 4246 538
rect 4280 504 4291 538
rect 4235 470 4291 504
rect 4235 436 4246 470
rect 4280 436 4291 470
rect 4235 402 4291 436
rect 4235 368 4246 402
rect 4280 368 4291 402
rect 4235 334 4291 368
rect 4235 300 4246 334
rect 4280 300 4291 334
rect 4235 266 4291 300
rect 4235 232 4246 266
rect 4280 232 4291 266
rect 4235 198 4291 232
rect 4235 164 4246 198
rect 4280 164 4291 198
rect 4235 130 4291 164
rect 4235 96 4246 130
rect 4280 96 4291 130
rect 4235 62 4291 96
rect 4235 28 4246 62
rect 4280 28 4291 62
rect 4235 16 4291 28
rect 4391 946 4447 1016
rect 4391 912 4402 946
rect 4436 912 4447 946
rect 4391 878 4447 912
rect 4391 844 4402 878
rect 4436 844 4447 878
rect 4391 810 4447 844
rect 4391 776 4402 810
rect 4436 776 4447 810
rect 4391 742 4447 776
rect 4391 708 4402 742
rect 4436 708 4447 742
rect 4391 674 4447 708
rect 4391 640 4402 674
rect 4436 640 4447 674
rect 4391 606 4447 640
rect 4391 572 4402 606
rect 4436 572 4447 606
rect 4391 538 4447 572
rect 4391 504 4402 538
rect 4436 504 4447 538
rect 4391 470 4447 504
rect 4391 436 4402 470
rect 4436 436 4447 470
rect 4391 402 4447 436
rect 4391 368 4402 402
rect 4436 368 4447 402
rect 4391 334 4447 368
rect 4391 300 4402 334
rect 4436 300 4447 334
rect 4391 266 4447 300
rect 4391 232 4402 266
rect 4436 232 4447 266
rect 4391 198 4447 232
rect 4391 164 4402 198
rect 4436 164 4447 198
rect 4391 130 4447 164
rect 4391 96 4402 130
rect 4436 96 4447 130
rect 4391 62 4447 96
rect 4391 28 4402 62
rect 4436 28 4447 62
rect 4391 16 4447 28
rect 4547 946 4603 1016
rect 4547 912 4558 946
rect 4592 912 4603 946
rect 4547 878 4603 912
rect 4547 844 4558 878
rect 4592 844 4603 878
rect 4547 810 4603 844
rect 4547 776 4558 810
rect 4592 776 4603 810
rect 4547 742 4603 776
rect 4547 708 4558 742
rect 4592 708 4603 742
rect 4547 674 4603 708
rect 4547 640 4558 674
rect 4592 640 4603 674
rect 4547 606 4603 640
rect 4547 572 4558 606
rect 4592 572 4603 606
rect 4547 538 4603 572
rect 4547 504 4558 538
rect 4592 504 4603 538
rect 4547 470 4603 504
rect 4547 436 4558 470
rect 4592 436 4603 470
rect 4547 402 4603 436
rect 4547 368 4558 402
rect 4592 368 4603 402
rect 4547 334 4603 368
rect 4547 300 4558 334
rect 4592 300 4603 334
rect 4547 266 4603 300
rect 4547 232 4558 266
rect 4592 232 4603 266
rect 4547 198 4603 232
rect 4547 164 4558 198
rect 4592 164 4603 198
rect 4547 130 4603 164
rect 4547 96 4558 130
rect 4592 96 4603 130
rect 4547 62 4603 96
rect 4547 28 4558 62
rect 4592 28 4603 62
rect 4547 16 4603 28
rect 4703 946 4759 1016
rect 4703 912 4714 946
rect 4748 912 4759 946
rect 4703 878 4759 912
rect 4703 844 4714 878
rect 4748 844 4759 878
rect 4703 810 4759 844
rect 4703 776 4714 810
rect 4748 776 4759 810
rect 4703 742 4759 776
rect 4703 708 4714 742
rect 4748 708 4759 742
rect 4703 674 4759 708
rect 4703 640 4714 674
rect 4748 640 4759 674
rect 4703 606 4759 640
rect 4703 572 4714 606
rect 4748 572 4759 606
rect 4703 538 4759 572
rect 4703 504 4714 538
rect 4748 504 4759 538
rect 4703 470 4759 504
rect 4703 436 4714 470
rect 4748 436 4759 470
rect 4703 402 4759 436
rect 4703 368 4714 402
rect 4748 368 4759 402
rect 4703 334 4759 368
rect 4703 300 4714 334
rect 4748 300 4759 334
rect 4703 266 4759 300
rect 4703 232 4714 266
rect 4748 232 4759 266
rect 4703 198 4759 232
rect 4703 164 4714 198
rect 4748 164 4759 198
rect 4703 130 4759 164
rect 4703 96 4714 130
rect 4748 96 4759 130
rect 4703 62 4759 96
rect 4703 28 4714 62
rect 4748 28 4759 62
rect 4703 16 4759 28
rect 4859 946 4915 1016
rect 4859 912 4870 946
rect 4904 912 4915 946
rect 4859 878 4915 912
rect 4859 844 4870 878
rect 4904 844 4915 878
rect 4859 810 4915 844
rect 4859 776 4870 810
rect 4904 776 4915 810
rect 4859 742 4915 776
rect 4859 708 4870 742
rect 4904 708 4915 742
rect 4859 674 4915 708
rect 4859 640 4870 674
rect 4904 640 4915 674
rect 4859 606 4915 640
rect 4859 572 4870 606
rect 4904 572 4915 606
rect 4859 538 4915 572
rect 4859 504 4870 538
rect 4904 504 4915 538
rect 4859 470 4915 504
rect 4859 436 4870 470
rect 4904 436 4915 470
rect 4859 402 4915 436
rect 4859 368 4870 402
rect 4904 368 4915 402
rect 4859 334 4915 368
rect 4859 300 4870 334
rect 4904 300 4915 334
rect 4859 266 4915 300
rect 4859 232 4870 266
rect 4904 232 4915 266
rect 4859 198 4915 232
rect 4859 164 4870 198
rect 4904 164 4915 198
rect 4859 130 4915 164
rect 4859 96 4870 130
rect 4904 96 4915 130
rect 4859 62 4915 96
rect 4859 28 4870 62
rect 4904 28 4915 62
rect 4859 16 4915 28
rect 5015 946 5071 1016
rect 5015 912 5026 946
rect 5060 912 5071 946
rect 5015 878 5071 912
rect 5015 844 5026 878
rect 5060 844 5071 878
rect 5015 810 5071 844
rect 5015 776 5026 810
rect 5060 776 5071 810
rect 5015 742 5071 776
rect 5015 708 5026 742
rect 5060 708 5071 742
rect 5015 674 5071 708
rect 5015 640 5026 674
rect 5060 640 5071 674
rect 5015 606 5071 640
rect 5015 572 5026 606
rect 5060 572 5071 606
rect 5015 538 5071 572
rect 5015 504 5026 538
rect 5060 504 5071 538
rect 5015 470 5071 504
rect 5015 436 5026 470
rect 5060 436 5071 470
rect 5015 402 5071 436
rect 5015 368 5026 402
rect 5060 368 5071 402
rect 5015 334 5071 368
rect 5015 300 5026 334
rect 5060 300 5071 334
rect 5015 266 5071 300
rect 5015 232 5026 266
rect 5060 232 5071 266
rect 5015 198 5071 232
rect 5015 164 5026 198
rect 5060 164 5071 198
rect 5015 130 5071 164
rect 5015 96 5026 130
rect 5060 96 5071 130
rect 5015 62 5071 96
rect 5015 28 5026 62
rect 5060 28 5071 62
rect 5015 16 5071 28
rect 5171 946 5227 1016
rect 5171 912 5182 946
rect 5216 912 5227 946
rect 5171 878 5227 912
rect 5171 844 5182 878
rect 5216 844 5227 878
rect 5171 810 5227 844
rect 5171 776 5182 810
rect 5216 776 5227 810
rect 5171 742 5227 776
rect 5171 708 5182 742
rect 5216 708 5227 742
rect 5171 674 5227 708
rect 5171 640 5182 674
rect 5216 640 5227 674
rect 5171 606 5227 640
rect 5171 572 5182 606
rect 5216 572 5227 606
rect 5171 538 5227 572
rect 5171 504 5182 538
rect 5216 504 5227 538
rect 5171 470 5227 504
rect 5171 436 5182 470
rect 5216 436 5227 470
rect 5171 402 5227 436
rect 5171 368 5182 402
rect 5216 368 5227 402
rect 5171 334 5227 368
rect 5171 300 5182 334
rect 5216 300 5227 334
rect 5171 266 5227 300
rect 5171 232 5182 266
rect 5216 232 5227 266
rect 5171 198 5227 232
rect 5171 164 5182 198
rect 5216 164 5227 198
rect 5171 130 5227 164
rect 5171 96 5182 130
rect 5216 96 5227 130
rect 5171 62 5227 96
rect 5171 28 5182 62
rect 5216 28 5227 62
rect 5171 16 5227 28
rect 5327 946 5383 1016
rect 5327 912 5338 946
rect 5372 912 5383 946
rect 5327 878 5383 912
rect 5327 844 5338 878
rect 5372 844 5383 878
rect 5327 810 5383 844
rect 5327 776 5338 810
rect 5372 776 5383 810
rect 5327 742 5383 776
rect 5327 708 5338 742
rect 5372 708 5383 742
rect 5327 674 5383 708
rect 5327 640 5338 674
rect 5372 640 5383 674
rect 5327 606 5383 640
rect 5327 572 5338 606
rect 5372 572 5383 606
rect 5327 538 5383 572
rect 5327 504 5338 538
rect 5372 504 5383 538
rect 5327 470 5383 504
rect 5327 436 5338 470
rect 5372 436 5383 470
rect 5327 402 5383 436
rect 5327 368 5338 402
rect 5372 368 5383 402
rect 5327 334 5383 368
rect 5327 300 5338 334
rect 5372 300 5383 334
rect 5327 266 5383 300
rect 5327 232 5338 266
rect 5372 232 5383 266
rect 5327 198 5383 232
rect 5327 164 5338 198
rect 5372 164 5383 198
rect 5327 130 5383 164
rect 5327 96 5338 130
rect 5372 96 5383 130
rect 5327 62 5383 96
rect 5327 28 5338 62
rect 5372 28 5383 62
rect 5327 16 5383 28
rect 5483 946 5536 1016
rect 5483 912 5494 946
rect 5528 912 5536 946
rect 5483 878 5536 912
rect 5483 844 5494 878
rect 5528 844 5536 878
rect 5483 810 5536 844
rect 5483 776 5494 810
rect 5528 776 5536 810
rect 5483 742 5536 776
rect 5483 708 5494 742
rect 5528 708 5536 742
rect 5483 674 5536 708
rect 5483 640 5494 674
rect 5528 640 5536 674
rect 5483 606 5536 640
rect 5483 572 5494 606
rect 5528 572 5536 606
rect 5483 538 5536 572
rect 5483 504 5494 538
rect 5528 504 5536 538
rect 5483 470 5536 504
rect 5483 436 5494 470
rect 5528 436 5536 470
rect 5483 402 5536 436
rect 5483 368 5494 402
rect 5528 368 5536 402
rect 5483 334 5536 368
rect 5483 300 5494 334
rect 5528 300 5536 334
rect 5483 266 5536 300
rect 5483 232 5494 266
rect 5528 232 5536 266
rect 5483 198 5536 232
rect 5483 164 5494 198
rect 5528 164 5536 198
rect 5483 130 5536 164
rect 5483 96 5494 130
rect 5528 96 5536 130
rect 5483 62 5536 96
rect 5483 28 5494 62
rect 5528 28 5536 62
rect 5483 16 5536 28
rect 5660 946 5713 1016
rect 5660 912 5668 946
rect 5702 912 5713 946
rect 5660 878 5713 912
rect 5660 844 5668 878
rect 5702 844 5713 878
rect 5660 810 5713 844
rect 5660 776 5668 810
rect 5702 776 5713 810
rect 5660 742 5713 776
rect 5660 708 5668 742
rect 5702 708 5713 742
rect 5660 674 5713 708
rect 5660 640 5668 674
rect 5702 640 5713 674
rect 5660 606 5713 640
rect 5660 572 5668 606
rect 5702 572 5713 606
rect 5660 538 5713 572
rect 5660 504 5668 538
rect 5702 504 5713 538
rect 5660 470 5713 504
rect 5660 436 5668 470
rect 5702 436 5713 470
rect 5660 402 5713 436
rect 5660 368 5668 402
rect 5702 368 5713 402
rect 5660 334 5713 368
rect 5660 300 5668 334
rect 5702 300 5713 334
rect 5660 266 5713 300
rect 5660 232 5668 266
rect 5702 232 5713 266
rect 5660 198 5713 232
rect 5660 164 5668 198
rect 5702 164 5713 198
rect 5660 130 5713 164
rect 5660 96 5668 130
rect 5702 96 5713 130
rect 5660 62 5713 96
rect 5660 28 5668 62
rect 5702 28 5713 62
rect 5660 16 5713 28
rect 5813 946 5869 1016
rect 5813 912 5824 946
rect 5858 912 5869 946
rect 5813 878 5869 912
rect 5813 844 5824 878
rect 5858 844 5869 878
rect 5813 810 5869 844
rect 5813 776 5824 810
rect 5858 776 5869 810
rect 5813 742 5869 776
rect 5813 708 5824 742
rect 5858 708 5869 742
rect 5813 674 5869 708
rect 5813 640 5824 674
rect 5858 640 5869 674
rect 5813 606 5869 640
rect 5813 572 5824 606
rect 5858 572 5869 606
rect 5813 538 5869 572
rect 5813 504 5824 538
rect 5858 504 5869 538
rect 5813 470 5869 504
rect 5813 436 5824 470
rect 5858 436 5869 470
rect 5813 402 5869 436
rect 5813 368 5824 402
rect 5858 368 5869 402
rect 5813 334 5869 368
rect 5813 300 5824 334
rect 5858 300 5869 334
rect 5813 266 5869 300
rect 5813 232 5824 266
rect 5858 232 5869 266
rect 5813 198 5869 232
rect 5813 164 5824 198
rect 5858 164 5869 198
rect 5813 130 5869 164
rect 5813 96 5824 130
rect 5858 96 5869 130
rect 5813 62 5869 96
rect 5813 28 5824 62
rect 5858 28 5869 62
rect 5813 16 5869 28
rect 5969 946 6025 1016
rect 5969 912 5980 946
rect 6014 912 6025 946
rect 5969 878 6025 912
rect 5969 844 5980 878
rect 6014 844 6025 878
rect 5969 810 6025 844
rect 5969 776 5980 810
rect 6014 776 6025 810
rect 5969 742 6025 776
rect 5969 708 5980 742
rect 6014 708 6025 742
rect 5969 674 6025 708
rect 5969 640 5980 674
rect 6014 640 6025 674
rect 5969 606 6025 640
rect 5969 572 5980 606
rect 6014 572 6025 606
rect 5969 538 6025 572
rect 5969 504 5980 538
rect 6014 504 6025 538
rect 5969 470 6025 504
rect 5969 436 5980 470
rect 6014 436 6025 470
rect 5969 402 6025 436
rect 5969 368 5980 402
rect 6014 368 6025 402
rect 5969 334 6025 368
rect 5969 300 5980 334
rect 6014 300 6025 334
rect 5969 266 6025 300
rect 5969 232 5980 266
rect 6014 232 6025 266
rect 5969 198 6025 232
rect 5969 164 5980 198
rect 6014 164 6025 198
rect 5969 130 6025 164
rect 5969 96 5980 130
rect 6014 96 6025 130
rect 5969 62 6025 96
rect 5969 28 5980 62
rect 6014 28 6025 62
rect 5969 16 6025 28
rect 6125 946 6181 1016
rect 6125 912 6136 946
rect 6170 912 6181 946
rect 6125 878 6181 912
rect 6125 844 6136 878
rect 6170 844 6181 878
rect 6125 810 6181 844
rect 6125 776 6136 810
rect 6170 776 6181 810
rect 6125 742 6181 776
rect 6125 708 6136 742
rect 6170 708 6181 742
rect 6125 674 6181 708
rect 6125 640 6136 674
rect 6170 640 6181 674
rect 6125 606 6181 640
rect 6125 572 6136 606
rect 6170 572 6181 606
rect 6125 538 6181 572
rect 6125 504 6136 538
rect 6170 504 6181 538
rect 6125 470 6181 504
rect 6125 436 6136 470
rect 6170 436 6181 470
rect 6125 402 6181 436
rect 6125 368 6136 402
rect 6170 368 6181 402
rect 6125 334 6181 368
rect 6125 300 6136 334
rect 6170 300 6181 334
rect 6125 266 6181 300
rect 6125 232 6136 266
rect 6170 232 6181 266
rect 6125 198 6181 232
rect 6125 164 6136 198
rect 6170 164 6181 198
rect 6125 130 6181 164
rect 6125 96 6136 130
rect 6170 96 6181 130
rect 6125 62 6181 96
rect 6125 28 6136 62
rect 6170 28 6181 62
rect 6125 16 6181 28
rect 6281 946 6334 1016
rect 6281 912 6292 946
rect 6326 912 6334 946
rect 6281 878 6334 912
rect 6281 844 6292 878
rect 6326 844 6334 878
rect 6281 810 6334 844
rect 6281 776 6292 810
rect 6326 776 6334 810
rect 6281 742 6334 776
rect 6281 708 6292 742
rect 6326 708 6334 742
rect 6281 674 6334 708
rect 6281 640 6292 674
rect 6326 640 6334 674
rect 6281 606 6334 640
rect 6281 572 6292 606
rect 6326 572 6334 606
rect 6281 538 6334 572
rect 6281 504 6292 538
rect 6326 504 6334 538
rect 6281 470 6334 504
rect 6281 436 6292 470
rect 6326 436 6334 470
rect 6281 402 6334 436
rect 6281 368 6292 402
rect 6326 368 6334 402
rect 6281 334 6334 368
rect 6281 300 6292 334
rect 6326 300 6334 334
rect 6281 266 6334 300
rect 6281 232 6292 266
rect 6326 232 6334 266
rect 6281 198 6334 232
rect 6281 164 6292 198
rect 6326 164 6334 198
rect 6281 130 6334 164
rect 6281 96 6292 130
rect 6326 96 6334 130
rect 6281 62 6334 96
rect 6281 28 6292 62
rect 6326 28 6334 62
rect 6281 16 6334 28
rect 6408 946 6461 1016
rect 6408 912 6416 946
rect 6450 912 6461 946
rect 6408 878 6461 912
rect 6408 844 6416 878
rect 6450 844 6461 878
rect 6408 810 6461 844
rect 6408 776 6416 810
rect 6450 776 6461 810
rect 6408 742 6461 776
rect 6408 708 6416 742
rect 6450 708 6461 742
rect 6408 674 6461 708
rect 6408 640 6416 674
rect 6450 640 6461 674
rect 6408 606 6461 640
rect 6408 572 6416 606
rect 6450 572 6461 606
rect 6408 538 6461 572
rect 6408 504 6416 538
rect 6450 504 6461 538
rect 6408 470 6461 504
rect 6408 436 6416 470
rect 6450 436 6461 470
rect 6408 402 6461 436
rect 6408 368 6416 402
rect 6450 368 6461 402
rect 6408 334 6461 368
rect 6408 300 6416 334
rect 6450 300 6461 334
rect 6408 266 6461 300
rect 6408 232 6416 266
rect 6450 232 6461 266
rect 6408 198 6461 232
rect 6408 164 6416 198
rect 6450 164 6461 198
rect 6408 130 6461 164
rect 6408 96 6416 130
rect 6450 96 6461 130
rect 6408 62 6461 96
rect 6408 28 6416 62
rect 6450 28 6461 62
rect 6408 16 6461 28
rect 6561 946 6614 1016
rect 6561 912 6572 946
rect 6606 912 6614 946
rect 6561 878 6614 912
rect 6561 844 6572 878
rect 6606 844 6614 878
rect 6561 810 6614 844
rect 6561 776 6572 810
rect 6606 776 6614 810
rect 6561 742 6614 776
rect 6561 708 6572 742
rect 6606 708 6614 742
rect 6561 674 6614 708
rect 6561 640 6572 674
rect 6606 640 6614 674
rect 6561 606 6614 640
rect 6561 572 6572 606
rect 6606 572 6614 606
rect 6561 538 6614 572
rect 6561 504 6572 538
rect 6606 504 6614 538
rect 6561 470 6614 504
rect 6561 436 6572 470
rect 6606 436 6614 470
rect 6561 402 6614 436
rect 6561 368 6572 402
rect 6606 368 6614 402
rect 6561 334 6614 368
rect 6561 300 6572 334
rect 6606 300 6614 334
rect 6561 266 6614 300
rect 6561 232 6572 266
rect 6606 232 6614 266
rect 6561 198 6614 232
rect 6561 164 6572 198
rect 6606 164 6614 198
rect 6561 130 6614 164
rect 6561 96 6572 130
rect 6606 96 6614 130
rect 6561 62 6614 96
rect 6561 28 6572 62
rect 6606 28 6614 62
rect 6561 16 6614 28
rect 6688 946 6741 1016
rect 6688 912 6696 946
rect 6730 912 6741 946
rect 6688 878 6741 912
rect 6688 844 6696 878
rect 6730 844 6741 878
rect 6688 810 6741 844
rect 6688 776 6696 810
rect 6730 776 6741 810
rect 6688 742 6741 776
rect 6688 708 6696 742
rect 6730 708 6741 742
rect 6688 674 6741 708
rect 6688 640 6696 674
rect 6730 640 6741 674
rect 6688 606 6741 640
rect 6688 572 6696 606
rect 6730 572 6741 606
rect 6688 538 6741 572
rect 6688 504 6696 538
rect 6730 504 6741 538
rect 6688 470 6741 504
rect 6688 436 6696 470
rect 6730 436 6741 470
rect 6688 402 6741 436
rect 6688 368 6696 402
rect 6730 368 6741 402
rect 6688 334 6741 368
rect 6688 300 6696 334
rect 6730 300 6741 334
rect 6688 266 6741 300
rect 6688 232 6696 266
rect 6730 232 6741 266
rect 6688 198 6741 232
rect 6688 164 6696 198
rect 6730 164 6741 198
rect 6688 130 6741 164
rect 6688 96 6696 130
rect 6730 96 6741 130
rect 6688 62 6741 96
rect 6688 28 6696 62
rect 6730 28 6741 62
rect 6688 16 6741 28
rect 6841 946 6897 1016
rect 6841 912 6852 946
rect 6886 912 6897 946
rect 6841 878 6897 912
rect 6841 844 6852 878
rect 6886 844 6897 878
rect 6841 810 6897 844
rect 6841 776 6852 810
rect 6886 776 6897 810
rect 6841 742 6897 776
rect 6841 708 6852 742
rect 6886 708 6897 742
rect 6841 674 6897 708
rect 6841 640 6852 674
rect 6886 640 6897 674
rect 6841 606 6897 640
rect 6841 572 6852 606
rect 6886 572 6897 606
rect 6841 538 6897 572
rect 6841 504 6852 538
rect 6886 504 6897 538
rect 6841 470 6897 504
rect 6841 436 6852 470
rect 6886 436 6897 470
rect 6841 402 6897 436
rect 6841 368 6852 402
rect 6886 368 6897 402
rect 6841 334 6897 368
rect 6841 300 6852 334
rect 6886 300 6897 334
rect 6841 266 6897 300
rect 6841 232 6852 266
rect 6886 232 6897 266
rect 6841 198 6897 232
rect 6841 164 6852 198
rect 6886 164 6897 198
rect 6841 130 6897 164
rect 6841 96 6852 130
rect 6886 96 6897 130
rect 6841 62 6897 96
rect 6841 28 6852 62
rect 6886 28 6897 62
rect 6841 16 6897 28
rect 6997 946 7050 1016
rect 6997 912 7008 946
rect 7042 912 7050 946
rect 6997 878 7050 912
rect 6997 844 7008 878
rect 7042 844 7050 878
rect 6997 810 7050 844
rect 6997 776 7008 810
rect 7042 776 7050 810
rect 6997 742 7050 776
rect 6997 708 7008 742
rect 7042 708 7050 742
rect 6997 674 7050 708
rect 6997 640 7008 674
rect 7042 640 7050 674
rect 6997 606 7050 640
rect 6997 572 7008 606
rect 7042 572 7050 606
rect 6997 538 7050 572
rect 6997 504 7008 538
rect 7042 504 7050 538
rect 6997 470 7050 504
rect 6997 436 7008 470
rect 7042 436 7050 470
rect 6997 402 7050 436
rect 6997 368 7008 402
rect 7042 368 7050 402
rect 6997 334 7050 368
rect 6997 300 7008 334
rect 7042 300 7050 334
rect 6997 266 7050 300
rect 6997 232 7008 266
rect 7042 232 7050 266
rect 6997 198 7050 232
rect 6997 164 7008 198
rect 7042 164 7050 198
rect 6997 130 7050 164
rect 6997 96 7008 130
rect 7042 96 7050 130
rect 6997 62 7050 96
rect 6997 28 7008 62
rect 7042 28 7050 62
rect 6997 16 7050 28
rect 13076 1069 15076 1077
rect 13076 1035 13088 1069
rect 13122 1035 13156 1069
rect 13190 1035 13224 1069
rect 13258 1035 13292 1069
rect 13326 1035 13360 1069
rect 13394 1035 13428 1069
rect 13462 1035 13496 1069
rect 13530 1035 13564 1069
rect 13598 1035 13632 1069
rect 13666 1035 13700 1069
rect 13734 1035 13768 1069
rect 13802 1035 13836 1069
rect 13870 1035 13904 1069
rect 13938 1035 13972 1069
rect 14006 1035 14040 1069
rect 14074 1035 14108 1069
rect 14142 1035 14176 1069
rect 14210 1035 14244 1069
rect 14278 1035 14312 1069
rect 14346 1035 14380 1069
rect 14414 1035 14448 1069
rect 14482 1035 14516 1069
rect 14550 1035 14584 1069
rect 14618 1035 14652 1069
rect 14686 1035 14720 1069
rect 14754 1035 14788 1069
rect 14822 1035 14856 1069
rect 14890 1035 14924 1069
rect 14958 1035 14992 1069
rect 15026 1035 15076 1069
rect 13076 1024 15076 1035
rect 8276 878 8329 948
rect 8276 844 8284 878
rect 8318 844 8329 878
rect 8276 810 8329 844
rect 8276 776 8284 810
rect 8318 776 8329 810
rect 8276 742 8329 776
rect 8276 708 8284 742
rect 8318 708 8329 742
rect 8276 674 8329 708
rect 8276 640 8284 674
rect 8318 640 8329 674
rect 8276 606 8329 640
rect 8276 572 8284 606
rect 8318 572 8329 606
rect 8276 538 8329 572
rect 8276 504 8284 538
rect 8318 504 8329 538
rect 8276 470 8329 504
rect 8276 436 8284 470
rect 8318 436 8329 470
rect 8276 402 8329 436
rect 8276 368 8284 402
rect 8318 368 8329 402
rect 8276 334 8329 368
rect 8276 300 8284 334
rect 8318 300 8329 334
rect 8276 266 8329 300
rect 8276 232 8284 266
rect 8318 232 8329 266
rect 8276 198 8329 232
rect 8276 164 8284 198
rect 8318 164 8329 198
rect 8276 130 8329 164
rect 8276 96 8284 130
rect 8318 96 8329 130
rect 8276 62 8329 96
rect 8276 28 8284 62
rect 8318 28 8329 62
rect 8276 -6 8329 28
rect 8276 -40 8284 -6
rect 8318 -40 8329 -6
rect 8276 -52 8329 -40
rect 8429 878 8485 948
rect 8429 844 8440 878
rect 8474 844 8485 878
rect 8429 810 8485 844
rect 8429 776 8440 810
rect 8474 776 8485 810
rect 8429 742 8485 776
rect 8429 708 8440 742
rect 8474 708 8485 742
rect 8429 674 8485 708
rect 8429 640 8440 674
rect 8474 640 8485 674
rect 8429 606 8485 640
rect 8429 572 8440 606
rect 8474 572 8485 606
rect 8429 538 8485 572
rect 8429 504 8440 538
rect 8474 504 8485 538
rect 8429 470 8485 504
rect 8429 436 8440 470
rect 8474 436 8485 470
rect 8429 402 8485 436
rect 8429 368 8440 402
rect 8474 368 8485 402
rect 8429 334 8485 368
rect 8429 300 8440 334
rect 8474 300 8485 334
rect 8429 266 8485 300
rect 8429 232 8440 266
rect 8474 232 8485 266
rect 8429 198 8485 232
rect 8429 164 8440 198
rect 8474 164 8485 198
rect 8429 130 8485 164
rect 8429 96 8440 130
rect 8474 96 8485 130
rect 8429 62 8485 96
rect 8429 28 8440 62
rect 8474 28 8485 62
rect 8429 -6 8485 28
rect 8429 -40 8440 -6
rect 8474 -40 8485 -6
rect 8429 -52 8485 -40
rect 8585 878 8641 948
rect 8585 844 8596 878
rect 8630 844 8641 878
rect 8585 810 8641 844
rect 8585 776 8596 810
rect 8630 776 8641 810
rect 8585 742 8641 776
rect 8585 708 8596 742
rect 8630 708 8641 742
rect 8585 674 8641 708
rect 8585 640 8596 674
rect 8630 640 8641 674
rect 8585 606 8641 640
rect 8585 572 8596 606
rect 8630 572 8641 606
rect 8585 538 8641 572
rect 8585 504 8596 538
rect 8630 504 8641 538
rect 8585 470 8641 504
rect 8585 436 8596 470
rect 8630 436 8641 470
rect 8585 402 8641 436
rect 8585 368 8596 402
rect 8630 368 8641 402
rect 8585 334 8641 368
rect 8585 300 8596 334
rect 8630 300 8641 334
rect 8585 266 8641 300
rect 8585 232 8596 266
rect 8630 232 8641 266
rect 8585 198 8641 232
rect 8585 164 8596 198
rect 8630 164 8641 198
rect 8585 130 8641 164
rect 8585 96 8596 130
rect 8630 96 8641 130
rect 8585 62 8641 96
rect 8585 28 8596 62
rect 8630 28 8641 62
rect 8585 -6 8641 28
rect 8585 -40 8596 -6
rect 8630 -40 8641 -6
rect 8585 -52 8641 -40
rect 8741 878 8797 948
rect 8741 844 8752 878
rect 8786 844 8797 878
rect 8741 810 8797 844
rect 8741 776 8752 810
rect 8786 776 8797 810
rect 8741 742 8797 776
rect 8741 708 8752 742
rect 8786 708 8797 742
rect 8741 674 8797 708
rect 8741 640 8752 674
rect 8786 640 8797 674
rect 8741 606 8797 640
rect 8741 572 8752 606
rect 8786 572 8797 606
rect 8741 538 8797 572
rect 8741 504 8752 538
rect 8786 504 8797 538
rect 8741 470 8797 504
rect 8741 436 8752 470
rect 8786 436 8797 470
rect 8741 402 8797 436
rect 8741 368 8752 402
rect 8786 368 8797 402
rect 8741 334 8797 368
rect 8741 300 8752 334
rect 8786 300 8797 334
rect 8741 266 8797 300
rect 8741 232 8752 266
rect 8786 232 8797 266
rect 8741 198 8797 232
rect 8741 164 8752 198
rect 8786 164 8797 198
rect 8741 130 8797 164
rect 8741 96 8752 130
rect 8786 96 8797 130
rect 8741 62 8797 96
rect 8741 28 8752 62
rect 8786 28 8797 62
rect 8741 -6 8797 28
rect 8741 -40 8752 -6
rect 8786 -40 8797 -6
rect 8741 -52 8797 -40
rect 8897 878 8953 948
rect 8897 844 8908 878
rect 8942 844 8953 878
rect 8897 810 8953 844
rect 8897 776 8908 810
rect 8942 776 8953 810
rect 8897 742 8953 776
rect 8897 708 8908 742
rect 8942 708 8953 742
rect 8897 674 8953 708
rect 8897 640 8908 674
rect 8942 640 8953 674
rect 8897 606 8953 640
rect 8897 572 8908 606
rect 8942 572 8953 606
rect 8897 538 8953 572
rect 8897 504 8908 538
rect 8942 504 8953 538
rect 8897 470 8953 504
rect 8897 436 8908 470
rect 8942 436 8953 470
rect 8897 402 8953 436
rect 8897 368 8908 402
rect 8942 368 8953 402
rect 8897 334 8953 368
rect 8897 300 8908 334
rect 8942 300 8953 334
rect 8897 266 8953 300
rect 8897 232 8908 266
rect 8942 232 8953 266
rect 8897 198 8953 232
rect 8897 164 8908 198
rect 8942 164 8953 198
rect 8897 130 8953 164
rect 8897 96 8908 130
rect 8942 96 8953 130
rect 8897 62 8953 96
rect 8897 28 8908 62
rect 8942 28 8953 62
rect 8897 -6 8953 28
rect 8897 -40 8908 -6
rect 8942 -40 8953 -6
rect 8897 -52 8953 -40
rect 9053 878 9109 948
rect 9053 844 9064 878
rect 9098 844 9109 878
rect 9053 810 9109 844
rect 9053 776 9064 810
rect 9098 776 9109 810
rect 9053 742 9109 776
rect 9053 708 9064 742
rect 9098 708 9109 742
rect 9053 674 9109 708
rect 9053 640 9064 674
rect 9098 640 9109 674
rect 9053 606 9109 640
rect 9053 572 9064 606
rect 9098 572 9109 606
rect 9053 538 9109 572
rect 9053 504 9064 538
rect 9098 504 9109 538
rect 9053 470 9109 504
rect 9053 436 9064 470
rect 9098 436 9109 470
rect 9053 402 9109 436
rect 9053 368 9064 402
rect 9098 368 9109 402
rect 9053 334 9109 368
rect 9053 300 9064 334
rect 9098 300 9109 334
rect 9053 266 9109 300
rect 9053 232 9064 266
rect 9098 232 9109 266
rect 9053 198 9109 232
rect 9053 164 9064 198
rect 9098 164 9109 198
rect 9053 130 9109 164
rect 9053 96 9064 130
rect 9098 96 9109 130
rect 9053 62 9109 96
rect 9053 28 9064 62
rect 9098 28 9109 62
rect 9053 -6 9109 28
rect 9053 -40 9064 -6
rect 9098 -40 9109 -6
rect 9053 -52 9109 -40
rect 9209 878 9265 948
rect 9209 844 9220 878
rect 9254 844 9265 878
rect 9209 810 9265 844
rect 9209 776 9220 810
rect 9254 776 9265 810
rect 9209 742 9265 776
rect 9209 708 9220 742
rect 9254 708 9265 742
rect 9209 674 9265 708
rect 9209 640 9220 674
rect 9254 640 9265 674
rect 9209 606 9265 640
rect 9209 572 9220 606
rect 9254 572 9265 606
rect 9209 538 9265 572
rect 9209 504 9220 538
rect 9254 504 9265 538
rect 9209 470 9265 504
rect 9209 436 9220 470
rect 9254 436 9265 470
rect 9209 402 9265 436
rect 9209 368 9220 402
rect 9254 368 9265 402
rect 9209 334 9265 368
rect 9209 300 9220 334
rect 9254 300 9265 334
rect 9209 266 9265 300
rect 9209 232 9220 266
rect 9254 232 9265 266
rect 9209 198 9265 232
rect 9209 164 9220 198
rect 9254 164 9265 198
rect 9209 130 9265 164
rect 9209 96 9220 130
rect 9254 96 9265 130
rect 9209 62 9265 96
rect 9209 28 9220 62
rect 9254 28 9265 62
rect 9209 -6 9265 28
rect 9209 -40 9220 -6
rect 9254 -40 9265 -6
rect 9209 -52 9265 -40
rect 9365 878 9421 948
rect 9365 844 9376 878
rect 9410 844 9421 878
rect 9365 810 9421 844
rect 9365 776 9376 810
rect 9410 776 9421 810
rect 9365 742 9421 776
rect 9365 708 9376 742
rect 9410 708 9421 742
rect 9365 674 9421 708
rect 9365 640 9376 674
rect 9410 640 9421 674
rect 9365 606 9421 640
rect 9365 572 9376 606
rect 9410 572 9421 606
rect 9365 538 9421 572
rect 9365 504 9376 538
rect 9410 504 9421 538
rect 9365 470 9421 504
rect 9365 436 9376 470
rect 9410 436 9421 470
rect 9365 402 9421 436
rect 9365 368 9376 402
rect 9410 368 9421 402
rect 9365 334 9421 368
rect 9365 300 9376 334
rect 9410 300 9421 334
rect 9365 266 9421 300
rect 9365 232 9376 266
rect 9410 232 9421 266
rect 9365 198 9421 232
rect 9365 164 9376 198
rect 9410 164 9421 198
rect 9365 130 9421 164
rect 9365 96 9376 130
rect 9410 96 9421 130
rect 9365 62 9421 96
rect 9365 28 9376 62
rect 9410 28 9421 62
rect 9365 -6 9421 28
rect 9365 -40 9376 -6
rect 9410 -40 9421 -6
rect 9365 -52 9421 -40
rect 9521 878 9577 948
rect 9521 844 9532 878
rect 9566 844 9577 878
rect 9521 810 9577 844
rect 9521 776 9532 810
rect 9566 776 9577 810
rect 9521 742 9577 776
rect 9521 708 9532 742
rect 9566 708 9577 742
rect 9521 674 9577 708
rect 9521 640 9532 674
rect 9566 640 9577 674
rect 9521 606 9577 640
rect 9521 572 9532 606
rect 9566 572 9577 606
rect 9521 538 9577 572
rect 9521 504 9532 538
rect 9566 504 9577 538
rect 9521 470 9577 504
rect 9521 436 9532 470
rect 9566 436 9577 470
rect 9521 402 9577 436
rect 9521 368 9532 402
rect 9566 368 9577 402
rect 9521 334 9577 368
rect 9521 300 9532 334
rect 9566 300 9577 334
rect 9521 266 9577 300
rect 9521 232 9532 266
rect 9566 232 9577 266
rect 9521 198 9577 232
rect 9521 164 9532 198
rect 9566 164 9577 198
rect 9521 130 9577 164
rect 9521 96 9532 130
rect 9566 96 9577 130
rect 9521 62 9577 96
rect 9521 28 9532 62
rect 9566 28 9577 62
rect 9521 -6 9577 28
rect 9521 -40 9532 -6
rect 9566 -40 9577 -6
rect 9521 -52 9577 -40
rect 9677 878 9733 948
rect 9677 844 9688 878
rect 9722 844 9733 878
rect 9677 810 9733 844
rect 9677 776 9688 810
rect 9722 776 9733 810
rect 9677 742 9733 776
rect 9677 708 9688 742
rect 9722 708 9733 742
rect 9677 674 9733 708
rect 9677 640 9688 674
rect 9722 640 9733 674
rect 9677 606 9733 640
rect 9677 572 9688 606
rect 9722 572 9733 606
rect 9677 538 9733 572
rect 9677 504 9688 538
rect 9722 504 9733 538
rect 9677 470 9733 504
rect 9677 436 9688 470
rect 9722 436 9733 470
rect 9677 402 9733 436
rect 9677 368 9688 402
rect 9722 368 9733 402
rect 9677 334 9733 368
rect 9677 300 9688 334
rect 9722 300 9733 334
rect 9677 266 9733 300
rect 9677 232 9688 266
rect 9722 232 9733 266
rect 9677 198 9733 232
rect 9677 164 9688 198
rect 9722 164 9733 198
rect 9677 130 9733 164
rect 9677 96 9688 130
rect 9722 96 9733 130
rect 9677 62 9733 96
rect 9677 28 9688 62
rect 9722 28 9733 62
rect 9677 -6 9733 28
rect 9677 -40 9688 -6
rect 9722 -40 9733 -6
rect 9677 -52 9733 -40
rect 9833 878 9889 948
rect 9833 844 9844 878
rect 9878 844 9889 878
rect 9833 810 9889 844
rect 9833 776 9844 810
rect 9878 776 9889 810
rect 9833 742 9889 776
rect 9833 708 9844 742
rect 9878 708 9889 742
rect 9833 674 9889 708
rect 9833 640 9844 674
rect 9878 640 9889 674
rect 9833 606 9889 640
rect 9833 572 9844 606
rect 9878 572 9889 606
rect 9833 538 9889 572
rect 9833 504 9844 538
rect 9878 504 9889 538
rect 9833 470 9889 504
rect 9833 436 9844 470
rect 9878 436 9889 470
rect 9833 402 9889 436
rect 9833 368 9844 402
rect 9878 368 9889 402
rect 9833 334 9889 368
rect 9833 300 9844 334
rect 9878 300 9889 334
rect 9833 266 9889 300
rect 9833 232 9844 266
rect 9878 232 9889 266
rect 9833 198 9889 232
rect 9833 164 9844 198
rect 9878 164 9889 198
rect 9833 130 9889 164
rect 9833 96 9844 130
rect 9878 96 9889 130
rect 9833 62 9889 96
rect 9833 28 9844 62
rect 9878 28 9889 62
rect 9833 -6 9889 28
rect 9833 -40 9844 -6
rect 9878 -40 9889 -6
rect 9833 -52 9889 -40
rect 9989 878 10045 948
rect 9989 844 10000 878
rect 10034 844 10045 878
rect 9989 810 10045 844
rect 9989 776 10000 810
rect 10034 776 10045 810
rect 9989 742 10045 776
rect 9989 708 10000 742
rect 10034 708 10045 742
rect 9989 674 10045 708
rect 9989 640 10000 674
rect 10034 640 10045 674
rect 9989 606 10045 640
rect 9989 572 10000 606
rect 10034 572 10045 606
rect 9989 538 10045 572
rect 9989 504 10000 538
rect 10034 504 10045 538
rect 9989 470 10045 504
rect 9989 436 10000 470
rect 10034 436 10045 470
rect 9989 402 10045 436
rect 9989 368 10000 402
rect 10034 368 10045 402
rect 9989 334 10045 368
rect 9989 300 10000 334
rect 10034 300 10045 334
rect 9989 266 10045 300
rect 9989 232 10000 266
rect 10034 232 10045 266
rect 9989 198 10045 232
rect 9989 164 10000 198
rect 10034 164 10045 198
rect 9989 130 10045 164
rect 9989 96 10000 130
rect 10034 96 10045 130
rect 9989 62 10045 96
rect 9989 28 10000 62
rect 10034 28 10045 62
rect 9989 -6 10045 28
rect 9989 -40 10000 -6
rect 10034 -40 10045 -6
rect 9989 -52 10045 -40
rect 10145 878 10201 948
rect 10145 844 10156 878
rect 10190 844 10201 878
rect 10145 810 10201 844
rect 10145 776 10156 810
rect 10190 776 10201 810
rect 10145 742 10201 776
rect 10145 708 10156 742
rect 10190 708 10201 742
rect 10145 674 10201 708
rect 10145 640 10156 674
rect 10190 640 10201 674
rect 10145 606 10201 640
rect 10145 572 10156 606
rect 10190 572 10201 606
rect 10145 538 10201 572
rect 10145 504 10156 538
rect 10190 504 10201 538
rect 10145 470 10201 504
rect 10145 436 10156 470
rect 10190 436 10201 470
rect 10145 402 10201 436
rect 10145 368 10156 402
rect 10190 368 10201 402
rect 10145 334 10201 368
rect 10145 300 10156 334
rect 10190 300 10201 334
rect 10145 266 10201 300
rect 10145 232 10156 266
rect 10190 232 10201 266
rect 10145 198 10201 232
rect 10145 164 10156 198
rect 10190 164 10201 198
rect 10145 130 10201 164
rect 10145 96 10156 130
rect 10190 96 10201 130
rect 10145 62 10201 96
rect 10145 28 10156 62
rect 10190 28 10201 62
rect 10145 -6 10201 28
rect 10145 -40 10156 -6
rect 10190 -40 10201 -6
rect 10145 -52 10201 -40
rect 10301 878 10357 948
rect 10301 844 10312 878
rect 10346 844 10357 878
rect 10301 810 10357 844
rect 10301 776 10312 810
rect 10346 776 10357 810
rect 10301 742 10357 776
rect 10301 708 10312 742
rect 10346 708 10357 742
rect 10301 674 10357 708
rect 10301 640 10312 674
rect 10346 640 10357 674
rect 10301 606 10357 640
rect 10301 572 10312 606
rect 10346 572 10357 606
rect 10301 538 10357 572
rect 10301 504 10312 538
rect 10346 504 10357 538
rect 10301 470 10357 504
rect 10301 436 10312 470
rect 10346 436 10357 470
rect 10301 402 10357 436
rect 10301 368 10312 402
rect 10346 368 10357 402
rect 10301 334 10357 368
rect 10301 300 10312 334
rect 10346 300 10357 334
rect 10301 266 10357 300
rect 10301 232 10312 266
rect 10346 232 10357 266
rect 10301 198 10357 232
rect 10301 164 10312 198
rect 10346 164 10357 198
rect 10301 130 10357 164
rect 10301 96 10312 130
rect 10346 96 10357 130
rect 10301 62 10357 96
rect 10301 28 10312 62
rect 10346 28 10357 62
rect 10301 -6 10357 28
rect 10301 -40 10312 -6
rect 10346 -40 10357 -6
rect 10301 -52 10357 -40
rect 10457 878 10510 948
rect 10457 844 10468 878
rect 10502 844 10510 878
rect 10457 810 10510 844
rect 10457 776 10468 810
rect 10502 776 10510 810
rect 10457 742 10510 776
rect 10457 708 10468 742
rect 10502 708 10510 742
rect 10457 674 10510 708
rect 10457 640 10468 674
rect 10502 640 10510 674
rect 10457 606 10510 640
rect 10457 572 10468 606
rect 10502 572 10510 606
rect 10457 538 10510 572
rect 10457 504 10468 538
rect 10502 504 10510 538
rect 10457 470 10510 504
rect 10457 436 10468 470
rect 10502 436 10510 470
rect 10457 402 10510 436
rect 10457 368 10468 402
rect 10502 368 10510 402
rect 10457 334 10510 368
rect 10457 300 10468 334
rect 10502 300 10510 334
rect 10457 266 10510 300
rect 10457 232 10468 266
rect 10502 232 10510 266
rect 10457 198 10510 232
rect 10457 164 10468 198
rect 10502 164 10510 198
rect 10457 130 10510 164
rect 10457 96 10468 130
rect 10502 96 10510 130
rect 10457 62 10510 96
rect 10457 28 10468 62
rect 10502 28 10510 62
rect 10457 -6 10510 28
rect 10457 -40 10468 -6
rect 10502 -40 10510 -6
rect 10457 -52 10510 -40
rect 10729 878 10782 948
rect 10729 844 10737 878
rect 10771 844 10782 878
rect 10729 810 10782 844
rect 10729 776 10737 810
rect 10771 776 10782 810
rect 10729 742 10782 776
rect 10729 708 10737 742
rect 10771 708 10782 742
rect 10729 674 10782 708
rect 10729 640 10737 674
rect 10771 640 10782 674
rect 10729 606 10782 640
rect 10729 572 10737 606
rect 10771 572 10782 606
rect 10729 538 10782 572
rect 10729 504 10737 538
rect 10771 504 10782 538
rect 10729 470 10782 504
rect 10729 436 10737 470
rect 10771 436 10782 470
rect 10729 402 10782 436
rect 10729 368 10737 402
rect 10771 368 10782 402
rect 10729 334 10782 368
rect 10729 300 10737 334
rect 10771 300 10782 334
rect 10729 266 10782 300
rect 10729 232 10737 266
rect 10771 232 10782 266
rect 10729 198 10782 232
rect 10729 164 10737 198
rect 10771 164 10782 198
rect 10729 130 10782 164
rect 10729 96 10737 130
rect 10771 96 10782 130
rect 10729 62 10782 96
rect 10729 28 10737 62
rect 10771 28 10782 62
rect 10729 -6 10782 28
rect 10729 -40 10737 -6
rect 10771 -40 10782 -6
rect 10729 -52 10782 -40
rect 11182 878 11238 948
rect 11182 844 11193 878
rect 11227 844 11238 878
rect 11182 810 11238 844
rect 11182 776 11193 810
rect 11227 776 11238 810
rect 11182 742 11238 776
rect 11182 708 11193 742
rect 11227 708 11238 742
rect 11182 674 11238 708
rect 11182 640 11193 674
rect 11227 640 11238 674
rect 11182 606 11238 640
rect 11182 572 11193 606
rect 11227 572 11238 606
rect 11182 538 11238 572
rect 11182 504 11193 538
rect 11227 504 11238 538
rect 11182 470 11238 504
rect 11182 436 11193 470
rect 11227 436 11238 470
rect 11182 402 11238 436
rect 11182 368 11193 402
rect 11227 368 11238 402
rect 11182 334 11238 368
rect 11182 300 11193 334
rect 11227 300 11238 334
rect 11182 266 11238 300
rect 11182 232 11193 266
rect 11227 232 11238 266
rect 11182 198 11238 232
rect 11182 164 11193 198
rect 11227 164 11238 198
rect 11182 130 11238 164
rect 11182 96 11193 130
rect 11227 96 11238 130
rect 11182 62 11238 96
rect 11182 28 11193 62
rect 11227 28 11238 62
rect 11182 -6 11238 28
rect 11182 -40 11193 -6
rect 11227 -40 11238 -6
rect 11182 -52 11238 -40
rect 11638 878 11694 948
rect 11638 844 11649 878
rect 11683 844 11694 878
rect 11638 810 11694 844
rect 11638 776 11649 810
rect 11683 776 11694 810
rect 11638 742 11694 776
rect 11638 708 11649 742
rect 11683 708 11694 742
rect 11638 674 11694 708
rect 11638 640 11649 674
rect 11683 640 11694 674
rect 11638 606 11694 640
rect 11638 572 11649 606
rect 11683 572 11694 606
rect 11638 538 11694 572
rect 11638 504 11649 538
rect 11683 504 11694 538
rect 11638 470 11694 504
rect 11638 436 11649 470
rect 11683 436 11694 470
rect 11638 402 11694 436
rect 11638 368 11649 402
rect 11683 368 11694 402
rect 11638 334 11694 368
rect 11638 300 11649 334
rect 11683 300 11694 334
rect 11638 266 11694 300
rect 11638 232 11649 266
rect 11683 232 11694 266
rect 11638 198 11694 232
rect 11638 164 11649 198
rect 11683 164 11694 198
rect 11638 130 11694 164
rect 11638 96 11649 130
rect 11683 96 11694 130
rect 11638 62 11694 96
rect 11638 28 11649 62
rect 11683 28 11694 62
rect 11638 -6 11694 28
rect 11638 -40 11649 -6
rect 11683 -40 11694 -6
rect 11638 -52 11694 -40
rect 12094 878 12150 948
rect 12094 844 12105 878
rect 12139 844 12150 878
rect 12094 810 12150 844
rect 12094 776 12105 810
rect 12139 776 12150 810
rect 12094 742 12150 776
rect 12094 708 12105 742
rect 12139 708 12150 742
rect 12094 674 12150 708
rect 12094 640 12105 674
rect 12139 640 12150 674
rect 12094 606 12150 640
rect 12094 572 12105 606
rect 12139 572 12150 606
rect 12094 538 12150 572
rect 12094 504 12105 538
rect 12139 504 12150 538
rect 12094 470 12150 504
rect 12094 436 12105 470
rect 12139 436 12150 470
rect 12094 402 12150 436
rect 12094 368 12105 402
rect 12139 368 12150 402
rect 12094 334 12150 368
rect 12094 300 12105 334
rect 12139 300 12150 334
rect 12094 266 12150 300
rect 12094 232 12105 266
rect 12139 232 12150 266
rect 12094 198 12150 232
rect 12094 164 12105 198
rect 12139 164 12150 198
rect 12094 130 12150 164
rect 12094 96 12105 130
rect 12139 96 12150 130
rect 12094 62 12150 96
rect 12094 28 12105 62
rect 12139 28 12150 62
rect 12094 -6 12150 28
rect 12094 -40 12105 -6
rect 12139 -40 12150 -6
rect 12094 -52 12150 -40
rect 12550 878 12603 948
rect 12550 844 12561 878
rect 12595 844 12603 878
rect 12550 810 12603 844
rect 12550 776 12561 810
rect 12595 776 12603 810
rect 12550 742 12603 776
rect 12775 930 12828 948
rect 12775 896 12783 930
rect 12817 896 12828 930
rect 12775 862 12828 896
rect 12775 828 12783 862
rect 12817 828 12828 862
rect 12775 794 12828 828
rect 12775 760 12783 794
rect 12817 760 12828 794
rect 12775 748 12828 760
rect 12948 930 13001 948
rect 12948 896 12959 930
rect 12993 896 13001 930
rect 12948 862 13001 896
rect 12948 828 12959 862
rect 12993 828 13001 862
rect 12948 794 13001 828
rect 12948 760 12959 794
rect 12993 760 13001 794
rect 13076 833 15076 844
rect 13076 799 13088 833
rect 13122 799 13156 833
rect 13190 799 13224 833
rect 13258 799 13292 833
rect 13326 799 13360 833
rect 13394 799 13428 833
rect 13462 799 13496 833
rect 13530 799 13564 833
rect 13598 799 13632 833
rect 13666 799 13700 833
rect 13734 799 13768 833
rect 13802 799 13836 833
rect 13870 799 13904 833
rect 13938 799 13972 833
rect 14006 799 14040 833
rect 14074 799 14108 833
rect 14142 799 14176 833
rect 14210 799 14244 833
rect 14278 799 14312 833
rect 14346 799 14380 833
rect 14414 799 14448 833
rect 14482 799 14516 833
rect 14550 799 14584 833
rect 14618 799 14652 833
rect 14686 799 14720 833
rect 14754 799 14788 833
rect 14822 799 14856 833
rect 14890 799 14924 833
rect 14958 799 14992 833
rect 15026 799 15076 833
rect 13076 788 15076 799
rect 15215 1022 15268 1034
rect 15215 988 15223 1022
rect 15257 988 15268 1022
rect 15215 954 15268 988
rect 15215 920 15223 954
rect 15257 920 15268 954
rect 15215 886 15268 920
rect 15215 852 15223 886
rect 15257 852 15268 886
rect 15215 834 15268 852
rect 15448 1022 15504 1034
rect 15448 988 15459 1022
rect 15493 988 15504 1022
rect 15448 954 15504 988
rect 15448 920 15459 954
rect 15493 920 15504 954
rect 15448 886 15504 920
rect 15448 852 15459 886
rect 15493 852 15504 886
rect 15448 834 15504 852
rect 15684 1022 15740 1034
rect 15684 988 15695 1022
rect 15729 988 15740 1022
rect 15684 954 15740 988
rect 15684 920 15695 954
rect 15729 920 15740 954
rect 15684 886 15740 920
rect 15684 852 15695 886
rect 15729 852 15740 886
rect 15684 834 15740 852
rect 15920 1022 15976 1034
rect 15920 988 15931 1022
rect 15965 988 15976 1022
rect 15920 954 15976 988
rect 15920 920 15931 954
rect 15965 920 15976 954
rect 15920 886 15976 920
rect 15920 852 15931 886
rect 15965 852 15976 886
rect 15920 834 15976 852
rect 16156 1022 16209 1034
rect 16156 988 16167 1022
rect 16201 988 16209 1022
rect 16156 954 16209 988
rect 16156 920 16167 954
rect 16201 920 16209 954
rect 16156 886 16209 920
rect 16156 852 16167 886
rect 16201 852 16209 886
rect 16156 834 16209 852
rect 12948 748 13001 760
rect 12550 708 12561 742
rect 12595 708 12603 742
rect 12550 674 12603 708
rect 12550 640 12561 674
rect 12595 640 12603 674
rect 12550 606 12603 640
rect 12550 572 12561 606
rect 12595 572 12603 606
rect 12550 538 12603 572
rect 12550 504 12561 538
rect 12595 504 12603 538
rect 12550 470 12603 504
rect 12550 436 12561 470
rect 12595 436 12603 470
rect 12550 402 12603 436
rect 12550 368 12561 402
rect 12595 368 12603 402
rect 12550 334 12603 368
rect 12550 300 12561 334
rect 12595 300 12603 334
rect 12550 266 12603 300
rect 12550 232 12561 266
rect 12595 232 12603 266
rect 12550 198 12603 232
rect 12550 164 12561 198
rect 12595 164 12603 198
rect 12550 130 12603 164
rect 12550 96 12561 130
rect 12595 96 12603 130
rect 12550 62 12603 96
rect 12550 28 12561 62
rect 12595 28 12603 62
rect 12550 -6 12603 28
rect 12550 -40 12561 -6
rect 12595 -40 12603 -6
rect 12550 -52 12603 -40
rect 13076 597 15076 608
rect 13076 563 13088 597
rect 13122 563 13156 597
rect 13190 563 13224 597
rect 13258 563 13292 597
rect 13326 563 13360 597
rect 13394 563 13428 597
rect 13462 563 13496 597
rect 13530 563 13564 597
rect 13598 563 13632 597
rect 13666 563 13700 597
rect 13734 563 13768 597
rect 13802 563 13836 597
rect 13870 563 13904 597
rect 13938 563 13972 597
rect 14006 563 14040 597
rect 14074 563 14108 597
rect 14142 563 14176 597
rect 14210 563 14244 597
rect 14278 563 14312 597
rect 14346 563 14380 597
rect 14414 563 14448 597
rect 14482 563 14516 597
rect 14550 563 14584 597
rect 14618 563 14652 597
rect 14686 563 14720 597
rect 14754 563 14788 597
rect 14822 563 14856 597
rect 14890 563 14924 597
rect 14958 563 14992 597
rect 15026 563 15076 597
rect 13076 552 15076 563
rect 15215 661 15268 679
rect 15215 627 15223 661
rect 15257 627 15268 661
rect 15215 593 15268 627
rect 15215 559 15223 593
rect 15257 559 15268 593
rect 15215 525 15268 559
rect 15215 491 15223 525
rect 15257 491 15268 525
rect 15215 479 15268 491
rect 15448 661 15504 679
rect 15448 627 15459 661
rect 15493 627 15504 661
rect 15448 593 15504 627
rect 15448 559 15459 593
rect 15493 559 15504 593
rect 15448 525 15504 559
rect 15448 491 15459 525
rect 15493 491 15504 525
rect 15448 479 15504 491
rect 15684 661 15740 679
rect 15684 627 15695 661
rect 15729 627 15740 661
rect 15684 593 15740 627
rect 15684 559 15695 593
rect 15729 559 15740 593
rect 15684 525 15740 559
rect 15684 491 15695 525
rect 15729 491 15740 525
rect 15684 479 15740 491
rect 15920 661 15976 679
rect 15920 627 15931 661
rect 15965 627 15976 661
rect 15920 593 15976 627
rect 15920 559 15931 593
rect 15965 559 15976 593
rect 15920 525 15976 559
rect 15920 491 15931 525
rect 15965 491 15976 525
rect 15920 479 15976 491
rect 16156 661 16209 679
rect 16156 627 16167 661
rect 16201 627 16209 661
rect 16156 593 16209 627
rect 16156 559 16167 593
rect 16201 559 16209 593
rect 16156 525 16209 559
rect 16156 491 16167 525
rect 16201 491 16209 525
rect 16156 479 16209 491
rect 13076 361 15076 372
rect 13076 327 13088 361
rect 13122 327 13156 361
rect 13190 327 13224 361
rect 13258 327 13292 361
rect 13326 327 13360 361
rect 13394 327 13428 361
rect 13462 327 13496 361
rect 13530 327 13564 361
rect 13598 327 13632 361
rect 13666 327 13700 361
rect 13734 327 13768 361
rect 13802 327 13836 361
rect 13870 327 13904 361
rect 13938 327 13972 361
rect 14006 327 14040 361
rect 14074 327 14108 361
rect 14142 327 14176 361
rect 14210 327 14244 361
rect 14278 327 14312 361
rect 14346 327 14380 361
rect 14414 327 14448 361
rect 14482 327 14516 361
rect 14550 327 14584 361
rect 14618 327 14652 361
rect 14686 327 14720 361
rect 14754 327 14788 361
rect 14822 327 14856 361
rect 14890 327 14924 361
rect 14958 327 14992 361
rect 15026 327 15076 361
rect 13076 316 15076 327
rect 13076 125 15076 136
rect 15215 282 15268 294
rect 15215 248 15223 282
rect 15257 248 15268 282
rect 15215 214 15268 248
rect 15215 180 15223 214
rect 15257 180 15268 214
rect 15215 146 15268 180
rect 13076 91 13088 125
rect 13122 91 13156 125
rect 13190 91 13224 125
rect 13258 91 13292 125
rect 13326 91 13360 125
rect 13394 91 13428 125
rect 13462 91 13496 125
rect 13530 91 13564 125
rect 13598 91 13632 125
rect 13666 91 13700 125
rect 13734 91 13768 125
rect 13802 91 13836 125
rect 13870 91 13904 125
rect 13938 91 13972 125
rect 14006 91 14040 125
rect 14074 91 14108 125
rect 14142 91 14176 125
rect 14210 91 14244 125
rect 14278 91 14312 125
rect 14346 91 14380 125
rect 14414 91 14448 125
rect 14482 91 14516 125
rect 14550 91 14584 125
rect 14618 91 14652 125
rect 14686 91 14720 125
rect 14754 91 14788 125
rect 14822 91 14856 125
rect 14890 91 14924 125
rect 14958 91 14992 125
rect 15026 91 15076 125
rect 15215 112 15223 146
rect 15257 112 15268 146
rect 15215 94 15268 112
rect 15448 282 15504 294
rect 15448 248 15459 282
rect 15493 248 15504 282
rect 15448 214 15504 248
rect 15448 180 15459 214
rect 15493 180 15504 214
rect 15448 146 15504 180
rect 15448 112 15459 146
rect 15493 112 15504 146
rect 15448 94 15504 112
rect 15684 282 15737 294
rect 15684 248 15695 282
rect 15729 248 15737 282
rect 18396 338 18596 346
rect 18396 304 18414 338
rect 18448 304 18482 338
rect 18516 304 18550 338
rect 18584 304 18596 338
rect 18396 293 18596 304
rect 15684 214 15737 248
rect 15684 180 15695 214
rect 15729 180 15737 214
rect 15684 146 15737 180
rect 15684 112 15695 146
rect 15729 112 15737 146
rect 15684 94 15737 112
rect 15876 107 15929 177
rect 13076 83 15076 91
rect 15876 73 15884 107
rect 15918 73 15929 107
rect 15876 39 15929 73
rect 15876 5 15884 39
rect 15918 5 15929 39
rect 15876 -29 15929 5
rect 15876 -63 15884 -29
rect 15918 -63 15929 -29
rect 15876 -97 15929 -63
rect 15876 -131 15884 -97
rect 15918 -131 15929 -97
rect 15876 -165 15929 -131
rect 15876 -199 15884 -165
rect 15918 -199 15929 -165
rect 15876 -233 15929 -199
rect 15876 -267 15884 -233
rect 15918 -267 15929 -233
rect 15876 -301 15929 -267
rect 15876 -335 15884 -301
rect 15918 -335 15929 -301
rect 15876 -369 15929 -335
rect 15876 -403 15884 -369
rect 15918 -403 15929 -369
rect 15876 -437 15929 -403
rect 15876 -471 15884 -437
rect 15918 -471 15929 -437
rect 15876 -505 15929 -471
rect 15876 -539 15884 -505
rect 15918 -539 15929 -505
rect 15876 -573 15929 -539
rect 15876 -607 15884 -573
rect 15918 -607 15929 -573
rect 15876 -641 15929 -607
rect 15876 -675 15884 -641
rect 15918 -675 15929 -641
rect 15876 -709 15929 -675
rect 15876 -743 15884 -709
rect 15918 -743 15929 -709
rect 15876 -777 15929 -743
rect 15876 -811 15884 -777
rect 15918 -811 15929 -777
rect 15876 -823 15929 -811
rect 16029 107 16085 177
rect 16029 73 16040 107
rect 16074 73 16085 107
rect 16029 39 16085 73
rect 16029 5 16040 39
rect 16074 5 16085 39
rect 16029 -29 16085 5
rect 16029 -63 16040 -29
rect 16074 -63 16085 -29
rect 16029 -97 16085 -63
rect 16029 -131 16040 -97
rect 16074 -131 16085 -97
rect 16029 -165 16085 -131
rect 16029 -199 16040 -165
rect 16074 -199 16085 -165
rect 16029 -233 16085 -199
rect 16029 -267 16040 -233
rect 16074 -267 16085 -233
rect 16029 -301 16085 -267
rect 16029 -335 16040 -301
rect 16074 -335 16085 -301
rect 16029 -369 16085 -335
rect 16029 -403 16040 -369
rect 16074 -403 16085 -369
rect 16029 -437 16085 -403
rect 16029 -471 16040 -437
rect 16074 -471 16085 -437
rect 16029 -505 16085 -471
rect 16029 -539 16040 -505
rect 16074 -539 16085 -505
rect 16029 -573 16085 -539
rect 16029 -607 16040 -573
rect 16074 -607 16085 -573
rect 16029 -641 16085 -607
rect 16029 -675 16040 -641
rect 16074 -675 16085 -641
rect 16029 -709 16085 -675
rect 16029 -743 16040 -709
rect 16074 -743 16085 -709
rect 16029 -777 16085 -743
rect 16029 -811 16040 -777
rect 16074 -811 16085 -777
rect 16029 -823 16085 -811
rect 16185 107 16238 177
rect 16185 73 16196 107
rect 16230 73 16238 107
rect 16185 39 16238 73
rect 16185 5 16196 39
rect 16230 5 16238 39
rect 16185 -29 16238 5
rect 16185 -63 16196 -29
rect 16230 -63 16238 -29
rect 16185 -97 16238 -63
rect 16185 -131 16196 -97
rect 16230 -131 16238 -97
rect 16185 -165 16238 -131
rect 16185 -199 16196 -165
rect 16230 -199 16238 -165
rect 16185 -233 16238 -199
rect 16185 -267 16196 -233
rect 16230 -267 16238 -233
rect 16185 -301 16238 -267
rect 16185 -335 16196 -301
rect 16230 -335 16238 -301
rect 16185 -369 16238 -335
rect 16185 -403 16196 -369
rect 16230 -403 16238 -369
rect 16185 -437 16238 -403
rect 16185 -471 16196 -437
rect 16230 -471 16238 -437
rect 16185 -505 16238 -471
rect 16185 -539 16196 -505
rect 16230 -539 16238 -505
rect 16185 -573 16238 -539
rect 16185 -607 16196 -573
rect 16230 -607 16238 -573
rect 16185 -641 16238 -607
rect 16185 -675 16196 -641
rect 16230 -675 16238 -641
rect 16185 -709 16238 -675
rect 16185 -743 16196 -709
rect 16230 -743 16238 -709
rect 16185 -777 16238 -743
rect 16185 -811 16196 -777
rect 16230 -811 16238 -777
rect 16185 -823 16238 -811
rect 18396 182 18596 193
rect 18396 148 18414 182
rect 18448 148 18482 182
rect 18516 148 18550 182
rect 18584 148 18596 182
rect 18396 137 18596 148
rect 18396 26 18596 37
rect 18396 -8 18414 26
rect 18448 -8 18482 26
rect 18516 -8 18550 26
rect 18584 -8 18596 26
rect 18396 -16 18596 -8
rect 515 -10956 548 -10922
rect 582 -10956 615 -10922
rect 515 -10964 615 -10956
rect 863 -3369 963 -3360
rect 863 -3403 896 -3369
rect 930 -3403 963 -3369
rect 2616 -9662 2669 -9584
rect 2616 -9696 2624 -9662
rect 2658 -9696 2669 -9662
rect 2616 -9730 2669 -9696
rect 2616 -9764 2624 -9730
rect 2658 -9764 2669 -9730
rect 2616 -9798 2669 -9764
rect 2616 -9832 2624 -9798
rect 2658 -9832 2669 -9798
rect 2616 -9866 2669 -9832
rect 2616 -9900 2624 -9866
rect 2658 -9900 2669 -9866
rect 2616 -9934 2669 -9900
rect 2616 -9968 2624 -9934
rect 2658 -9968 2669 -9934
rect 2616 -10002 2669 -9968
rect 2616 -10036 2624 -10002
rect 2658 -10036 2669 -10002
rect 2616 -10070 2669 -10036
rect 2616 -10104 2624 -10070
rect 2658 -10104 2669 -10070
rect 2616 -10138 2669 -10104
rect 2616 -10172 2624 -10138
rect 2658 -10172 2669 -10138
rect 2616 -10184 2669 -10172
rect 2769 -9662 2825 -9584
rect 2769 -9696 2780 -9662
rect 2814 -9696 2825 -9662
rect 2769 -9730 2825 -9696
rect 2769 -9764 2780 -9730
rect 2814 -9764 2825 -9730
rect 2769 -9798 2825 -9764
rect 2769 -9832 2780 -9798
rect 2814 -9832 2825 -9798
rect 2769 -9866 2825 -9832
rect 2769 -9900 2780 -9866
rect 2814 -9900 2825 -9866
rect 2769 -9934 2825 -9900
rect 2769 -9968 2780 -9934
rect 2814 -9968 2825 -9934
rect 2769 -10002 2825 -9968
rect 2769 -10036 2780 -10002
rect 2814 -10036 2825 -10002
rect 2769 -10070 2825 -10036
rect 2769 -10104 2780 -10070
rect 2814 -10104 2825 -10070
rect 2769 -10138 2825 -10104
rect 2769 -10172 2780 -10138
rect 2814 -10172 2825 -10138
rect 2769 -10184 2825 -10172
rect 2925 -9662 2978 -9584
rect 2925 -9696 2936 -9662
rect 2970 -9696 2978 -9662
rect 2925 -9730 2978 -9696
rect 2925 -9764 2936 -9730
rect 2970 -9764 2978 -9730
rect 2925 -9798 2978 -9764
rect 2925 -9832 2936 -9798
rect 2970 -9832 2978 -9798
rect 2925 -9866 2978 -9832
rect 2925 -9900 2936 -9866
rect 2970 -9900 2978 -9866
rect 2925 -9934 2978 -9900
rect 2925 -9968 2936 -9934
rect 2970 -9968 2978 -9934
rect 2925 -10002 2978 -9968
rect 2925 -10036 2936 -10002
rect 2970 -10036 2978 -10002
rect 2925 -10070 2978 -10036
rect 2925 -10104 2936 -10070
rect 2970 -10104 2978 -10070
rect 2925 -10138 2978 -10104
rect 2925 -10172 2936 -10138
rect 2970 -10172 2978 -10138
rect 2925 -10184 2978 -10172
<< mvpdiff >>
rect 8706 4792 8759 4804
rect 8706 4758 8714 4792
rect 8748 4758 8759 4792
rect 8706 4724 8759 4758
rect 8706 4690 8714 4724
rect 8748 4690 8759 4724
rect 8706 4656 8759 4690
rect 8706 4622 8714 4656
rect 8748 4622 8759 4656
rect 8706 4588 8759 4622
rect 8706 4554 8714 4588
rect 8748 4554 8759 4588
rect 8706 4520 8759 4554
rect 8706 4486 8714 4520
rect 8748 4486 8759 4520
rect 8706 4452 8759 4486
rect 8706 4418 8714 4452
rect 8748 4418 8759 4452
rect 8706 4384 8759 4418
rect 8706 4350 8714 4384
rect 8748 4350 8759 4384
rect 8706 4316 8759 4350
rect 8706 4282 8714 4316
rect 8748 4282 8759 4316
rect 8706 4248 8759 4282
rect 8706 4214 8714 4248
rect 8748 4214 8759 4248
rect 8706 4180 8759 4214
rect 8706 4146 8714 4180
rect 8748 4146 8759 4180
rect 8706 4112 8759 4146
rect 8706 4078 8714 4112
rect 8748 4078 8759 4112
rect 8706 4044 8759 4078
rect 8706 4010 8714 4044
rect 8748 4010 8759 4044
rect 8706 3976 8759 4010
rect 8706 3942 8714 3976
rect 8748 3942 8759 3976
rect 8706 3908 8759 3942
rect 8706 3874 8714 3908
rect 8748 3874 8759 3908
rect 8706 3804 8759 3874
rect 8859 4792 8915 4804
rect 8859 4758 8870 4792
rect 8904 4758 8915 4792
rect 8859 4724 8915 4758
rect 8859 4690 8870 4724
rect 8904 4690 8915 4724
rect 8859 4656 8915 4690
rect 8859 4622 8870 4656
rect 8904 4622 8915 4656
rect 8859 4588 8915 4622
rect 8859 4554 8870 4588
rect 8904 4554 8915 4588
rect 8859 4520 8915 4554
rect 8859 4486 8870 4520
rect 8904 4486 8915 4520
rect 8859 4452 8915 4486
rect 8859 4418 8870 4452
rect 8904 4418 8915 4452
rect 8859 4384 8915 4418
rect 8859 4350 8870 4384
rect 8904 4350 8915 4384
rect 8859 4316 8915 4350
rect 8859 4282 8870 4316
rect 8904 4282 8915 4316
rect 8859 4248 8915 4282
rect 8859 4214 8870 4248
rect 8904 4214 8915 4248
rect 8859 4180 8915 4214
rect 8859 4146 8870 4180
rect 8904 4146 8915 4180
rect 8859 4112 8915 4146
rect 8859 4078 8870 4112
rect 8904 4078 8915 4112
rect 8859 4044 8915 4078
rect 8859 4010 8870 4044
rect 8904 4010 8915 4044
rect 8859 3976 8915 4010
rect 8859 3942 8870 3976
rect 8904 3942 8915 3976
rect 8859 3908 8915 3942
rect 8859 3874 8870 3908
rect 8904 3874 8915 3908
rect 8859 3804 8915 3874
rect 9015 4792 9071 4804
rect 9015 4758 9026 4792
rect 9060 4758 9071 4792
rect 9015 4724 9071 4758
rect 9015 4690 9026 4724
rect 9060 4690 9071 4724
rect 9015 4656 9071 4690
rect 9015 4622 9026 4656
rect 9060 4622 9071 4656
rect 9015 4588 9071 4622
rect 9015 4554 9026 4588
rect 9060 4554 9071 4588
rect 9015 4520 9071 4554
rect 9015 4486 9026 4520
rect 9060 4486 9071 4520
rect 9015 4452 9071 4486
rect 9015 4418 9026 4452
rect 9060 4418 9071 4452
rect 9015 4384 9071 4418
rect 9015 4350 9026 4384
rect 9060 4350 9071 4384
rect 9015 4316 9071 4350
rect 9015 4282 9026 4316
rect 9060 4282 9071 4316
rect 9015 4248 9071 4282
rect 9015 4214 9026 4248
rect 9060 4214 9071 4248
rect 9015 4180 9071 4214
rect 9015 4146 9026 4180
rect 9060 4146 9071 4180
rect 9015 4112 9071 4146
rect 9015 4078 9026 4112
rect 9060 4078 9071 4112
rect 9015 4044 9071 4078
rect 9015 4010 9026 4044
rect 9060 4010 9071 4044
rect 9015 3976 9071 4010
rect 9015 3942 9026 3976
rect 9060 3942 9071 3976
rect 9015 3908 9071 3942
rect 9015 3874 9026 3908
rect 9060 3874 9071 3908
rect 9015 3804 9071 3874
rect 9171 4792 9227 4804
rect 9171 4758 9182 4792
rect 9216 4758 9227 4792
rect 9171 4724 9227 4758
rect 9171 4690 9182 4724
rect 9216 4690 9227 4724
rect 9171 4656 9227 4690
rect 9171 4622 9182 4656
rect 9216 4622 9227 4656
rect 9171 4588 9227 4622
rect 9171 4554 9182 4588
rect 9216 4554 9227 4588
rect 9171 4520 9227 4554
rect 9171 4486 9182 4520
rect 9216 4486 9227 4520
rect 9171 4452 9227 4486
rect 9171 4418 9182 4452
rect 9216 4418 9227 4452
rect 9171 4384 9227 4418
rect 9171 4350 9182 4384
rect 9216 4350 9227 4384
rect 9171 4316 9227 4350
rect 9171 4282 9182 4316
rect 9216 4282 9227 4316
rect 9171 4248 9227 4282
rect 9171 4214 9182 4248
rect 9216 4214 9227 4248
rect 9171 4180 9227 4214
rect 9171 4146 9182 4180
rect 9216 4146 9227 4180
rect 9171 4112 9227 4146
rect 9171 4078 9182 4112
rect 9216 4078 9227 4112
rect 9171 4044 9227 4078
rect 9171 4010 9182 4044
rect 9216 4010 9227 4044
rect 9171 3976 9227 4010
rect 9171 3942 9182 3976
rect 9216 3942 9227 3976
rect 9171 3908 9227 3942
rect 9171 3874 9182 3908
rect 9216 3874 9227 3908
rect 9171 3804 9227 3874
rect 9327 4792 9380 4804
rect 9327 4758 9338 4792
rect 9372 4758 9380 4792
rect 9327 4724 9380 4758
rect 9327 4690 9338 4724
rect 9372 4690 9380 4724
rect 9327 4656 9380 4690
rect 9327 4622 9338 4656
rect 9372 4622 9380 4656
rect 9327 4588 9380 4622
rect 9327 4554 9338 4588
rect 9372 4554 9380 4588
rect 9327 4520 9380 4554
rect 9327 4486 9338 4520
rect 9372 4486 9380 4520
rect 9327 4452 9380 4486
rect 9327 4418 9338 4452
rect 9372 4418 9380 4452
rect 9327 4384 9380 4418
rect 9327 4350 9338 4384
rect 9372 4350 9380 4384
rect 9327 4316 9380 4350
rect 9327 4282 9338 4316
rect 9372 4282 9380 4316
rect 9327 4248 9380 4282
rect 9327 4214 9338 4248
rect 9372 4214 9380 4248
rect 9327 4180 9380 4214
rect 9327 4146 9338 4180
rect 9372 4146 9380 4180
rect 9327 4112 9380 4146
rect 9327 4078 9338 4112
rect 9372 4078 9380 4112
rect 9327 4044 9380 4078
rect 9327 4010 9338 4044
rect 9372 4010 9380 4044
rect 9327 3976 9380 4010
rect 9327 3942 9338 3976
rect 9372 3942 9380 3976
rect 9327 3908 9380 3942
rect 9327 3874 9338 3908
rect 9372 3874 9380 3908
rect 9327 3804 9380 3874
rect 9454 4792 9507 4804
rect 9454 4758 9462 4792
rect 9496 4758 9507 4792
rect 9454 4724 9507 4758
rect 9454 4690 9462 4724
rect 9496 4690 9507 4724
rect 9454 4656 9507 4690
rect 9454 4622 9462 4656
rect 9496 4622 9507 4656
rect 9454 4588 9507 4622
rect 9454 4554 9462 4588
rect 9496 4554 9507 4588
rect 9454 4520 9507 4554
rect 9454 4486 9462 4520
rect 9496 4486 9507 4520
rect 9454 4452 9507 4486
rect 9454 4418 9462 4452
rect 9496 4418 9507 4452
rect 9454 4384 9507 4418
rect 9454 4350 9462 4384
rect 9496 4350 9507 4384
rect 9454 4316 9507 4350
rect 9454 4282 9462 4316
rect 9496 4282 9507 4316
rect 9454 4248 9507 4282
rect 9454 4214 9462 4248
rect 9496 4214 9507 4248
rect 9454 4180 9507 4214
rect 9454 4146 9462 4180
rect 9496 4146 9507 4180
rect 9454 4112 9507 4146
rect 9454 4078 9462 4112
rect 9496 4078 9507 4112
rect 9454 4044 9507 4078
rect 9454 4010 9462 4044
rect 9496 4010 9507 4044
rect 9454 3976 9507 4010
rect 9454 3942 9462 3976
rect 9496 3942 9507 3976
rect 9454 3908 9507 3942
rect 9454 3874 9462 3908
rect 9496 3874 9507 3908
rect 9454 3804 9507 3874
rect 9607 4792 9660 4804
rect 9607 4758 9618 4792
rect 9652 4758 9660 4792
rect 9607 4724 9660 4758
rect 9607 4690 9618 4724
rect 9652 4690 9660 4724
rect 9607 4656 9660 4690
rect 9607 4622 9618 4656
rect 9652 4622 9660 4656
rect 9607 4588 9660 4622
rect 9607 4554 9618 4588
rect 9652 4554 9660 4588
rect 9607 4520 9660 4554
rect 9607 4486 9618 4520
rect 9652 4486 9660 4520
rect 9607 4452 9660 4486
rect 9607 4418 9618 4452
rect 9652 4418 9660 4452
rect 9607 4384 9660 4418
rect 9607 4350 9618 4384
rect 9652 4350 9660 4384
rect 9607 4316 9660 4350
rect 9607 4282 9618 4316
rect 9652 4282 9660 4316
rect 9607 4248 9660 4282
rect 9607 4214 9618 4248
rect 9652 4214 9660 4248
rect 9607 4180 9660 4214
rect 9607 4146 9618 4180
rect 9652 4146 9660 4180
rect 9607 4112 9660 4146
rect 9607 4078 9618 4112
rect 9652 4078 9660 4112
rect 9607 4044 9660 4078
rect 9607 4010 9618 4044
rect 9652 4010 9660 4044
rect 9607 3976 9660 4010
rect 9607 3942 9618 3976
rect 9652 3942 9660 3976
rect 9607 3908 9660 3942
rect 9607 3874 9618 3908
rect 9652 3874 9660 3908
rect 9607 3804 9660 3874
rect 9734 4792 9787 4804
rect 9734 4758 9742 4792
rect 9776 4758 9787 4792
rect 9734 4724 9787 4758
rect 9734 4690 9742 4724
rect 9776 4690 9787 4724
rect 9734 4656 9787 4690
rect 9734 4622 9742 4656
rect 9776 4622 9787 4656
rect 9734 4588 9787 4622
rect 9734 4554 9742 4588
rect 9776 4554 9787 4588
rect 9734 4520 9787 4554
rect 9734 4486 9742 4520
rect 9776 4486 9787 4520
rect 9734 4452 9787 4486
rect 9734 4418 9742 4452
rect 9776 4418 9787 4452
rect 9734 4384 9787 4418
rect 9734 4350 9742 4384
rect 9776 4350 9787 4384
rect 9734 4316 9787 4350
rect 9734 4282 9742 4316
rect 9776 4282 9787 4316
rect 9734 4248 9787 4282
rect 9734 4214 9742 4248
rect 9776 4214 9787 4248
rect 9734 4180 9787 4214
rect 9734 4146 9742 4180
rect 9776 4146 9787 4180
rect 9734 4112 9787 4146
rect 9734 4078 9742 4112
rect 9776 4078 9787 4112
rect 9734 4044 9787 4078
rect 9734 4010 9742 4044
rect 9776 4010 9787 4044
rect 9734 3976 9787 4010
rect 9734 3942 9742 3976
rect 9776 3942 9787 3976
rect 9734 3908 9787 3942
rect 9734 3874 9742 3908
rect 9776 3874 9787 3908
rect 9734 3804 9787 3874
rect 9887 4792 9943 4804
rect 9887 4758 9898 4792
rect 9932 4758 9943 4792
rect 9887 4724 9943 4758
rect 9887 4690 9898 4724
rect 9932 4690 9943 4724
rect 9887 4656 9943 4690
rect 9887 4622 9898 4656
rect 9932 4622 9943 4656
rect 9887 4588 9943 4622
rect 9887 4554 9898 4588
rect 9932 4554 9943 4588
rect 9887 4520 9943 4554
rect 9887 4486 9898 4520
rect 9932 4486 9943 4520
rect 9887 4452 9943 4486
rect 9887 4418 9898 4452
rect 9932 4418 9943 4452
rect 9887 4384 9943 4418
rect 9887 4350 9898 4384
rect 9932 4350 9943 4384
rect 9887 4316 9943 4350
rect 9887 4282 9898 4316
rect 9932 4282 9943 4316
rect 9887 4248 9943 4282
rect 9887 4214 9898 4248
rect 9932 4214 9943 4248
rect 9887 4180 9943 4214
rect 9887 4146 9898 4180
rect 9932 4146 9943 4180
rect 9887 4112 9943 4146
rect 9887 4078 9898 4112
rect 9932 4078 9943 4112
rect 9887 4044 9943 4078
rect 9887 4010 9898 4044
rect 9932 4010 9943 4044
rect 9887 3976 9943 4010
rect 9887 3942 9898 3976
rect 9932 3942 9943 3976
rect 9887 3908 9943 3942
rect 9887 3874 9898 3908
rect 9932 3874 9943 3908
rect 9887 3804 9943 3874
rect 10043 4792 10096 4804
rect 10043 4758 10054 4792
rect 10088 4758 10096 4792
rect 10043 4724 10096 4758
rect 10043 4690 10054 4724
rect 10088 4690 10096 4724
rect 10043 4656 10096 4690
rect 10043 4622 10054 4656
rect 10088 4622 10096 4656
rect 10043 4588 10096 4622
rect 10043 4554 10054 4588
rect 10088 4554 10096 4588
rect 10043 4520 10096 4554
rect 10043 4486 10054 4520
rect 10088 4486 10096 4520
rect 10043 4452 10096 4486
rect 10043 4418 10054 4452
rect 10088 4418 10096 4452
rect 10043 4384 10096 4418
rect 10043 4350 10054 4384
rect 10088 4350 10096 4384
rect 10043 4316 10096 4350
rect 10043 4282 10054 4316
rect 10088 4282 10096 4316
rect 10043 4248 10096 4282
rect 10043 4214 10054 4248
rect 10088 4214 10096 4248
rect 10043 4180 10096 4214
rect 10043 4146 10054 4180
rect 10088 4146 10096 4180
rect 10043 4112 10096 4146
rect 10043 4078 10054 4112
rect 10088 4078 10096 4112
rect 10043 4044 10096 4078
rect 10043 4010 10054 4044
rect 10088 4010 10096 4044
rect 10043 3976 10096 4010
rect 10043 3942 10054 3976
rect 10088 3942 10096 3976
rect 10043 3908 10096 3942
rect 10043 3874 10054 3908
rect 10088 3874 10096 3908
rect 10043 3804 10096 3874
rect 10323 4792 10376 4804
rect 10323 4758 10331 4792
rect 10365 4758 10376 4792
rect 10323 4724 10376 4758
rect 10323 4690 10331 4724
rect 10365 4690 10376 4724
rect 10323 4656 10376 4690
rect 10323 4622 10331 4656
rect 10365 4622 10376 4656
rect 10323 4588 10376 4622
rect 10323 4554 10331 4588
rect 10365 4554 10376 4588
rect 10323 4520 10376 4554
rect 10323 4486 10331 4520
rect 10365 4486 10376 4520
rect 10323 4452 10376 4486
rect 10323 4418 10331 4452
rect 10365 4418 10376 4452
rect 10323 4384 10376 4418
rect 10323 4350 10331 4384
rect 10365 4350 10376 4384
rect 10323 4316 10376 4350
rect 10323 4282 10331 4316
rect 10365 4282 10376 4316
rect 10323 4248 10376 4282
rect 10323 4214 10331 4248
rect 10365 4214 10376 4248
rect 10323 4180 10376 4214
rect 10323 4146 10331 4180
rect 10365 4146 10376 4180
rect 10323 4112 10376 4146
rect 10323 4078 10331 4112
rect 10365 4078 10376 4112
rect 10323 4044 10376 4078
rect 10323 4010 10331 4044
rect 10365 4010 10376 4044
rect 10323 3976 10376 4010
rect 10323 3942 10331 3976
rect 10365 3942 10376 3976
rect 10323 3908 10376 3942
rect 10323 3874 10331 3908
rect 10365 3874 10376 3908
rect 10323 3804 10376 3874
rect 10476 4792 10532 4804
rect 10476 4758 10487 4792
rect 10521 4758 10532 4792
rect 10476 4724 10532 4758
rect 10476 4690 10487 4724
rect 10521 4690 10532 4724
rect 10476 4656 10532 4690
rect 10476 4622 10487 4656
rect 10521 4622 10532 4656
rect 10476 4588 10532 4622
rect 10476 4554 10487 4588
rect 10521 4554 10532 4588
rect 10476 4520 10532 4554
rect 10476 4486 10487 4520
rect 10521 4486 10532 4520
rect 10476 4452 10532 4486
rect 10476 4418 10487 4452
rect 10521 4418 10532 4452
rect 10476 4384 10532 4418
rect 10476 4350 10487 4384
rect 10521 4350 10532 4384
rect 10476 4316 10532 4350
rect 10476 4282 10487 4316
rect 10521 4282 10532 4316
rect 10476 4248 10532 4282
rect 10476 4214 10487 4248
rect 10521 4214 10532 4248
rect 10476 4180 10532 4214
rect 10476 4146 10487 4180
rect 10521 4146 10532 4180
rect 10476 4112 10532 4146
rect 10476 4078 10487 4112
rect 10521 4078 10532 4112
rect 10476 4044 10532 4078
rect 10476 4010 10487 4044
rect 10521 4010 10532 4044
rect 10476 3976 10532 4010
rect 10476 3942 10487 3976
rect 10521 3942 10532 3976
rect 10476 3908 10532 3942
rect 10476 3874 10487 3908
rect 10521 3874 10532 3908
rect 10476 3804 10532 3874
rect 10632 4792 10688 4804
rect 10632 4758 10643 4792
rect 10677 4758 10688 4792
rect 10632 4724 10688 4758
rect 10632 4690 10643 4724
rect 10677 4690 10688 4724
rect 10632 4656 10688 4690
rect 10632 4622 10643 4656
rect 10677 4622 10688 4656
rect 10632 4588 10688 4622
rect 10632 4554 10643 4588
rect 10677 4554 10688 4588
rect 10632 4520 10688 4554
rect 10632 4486 10643 4520
rect 10677 4486 10688 4520
rect 10632 4452 10688 4486
rect 10632 4418 10643 4452
rect 10677 4418 10688 4452
rect 10632 4384 10688 4418
rect 10632 4350 10643 4384
rect 10677 4350 10688 4384
rect 10632 4316 10688 4350
rect 10632 4282 10643 4316
rect 10677 4282 10688 4316
rect 10632 4248 10688 4282
rect 10632 4214 10643 4248
rect 10677 4214 10688 4248
rect 10632 4180 10688 4214
rect 10632 4146 10643 4180
rect 10677 4146 10688 4180
rect 10632 4112 10688 4146
rect 10632 4078 10643 4112
rect 10677 4078 10688 4112
rect 10632 4044 10688 4078
rect 10632 4010 10643 4044
rect 10677 4010 10688 4044
rect 10632 3976 10688 4010
rect 10632 3942 10643 3976
rect 10677 3942 10688 3976
rect 10632 3908 10688 3942
rect 10632 3874 10643 3908
rect 10677 3874 10688 3908
rect 10632 3804 10688 3874
rect 10788 4792 10844 4804
rect 10788 4758 10799 4792
rect 10833 4758 10844 4792
rect 10788 4724 10844 4758
rect 10788 4690 10799 4724
rect 10833 4690 10844 4724
rect 10788 4656 10844 4690
rect 10788 4622 10799 4656
rect 10833 4622 10844 4656
rect 10788 4588 10844 4622
rect 10788 4554 10799 4588
rect 10833 4554 10844 4588
rect 10788 4520 10844 4554
rect 10788 4486 10799 4520
rect 10833 4486 10844 4520
rect 10788 4452 10844 4486
rect 10788 4418 10799 4452
rect 10833 4418 10844 4452
rect 10788 4384 10844 4418
rect 10788 4350 10799 4384
rect 10833 4350 10844 4384
rect 10788 4316 10844 4350
rect 10788 4282 10799 4316
rect 10833 4282 10844 4316
rect 10788 4248 10844 4282
rect 10788 4214 10799 4248
rect 10833 4214 10844 4248
rect 10788 4180 10844 4214
rect 10788 4146 10799 4180
rect 10833 4146 10844 4180
rect 10788 4112 10844 4146
rect 10788 4078 10799 4112
rect 10833 4078 10844 4112
rect 10788 4044 10844 4078
rect 10788 4010 10799 4044
rect 10833 4010 10844 4044
rect 10788 3976 10844 4010
rect 10788 3942 10799 3976
rect 10833 3942 10844 3976
rect 10788 3908 10844 3942
rect 10788 3874 10799 3908
rect 10833 3874 10844 3908
rect 10788 3804 10844 3874
rect 10944 4792 11000 4804
rect 10944 4758 10955 4792
rect 10989 4758 11000 4792
rect 10944 4724 11000 4758
rect 10944 4690 10955 4724
rect 10989 4690 11000 4724
rect 10944 4656 11000 4690
rect 10944 4622 10955 4656
rect 10989 4622 11000 4656
rect 10944 4588 11000 4622
rect 10944 4554 10955 4588
rect 10989 4554 11000 4588
rect 10944 4520 11000 4554
rect 10944 4486 10955 4520
rect 10989 4486 11000 4520
rect 10944 4452 11000 4486
rect 10944 4418 10955 4452
rect 10989 4418 11000 4452
rect 10944 4384 11000 4418
rect 10944 4350 10955 4384
rect 10989 4350 11000 4384
rect 10944 4316 11000 4350
rect 10944 4282 10955 4316
rect 10989 4282 11000 4316
rect 10944 4248 11000 4282
rect 10944 4214 10955 4248
rect 10989 4214 11000 4248
rect 10944 4180 11000 4214
rect 10944 4146 10955 4180
rect 10989 4146 11000 4180
rect 10944 4112 11000 4146
rect 10944 4078 10955 4112
rect 10989 4078 11000 4112
rect 10944 4044 11000 4078
rect 10944 4010 10955 4044
rect 10989 4010 11000 4044
rect 10944 3976 11000 4010
rect 10944 3942 10955 3976
rect 10989 3942 11000 3976
rect 10944 3908 11000 3942
rect 10944 3874 10955 3908
rect 10989 3874 11000 3908
rect 10944 3804 11000 3874
rect 11100 4792 11153 4804
rect 11100 4758 11111 4792
rect 11145 4758 11153 4792
rect 11100 4724 11153 4758
rect 11100 4690 11111 4724
rect 11145 4690 11153 4724
rect 11100 4656 11153 4690
rect 11100 4622 11111 4656
rect 11145 4622 11153 4656
rect 11100 4588 11153 4622
rect 11100 4554 11111 4588
rect 11145 4554 11153 4588
rect 11100 4520 11153 4554
rect 11100 4486 11111 4520
rect 11145 4486 11153 4520
rect 11100 4452 11153 4486
rect 11100 4418 11111 4452
rect 11145 4418 11153 4452
rect 11100 4384 11153 4418
rect 11100 4350 11111 4384
rect 11145 4350 11153 4384
rect 11100 4316 11153 4350
rect 11100 4282 11111 4316
rect 11145 4282 11153 4316
rect 11100 4248 11153 4282
rect 11100 4214 11111 4248
rect 11145 4214 11153 4248
rect 11100 4180 11153 4214
rect 11100 4146 11111 4180
rect 11145 4146 11153 4180
rect 11100 4112 11153 4146
rect 11100 4078 11111 4112
rect 11145 4078 11153 4112
rect 11100 4044 11153 4078
rect 11100 4010 11111 4044
rect 11145 4010 11153 4044
rect 11100 3976 11153 4010
rect 11100 3942 11111 3976
rect 11145 3942 11153 3976
rect 11100 3908 11153 3942
rect 11100 3874 11111 3908
rect 11145 3874 11153 3908
rect 11100 3804 11153 3874
rect 10571 3523 10624 3561
rect 8893 3509 9893 3517
rect 8893 3475 8905 3509
rect 8939 3475 8973 3509
rect 9007 3475 9041 3509
rect 9075 3475 9109 3509
rect 9143 3475 9177 3509
rect 9211 3475 9245 3509
rect 9279 3475 9313 3509
rect 9347 3475 9381 3509
rect 9415 3475 9449 3509
rect 9483 3475 9517 3509
rect 9551 3475 9585 3509
rect 9619 3475 9653 3509
rect 9687 3475 9721 3509
rect 9755 3475 9789 3509
rect 9823 3475 9893 3509
rect 10571 3489 10579 3523
rect 10613 3489 10624 3523
rect 10571 3477 10624 3489
rect 10824 3523 10877 3561
rect 10824 3489 10835 3523
rect 10869 3489 10877 3523
rect 10824 3477 10877 3489
rect 8893 3464 9893 3475
rect 8893 3353 9893 3364
rect 8893 3319 8905 3353
rect 8939 3319 8973 3353
rect 9007 3319 9041 3353
rect 9075 3319 9109 3353
rect 9143 3319 9177 3353
rect 9211 3319 9245 3353
rect 9279 3319 9313 3353
rect 9347 3319 9381 3353
rect 9415 3319 9449 3353
rect 9483 3319 9517 3353
rect 9551 3319 9585 3353
rect 9619 3319 9653 3353
rect 9687 3319 9721 3353
rect 9755 3319 9789 3353
rect 9823 3319 9893 3353
rect 8893 3308 9893 3319
rect 10152 3370 11152 3378
rect 10152 3336 10222 3370
rect 10256 3336 10290 3370
rect 10324 3336 10358 3370
rect 10392 3336 10426 3370
rect 10460 3336 10494 3370
rect 10528 3336 10562 3370
rect 10596 3336 10630 3370
rect 10664 3336 10698 3370
rect 10732 3336 10766 3370
rect 10800 3336 10834 3370
rect 10868 3336 10902 3370
rect 10936 3336 10970 3370
rect 11004 3336 11038 3370
rect 11072 3336 11106 3370
rect 11140 3336 11152 3370
rect 10152 3325 11152 3336
rect 10152 3214 11152 3225
rect 8893 3197 9893 3208
rect 8893 3163 8905 3197
rect 8939 3163 8973 3197
rect 9007 3163 9041 3197
rect 9075 3163 9109 3197
rect 9143 3163 9177 3197
rect 9211 3163 9245 3197
rect 9279 3163 9313 3197
rect 9347 3163 9381 3197
rect 9415 3163 9449 3197
rect 9483 3163 9517 3197
rect 9551 3163 9585 3197
rect 9619 3163 9653 3197
rect 9687 3163 9721 3197
rect 9755 3163 9789 3197
rect 9823 3163 9893 3197
rect 10152 3180 10222 3214
rect 10256 3180 10290 3214
rect 10324 3180 10358 3214
rect 10392 3180 10426 3214
rect 10460 3180 10494 3214
rect 10528 3180 10562 3214
rect 10596 3180 10630 3214
rect 10664 3180 10698 3214
rect 10732 3180 10766 3214
rect 10800 3180 10834 3214
rect 10868 3180 10902 3214
rect 10936 3180 10970 3214
rect 11004 3180 11038 3214
rect 11072 3180 11106 3214
rect 11140 3180 11152 3214
rect 10152 3172 11152 3180
rect 8893 3155 9893 3163
rect 16971 3229 17571 3237
rect 16971 3195 17049 3229
rect 17083 3195 17117 3229
rect 17151 3195 17185 3229
rect 17219 3195 17253 3229
rect 17287 3195 17321 3229
rect 17355 3195 17389 3229
rect 17423 3195 17457 3229
rect 17491 3195 17525 3229
rect 17559 3195 17571 3229
rect 16971 3184 17571 3195
rect 17790 3216 17843 3234
rect 16971 3053 17571 3064
rect 16971 3019 17049 3053
rect 17083 3019 17117 3053
rect 17151 3019 17185 3053
rect 17219 3019 17253 3053
rect 17287 3019 17321 3053
rect 17355 3019 17389 3053
rect 17423 3019 17457 3053
rect 17491 3019 17525 3053
rect 17559 3019 17571 3053
rect 17790 3182 17798 3216
rect 17832 3182 17843 3216
rect 17790 3148 17843 3182
rect 17790 3114 17798 3148
rect 17832 3114 17843 3148
rect 17790 3080 17843 3114
rect 17790 3046 17798 3080
rect 17832 3046 17843 3080
rect 17790 3034 17843 3046
rect 17943 3216 17999 3234
rect 17943 3182 17954 3216
rect 17988 3182 17999 3216
rect 17943 3148 17999 3182
rect 17943 3114 17954 3148
rect 17988 3114 17999 3148
rect 17943 3080 17999 3114
rect 17943 3046 17954 3080
rect 17988 3046 17999 3080
rect 17943 3034 17999 3046
rect 18099 3216 18152 3234
rect 18099 3182 18110 3216
rect 18144 3182 18152 3216
rect 18099 3148 18152 3182
rect 18099 3114 18110 3148
rect 18144 3114 18152 3148
rect 18099 3080 18152 3114
rect 18099 3046 18110 3080
rect 18144 3046 18152 3080
rect 18099 3034 18152 3046
rect 18274 3216 18327 3234
rect 18274 3182 18282 3216
rect 18316 3182 18327 3216
rect 18274 3148 18327 3182
rect 18274 3114 18282 3148
rect 18316 3114 18327 3148
rect 18274 3080 18327 3114
rect 18274 3046 18282 3080
rect 18316 3046 18327 3080
rect 18274 3034 18327 3046
rect 18427 3216 18483 3234
rect 18427 3182 18438 3216
rect 18472 3182 18483 3216
rect 18427 3148 18483 3182
rect 18427 3114 18438 3148
rect 18472 3114 18483 3148
rect 18427 3080 18483 3114
rect 18427 3046 18438 3080
rect 18472 3046 18483 3080
rect 18427 3034 18483 3046
rect 18583 3216 18636 3234
rect 18583 3182 18594 3216
rect 18628 3182 18636 3216
rect 18583 3148 18636 3182
rect 18583 3114 18594 3148
rect 18628 3114 18636 3148
rect 18583 3080 18636 3114
rect 18583 3046 18594 3080
rect 18628 3046 18636 3080
rect 18583 3034 18636 3046
rect 18736 3216 18789 3234
rect 18736 3182 18744 3216
rect 18778 3182 18789 3216
rect 18736 3148 18789 3182
rect 18736 3114 18744 3148
rect 18778 3114 18789 3148
rect 18736 3080 18789 3114
rect 18736 3046 18744 3080
rect 18778 3046 18789 3080
rect 18736 3034 18789 3046
rect 18889 3216 18945 3234
rect 18889 3182 18900 3216
rect 18934 3182 18945 3216
rect 18889 3148 18945 3182
rect 18889 3114 18900 3148
rect 18934 3114 18945 3148
rect 18889 3080 18945 3114
rect 18889 3046 18900 3080
rect 18934 3046 18945 3080
rect 18889 3034 18945 3046
rect 19045 3216 19098 3234
rect 19045 3182 19056 3216
rect 19090 3182 19098 3216
rect 19045 3148 19098 3182
rect 19045 3114 19056 3148
rect 19090 3114 19098 3148
rect 19045 3080 19098 3114
rect 19045 3046 19056 3080
rect 19090 3046 19098 3080
rect 19045 3034 19098 3046
rect 16971 3011 17571 3019
rect 18086 2883 19086 2891
rect 18086 2849 18156 2883
rect 18190 2849 18224 2883
rect 18258 2849 18292 2883
rect 18326 2849 18360 2883
rect 18394 2849 18428 2883
rect 18462 2849 18496 2883
rect 18530 2849 18564 2883
rect 18598 2849 18632 2883
rect 18666 2849 18700 2883
rect 18734 2849 18768 2883
rect 18802 2849 18836 2883
rect 18870 2849 18904 2883
rect 18938 2849 18972 2883
rect 19006 2849 19040 2883
rect 19074 2849 19086 2883
rect 18086 2838 19086 2849
rect 574 2433 1574 2441
rect 574 2399 586 2433
rect 620 2399 654 2433
rect 688 2399 722 2433
rect 756 2399 790 2433
rect 824 2399 858 2433
rect 892 2399 926 2433
rect 960 2399 994 2433
rect 1028 2399 1062 2433
rect 1096 2399 1130 2433
rect 1164 2399 1198 2433
rect 1232 2399 1266 2433
rect 1300 2399 1334 2433
rect 1368 2399 1402 2433
rect 1436 2399 1470 2433
rect 1504 2399 1574 2433
rect 574 2388 1574 2399
rect 574 2277 1574 2288
rect 574 2243 586 2277
rect 620 2243 654 2277
rect 688 2243 722 2277
rect 756 2243 790 2277
rect 824 2243 858 2277
rect 892 2243 926 2277
rect 960 2243 994 2277
rect 1028 2243 1062 2277
rect 1096 2243 1130 2277
rect 1164 2243 1198 2277
rect 1232 2243 1266 2277
rect 1300 2243 1334 2277
rect 1368 2243 1402 2277
rect 1436 2243 1470 2277
rect 1504 2243 1574 2277
rect 574 2235 1574 2243
rect 574 1841 1574 1849
rect 574 1807 586 1841
rect 620 1807 654 1841
rect 688 1807 722 1841
rect 756 1807 790 1841
rect 824 1807 858 1841
rect 892 1807 926 1841
rect 960 1807 994 1841
rect 1028 1807 1062 1841
rect 1096 1807 1130 1841
rect 1164 1807 1198 1841
rect 1232 1807 1266 1841
rect 1300 1807 1334 1841
rect 1368 1807 1402 1841
rect 1436 1807 1470 1841
rect 1504 1807 1574 1841
rect 574 1796 1574 1807
rect 574 1685 1574 1696
rect 574 1651 586 1685
rect 620 1651 654 1685
rect 688 1651 722 1685
rect 756 1651 790 1685
rect 824 1651 858 1685
rect 892 1651 926 1685
rect 960 1651 994 1685
rect 1028 1651 1062 1685
rect 1096 1651 1130 1685
rect 1164 1651 1198 1685
rect 1232 1651 1266 1685
rect 1300 1651 1334 1685
rect 1368 1651 1402 1685
rect 1436 1651 1470 1685
rect 1504 1651 1574 1685
rect 574 1640 1574 1651
rect 574 1529 1574 1540
rect 574 1495 586 1529
rect 620 1495 654 1529
rect 688 1495 722 1529
rect 756 1495 790 1529
rect 824 1495 858 1529
rect 892 1495 926 1529
rect 960 1495 994 1529
rect 1028 1495 1062 1529
rect 1096 1495 1130 1529
rect 1164 1495 1198 1529
rect 1232 1495 1266 1529
rect 1300 1495 1334 1529
rect 1368 1495 1402 1529
rect 1436 1495 1470 1529
rect 1504 1495 1574 1529
rect 574 1487 1574 1495
rect 18086 2727 19086 2738
rect 18086 2693 18156 2727
rect 18190 2693 18224 2727
rect 18258 2693 18292 2727
rect 18326 2693 18360 2727
rect 18394 2693 18428 2727
rect 18462 2693 18496 2727
rect 18530 2693 18564 2727
rect 18598 2693 18632 2727
rect 18666 2693 18700 2727
rect 18734 2693 18768 2727
rect 18802 2693 18836 2727
rect 18870 2693 18904 2727
rect 18938 2693 18972 2727
rect 19006 2693 19040 2727
rect 19074 2693 19086 2727
rect 18086 2685 19086 2693
rect 574 1279 1574 1287
rect 574 1245 586 1279
rect 620 1245 654 1279
rect 688 1245 722 1279
rect 756 1245 790 1279
rect 824 1245 858 1279
rect 892 1245 926 1279
rect 960 1245 994 1279
rect 1028 1245 1062 1279
rect 1096 1245 1130 1279
rect 1164 1245 1198 1279
rect 1232 1245 1266 1279
rect 1300 1245 1334 1279
rect 1368 1245 1402 1279
rect 1436 1245 1470 1279
rect 1504 1245 1574 1279
rect 574 1234 1574 1245
rect 574 1123 1574 1134
rect 574 1089 586 1123
rect 620 1089 654 1123
rect 688 1089 722 1123
rect 756 1089 790 1123
rect 824 1089 858 1123
rect 892 1089 926 1123
rect 960 1089 994 1123
rect 1028 1089 1062 1123
rect 1096 1089 1130 1123
rect 1164 1089 1198 1123
rect 1232 1089 1266 1123
rect 1300 1089 1334 1123
rect 1368 1089 1402 1123
rect 1436 1089 1470 1123
rect 1504 1089 1574 1123
rect 574 1078 1574 1089
rect 574 967 1574 978
rect 574 933 586 967
rect 620 933 654 967
rect 688 933 722 967
rect 756 933 790 967
rect 824 933 858 967
rect 892 933 926 967
rect 960 933 994 967
rect 1028 933 1062 967
rect 1096 933 1130 967
rect 1164 933 1198 967
rect 1232 933 1266 967
rect 1300 933 1334 967
rect 1368 933 1402 967
rect 1436 933 1470 967
rect 1504 933 1574 967
rect 574 922 1574 933
rect 574 811 1574 822
rect 574 777 586 811
rect 620 777 654 811
rect 688 777 722 811
rect 756 777 790 811
rect 824 777 858 811
rect 892 777 926 811
rect 960 777 994 811
rect 1028 777 1062 811
rect 1096 777 1130 811
rect 1164 777 1198 811
rect 1232 777 1266 811
rect 1300 777 1334 811
rect 1368 777 1402 811
rect 1436 777 1470 811
rect 1504 777 1574 811
rect 574 766 1574 777
rect 574 655 1574 666
rect 574 621 586 655
rect 620 621 654 655
rect 688 621 722 655
rect 756 621 790 655
rect 824 621 858 655
rect 892 621 926 655
rect 960 621 994 655
rect 1028 621 1062 655
rect 1096 621 1130 655
rect 1164 621 1198 655
rect 1232 621 1266 655
rect 1300 621 1334 655
rect 1368 621 1402 655
rect 1436 621 1470 655
rect 1504 621 1574 655
rect 574 610 1574 621
rect 574 499 1574 510
rect 574 465 586 499
rect 620 465 654 499
rect 688 465 722 499
rect 756 465 790 499
rect 824 465 858 499
rect 892 465 926 499
rect 960 465 994 499
rect 1028 465 1062 499
rect 1096 465 1130 499
rect 1164 465 1198 499
rect 1232 465 1266 499
rect 1300 465 1334 499
rect 1368 465 1402 499
rect 1436 465 1470 499
rect 1504 465 1574 499
rect 574 454 1574 465
rect 574 343 1574 354
rect 574 309 586 343
rect 620 309 654 343
rect 688 309 722 343
rect 756 309 790 343
rect 824 309 858 343
rect 892 309 926 343
rect 960 309 994 343
rect 1028 309 1062 343
rect 1096 309 1130 343
rect 1164 309 1198 343
rect 1232 309 1266 343
rect 1300 309 1334 343
rect 1368 309 1402 343
rect 1436 309 1470 343
rect 1504 309 1574 343
rect 574 298 1574 309
rect 574 187 1574 198
rect 574 153 586 187
rect 620 153 654 187
rect 688 153 722 187
rect 756 153 790 187
rect 824 153 858 187
rect 892 153 926 187
rect 960 153 994 187
rect 1028 153 1062 187
rect 1096 153 1130 187
rect 1164 153 1198 187
rect 1232 153 1266 187
rect 1300 153 1334 187
rect 1368 153 1402 187
rect 1436 153 1470 187
rect 1504 153 1574 187
rect 574 142 1574 153
rect 574 31 1574 42
rect 574 -3 586 31
rect 620 -3 654 31
rect 688 -3 722 31
rect 756 -3 790 31
rect 824 -3 858 31
rect 892 -3 926 31
rect 960 -3 994 31
rect 1028 -3 1062 31
rect 1096 -3 1130 31
rect 1164 -3 1198 31
rect 1232 -3 1266 31
rect 1300 -3 1334 31
rect 1368 -3 1402 31
rect 1436 -3 1470 31
rect 1504 -3 1574 31
rect 574 -14 1574 -3
rect 574 -125 1574 -114
rect 574 -159 586 -125
rect 620 -159 654 -125
rect 688 -159 722 -125
rect 756 -159 790 -125
rect 824 -159 858 -125
rect 892 -159 926 -125
rect 960 -159 994 -125
rect 1028 -159 1062 -125
rect 1096 -159 1130 -125
rect 1164 -159 1198 -125
rect 1232 -159 1266 -125
rect 1300 -159 1334 -125
rect 1368 -159 1402 -125
rect 1436 -159 1470 -125
rect 1504 -159 1574 -125
rect 574 -170 1574 -159
rect 574 -281 1574 -270
rect 574 -315 586 -281
rect 620 -315 654 -281
rect 688 -315 722 -281
rect 756 -315 790 -281
rect 824 -315 858 -281
rect 892 -315 926 -281
rect 960 -315 994 -281
rect 1028 -315 1062 -281
rect 1096 -315 1130 -281
rect 1164 -315 1198 -281
rect 1232 -315 1266 -281
rect 1300 -315 1334 -281
rect 1368 -315 1402 -281
rect 1436 -315 1470 -281
rect 1504 -315 1574 -281
rect 574 -326 1574 -315
rect 574 -437 1574 -426
rect 574 -471 586 -437
rect 620 -471 654 -437
rect 688 -471 722 -437
rect 756 -471 790 -437
rect 824 -471 858 -437
rect 892 -471 926 -437
rect 960 -471 994 -437
rect 1028 -471 1062 -437
rect 1096 -471 1130 -437
rect 1164 -471 1198 -437
rect 1232 -471 1266 -437
rect 1300 -471 1334 -437
rect 1368 -471 1402 -437
rect 1436 -471 1470 -437
rect 1504 -471 1574 -437
rect 574 -482 1574 -471
rect 574 -593 1574 -582
rect 574 -627 586 -593
rect 620 -627 654 -593
rect 688 -627 722 -593
rect 756 -627 790 -593
rect 824 -627 858 -593
rect 892 -627 926 -593
rect 960 -627 994 -593
rect 1028 -627 1062 -593
rect 1096 -627 1130 -593
rect 1164 -627 1198 -593
rect 1232 -627 1266 -593
rect 1300 -627 1334 -593
rect 1368 -627 1402 -593
rect 1436 -627 1470 -593
rect 1504 -627 1574 -593
rect 574 -638 1574 -627
rect 574 -749 1574 -738
rect 574 -783 586 -749
rect 620 -783 654 -749
rect 688 -783 722 -749
rect 756 -783 790 -749
rect 824 -783 858 -749
rect 892 -783 926 -749
rect 960 -783 994 -749
rect 1028 -783 1062 -749
rect 1096 -783 1130 -749
rect 1164 -783 1198 -749
rect 1232 -783 1266 -749
rect 1300 -783 1334 -749
rect 1368 -783 1402 -749
rect 1436 -783 1470 -749
rect 1504 -783 1574 -749
rect 574 -791 1574 -783
rect 574 -1034 1574 -1026
rect 574 -1068 586 -1034
rect 620 -1068 654 -1034
rect 688 -1068 722 -1034
rect 756 -1068 790 -1034
rect 824 -1068 858 -1034
rect 892 -1068 926 -1034
rect 960 -1068 994 -1034
rect 1028 -1068 1062 -1034
rect 1096 -1068 1130 -1034
rect 1164 -1068 1198 -1034
rect 1232 -1068 1266 -1034
rect 1300 -1068 1334 -1034
rect 1368 -1068 1402 -1034
rect 1436 -1068 1470 -1034
rect 1504 -1068 1574 -1034
rect 574 -1079 1574 -1068
rect 574 -1190 1574 -1179
rect 574 -1224 586 -1190
rect 620 -1224 654 -1190
rect 688 -1224 722 -1190
rect 756 -1224 790 -1190
rect 824 -1224 858 -1190
rect 892 -1224 926 -1190
rect 960 -1224 994 -1190
rect 1028 -1224 1062 -1190
rect 1096 -1224 1130 -1190
rect 1164 -1224 1198 -1190
rect 1232 -1224 1266 -1190
rect 1300 -1224 1334 -1190
rect 1368 -1224 1402 -1190
rect 1436 -1224 1470 -1190
rect 1504 -1224 1574 -1190
rect 574 -1235 1574 -1224
rect 574 -1346 1574 -1335
rect 574 -1380 586 -1346
rect 620 -1380 654 -1346
rect 688 -1380 722 -1346
rect 756 -1380 790 -1346
rect 824 -1380 858 -1346
rect 892 -1380 926 -1346
rect 960 -1380 994 -1346
rect 1028 -1380 1062 -1346
rect 1096 -1380 1130 -1346
rect 1164 -1380 1198 -1346
rect 1232 -1380 1266 -1346
rect 1300 -1380 1334 -1346
rect 1368 -1380 1402 -1346
rect 1436 -1380 1470 -1346
rect 1504 -1380 1574 -1346
rect 574 -1391 1574 -1380
rect 574 -1502 1574 -1491
rect 574 -1536 586 -1502
rect 620 -1536 654 -1502
rect 688 -1536 722 -1502
rect 756 -1536 790 -1502
rect 824 -1536 858 -1502
rect 892 -1536 926 -1502
rect 960 -1536 994 -1502
rect 1028 -1536 1062 -1502
rect 1096 -1536 1130 -1502
rect 1164 -1536 1198 -1502
rect 1232 -1536 1266 -1502
rect 1300 -1536 1334 -1502
rect 1368 -1536 1402 -1502
rect 1436 -1536 1470 -1502
rect 1504 -1536 1574 -1502
rect 574 -1547 1574 -1536
rect 574 -1658 1574 -1647
rect 574 -1692 586 -1658
rect 620 -1692 654 -1658
rect 688 -1692 722 -1658
rect 756 -1692 790 -1658
rect 824 -1692 858 -1658
rect 892 -1692 926 -1658
rect 960 -1692 994 -1658
rect 1028 -1692 1062 -1658
rect 1096 -1692 1130 -1658
rect 1164 -1692 1198 -1658
rect 1232 -1692 1266 -1658
rect 1300 -1692 1334 -1658
rect 1368 -1692 1402 -1658
rect 1436 -1692 1470 -1658
rect 1504 -1692 1574 -1658
rect 574 -1703 1574 -1692
rect 574 -1814 1574 -1803
rect 574 -1848 586 -1814
rect 620 -1848 654 -1814
rect 688 -1848 722 -1814
rect 756 -1848 790 -1814
rect 824 -1848 858 -1814
rect 892 -1848 926 -1814
rect 960 -1848 994 -1814
rect 1028 -1848 1062 -1814
rect 1096 -1848 1130 -1814
rect 1164 -1848 1198 -1814
rect 1232 -1848 1266 -1814
rect 1300 -1848 1334 -1814
rect 1368 -1848 1402 -1814
rect 1436 -1848 1470 -1814
rect 1504 -1848 1574 -1814
rect 574 -1859 1574 -1848
rect 574 -1970 1574 -1959
rect 574 -2004 586 -1970
rect 620 -2004 654 -1970
rect 688 -2004 722 -1970
rect 756 -2004 790 -1970
rect 824 -2004 858 -1970
rect 892 -2004 926 -1970
rect 960 -2004 994 -1970
rect 1028 -2004 1062 -1970
rect 1096 -2004 1130 -1970
rect 1164 -2004 1198 -1970
rect 1232 -2004 1266 -1970
rect 1300 -2004 1334 -1970
rect 1368 -2004 1402 -1970
rect 1436 -2004 1470 -1970
rect 1504 -2004 1574 -1970
rect 574 -2015 1574 -2004
rect 574 -2126 1574 -2115
rect 574 -2160 586 -2126
rect 620 -2160 654 -2126
rect 688 -2160 722 -2126
rect 756 -2160 790 -2126
rect 824 -2160 858 -2126
rect 892 -2160 926 -2126
rect 960 -2160 994 -2126
rect 1028 -2160 1062 -2126
rect 1096 -2160 1130 -2126
rect 1164 -2160 1198 -2126
rect 1232 -2160 1266 -2126
rect 1300 -2160 1334 -2126
rect 1368 -2160 1402 -2126
rect 1436 -2160 1470 -2126
rect 1504 -2160 1574 -2126
rect 574 -2171 1574 -2160
rect 574 -2282 1574 -2271
rect 574 -2316 586 -2282
rect 620 -2316 654 -2282
rect 688 -2316 722 -2282
rect 756 -2316 790 -2282
rect 824 -2316 858 -2282
rect 892 -2316 926 -2282
rect 960 -2316 994 -2282
rect 1028 -2316 1062 -2282
rect 1096 -2316 1130 -2282
rect 1164 -2316 1198 -2282
rect 1232 -2316 1266 -2282
rect 1300 -2316 1334 -2282
rect 1368 -2316 1402 -2282
rect 1436 -2316 1470 -2282
rect 1504 -2316 1574 -2282
rect 574 -2324 1574 -2316
rect 3015 -17112 3068 -17100
rect 3015 -17146 3023 -17112
rect 3057 -17146 3068 -17112
rect 3015 -17180 3068 -17146
rect 3015 -17214 3023 -17180
rect 3057 -17214 3068 -17180
rect 3015 -17248 3068 -17214
rect 3015 -17282 3023 -17248
rect 3057 -17282 3068 -17248
rect 3015 -17316 3068 -17282
rect 3015 -17350 3023 -17316
rect 3057 -17350 3068 -17316
rect 3015 -17384 3068 -17350
rect 3015 -17418 3023 -17384
rect 3057 -17418 3068 -17384
rect 3015 -17452 3068 -17418
rect 3015 -17486 3023 -17452
rect 3057 -17486 3068 -17452
rect 3015 -17520 3068 -17486
rect 3015 -17554 3023 -17520
rect 3057 -17554 3068 -17520
rect 3015 -17588 3068 -17554
rect 3015 -17622 3023 -17588
rect 3057 -17622 3068 -17588
rect 3015 -17700 3068 -17622
rect 3168 -17112 3224 -17100
rect 3168 -17146 3179 -17112
rect 3213 -17146 3224 -17112
rect 3168 -17180 3224 -17146
rect 3168 -17214 3179 -17180
rect 3213 -17214 3224 -17180
rect 3168 -17248 3224 -17214
rect 3168 -17282 3179 -17248
rect 3213 -17282 3224 -17248
rect 3168 -17316 3224 -17282
rect 3168 -17350 3179 -17316
rect 3213 -17350 3224 -17316
rect 3168 -17384 3224 -17350
rect 3168 -17418 3179 -17384
rect 3213 -17418 3224 -17384
rect 3168 -17452 3224 -17418
rect 3168 -17486 3179 -17452
rect 3213 -17486 3224 -17452
rect 3168 -17520 3224 -17486
rect 3168 -17554 3179 -17520
rect 3213 -17554 3224 -17520
rect 3168 -17588 3224 -17554
rect 3168 -17622 3179 -17588
rect 3213 -17622 3224 -17588
rect 3168 -17700 3224 -17622
rect 3324 -17112 3377 -17100
rect 3324 -17146 3335 -17112
rect 3369 -17146 3377 -17112
rect 3324 -17180 3377 -17146
rect 3324 -17214 3335 -17180
rect 3369 -17214 3377 -17180
rect 3324 -17248 3377 -17214
rect 3324 -17282 3335 -17248
rect 3369 -17282 3377 -17248
rect 3324 -17316 3377 -17282
rect 3324 -17350 3335 -17316
rect 3369 -17350 3377 -17316
rect 3324 -17384 3377 -17350
rect 3324 -17418 3335 -17384
rect 3369 -17418 3377 -17384
rect 3324 -17452 3377 -17418
rect 3324 -17486 3335 -17452
rect 3369 -17486 3377 -17452
rect 3324 -17520 3377 -17486
rect 3324 -17554 3335 -17520
rect 3369 -17554 3377 -17520
rect 3324 -17588 3377 -17554
rect 3324 -17622 3335 -17588
rect 3369 -17622 3377 -17588
rect 3324 -17700 3377 -17622
rect 2572 -17985 2625 -17915
rect 2572 -18019 2580 -17985
rect 2614 -18019 2625 -17985
rect 2572 -18053 2625 -18019
rect 2572 -18087 2580 -18053
rect 2614 -18087 2625 -18053
rect 2572 -18121 2625 -18087
rect 2572 -18155 2580 -18121
rect 2614 -18155 2625 -18121
rect 2572 -18189 2625 -18155
rect 2572 -18223 2580 -18189
rect 2614 -18223 2625 -18189
rect 2572 -18257 2625 -18223
rect 2572 -18291 2580 -18257
rect 2614 -18291 2625 -18257
rect 2572 -18325 2625 -18291
rect 2572 -18359 2580 -18325
rect 2614 -18359 2625 -18325
rect 2572 -18393 2625 -18359
rect 2572 -18427 2580 -18393
rect 2614 -18427 2625 -18393
rect 2572 -18461 2625 -18427
rect 2572 -18495 2580 -18461
rect 2614 -18495 2625 -18461
rect 2572 -18529 2625 -18495
rect 2572 -18563 2580 -18529
rect 2614 -18563 2625 -18529
rect 2572 -18597 2625 -18563
rect 2572 -18631 2580 -18597
rect 2614 -18631 2625 -18597
rect 2572 -18665 2625 -18631
rect 2572 -18699 2580 -18665
rect 2614 -18699 2625 -18665
rect 2572 -18733 2625 -18699
rect 2572 -18767 2580 -18733
rect 2614 -18767 2625 -18733
rect 2572 -18801 2625 -18767
rect 2572 -18835 2580 -18801
rect 2614 -18835 2625 -18801
rect 2572 -18869 2625 -18835
rect 2572 -18903 2580 -18869
rect 2614 -18903 2625 -18869
rect 2572 -18915 2625 -18903
rect 2725 -17985 2781 -17915
rect 2725 -18019 2736 -17985
rect 2770 -18019 2781 -17985
rect 2725 -18053 2781 -18019
rect 2725 -18087 2736 -18053
rect 2770 -18087 2781 -18053
rect 2725 -18121 2781 -18087
rect 2725 -18155 2736 -18121
rect 2770 -18155 2781 -18121
rect 2725 -18189 2781 -18155
rect 2725 -18223 2736 -18189
rect 2770 -18223 2781 -18189
rect 2725 -18257 2781 -18223
rect 2725 -18291 2736 -18257
rect 2770 -18291 2781 -18257
rect 2725 -18325 2781 -18291
rect 2725 -18359 2736 -18325
rect 2770 -18359 2781 -18325
rect 2725 -18393 2781 -18359
rect 2725 -18427 2736 -18393
rect 2770 -18427 2781 -18393
rect 2725 -18461 2781 -18427
rect 2725 -18495 2736 -18461
rect 2770 -18495 2781 -18461
rect 2725 -18529 2781 -18495
rect 2725 -18563 2736 -18529
rect 2770 -18563 2781 -18529
rect 2725 -18597 2781 -18563
rect 2725 -18631 2736 -18597
rect 2770 -18631 2781 -18597
rect 2725 -18665 2781 -18631
rect 2725 -18699 2736 -18665
rect 2770 -18699 2781 -18665
rect 2725 -18733 2781 -18699
rect 2725 -18767 2736 -18733
rect 2770 -18767 2781 -18733
rect 2725 -18801 2781 -18767
rect 2725 -18835 2736 -18801
rect 2770 -18835 2781 -18801
rect 2725 -18869 2781 -18835
rect 2725 -18903 2736 -18869
rect 2770 -18903 2781 -18869
rect 2725 -18915 2781 -18903
rect 2881 -17985 2934 -17915
rect 2881 -18019 2892 -17985
rect 2926 -18019 2934 -17985
rect 2881 -18053 2934 -18019
rect 2881 -18087 2892 -18053
rect 2926 -18087 2934 -18053
rect 2881 -18121 2934 -18087
rect 2881 -18155 2892 -18121
rect 2926 -18155 2934 -18121
rect 2881 -18189 2934 -18155
rect 2881 -18223 2892 -18189
rect 2926 -18223 2934 -18189
rect 2881 -18257 2934 -18223
rect 2881 -18291 2892 -18257
rect 2926 -18291 2934 -18257
rect 2881 -18325 2934 -18291
rect 2881 -18359 2892 -18325
rect 2926 -18359 2934 -18325
rect 2881 -18393 2934 -18359
rect 2881 -18427 2892 -18393
rect 2926 -18427 2934 -18393
rect 2881 -18461 2934 -18427
rect 2881 -18495 2892 -18461
rect 2926 -18495 2934 -18461
rect 2881 -18529 2934 -18495
rect 2881 -18563 2892 -18529
rect 2926 -18563 2934 -18529
rect 2881 -18597 2934 -18563
rect 2881 -18631 2892 -18597
rect 2926 -18631 2934 -18597
rect 2881 -18665 2934 -18631
rect 2881 -18699 2892 -18665
rect 2926 -18699 2934 -18665
rect 2881 -18733 2934 -18699
rect 2881 -18767 2892 -18733
rect 2926 -18767 2934 -18733
rect 2881 -18801 2934 -18767
rect 2881 -18835 2892 -18801
rect 2926 -18835 2934 -18801
rect 2881 -18869 2934 -18835
rect 2881 -18903 2892 -18869
rect 2926 -18903 2934 -18869
rect 2881 -18915 2934 -18903
<< ndiffc >>
rect 7424 1295 7458 1329
rect 7424 1227 7458 1261
rect 7424 1159 7458 1193
rect 7424 1091 7458 1125
rect 7424 1023 7458 1057
rect 7424 955 7458 989
rect 7424 887 7458 921
rect 7424 819 7458 853
rect 7424 751 7458 785
rect 7424 683 7458 717
rect 7424 615 7458 649
rect 7424 547 7458 581
rect 7424 479 7458 513
rect 7424 411 7458 445
rect 7424 343 7458 377
rect 7424 275 7458 309
rect 7424 207 7458 241
rect 7424 139 7458 173
rect 7424 71 7458 105
rect 7424 3 7458 37
rect 7510 1295 7544 1329
rect 7510 1227 7544 1261
rect 7510 1159 7544 1193
rect 7510 1091 7544 1125
rect 7510 1023 7544 1057
rect 7510 955 7544 989
rect 7510 887 7544 921
rect 7510 819 7544 853
rect 7510 751 7544 785
rect 7510 683 7544 717
rect 7510 615 7544 649
rect 7510 547 7544 581
rect 7510 479 7544 513
rect 7510 411 7544 445
rect 7510 343 7544 377
rect 7510 275 7544 309
rect 7510 207 7544 241
rect 7510 139 7544 173
rect 7510 71 7544 105
rect 7510 3 7544 37
rect 7596 1295 7630 1329
rect 7596 1227 7630 1261
rect 7596 1159 7630 1193
rect 7596 1091 7630 1125
rect 7596 1023 7630 1057
rect 7596 955 7630 989
rect 7596 887 7630 921
rect 7596 819 7630 853
rect 7596 751 7630 785
rect 7596 683 7630 717
rect 7596 615 7630 649
rect 7596 547 7630 581
rect 7596 479 7630 513
rect 7596 411 7630 445
rect 7596 343 7630 377
rect 7596 275 7630 309
rect 7596 207 7630 241
rect 7596 139 7630 173
rect 7596 71 7630 105
rect 7596 3 7630 37
rect 7682 1295 7716 1329
rect 7682 1227 7716 1261
rect 7682 1159 7716 1193
rect 7682 1091 7716 1125
rect 7682 1023 7716 1057
rect 7682 955 7716 989
rect 7682 887 7716 921
rect 7682 819 7716 853
rect 7682 751 7716 785
rect 7682 683 7716 717
rect 7682 615 7716 649
rect 7682 547 7716 581
rect 7682 479 7716 513
rect 7682 411 7716 445
rect 7682 343 7716 377
rect 7682 275 7716 309
rect 7682 207 7716 241
rect 7682 139 7716 173
rect 7682 71 7716 105
rect 7682 3 7716 37
rect 7768 1295 7802 1329
rect 7768 1227 7802 1261
rect 7768 1159 7802 1193
rect 7768 1091 7802 1125
rect 7768 1023 7802 1057
rect 7768 955 7802 989
rect 7768 887 7802 921
rect 7768 819 7802 853
rect 7768 751 7802 785
rect 7768 683 7802 717
rect 7768 615 7802 649
rect 7768 547 7802 581
rect 7768 479 7802 513
rect 7768 411 7802 445
rect 7768 343 7802 377
rect 7768 275 7802 309
rect 7768 207 7802 241
rect 7768 139 7802 173
rect 7768 71 7802 105
rect 7768 3 7802 37
rect 7854 1295 7888 1329
rect 7854 1227 7888 1261
rect 7854 1159 7888 1193
rect 7854 1091 7888 1125
rect 7854 1023 7888 1057
rect 7854 955 7888 989
rect 7854 887 7888 921
rect 7854 819 7888 853
rect 7854 751 7888 785
rect 7854 683 7888 717
rect 7854 615 7888 649
rect 7854 547 7888 581
rect 7854 479 7888 513
rect 7854 411 7888 445
rect 7854 343 7888 377
rect 7854 275 7888 309
rect 7854 207 7888 241
rect 7854 139 7888 173
rect 7854 71 7888 105
rect 7854 3 7888 37
<< pdiffc >>
rect 871 4773 905 4807
rect 1727 4773 1761 4807
rect 1983 4773 2017 4807
rect 2239 4773 2273 4807
rect 2495 4773 2529 4807
rect 2751 4773 2785 4807
rect 3007 4773 3041 4807
rect 3263 4773 3297 4807
rect 3519 4773 3553 4807
rect 3775 4773 3809 4807
rect 4031 4773 4065 4807
rect 4287 4773 4321 4807
rect 4543 4773 4577 4807
rect 4799 4773 4833 4807
rect 5055 4773 5089 4807
rect 5311 4773 5345 4807
rect 5567 4773 5601 4807
rect 5823 4773 5857 4807
rect 6079 4773 6113 4807
rect 6335 4773 6369 4807
rect 6591 4773 6625 4807
rect 6847 4773 6881 4807
rect 7703 4773 7737 4807
rect 871 4303 905 4337
rect 1727 4303 1761 4337
rect 1983 4303 2017 4337
rect 2239 4303 2273 4337
rect 2495 4303 2529 4337
rect 2751 4303 2785 4337
rect 3007 4303 3041 4337
rect 3263 4303 3297 4337
rect 3519 4303 3553 4337
rect 3775 4303 3809 4337
rect 4031 4303 4065 4337
rect 4287 4303 4321 4337
rect 4543 4303 4577 4337
rect 4799 4303 4833 4337
rect 5055 4303 5089 4337
rect 5311 4303 5345 4337
rect 5567 4303 5601 4337
rect 5823 4303 5857 4337
rect 6079 4303 6113 4337
rect 6335 4303 6369 4337
rect 6591 4303 6625 4337
rect 6847 4303 6881 4337
rect 7703 4303 7737 4337
rect 871 3763 905 3797
rect 1727 3763 1761 3797
rect 1983 3763 2017 3797
rect 2239 3763 2273 3797
rect 2495 3763 2529 3797
rect 2751 3763 2785 3797
rect 3007 3763 3041 3797
rect 3263 3763 3297 3797
rect 3519 3763 3553 3797
rect 3775 3763 3809 3797
rect 4031 3763 4065 3797
rect 4287 3763 4321 3797
rect 4543 3763 4577 3797
rect 4799 3763 4833 3797
rect 5055 3763 5089 3797
rect 5311 3763 5345 3797
rect 5567 3763 5601 3797
rect 5823 3763 5857 3797
rect 6079 3763 6113 3797
rect 6335 3763 6369 3797
rect 6591 3763 6625 3797
rect 6847 3763 6881 3797
rect 7703 3763 7737 3797
rect 871 3293 905 3327
rect 1727 3293 1761 3327
rect 1983 3293 2017 3327
rect 2239 3293 2273 3327
rect 2495 3293 2529 3327
rect 2751 3293 2785 3327
rect 3007 3293 3041 3327
rect 3263 3293 3297 3327
rect 3519 3293 3553 3327
rect 3775 3293 3809 3327
rect 4031 3293 4065 3327
rect 4287 3293 4321 3327
rect 4543 3293 4577 3327
rect 4799 3293 4833 3327
rect 5055 3293 5089 3327
rect 5311 3293 5345 3327
rect 5567 3293 5601 3327
rect 5823 3293 5857 3327
rect 6079 3293 6113 3327
rect 6335 3293 6369 3327
rect 6591 3293 6625 3327
rect 6847 3293 6881 3327
rect 7703 3293 7737 3327
<< mvndiffc >>
rect 7515 2203 7549 2237
rect 7583 2203 7617 2237
rect 7651 2203 7685 2237
rect 7719 2203 7753 2237
rect 7787 2203 7821 2237
rect 7855 2203 7889 2237
rect 7923 2203 7957 2237
rect 7991 2203 8025 2237
rect 8059 2203 8093 2237
rect 8127 2203 8161 2237
rect 8195 2203 8229 2237
rect 8263 2203 8297 2237
rect 8331 2203 8365 2237
rect 8399 2203 8433 2237
rect 2436 2103 2470 2137
rect 2504 2103 2538 2137
rect 2572 2103 2606 2137
rect 2640 2103 2674 2137
rect 2708 2103 2742 2137
rect 2776 2103 2810 2137
rect 2844 2103 2878 2137
rect 2912 2103 2946 2137
rect 2980 2103 3014 2137
rect 3048 2103 3082 2137
rect 3116 2103 3150 2137
rect 3184 2103 3218 2137
rect 3252 2103 3286 2137
rect 3320 2103 3354 2137
rect 3388 2103 3422 2137
rect 3456 2103 3490 2137
rect 3524 2103 3558 2137
rect 3592 2103 3626 2137
rect 3660 2103 3694 2137
rect 3728 2103 3762 2137
rect 3796 2103 3830 2137
rect 3864 2103 3898 2137
rect 3932 2103 3966 2137
rect 4000 2103 4034 2137
rect 4068 2103 4102 2137
rect 4136 2103 4170 2137
rect 4204 2103 4238 2137
rect 4272 2103 4306 2137
rect 4340 2103 4374 2137
rect 4712 2103 4746 2137
rect 4780 2103 4814 2137
rect 4848 2103 4882 2137
rect 4916 2103 4950 2137
rect 4984 2103 5018 2137
rect 5052 2103 5086 2137
rect 5120 2103 5154 2137
rect 5188 2103 5222 2137
rect 5256 2103 5290 2137
rect 5324 2103 5358 2137
rect 5392 2103 5426 2137
rect 5460 2103 5494 2137
rect 5528 2103 5562 2137
rect 5596 2103 5630 2137
rect 5664 2103 5698 2137
rect 5732 2103 5766 2137
rect 5800 2103 5834 2137
rect 5868 2103 5902 2137
rect 5936 2103 5970 2137
rect 6004 2103 6038 2137
rect 6072 2103 6106 2137
rect 6140 2103 6174 2137
rect 6208 2103 6242 2137
rect 6276 2103 6310 2137
rect 6344 2103 6378 2137
rect 6412 2103 6446 2137
rect 6480 2103 6514 2137
rect 6548 2103 6582 2137
rect 6616 2103 6650 2137
rect 2436 1867 2470 1901
rect 2504 1867 2538 1901
rect 2572 1867 2606 1901
rect 2640 1867 2674 1901
rect 2708 1867 2742 1901
rect 2776 1867 2810 1901
rect 2844 1867 2878 1901
rect 2912 1867 2946 1901
rect 2980 1867 3014 1901
rect 3048 1867 3082 1901
rect 3116 1867 3150 1901
rect 3184 1867 3218 1901
rect 3252 1867 3286 1901
rect 3320 1867 3354 1901
rect 3388 1867 3422 1901
rect 3456 1867 3490 1901
rect 3524 1867 3558 1901
rect 3592 1867 3626 1901
rect 3660 1867 3694 1901
rect 3728 1867 3762 1901
rect 3796 1867 3830 1901
rect 3864 1867 3898 1901
rect 3932 1867 3966 1901
rect 4000 1867 4034 1901
rect 4068 1867 4102 1901
rect 4136 1867 4170 1901
rect 4204 1867 4238 1901
rect 4272 1867 4306 1901
rect 4340 1867 4374 1901
rect 7515 2047 7549 2081
rect 7583 2047 7617 2081
rect 7651 2047 7685 2081
rect 7719 2047 7753 2081
rect 7787 2047 7821 2081
rect 7855 2047 7889 2081
rect 7923 2047 7957 2081
rect 7991 2047 8025 2081
rect 8059 2047 8093 2081
rect 8127 2047 8161 2081
rect 8195 2047 8229 2081
rect 8263 2047 8297 2081
rect 8331 2047 8365 2081
rect 8399 2047 8433 2081
rect 4712 1867 4746 1901
rect 4780 1867 4814 1901
rect 4848 1867 4882 1901
rect 4916 1867 4950 1901
rect 4984 1867 5018 1901
rect 5052 1867 5086 1901
rect 5120 1867 5154 1901
rect 5188 1867 5222 1901
rect 5256 1867 5290 1901
rect 5324 1867 5358 1901
rect 5392 1867 5426 1901
rect 5460 1867 5494 1901
rect 5528 1867 5562 1901
rect 5596 1867 5630 1901
rect 5664 1867 5698 1901
rect 5732 1867 5766 1901
rect 5800 1867 5834 1901
rect 5868 1867 5902 1901
rect 5936 1867 5970 1901
rect 6004 1867 6038 1901
rect 6072 1867 6106 1901
rect 6140 1867 6174 1901
rect 6208 1867 6242 1901
rect 6276 1867 6310 1901
rect 6344 1867 6378 1901
rect 6412 1867 6446 1901
rect 6480 1867 6514 1901
rect 6548 1867 6582 1901
rect 6616 1867 6650 1901
rect 6829 1908 6863 1942
rect 8485 1908 8519 1942
rect 2436 1631 2470 1665
rect 2504 1631 2538 1665
rect 2572 1631 2606 1665
rect 2640 1631 2674 1665
rect 2708 1631 2742 1665
rect 2776 1631 2810 1665
rect 2844 1631 2878 1665
rect 2912 1631 2946 1665
rect 2980 1631 3014 1665
rect 3048 1631 3082 1665
rect 3116 1631 3150 1665
rect 3184 1631 3218 1665
rect 3252 1631 3286 1665
rect 3320 1631 3354 1665
rect 3388 1631 3422 1665
rect 3456 1631 3490 1665
rect 3524 1631 3558 1665
rect 3592 1631 3626 1665
rect 3660 1631 3694 1665
rect 3728 1631 3762 1665
rect 3796 1631 3830 1665
rect 3864 1631 3898 1665
rect 3932 1631 3966 1665
rect 4000 1631 4034 1665
rect 4068 1631 4102 1665
rect 4136 1631 4170 1665
rect 4204 1631 4238 1665
rect 4272 1631 4306 1665
rect 4340 1631 4374 1665
rect 4712 1631 4746 1665
rect 4780 1631 4814 1665
rect 4848 1631 4882 1665
rect 4916 1631 4950 1665
rect 4984 1631 5018 1665
rect 5052 1631 5086 1665
rect 5120 1631 5154 1665
rect 5188 1631 5222 1665
rect 5256 1631 5290 1665
rect 5324 1631 5358 1665
rect 5392 1631 5426 1665
rect 5460 1631 5494 1665
rect 5528 1631 5562 1665
rect 5596 1631 5630 1665
rect 5664 1631 5698 1665
rect 5732 1631 5766 1665
rect 5800 1631 5834 1665
rect 5868 1631 5902 1665
rect 5936 1631 5970 1665
rect 6004 1631 6038 1665
rect 6072 1631 6106 1665
rect 6140 1631 6174 1665
rect 6208 1631 6242 1665
rect 6276 1631 6310 1665
rect 6344 1631 6378 1665
rect 6412 1631 6446 1665
rect 6480 1631 6514 1665
rect 6548 1631 6582 1665
rect 6616 1631 6650 1665
rect 6829 1668 6863 1702
rect 8485 1668 8519 1702
rect 10637 2676 10671 2710
rect 10634 2154 10668 2188
rect 2436 1395 2470 1429
rect 2504 1395 2538 1429
rect 2572 1395 2606 1429
rect 2640 1395 2674 1429
rect 2708 1395 2742 1429
rect 2776 1395 2810 1429
rect 2844 1395 2878 1429
rect 2912 1395 2946 1429
rect 2980 1395 3014 1429
rect 3048 1395 3082 1429
rect 3116 1395 3150 1429
rect 3184 1395 3218 1429
rect 3252 1395 3286 1429
rect 3320 1395 3354 1429
rect 3388 1395 3422 1429
rect 3456 1395 3490 1429
rect 3524 1395 3558 1429
rect 3592 1395 3626 1429
rect 3660 1395 3694 1429
rect 3728 1395 3762 1429
rect 3796 1395 3830 1429
rect 3864 1395 3898 1429
rect 3932 1395 3966 1429
rect 4000 1395 4034 1429
rect 4068 1395 4102 1429
rect 4136 1395 4170 1429
rect 4204 1395 4238 1429
rect 4272 1395 4306 1429
rect 4340 1395 4374 1429
rect 4712 1395 4746 1429
rect 4780 1395 4814 1429
rect 4848 1395 4882 1429
rect 4916 1395 4950 1429
rect 4984 1395 5018 1429
rect 5052 1395 5086 1429
rect 5120 1395 5154 1429
rect 5188 1395 5222 1429
rect 5256 1395 5290 1429
rect 5324 1395 5358 1429
rect 5392 1395 5426 1429
rect 5460 1395 5494 1429
rect 5528 1395 5562 1429
rect 5596 1395 5630 1429
rect 5664 1395 5698 1429
rect 5732 1395 5766 1429
rect 5800 1395 5834 1429
rect 5868 1395 5902 1429
rect 5936 1395 5970 1429
rect 6004 1395 6038 1429
rect 6072 1395 6106 1429
rect 6140 1395 6174 1429
rect 6208 1395 6242 1429
rect 6276 1395 6310 1429
rect 6344 1395 6378 1429
rect 6412 1395 6446 1429
rect 6480 1395 6514 1429
rect 6548 1395 6582 1429
rect 6616 1395 6650 1429
rect 2436 1159 2470 1193
rect 2504 1159 2538 1193
rect 2572 1159 2606 1193
rect 2640 1159 2674 1193
rect 2708 1159 2742 1193
rect 2776 1159 2810 1193
rect 2844 1159 2878 1193
rect 2912 1159 2946 1193
rect 2980 1159 3014 1193
rect 3048 1159 3082 1193
rect 3116 1159 3150 1193
rect 3184 1159 3218 1193
rect 3252 1159 3286 1193
rect 3320 1159 3354 1193
rect 3388 1159 3422 1193
rect 3456 1159 3490 1193
rect 3524 1159 3558 1193
rect 3592 1159 3626 1193
rect 3660 1159 3694 1193
rect 3728 1159 3762 1193
rect 3796 1159 3830 1193
rect 3864 1159 3898 1193
rect 3932 1159 3966 1193
rect 4000 1159 4034 1193
rect 4068 1159 4102 1193
rect 4136 1159 4170 1193
rect 4204 1159 4238 1193
rect 4272 1159 4306 1193
rect 4340 1159 4374 1193
rect 4712 1159 4746 1193
rect 4780 1159 4814 1193
rect 4848 1159 4882 1193
rect 4916 1159 4950 1193
rect 4984 1159 5018 1193
rect 5052 1159 5086 1193
rect 5120 1159 5154 1193
rect 5188 1159 5222 1193
rect 5256 1159 5290 1193
rect 5324 1159 5358 1193
rect 5392 1159 5426 1193
rect 5460 1159 5494 1193
rect 5528 1159 5562 1193
rect 5596 1159 5630 1193
rect 5664 1159 5698 1193
rect 5732 1159 5766 1193
rect 5800 1159 5834 1193
rect 5868 1159 5902 1193
rect 5936 1159 5970 1193
rect 6004 1159 6038 1193
rect 6072 1159 6106 1193
rect 6140 1159 6174 1193
rect 6208 1159 6242 1193
rect 6276 1159 6310 1193
rect 6344 1159 6378 1193
rect 6412 1159 6446 1193
rect 6480 1159 6514 1193
rect 6548 1159 6582 1193
rect 6616 1159 6650 1193
rect 2406 912 2440 946
rect 2406 844 2440 878
rect 2406 776 2440 810
rect 2406 708 2440 742
rect 2406 640 2440 674
rect 2406 572 2440 606
rect 2406 504 2440 538
rect 2406 436 2440 470
rect 2406 368 2440 402
rect 2406 300 2440 334
rect 2406 232 2440 266
rect 2406 164 2440 198
rect 2406 96 2440 130
rect 2406 28 2440 62
rect 2562 912 2596 946
rect 2562 844 2596 878
rect 2562 776 2596 810
rect 2562 708 2596 742
rect 2562 640 2596 674
rect 2562 572 2596 606
rect 2562 504 2596 538
rect 2562 436 2596 470
rect 2562 368 2596 402
rect 2562 300 2596 334
rect 2562 232 2596 266
rect 2562 164 2596 198
rect 2562 96 2596 130
rect 2562 28 2596 62
rect 2718 912 2752 946
rect 2718 844 2752 878
rect 2718 776 2752 810
rect 2718 708 2752 742
rect 2718 640 2752 674
rect 2718 572 2752 606
rect 2718 504 2752 538
rect 2718 436 2752 470
rect 2718 368 2752 402
rect 2718 300 2752 334
rect 2718 232 2752 266
rect 2718 164 2752 198
rect 2718 96 2752 130
rect 2718 28 2752 62
rect 2874 912 2908 946
rect 2874 844 2908 878
rect 2874 776 2908 810
rect 2874 708 2908 742
rect 2874 640 2908 674
rect 2874 572 2908 606
rect 2874 504 2908 538
rect 2874 436 2908 470
rect 2874 368 2908 402
rect 2874 300 2908 334
rect 2874 232 2908 266
rect 2874 164 2908 198
rect 2874 96 2908 130
rect 2874 28 2908 62
rect 3030 912 3064 946
rect 3030 844 3064 878
rect 3030 776 3064 810
rect 3030 708 3064 742
rect 3030 640 3064 674
rect 3030 572 3064 606
rect 3030 504 3064 538
rect 3030 436 3064 470
rect 3030 368 3064 402
rect 3030 300 3064 334
rect 3030 232 3064 266
rect 3030 164 3064 198
rect 3030 96 3064 130
rect 3030 28 3064 62
rect 3186 912 3220 946
rect 3186 844 3220 878
rect 3186 776 3220 810
rect 3186 708 3220 742
rect 3186 640 3220 674
rect 3186 572 3220 606
rect 3186 504 3220 538
rect 3186 436 3220 470
rect 3186 368 3220 402
rect 3186 300 3220 334
rect 3186 232 3220 266
rect 3186 164 3220 198
rect 3186 96 3220 130
rect 3186 28 3220 62
rect 3342 912 3376 946
rect 3342 844 3376 878
rect 3342 776 3376 810
rect 3342 708 3376 742
rect 3342 640 3376 674
rect 3342 572 3376 606
rect 3342 504 3376 538
rect 3342 436 3376 470
rect 3342 368 3376 402
rect 3342 300 3376 334
rect 3342 232 3376 266
rect 3342 164 3376 198
rect 3342 96 3376 130
rect 3342 28 3376 62
rect 3498 912 3532 946
rect 3498 844 3532 878
rect 3498 776 3532 810
rect 3498 708 3532 742
rect 3498 640 3532 674
rect 3498 572 3532 606
rect 3498 504 3532 538
rect 3498 436 3532 470
rect 3498 368 3532 402
rect 3498 300 3532 334
rect 3498 232 3532 266
rect 3498 164 3532 198
rect 3498 96 3532 130
rect 3498 28 3532 62
rect 3654 912 3688 946
rect 3654 844 3688 878
rect 3654 776 3688 810
rect 3654 708 3688 742
rect 3654 640 3688 674
rect 3654 572 3688 606
rect 3654 504 3688 538
rect 3654 436 3688 470
rect 3654 368 3688 402
rect 3654 300 3688 334
rect 3654 232 3688 266
rect 3654 164 3688 198
rect 3654 96 3688 130
rect 3654 28 3688 62
rect 3778 912 3812 946
rect 3778 844 3812 878
rect 3778 776 3812 810
rect 3778 708 3812 742
rect 3778 640 3812 674
rect 3778 572 3812 606
rect 3778 504 3812 538
rect 3778 436 3812 470
rect 3778 368 3812 402
rect 3778 300 3812 334
rect 3778 232 3812 266
rect 3778 164 3812 198
rect 3778 96 3812 130
rect 3778 28 3812 62
rect 3934 912 3968 946
rect 3934 844 3968 878
rect 3934 776 3968 810
rect 3934 708 3968 742
rect 3934 640 3968 674
rect 3934 572 3968 606
rect 3934 504 3968 538
rect 3934 436 3968 470
rect 3934 368 3968 402
rect 3934 300 3968 334
rect 3934 232 3968 266
rect 3934 164 3968 198
rect 3934 96 3968 130
rect 3934 28 3968 62
rect 4090 912 4124 946
rect 4090 844 4124 878
rect 4090 776 4124 810
rect 4090 708 4124 742
rect 4090 640 4124 674
rect 4090 572 4124 606
rect 4090 504 4124 538
rect 4090 436 4124 470
rect 4090 368 4124 402
rect 4090 300 4124 334
rect 4090 232 4124 266
rect 4090 164 4124 198
rect 4090 96 4124 130
rect 4090 28 4124 62
rect 4246 912 4280 946
rect 4246 844 4280 878
rect 4246 776 4280 810
rect 4246 708 4280 742
rect 4246 640 4280 674
rect 4246 572 4280 606
rect 4246 504 4280 538
rect 4246 436 4280 470
rect 4246 368 4280 402
rect 4246 300 4280 334
rect 4246 232 4280 266
rect 4246 164 4280 198
rect 4246 96 4280 130
rect 4246 28 4280 62
rect 4402 912 4436 946
rect 4402 844 4436 878
rect 4402 776 4436 810
rect 4402 708 4436 742
rect 4402 640 4436 674
rect 4402 572 4436 606
rect 4402 504 4436 538
rect 4402 436 4436 470
rect 4402 368 4436 402
rect 4402 300 4436 334
rect 4402 232 4436 266
rect 4402 164 4436 198
rect 4402 96 4436 130
rect 4402 28 4436 62
rect 4558 912 4592 946
rect 4558 844 4592 878
rect 4558 776 4592 810
rect 4558 708 4592 742
rect 4558 640 4592 674
rect 4558 572 4592 606
rect 4558 504 4592 538
rect 4558 436 4592 470
rect 4558 368 4592 402
rect 4558 300 4592 334
rect 4558 232 4592 266
rect 4558 164 4592 198
rect 4558 96 4592 130
rect 4558 28 4592 62
rect 4714 912 4748 946
rect 4714 844 4748 878
rect 4714 776 4748 810
rect 4714 708 4748 742
rect 4714 640 4748 674
rect 4714 572 4748 606
rect 4714 504 4748 538
rect 4714 436 4748 470
rect 4714 368 4748 402
rect 4714 300 4748 334
rect 4714 232 4748 266
rect 4714 164 4748 198
rect 4714 96 4748 130
rect 4714 28 4748 62
rect 4870 912 4904 946
rect 4870 844 4904 878
rect 4870 776 4904 810
rect 4870 708 4904 742
rect 4870 640 4904 674
rect 4870 572 4904 606
rect 4870 504 4904 538
rect 4870 436 4904 470
rect 4870 368 4904 402
rect 4870 300 4904 334
rect 4870 232 4904 266
rect 4870 164 4904 198
rect 4870 96 4904 130
rect 4870 28 4904 62
rect 5026 912 5060 946
rect 5026 844 5060 878
rect 5026 776 5060 810
rect 5026 708 5060 742
rect 5026 640 5060 674
rect 5026 572 5060 606
rect 5026 504 5060 538
rect 5026 436 5060 470
rect 5026 368 5060 402
rect 5026 300 5060 334
rect 5026 232 5060 266
rect 5026 164 5060 198
rect 5026 96 5060 130
rect 5026 28 5060 62
rect 5182 912 5216 946
rect 5182 844 5216 878
rect 5182 776 5216 810
rect 5182 708 5216 742
rect 5182 640 5216 674
rect 5182 572 5216 606
rect 5182 504 5216 538
rect 5182 436 5216 470
rect 5182 368 5216 402
rect 5182 300 5216 334
rect 5182 232 5216 266
rect 5182 164 5216 198
rect 5182 96 5216 130
rect 5182 28 5216 62
rect 5338 912 5372 946
rect 5338 844 5372 878
rect 5338 776 5372 810
rect 5338 708 5372 742
rect 5338 640 5372 674
rect 5338 572 5372 606
rect 5338 504 5372 538
rect 5338 436 5372 470
rect 5338 368 5372 402
rect 5338 300 5372 334
rect 5338 232 5372 266
rect 5338 164 5372 198
rect 5338 96 5372 130
rect 5338 28 5372 62
rect 5494 912 5528 946
rect 5494 844 5528 878
rect 5494 776 5528 810
rect 5494 708 5528 742
rect 5494 640 5528 674
rect 5494 572 5528 606
rect 5494 504 5528 538
rect 5494 436 5528 470
rect 5494 368 5528 402
rect 5494 300 5528 334
rect 5494 232 5528 266
rect 5494 164 5528 198
rect 5494 96 5528 130
rect 5494 28 5528 62
rect 5668 912 5702 946
rect 5668 844 5702 878
rect 5668 776 5702 810
rect 5668 708 5702 742
rect 5668 640 5702 674
rect 5668 572 5702 606
rect 5668 504 5702 538
rect 5668 436 5702 470
rect 5668 368 5702 402
rect 5668 300 5702 334
rect 5668 232 5702 266
rect 5668 164 5702 198
rect 5668 96 5702 130
rect 5668 28 5702 62
rect 5824 912 5858 946
rect 5824 844 5858 878
rect 5824 776 5858 810
rect 5824 708 5858 742
rect 5824 640 5858 674
rect 5824 572 5858 606
rect 5824 504 5858 538
rect 5824 436 5858 470
rect 5824 368 5858 402
rect 5824 300 5858 334
rect 5824 232 5858 266
rect 5824 164 5858 198
rect 5824 96 5858 130
rect 5824 28 5858 62
rect 5980 912 6014 946
rect 5980 844 6014 878
rect 5980 776 6014 810
rect 5980 708 6014 742
rect 5980 640 6014 674
rect 5980 572 6014 606
rect 5980 504 6014 538
rect 5980 436 6014 470
rect 5980 368 6014 402
rect 5980 300 6014 334
rect 5980 232 6014 266
rect 5980 164 6014 198
rect 5980 96 6014 130
rect 5980 28 6014 62
rect 6136 912 6170 946
rect 6136 844 6170 878
rect 6136 776 6170 810
rect 6136 708 6170 742
rect 6136 640 6170 674
rect 6136 572 6170 606
rect 6136 504 6170 538
rect 6136 436 6170 470
rect 6136 368 6170 402
rect 6136 300 6170 334
rect 6136 232 6170 266
rect 6136 164 6170 198
rect 6136 96 6170 130
rect 6136 28 6170 62
rect 6292 912 6326 946
rect 6292 844 6326 878
rect 6292 776 6326 810
rect 6292 708 6326 742
rect 6292 640 6326 674
rect 6292 572 6326 606
rect 6292 504 6326 538
rect 6292 436 6326 470
rect 6292 368 6326 402
rect 6292 300 6326 334
rect 6292 232 6326 266
rect 6292 164 6326 198
rect 6292 96 6326 130
rect 6292 28 6326 62
rect 6416 912 6450 946
rect 6416 844 6450 878
rect 6416 776 6450 810
rect 6416 708 6450 742
rect 6416 640 6450 674
rect 6416 572 6450 606
rect 6416 504 6450 538
rect 6416 436 6450 470
rect 6416 368 6450 402
rect 6416 300 6450 334
rect 6416 232 6450 266
rect 6416 164 6450 198
rect 6416 96 6450 130
rect 6416 28 6450 62
rect 6572 912 6606 946
rect 6572 844 6606 878
rect 6572 776 6606 810
rect 6572 708 6606 742
rect 6572 640 6606 674
rect 6572 572 6606 606
rect 6572 504 6606 538
rect 6572 436 6606 470
rect 6572 368 6606 402
rect 6572 300 6606 334
rect 6572 232 6606 266
rect 6572 164 6606 198
rect 6572 96 6606 130
rect 6572 28 6606 62
rect 6696 912 6730 946
rect 6696 844 6730 878
rect 6696 776 6730 810
rect 6696 708 6730 742
rect 6696 640 6730 674
rect 6696 572 6730 606
rect 6696 504 6730 538
rect 6696 436 6730 470
rect 6696 368 6730 402
rect 6696 300 6730 334
rect 6696 232 6730 266
rect 6696 164 6730 198
rect 6696 96 6730 130
rect 6696 28 6730 62
rect 6852 912 6886 946
rect 6852 844 6886 878
rect 6852 776 6886 810
rect 6852 708 6886 742
rect 6852 640 6886 674
rect 6852 572 6886 606
rect 6852 504 6886 538
rect 6852 436 6886 470
rect 6852 368 6886 402
rect 6852 300 6886 334
rect 6852 232 6886 266
rect 6852 164 6886 198
rect 6852 96 6886 130
rect 6852 28 6886 62
rect 7008 912 7042 946
rect 7008 844 7042 878
rect 7008 776 7042 810
rect 7008 708 7042 742
rect 7008 640 7042 674
rect 7008 572 7042 606
rect 7008 504 7042 538
rect 7008 436 7042 470
rect 7008 368 7042 402
rect 7008 300 7042 334
rect 7008 232 7042 266
rect 7008 164 7042 198
rect 7008 96 7042 130
rect 7008 28 7042 62
rect 13088 1035 13122 1069
rect 13156 1035 13190 1069
rect 13224 1035 13258 1069
rect 13292 1035 13326 1069
rect 13360 1035 13394 1069
rect 13428 1035 13462 1069
rect 13496 1035 13530 1069
rect 13564 1035 13598 1069
rect 13632 1035 13666 1069
rect 13700 1035 13734 1069
rect 13768 1035 13802 1069
rect 13836 1035 13870 1069
rect 13904 1035 13938 1069
rect 13972 1035 14006 1069
rect 14040 1035 14074 1069
rect 14108 1035 14142 1069
rect 14176 1035 14210 1069
rect 14244 1035 14278 1069
rect 14312 1035 14346 1069
rect 14380 1035 14414 1069
rect 14448 1035 14482 1069
rect 14516 1035 14550 1069
rect 14584 1035 14618 1069
rect 14652 1035 14686 1069
rect 14720 1035 14754 1069
rect 14788 1035 14822 1069
rect 14856 1035 14890 1069
rect 14924 1035 14958 1069
rect 14992 1035 15026 1069
rect 8284 844 8318 878
rect 8284 776 8318 810
rect 8284 708 8318 742
rect 8284 640 8318 674
rect 8284 572 8318 606
rect 8284 504 8318 538
rect 8284 436 8318 470
rect 8284 368 8318 402
rect 8284 300 8318 334
rect 8284 232 8318 266
rect 8284 164 8318 198
rect 8284 96 8318 130
rect 8284 28 8318 62
rect 8284 -40 8318 -6
rect 8440 844 8474 878
rect 8440 776 8474 810
rect 8440 708 8474 742
rect 8440 640 8474 674
rect 8440 572 8474 606
rect 8440 504 8474 538
rect 8440 436 8474 470
rect 8440 368 8474 402
rect 8440 300 8474 334
rect 8440 232 8474 266
rect 8440 164 8474 198
rect 8440 96 8474 130
rect 8440 28 8474 62
rect 8440 -40 8474 -6
rect 8596 844 8630 878
rect 8596 776 8630 810
rect 8596 708 8630 742
rect 8596 640 8630 674
rect 8596 572 8630 606
rect 8596 504 8630 538
rect 8596 436 8630 470
rect 8596 368 8630 402
rect 8596 300 8630 334
rect 8596 232 8630 266
rect 8596 164 8630 198
rect 8596 96 8630 130
rect 8596 28 8630 62
rect 8596 -40 8630 -6
rect 8752 844 8786 878
rect 8752 776 8786 810
rect 8752 708 8786 742
rect 8752 640 8786 674
rect 8752 572 8786 606
rect 8752 504 8786 538
rect 8752 436 8786 470
rect 8752 368 8786 402
rect 8752 300 8786 334
rect 8752 232 8786 266
rect 8752 164 8786 198
rect 8752 96 8786 130
rect 8752 28 8786 62
rect 8752 -40 8786 -6
rect 8908 844 8942 878
rect 8908 776 8942 810
rect 8908 708 8942 742
rect 8908 640 8942 674
rect 8908 572 8942 606
rect 8908 504 8942 538
rect 8908 436 8942 470
rect 8908 368 8942 402
rect 8908 300 8942 334
rect 8908 232 8942 266
rect 8908 164 8942 198
rect 8908 96 8942 130
rect 8908 28 8942 62
rect 8908 -40 8942 -6
rect 9064 844 9098 878
rect 9064 776 9098 810
rect 9064 708 9098 742
rect 9064 640 9098 674
rect 9064 572 9098 606
rect 9064 504 9098 538
rect 9064 436 9098 470
rect 9064 368 9098 402
rect 9064 300 9098 334
rect 9064 232 9098 266
rect 9064 164 9098 198
rect 9064 96 9098 130
rect 9064 28 9098 62
rect 9064 -40 9098 -6
rect 9220 844 9254 878
rect 9220 776 9254 810
rect 9220 708 9254 742
rect 9220 640 9254 674
rect 9220 572 9254 606
rect 9220 504 9254 538
rect 9220 436 9254 470
rect 9220 368 9254 402
rect 9220 300 9254 334
rect 9220 232 9254 266
rect 9220 164 9254 198
rect 9220 96 9254 130
rect 9220 28 9254 62
rect 9220 -40 9254 -6
rect 9376 844 9410 878
rect 9376 776 9410 810
rect 9376 708 9410 742
rect 9376 640 9410 674
rect 9376 572 9410 606
rect 9376 504 9410 538
rect 9376 436 9410 470
rect 9376 368 9410 402
rect 9376 300 9410 334
rect 9376 232 9410 266
rect 9376 164 9410 198
rect 9376 96 9410 130
rect 9376 28 9410 62
rect 9376 -40 9410 -6
rect 9532 844 9566 878
rect 9532 776 9566 810
rect 9532 708 9566 742
rect 9532 640 9566 674
rect 9532 572 9566 606
rect 9532 504 9566 538
rect 9532 436 9566 470
rect 9532 368 9566 402
rect 9532 300 9566 334
rect 9532 232 9566 266
rect 9532 164 9566 198
rect 9532 96 9566 130
rect 9532 28 9566 62
rect 9532 -40 9566 -6
rect 9688 844 9722 878
rect 9688 776 9722 810
rect 9688 708 9722 742
rect 9688 640 9722 674
rect 9688 572 9722 606
rect 9688 504 9722 538
rect 9688 436 9722 470
rect 9688 368 9722 402
rect 9688 300 9722 334
rect 9688 232 9722 266
rect 9688 164 9722 198
rect 9688 96 9722 130
rect 9688 28 9722 62
rect 9688 -40 9722 -6
rect 9844 844 9878 878
rect 9844 776 9878 810
rect 9844 708 9878 742
rect 9844 640 9878 674
rect 9844 572 9878 606
rect 9844 504 9878 538
rect 9844 436 9878 470
rect 9844 368 9878 402
rect 9844 300 9878 334
rect 9844 232 9878 266
rect 9844 164 9878 198
rect 9844 96 9878 130
rect 9844 28 9878 62
rect 9844 -40 9878 -6
rect 10000 844 10034 878
rect 10000 776 10034 810
rect 10000 708 10034 742
rect 10000 640 10034 674
rect 10000 572 10034 606
rect 10000 504 10034 538
rect 10000 436 10034 470
rect 10000 368 10034 402
rect 10000 300 10034 334
rect 10000 232 10034 266
rect 10000 164 10034 198
rect 10000 96 10034 130
rect 10000 28 10034 62
rect 10000 -40 10034 -6
rect 10156 844 10190 878
rect 10156 776 10190 810
rect 10156 708 10190 742
rect 10156 640 10190 674
rect 10156 572 10190 606
rect 10156 504 10190 538
rect 10156 436 10190 470
rect 10156 368 10190 402
rect 10156 300 10190 334
rect 10156 232 10190 266
rect 10156 164 10190 198
rect 10156 96 10190 130
rect 10156 28 10190 62
rect 10156 -40 10190 -6
rect 10312 844 10346 878
rect 10312 776 10346 810
rect 10312 708 10346 742
rect 10312 640 10346 674
rect 10312 572 10346 606
rect 10312 504 10346 538
rect 10312 436 10346 470
rect 10312 368 10346 402
rect 10312 300 10346 334
rect 10312 232 10346 266
rect 10312 164 10346 198
rect 10312 96 10346 130
rect 10312 28 10346 62
rect 10312 -40 10346 -6
rect 10468 844 10502 878
rect 10468 776 10502 810
rect 10468 708 10502 742
rect 10468 640 10502 674
rect 10468 572 10502 606
rect 10468 504 10502 538
rect 10468 436 10502 470
rect 10468 368 10502 402
rect 10468 300 10502 334
rect 10468 232 10502 266
rect 10468 164 10502 198
rect 10468 96 10502 130
rect 10468 28 10502 62
rect 10468 -40 10502 -6
rect 10737 844 10771 878
rect 10737 776 10771 810
rect 10737 708 10771 742
rect 10737 640 10771 674
rect 10737 572 10771 606
rect 10737 504 10771 538
rect 10737 436 10771 470
rect 10737 368 10771 402
rect 10737 300 10771 334
rect 10737 232 10771 266
rect 10737 164 10771 198
rect 10737 96 10771 130
rect 10737 28 10771 62
rect 10737 -40 10771 -6
rect 11193 844 11227 878
rect 11193 776 11227 810
rect 11193 708 11227 742
rect 11193 640 11227 674
rect 11193 572 11227 606
rect 11193 504 11227 538
rect 11193 436 11227 470
rect 11193 368 11227 402
rect 11193 300 11227 334
rect 11193 232 11227 266
rect 11193 164 11227 198
rect 11193 96 11227 130
rect 11193 28 11227 62
rect 11193 -40 11227 -6
rect 11649 844 11683 878
rect 11649 776 11683 810
rect 11649 708 11683 742
rect 11649 640 11683 674
rect 11649 572 11683 606
rect 11649 504 11683 538
rect 11649 436 11683 470
rect 11649 368 11683 402
rect 11649 300 11683 334
rect 11649 232 11683 266
rect 11649 164 11683 198
rect 11649 96 11683 130
rect 11649 28 11683 62
rect 11649 -40 11683 -6
rect 12105 844 12139 878
rect 12105 776 12139 810
rect 12105 708 12139 742
rect 12105 640 12139 674
rect 12105 572 12139 606
rect 12105 504 12139 538
rect 12105 436 12139 470
rect 12105 368 12139 402
rect 12105 300 12139 334
rect 12105 232 12139 266
rect 12105 164 12139 198
rect 12105 96 12139 130
rect 12105 28 12139 62
rect 12105 -40 12139 -6
rect 12561 844 12595 878
rect 12561 776 12595 810
rect 12783 896 12817 930
rect 12783 828 12817 862
rect 12783 760 12817 794
rect 12959 896 12993 930
rect 12959 828 12993 862
rect 12959 760 12993 794
rect 13088 799 13122 833
rect 13156 799 13190 833
rect 13224 799 13258 833
rect 13292 799 13326 833
rect 13360 799 13394 833
rect 13428 799 13462 833
rect 13496 799 13530 833
rect 13564 799 13598 833
rect 13632 799 13666 833
rect 13700 799 13734 833
rect 13768 799 13802 833
rect 13836 799 13870 833
rect 13904 799 13938 833
rect 13972 799 14006 833
rect 14040 799 14074 833
rect 14108 799 14142 833
rect 14176 799 14210 833
rect 14244 799 14278 833
rect 14312 799 14346 833
rect 14380 799 14414 833
rect 14448 799 14482 833
rect 14516 799 14550 833
rect 14584 799 14618 833
rect 14652 799 14686 833
rect 14720 799 14754 833
rect 14788 799 14822 833
rect 14856 799 14890 833
rect 14924 799 14958 833
rect 14992 799 15026 833
rect 15223 988 15257 1022
rect 15223 920 15257 954
rect 15223 852 15257 886
rect 15459 988 15493 1022
rect 15459 920 15493 954
rect 15459 852 15493 886
rect 15695 988 15729 1022
rect 15695 920 15729 954
rect 15695 852 15729 886
rect 15931 988 15965 1022
rect 15931 920 15965 954
rect 15931 852 15965 886
rect 16167 988 16201 1022
rect 16167 920 16201 954
rect 16167 852 16201 886
rect 12561 708 12595 742
rect 12561 640 12595 674
rect 12561 572 12595 606
rect 12561 504 12595 538
rect 12561 436 12595 470
rect 12561 368 12595 402
rect 12561 300 12595 334
rect 12561 232 12595 266
rect 12561 164 12595 198
rect 12561 96 12595 130
rect 12561 28 12595 62
rect 12561 -40 12595 -6
rect 13088 563 13122 597
rect 13156 563 13190 597
rect 13224 563 13258 597
rect 13292 563 13326 597
rect 13360 563 13394 597
rect 13428 563 13462 597
rect 13496 563 13530 597
rect 13564 563 13598 597
rect 13632 563 13666 597
rect 13700 563 13734 597
rect 13768 563 13802 597
rect 13836 563 13870 597
rect 13904 563 13938 597
rect 13972 563 14006 597
rect 14040 563 14074 597
rect 14108 563 14142 597
rect 14176 563 14210 597
rect 14244 563 14278 597
rect 14312 563 14346 597
rect 14380 563 14414 597
rect 14448 563 14482 597
rect 14516 563 14550 597
rect 14584 563 14618 597
rect 14652 563 14686 597
rect 14720 563 14754 597
rect 14788 563 14822 597
rect 14856 563 14890 597
rect 14924 563 14958 597
rect 14992 563 15026 597
rect 15223 627 15257 661
rect 15223 559 15257 593
rect 15223 491 15257 525
rect 15459 627 15493 661
rect 15459 559 15493 593
rect 15459 491 15493 525
rect 15695 627 15729 661
rect 15695 559 15729 593
rect 15695 491 15729 525
rect 15931 627 15965 661
rect 15931 559 15965 593
rect 15931 491 15965 525
rect 16167 627 16201 661
rect 16167 559 16201 593
rect 16167 491 16201 525
rect 13088 327 13122 361
rect 13156 327 13190 361
rect 13224 327 13258 361
rect 13292 327 13326 361
rect 13360 327 13394 361
rect 13428 327 13462 361
rect 13496 327 13530 361
rect 13564 327 13598 361
rect 13632 327 13666 361
rect 13700 327 13734 361
rect 13768 327 13802 361
rect 13836 327 13870 361
rect 13904 327 13938 361
rect 13972 327 14006 361
rect 14040 327 14074 361
rect 14108 327 14142 361
rect 14176 327 14210 361
rect 14244 327 14278 361
rect 14312 327 14346 361
rect 14380 327 14414 361
rect 14448 327 14482 361
rect 14516 327 14550 361
rect 14584 327 14618 361
rect 14652 327 14686 361
rect 14720 327 14754 361
rect 14788 327 14822 361
rect 14856 327 14890 361
rect 14924 327 14958 361
rect 14992 327 15026 361
rect 15223 248 15257 282
rect 15223 180 15257 214
rect 13088 91 13122 125
rect 13156 91 13190 125
rect 13224 91 13258 125
rect 13292 91 13326 125
rect 13360 91 13394 125
rect 13428 91 13462 125
rect 13496 91 13530 125
rect 13564 91 13598 125
rect 13632 91 13666 125
rect 13700 91 13734 125
rect 13768 91 13802 125
rect 13836 91 13870 125
rect 13904 91 13938 125
rect 13972 91 14006 125
rect 14040 91 14074 125
rect 14108 91 14142 125
rect 14176 91 14210 125
rect 14244 91 14278 125
rect 14312 91 14346 125
rect 14380 91 14414 125
rect 14448 91 14482 125
rect 14516 91 14550 125
rect 14584 91 14618 125
rect 14652 91 14686 125
rect 14720 91 14754 125
rect 14788 91 14822 125
rect 14856 91 14890 125
rect 14924 91 14958 125
rect 14992 91 15026 125
rect 15223 112 15257 146
rect 15459 248 15493 282
rect 15459 180 15493 214
rect 15459 112 15493 146
rect 15695 248 15729 282
rect 18414 304 18448 338
rect 18482 304 18516 338
rect 18550 304 18584 338
rect 15695 180 15729 214
rect 15695 112 15729 146
rect 15884 73 15918 107
rect 15884 5 15918 39
rect 15884 -63 15918 -29
rect 15884 -131 15918 -97
rect 15884 -199 15918 -165
rect 15884 -267 15918 -233
rect 15884 -335 15918 -301
rect 15884 -403 15918 -369
rect 15884 -471 15918 -437
rect 15884 -539 15918 -505
rect 15884 -607 15918 -573
rect 15884 -675 15918 -641
rect 15884 -743 15918 -709
rect 15884 -811 15918 -777
rect 16040 73 16074 107
rect 16040 5 16074 39
rect 16040 -63 16074 -29
rect 16040 -131 16074 -97
rect 16040 -199 16074 -165
rect 16040 -267 16074 -233
rect 16040 -335 16074 -301
rect 16040 -403 16074 -369
rect 16040 -471 16074 -437
rect 16040 -539 16074 -505
rect 16040 -607 16074 -573
rect 16040 -675 16074 -641
rect 16040 -743 16074 -709
rect 16040 -811 16074 -777
rect 16196 73 16230 107
rect 16196 5 16230 39
rect 16196 -63 16230 -29
rect 16196 -131 16230 -97
rect 16196 -199 16230 -165
rect 16196 -267 16230 -233
rect 16196 -335 16230 -301
rect 16196 -403 16230 -369
rect 16196 -471 16230 -437
rect 16196 -539 16230 -505
rect 16196 -607 16230 -573
rect 16196 -675 16230 -641
rect 16196 -743 16230 -709
rect 16196 -811 16230 -777
rect 18414 148 18448 182
rect 18482 148 18516 182
rect 18550 148 18584 182
rect 18414 -8 18448 26
rect 18482 -8 18516 26
rect 18550 -8 18584 26
rect 548 -10956 582 -10922
rect 896 -3403 930 -3369
rect 2624 -9696 2658 -9662
rect 2624 -9764 2658 -9730
rect 2624 -9832 2658 -9798
rect 2624 -9900 2658 -9866
rect 2624 -9968 2658 -9934
rect 2624 -10036 2658 -10002
rect 2624 -10104 2658 -10070
rect 2624 -10172 2658 -10138
rect 2780 -9696 2814 -9662
rect 2780 -9764 2814 -9730
rect 2780 -9832 2814 -9798
rect 2780 -9900 2814 -9866
rect 2780 -9968 2814 -9934
rect 2780 -10036 2814 -10002
rect 2780 -10104 2814 -10070
rect 2780 -10172 2814 -10138
rect 2936 -9696 2970 -9662
rect 2936 -9764 2970 -9730
rect 2936 -9832 2970 -9798
rect 2936 -9900 2970 -9866
rect 2936 -9968 2970 -9934
rect 2936 -10036 2970 -10002
rect 2936 -10104 2970 -10070
rect 2936 -10172 2970 -10138
<< mvpdiffc >>
rect 8714 4758 8748 4792
rect 8714 4690 8748 4724
rect 8714 4622 8748 4656
rect 8714 4554 8748 4588
rect 8714 4486 8748 4520
rect 8714 4418 8748 4452
rect 8714 4350 8748 4384
rect 8714 4282 8748 4316
rect 8714 4214 8748 4248
rect 8714 4146 8748 4180
rect 8714 4078 8748 4112
rect 8714 4010 8748 4044
rect 8714 3942 8748 3976
rect 8714 3874 8748 3908
rect 8870 4758 8904 4792
rect 8870 4690 8904 4724
rect 8870 4622 8904 4656
rect 8870 4554 8904 4588
rect 8870 4486 8904 4520
rect 8870 4418 8904 4452
rect 8870 4350 8904 4384
rect 8870 4282 8904 4316
rect 8870 4214 8904 4248
rect 8870 4146 8904 4180
rect 8870 4078 8904 4112
rect 8870 4010 8904 4044
rect 8870 3942 8904 3976
rect 8870 3874 8904 3908
rect 9026 4758 9060 4792
rect 9026 4690 9060 4724
rect 9026 4622 9060 4656
rect 9026 4554 9060 4588
rect 9026 4486 9060 4520
rect 9026 4418 9060 4452
rect 9026 4350 9060 4384
rect 9026 4282 9060 4316
rect 9026 4214 9060 4248
rect 9026 4146 9060 4180
rect 9026 4078 9060 4112
rect 9026 4010 9060 4044
rect 9026 3942 9060 3976
rect 9026 3874 9060 3908
rect 9182 4758 9216 4792
rect 9182 4690 9216 4724
rect 9182 4622 9216 4656
rect 9182 4554 9216 4588
rect 9182 4486 9216 4520
rect 9182 4418 9216 4452
rect 9182 4350 9216 4384
rect 9182 4282 9216 4316
rect 9182 4214 9216 4248
rect 9182 4146 9216 4180
rect 9182 4078 9216 4112
rect 9182 4010 9216 4044
rect 9182 3942 9216 3976
rect 9182 3874 9216 3908
rect 9338 4758 9372 4792
rect 9338 4690 9372 4724
rect 9338 4622 9372 4656
rect 9338 4554 9372 4588
rect 9338 4486 9372 4520
rect 9338 4418 9372 4452
rect 9338 4350 9372 4384
rect 9338 4282 9372 4316
rect 9338 4214 9372 4248
rect 9338 4146 9372 4180
rect 9338 4078 9372 4112
rect 9338 4010 9372 4044
rect 9338 3942 9372 3976
rect 9338 3874 9372 3908
rect 9462 4758 9496 4792
rect 9462 4690 9496 4724
rect 9462 4622 9496 4656
rect 9462 4554 9496 4588
rect 9462 4486 9496 4520
rect 9462 4418 9496 4452
rect 9462 4350 9496 4384
rect 9462 4282 9496 4316
rect 9462 4214 9496 4248
rect 9462 4146 9496 4180
rect 9462 4078 9496 4112
rect 9462 4010 9496 4044
rect 9462 3942 9496 3976
rect 9462 3874 9496 3908
rect 9618 4758 9652 4792
rect 9618 4690 9652 4724
rect 9618 4622 9652 4656
rect 9618 4554 9652 4588
rect 9618 4486 9652 4520
rect 9618 4418 9652 4452
rect 9618 4350 9652 4384
rect 9618 4282 9652 4316
rect 9618 4214 9652 4248
rect 9618 4146 9652 4180
rect 9618 4078 9652 4112
rect 9618 4010 9652 4044
rect 9618 3942 9652 3976
rect 9618 3874 9652 3908
rect 9742 4758 9776 4792
rect 9742 4690 9776 4724
rect 9742 4622 9776 4656
rect 9742 4554 9776 4588
rect 9742 4486 9776 4520
rect 9742 4418 9776 4452
rect 9742 4350 9776 4384
rect 9742 4282 9776 4316
rect 9742 4214 9776 4248
rect 9742 4146 9776 4180
rect 9742 4078 9776 4112
rect 9742 4010 9776 4044
rect 9742 3942 9776 3976
rect 9742 3874 9776 3908
rect 9898 4758 9932 4792
rect 9898 4690 9932 4724
rect 9898 4622 9932 4656
rect 9898 4554 9932 4588
rect 9898 4486 9932 4520
rect 9898 4418 9932 4452
rect 9898 4350 9932 4384
rect 9898 4282 9932 4316
rect 9898 4214 9932 4248
rect 9898 4146 9932 4180
rect 9898 4078 9932 4112
rect 9898 4010 9932 4044
rect 9898 3942 9932 3976
rect 9898 3874 9932 3908
rect 10054 4758 10088 4792
rect 10054 4690 10088 4724
rect 10054 4622 10088 4656
rect 10054 4554 10088 4588
rect 10054 4486 10088 4520
rect 10054 4418 10088 4452
rect 10054 4350 10088 4384
rect 10054 4282 10088 4316
rect 10054 4214 10088 4248
rect 10054 4146 10088 4180
rect 10054 4078 10088 4112
rect 10054 4010 10088 4044
rect 10054 3942 10088 3976
rect 10054 3874 10088 3908
rect 10331 4758 10365 4792
rect 10331 4690 10365 4724
rect 10331 4622 10365 4656
rect 10331 4554 10365 4588
rect 10331 4486 10365 4520
rect 10331 4418 10365 4452
rect 10331 4350 10365 4384
rect 10331 4282 10365 4316
rect 10331 4214 10365 4248
rect 10331 4146 10365 4180
rect 10331 4078 10365 4112
rect 10331 4010 10365 4044
rect 10331 3942 10365 3976
rect 10331 3874 10365 3908
rect 10487 4758 10521 4792
rect 10487 4690 10521 4724
rect 10487 4622 10521 4656
rect 10487 4554 10521 4588
rect 10487 4486 10521 4520
rect 10487 4418 10521 4452
rect 10487 4350 10521 4384
rect 10487 4282 10521 4316
rect 10487 4214 10521 4248
rect 10487 4146 10521 4180
rect 10487 4078 10521 4112
rect 10487 4010 10521 4044
rect 10487 3942 10521 3976
rect 10487 3874 10521 3908
rect 10643 4758 10677 4792
rect 10643 4690 10677 4724
rect 10643 4622 10677 4656
rect 10643 4554 10677 4588
rect 10643 4486 10677 4520
rect 10643 4418 10677 4452
rect 10643 4350 10677 4384
rect 10643 4282 10677 4316
rect 10643 4214 10677 4248
rect 10643 4146 10677 4180
rect 10643 4078 10677 4112
rect 10643 4010 10677 4044
rect 10643 3942 10677 3976
rect 10643 3874 10677 3908
rect 10799 4758 10833 4792
rect 10799 4690 10833 4724
rect 10799 4622 10833 4656
rect 10799 4554 10833 4588
rect 10799 4486 10833 4520
rect 10799 4418 10833 4452
rect 10799 4350 10833 4384
rect 10799 4282 10833 4316
rect 10799 4214 10833 4248
rect 10799 4146 10833 4180
rect 10799 4078 10833 4112
rect 10799 4010 10833 4044
rect 10799 3942 10833 3976
rect 10799 3874 10833 3908
rect 10955 4758 10989 4792
rect 10955 4690 10989 4724
rect 10955 4622 10989 4656
rect 10955 4554 10989 4588
rect 10955 4486 10989 4520
rect 10955 4418 10989 4452
rect 10955 4350 10989 4384
rect 10955 4282 10989 4316
rect 10955 4214 10989 4248
rect 10955 4146 10989 4180
rect 10955 4078 10989 4112
rect 10955 4010 10989 4044
rect 10955 3942 10989 3976
rect 10955 3874 10989 3908
rect 11111 4758 11145 4792
rect 11111 4690 11145 4724
rect 11111 4622 11145 4656
rect 11111 4554 11145 4588
rect 11111 4486 11145 4520
rect 11111 4418 11145 4452
rect 11111 4350 11145 4384
rect 11111 4282 11145 4316
rect 11111 4214 11145 4248
rect 11111 4146 11145 4180
rect 11111 4078 11145 4112
rect 11111 4010 11145 4044
rect 11111 3942 11145 3976
rect 11111 3874 11145 3908
rect 8905 3475 8939 3509
rect 8973 3475 9007 3509
rect 9041 3475 9075 3509
rect 9109 3475 9143 3509
rect 9177 3475 9211 3509
rect 9245 3475 9279 3509
rect 9313 3475 9347 3509
rect 9381 3475 9415 3509
rect 9449 3475 9483 3509
rect 9517 3475 9551 3509
rect 9585 3475 9619 3509
rect 9653 3475 9687 3509
rect 9721 3475 9755 3509
rect 9789 3475 9823 3509
rect 10579 3489 10613 3523
rect 10835 3489 10869 3523
rect 8905 3319 8939 3353
rect 8973 3319 9007 3353
rect 9041 3319 9075 3353
rect 9109 3319 9143 3353
rect 9177 3319 9211 3353
rect 9245 3319 9279 3353
rect 9313 3319 9347 3353
rect 9381 3319 9415 3353
rect 9449 3319 9483 3353
rect 9517 3319 9551 3353
rect 9585 3319 9619 3353
rect 9653 3319 9687 3353
rect 9721 3319 9755 3353
rect 9789 3319 9823 3353
rect 10222 3336 10256 3370
rect 10290 3336 10324 3370
rect 10358 3336 10392 3370
rect 10426 3336 10460 3370
rect 10494 3336 10528 3370
rect 10562 3336 10596 3370
rect 10630 3336 10664 3370
rect 10698 3336 10732 3370
rect 10766 3336 10800 3370
rect 10834 3336 10868 3370
rect 10902 3336 10936 3370
rect 10970 3336 11004 3370
rect 11038 3336 11072 3370
rect 11106 3336 11140 3370
rect 8905 3163 8939 3197
rect 8973 3163 9007 3197
rect 9041 3163 9075 3197
rect 9109 3163 9143 3197
rect 9177 3163 9211 3197
rect 9245 3163 9279 3197
rect 9313 3163 9347 3197
rect 9381 3163 9415 3197
rect 9449 3163 9483 3197
rect 9517 3163 9551 3197
rect 9585 3163 9619 3197
rect 9653 3163 9687 3197
rect 9721 3163 9755 3197
rect 9789 3163 9823 3197
rect 10222 3180 10256 3214
rect 10290 3180 10324 3214
rect 10358 3180 10392 3214
rect 10426 3180 10460 3214
rect 10494 3180 10528 3214
rect 10562 3180 10596 3214
rect 10630 3180 10664 3214
rect 10698 3180 10732 3214
rect 10766 3180 10800 3214
rect 10834 3180 10868 3214
rect 10902 3180 10936 3214
rect 10970 3180 11004 3214
rect 11038 3180 11072 3214
rect 11106 3180 11140 3214
rect 17049 3195 17083 3229
rect 17117 3195 17151 3229
rect 17185 3195 17219 3229
rect 17253 3195 17287 3229
rect 17321 3195 17355 3229
rect 17389 3195 17423 3229
rect 17457 3195 17491 3229
rect 17525 3195 17559 3229
rect 17049 3019 17083 3053
rect 17117 3019 17151 3053
rect 17185 3019 17219 3053
rect 17253 3019 17287 3053
rect 17321 3019 17355 3053
rect 17389 3019 17423 3053
rect 17457 3019 17491 3053
rect 17525 3019 17559 3053
rect 17798 3182 17832 3216
rect 17798 3114 17832 3148
rect 17798 3046 17832 3080
rect 17954 3182 17988 3216
rect 17954 3114 17988 3148
rect 17954 3046 17988 3080
rect 18110 3182 18144 3216
rect 18110 3114 18144 3148
rect 18110 3046 18144 3080
rect 18282 3182 18316 3216
rect 18282 3114 18316 3148
rect 18282 3046 18316 3080
rect 18438 3182 18472 3216
rect 18438 3114 18472 3148
rect 18438 3046 18472 3080
rect 18594 3182 18628 3216
rect 18594 3114 18628 3148
rect 18594 3046 18628 3080
rect 18744 3182 18778 3216
rect 18744 3114 18778 3148
rect 18744 3046 18778 3080
rect 18900 3182 18934 3216
rect 18900 3114 18934 3148
rect 18900 3046 18934 3080
rect 19056 3182 19090 3216
rect 19056 3114 19090 3148
rect 19056 3046 19090 3080
rect 18156 2849 18190 2883
rect 18224 2849 18258 2883
rect 18292 2849 18326 2883
rect 18360 2849 18394 2883
rect 18428 2849 18462 2883
rect 18496 2849 18530 2883
rect 18564 2849 18598 2883
rect 18632 2849 18666 2883
rect 18700 2849 18734 2883
rect 18768 2849 18802 2883
rect 18836 2849 18870 2883
rect 18904 2849 18938 2883
rect 18972 2849 19006 2883
rect 19040 2849 19074 2883
rect 586 2399 620 2433
rect 654 2399 688 2433
rect 722 2399 756 2433
rect 790 2399 824 2433
rect 858 2399 892 2433
rect 926 2399 960 2433
rect 994 2399 1028 2433
rect 1062 2399 1096 2433
rect 1130 2399 1164 2433
rect 1198 2399 1232 2433
rect 1266 2399 1300 2433
rect 1334 2399 1368 2433
rect 1402 2399 1436 2433
rect 1470 2399 1504 2433
rect 586 2243 620 2277
rect 654 2243 688 2277
rect 722 2243 756 2277
rect 790 2243 824 2277
rect 858 2243 892 2277
rect 926 2243 960 2277
rect 994 2243 1028 2277
rect 1062 2243 1096 2277
rect 1130 2243 1164 2277
rect 1198 2243 1232 2277
rect 1266 2243 1300 2277
rect 1334 2243 1368 2277
rect 1402 2243 1436 2277
rect 1470 2243 1504 2277
rect 586 1807 620 1841
rect 654 1807 688 1841
rect 722 1807 756 1841
rect 790 1807 824 1841
rect 858 1807 892 1841
rect 926 1807 960 1841
rect 994 1807 1028 1841
rect 1062 1807 1096 1841
rect 1130 1807 1164 1841
rect 1198 1807 1232 1841
rect 1266 1807 1300 1841
rect 1334 1807 1368 1841
rect 1402 1807 1436 1841
rect 1470 1807 1504 1841
rect 586 1651 620 1685
rect 654 1651 688 1685
rect 722 1651 756 1685
rect 790 1651 824 1685
rect 858 1651 892 1685
rect 926 1651 960 1685
rect 994 1651 1028 1685
rect 1062 1651 1096 1685
rect 1130 1651 1164 1685
rect 1198 1651 1232 1685
rect 1266 1651 1300 1685
rect 1334 1651 1368 1685
rect 1402 1651 1436 1685
rect 1470 1651 1504 1685
rect 586 1495 620 1529
rect 654 1495 688 1529
rect 722 1495 756 1529
rect 790 1495 824 1529
rect 858 1495 892 1529
rect 926 1495 960 1529
rect 994 1495 1028 1529
rect 1062 1495 1096 1529
rect 1130 1495 1164 1529
rect 1198 1495 1232 1529
rect 1266 1495 1300 1529
rect 1334 1495 1368 1529
rect 1402 1495 1436 1529
rect 1470 1495 1504 1529
rect 18156 2693 18190 2727
rect 18224 2693 18258 2727
rect 18292 2693 18326 2727
rect 18360 2693 18394 2727
rect 18428 2693 18462 2727
rect 18496 2693 18530 2727
rect 18564 2693 18598 2727
rect 18632 2693 18666 2727
rect 18700 2693 18734 2727
rect 18768 2693 18802 2727
rect 18836 2693 18870 2727
rect 18904 2693 18938 2727
rect 18972 2693 19006 2727
rect 19040 2693 19074 2727
rect 586 1245 620 1279
rect 654 1245 688 1279
rect 722 1245 756 1279
rect 790 1245 824 1279
rect 858 1245 892 1279
rect 926 1245 960 1279
rect 994 1245 1028 1279
rect 1062 1245 1096 1279
rect 1130 1245 1164 1279
rect 1198 1245 1232 1279
rect 1266 1245 1300 1279
rect 1334 1245 1368 1279
rect 1402 1245 1436 1279
rect 1470 1245 1504 1279
rect 586 1089 620 1123
rect 654 1089 688 1123
rect 722 1089 756 1123
rect 790 1089 824 1123
rect 858 1089 892 1123
rect 926 1089 960 1123
rect 994 1089 1028 1123
rect 1062 1089 1096 1123
rect 1130 1089 1164 1123
rect 1198 1089 1232 1123
rect 1266 1089 1300 1123
rect 1334 1089 1368 1123
rect 1402 1089 1436 1123
rect 1470 1089 1504 1123
rect 586 933 620 967
rect 654 933 688 967
rect 722 933 756 967
rect 790 933 824 967
rect 858 933 892 967
rect 926 933 960 967
rect 994 933 1028 967
rect 1062 933 1096 967
rect 1130 933 1164 967
rect 1198 933 1232 967
rect 1266 933 1300 967
rect 1334 933 1368 967
rect 1402 933 1436 967
rect 1470 933 1504 967
rect 586 777 620 811
rect 654 777 688 811
rect 722 777 756 811
rect 790 777 824 811
rect 858 777 892 811
rect 926 777 960 811
rect 994 777 1028 811
rect 1062 777 1096 811
rect 1130 777 1164 811
rect 1198 777 1232 811
rect 1266 777 1300 811
rect 1334 777 1368 811
rect 1402 777 1436 811
rect 1470 777 1504 811
rect 586 621 620 655
rect 654 621 688 655
rect 722 621 756 655
rect 790 621 824 655
rect 858 621 892 655
rect 926 621 960 655
rect 994 621 1028 655
rect 1062 621 1096 655
rect 1130 621 1164 655
rect 1198 621 1232 655
rect 1266 621 1300 655
rect 1334 621 1368 655
rect 1402 621 1436 655
rect 1470 621 1504 655
rect 586 465 620 499
rect 654 465 688 499
rect 722 465 756 499
rect 790 465 824 499
rect 858 465 892 499
rect 926 465 960 499
rect 994 465 1028 499
rect 1062 465 1096 499
rect 1130 465 1164 499
rect 1198 465 1232 499
rect 1266 465 1300 499
rect 1334 465 1368 499
rect 1402 465 1436 499
rect 1470 465 1504 499
rect 586 309 620 343
rect 654 309 688 343
rect 722 309 756 343
rect 790 309 824 343
rect 858 309 892 343
rect 926 309 960 343
rect 994 309 1028 343
rect 1062 309 1096 343
rect 1130 309 1164 343
rect 1198 309 1232 343
rect 1266 309 1300 343
rect 1334 309 1368 343
rect 1402 309 1436 343
rect 1470 309 1504 343
rect 586 153 620 187
rect 654 153 688 187
rect 722 153 756 187
rect 790 153 824 187
rect 858 153 892 187
rect 926 153 960 187
rect 994 153 1028 187
rect 1062 153 1096 187
rect 1130 153 1164 187
rect 1198 153 1232 187
rect 1266 153 1300 187
rect 1334 153 1368 187
rect 1402 153 1436 187
rect 1470 153 1504 187
rect 586 -3 620 31
rect 654 -3 688 31
rect 722 -3 756 31
rect 790 -3 824 31
rect 858 -3 892 31
rect 926 -3 960 31
rect 994 -3 1028 31
rect 1062 -3 1096 31
rect 1130 -3 1164 31
rect 1198 -3 1232 31
rect 1266 -3 1300 31
rect 1334 -3 1368 31
rect 1402 -3 1436 31
rect 1470 -3 1504 31
rect 586 -159 620 -125
rect 654 -159 688 -125
rect 722 -159 756 -125
rect 790 -159 824 -125
rect 858 -159 892 -125
rect 926 -159 960 -125
rect 994 -159 1028 -125
rect 1062 -159 1096 -125
rect 1130 -159 1164 -125
rect 1198 -159 1232 -125
rect 1266 -159 1300 -125
rect 1334 -159 1368 -125
rect 1402 -159 1436 -125
rect 1470 -159 1504 -125
rect 586 -315 620 -281
rect 654 -315 688 -281
rect 722 -315 756 -281
rect 790 -315 824 -281
rect 858 -315 892 -281
rect 926 -315 960 -281
rect 994 -315 1028 -281
rect 1062 -315 1096 -281
rect 1130 -315 1164 -281
rect 1198 -315 1232 -281
rect 1266 -315 1300 -281
rect 1334 -315 1368 -281
rect 1402 -315 1436 -281
rect 1470 -315 1504 -281
rect 586 -471 620 -437
rect 654 -471 688 -437
rect 722 -471 756 -437
rect 790 -471 824 -437
rect 858 -471 892 -437
rect 926 -471 960 -437
rect 994 -471 1028 -437
rect 1062 -471 1096 -437
rect 1130 -471 1164 -437
rect 1198 -471 1232 -437
rect 1266 -471 1300 -437
rect 1334 -471 1368 -437
rect 1402 -471 1436 -437
rect 1470 -471 1504 -437
rect 586 -627 620 -593
rect 654 -627 688 -593
rect 722 -627 756 -593
rect 790 -627 824 -593
rect 858 -627 892 -593
rect 926 -627 960 -593
rect 994 -627 1028 -593
rect 1062 -627 1096 -593
rect 1130 -627 1164 -593
rect 1198 -627 1232 -593
rect 1266 -627 1300 -593
rect 1334 -627 1368 -593
rect 1402 -627 1436 -593
rect 1470 -627 1504 -593
rect 586 -783 620 -749
rect 654 -783 688 -749
rect 722 -783 756 -749
rect 790 -783 824 -749
rect 858 -783 892 -749
rect 926 -783 960 -749
rect 994 -783 1028 -749
rect 1062 -783 1096 -749
rect 1130 -783 1164 -749
rect 1198 -783 1232 -749
rect 1266 -783 1300 -749
rect 1334 -783 1368 -749
rect 1402 -783 1436 -749
rect 1470 -783 1504 -749
rect 586 -1068 620 -1034
rect 654 -1068 688 -1034
rect 722 -1068 756 -1034
rect 790 -1068 824 -1034
rect 858 -1068 892 -1034
rect 926 -1068 960 -1034
rect 994 -1068 1028 -1034
rect 1062 -1068 1096 -1034
rect 1130 -1068 1164 -1034
rect 1198 -1068 1232 -1034
rect 1266 -1068 1300 -1034
rect 1334 -1068 1368 -1034
rect 1402 -1068 1436 -1034
rect 1470 -1068 1504 -1034
rect 586 -1224 620 -1190
rect 654 -1224 688 -1190
rect 722 -1224 756 -1190
rect 790 -1224 824 -1190
rect 858 -1224 892 -1190
rect 926 -1224 960 -1190
rect 994 -1224 1028 -1190
rect 1062 -1224 1096 -1190
rect 1130 -1224 1164 -1190
rect 1198 -1224 1232 -1190
rect 1266 -1224 1300 -1190
rect 1334 -1224 1368 -1190
rect 1402 -1224 1436 -1190
rect 1470 -1224 1504 -1190
rect 586 -1380 620 -1346
rect 654 -1380 688 -1346
rect 722 -1380 756 -1346
rect 790 -1380 824 -1346
rect 858 -1380 892 -1346
rect 926 -1380 960 -1346
rect 994 -1380 1028 -1346
rect 1062 -1380 1096 -1346
rect 1130 -1380 1164 -1346
rect 1198 -1380 1232 -1346
rect 1266 -1380 1300 -1346
rect 1334 -1380 1368 -1346
rect 1402 -1380 1436 -1346
rect 1470 -1380 1504 -1346
rect 586 -1536 620 -1502
rect 654 -1536 688 -1502
rect 722 -1536 756 -1502
rect 790 -1536 824 -1502
rect 858 -1536 892 -1502
rect 926 -1536 960 -1502
rect 994 -1536 1028 -1502
rect 1062 -1536 1096 -1502
rect 1130 -1536 1164 -1502
rect 1198 -1536 1232 -1502
rect 1266 -1536 1300 -1502
rect 1334 -1536 1368 -1502
rect 1402 -1536 1436 -1502
rect 1470 -1536 1504 -1502
rect 586 -1692 620 -1658
rect 654 -1692 688 -1658
rect 722 -1692 756 -1658
rect 790 -1692 824 -1658
rect 858 -1692 892 -1658
rect 926 -1692 960 -1658
rect 994 -1692 1028 -1658
rect 1062 -1692 1096 -1658
rect 1130 -1692 1164 -1658
rect 1198 -1692 1232 -1658
rect 1266 -1692 1300 -1658
rect 1334 -1692 1368 -1658
rect 1402 -1692 1436 -1658
rect 1470 -1692 1504 -1658
rect 586 -1848 620 -1814
rect 654 -1848 688 -1814
rect 722 -1848 756 -1814
rect 790 -1848 824 -1814
rect 858 -1848 892 -1814
rect 926 -1848 960 -1814
rect 994 -1848 1028 -1814
rect 1062 -1848 1096 -1814
rect 1130 -1848 1164 -1814
rect 1198 -1848 1232 -1814
rect 1266 -1848 1300 -1814
rect 1334 -1848 1368 -1814
rect 1402 -1848 1436 -1814
rect 1470 -1848 1504 -1814
rect 586 -2004 620 -1970
rect 654 -2004 688 -1970
rect 722 -2004 756 -1970
rect 790 -2004 824 -1970
rect 858 -2004 892 -1970
rect 926 -2004 960 -1970
rect 994 -2004 1028 -1970
rect 1062 -2004 1096 -1970
rect 1130 -2004 1164 -1970
rect 1198 -2004 1232 -1970
rect 1266 -2004 1300 -1970
rect 1334 -2004 1368 -1970
rect 1402 -2004 1436 -1970
rect 1470 -2004 1504 -1970
rect 586 -2160 620 -2126
rect 654 -2160 688 -2126
rect 722 -2160 756 -2126
rect 790 -2160 824 -2126
rect 858 -2160 892 -2126
rect 926 -2160 960 -2126
rect 994 -2160 1028 -2126
rect 1062 -2160 1096 -2126
rect 1130 -2160 1164 -2126
rect 1198 -2160 1232 -2126
rect 1266 -2160 1300 -2126
rect 1334 -2160 1368 -2126
rect 1402 -2160 1436 -2126
rect 1470 -2160 1504 -2126
rect 586 -2316 620 -2282
rect 654 -2316 688 -2282
rect 722 -2316 756 -2282
rect 790 -2316 824 -2282
rect 858 -2316 892 -2282
rect 926 -2316 960 -2282
rect 994 -2316 1028 -2282
rect 1062 -2316 1096 -2282
rect 1130 -2316 1164 -2282
rect 1198 -2316 1232 -2282
rect 1266 -2316 1300 -2282
rect 1334 -2316 1368 -2282
rect 1402 -2316 1436 -2282
rect 1470 -2316 1504 -2282
rect 3023 -17146 3057 -17112
rect 3023 -17214 3057 -17180
rect 3023 -17282 3057 -17248
rect 3023 -17350 3057 -17316
rect 3023 -17418 3057 -17384
rect 3023 -17486 3057 -17452
rect 3023 -17554 3057 -17520
rect 3023 -17622 3057 -17588
rect 3179 -17146 3213 -17112
rect 3179 -17214 3213 -17180
rect 3179 -17282 3213 -17248
rect 3179 -17350 3213 -17316
rect 3179 -17418 3213 -17384
rect 3179 -17486 3213 -17452
rect 3179 -17554 3213 -17520
rect 3179 -17622 3213 -17588
rect 3335 -17146 3369 -17112
rect 3335 -17214 3369 -17180
rect 3335 -17282 3369 -17248
rect 3335 -17350 3369 -17316
rect 3335 -17418 3369 -17384
rect 3335 -17486 3369 -17452
rect 3335 -17554 3369 -17520
rect 3335 -17622 3369 -17588
rect 2580 -18019 2614 -17985
rect 2580 -18087 2614 -18053
rect 2580 -18155 2614 -18121
rect 2580 -18223 2614 -18189
rect 2580 -18291 2614 -18257
rect 2580 -18359 2614 -18325
rect 2580 -18427 2614 -18393
rect 2580 -18495 2614 -18461
rect 2580 -18563 2614 -18529
rect 2580 -18631 2614 -18597
rect 2580 -18699 2614 -18665
rect 2580 -18767 2614 -18733
rect 2580 -18835 2614 -18801
rect 2580 -18903 2614 -18869
rect 2736 -18019 2770 -17985
rect 2736 -18087 2770 -18053
rect 2736 -18155 2770 -18121
rect 2736 -18223 2770 -18189
rect 2736 -18291 2770 -18257
rect 2736 -18359 2770 -18325
rect 2736 -18427 2770 -18393
rect 2736 -18495 2770 -18461
rect 2736 -18563 2770 -18529
rect 2736 -18631 2770 -18597
rect 2736 -18699 2770 -18665
rect 2736 -18767 2770 -18733
rect 2736 -18835 2770 -18801
rect 2736 -18903 2770 -18869
rect 2892 -18019 2926 -17985
rect 2892 -18087 2926 -18053
rect 2892 -18155 2926 -18121
rect 2892 -18223 2926 -18189
rect 2892 -18291 2926 -18257
rect 2892 -18359 2926 -18325
rect 2892 -18427 2926 -18393
rect 2892 -18495 2926 -18461
rect 2892 -18563 2926 -18529
rect 2892 -18631 2926 -18597
rect 2892 -18699 2926 -18665
rect 2892 -18767 2926 -18733
rect 2892 -18835 2926 -18801
rect 2892 -18903 2926 -18869
<< psubdiff >>
rect 20252 1428 20286 1452
rect 20252 1310 20286 1394
rect 20252 1252 20286 1276
<< nsubdiff >>
rect 522 4937 590 4971
rect 624 4937 658 4971
rect 692 4937 726 4971
rect 760 4937 794 4971
rect 828 4937 862 4971
rect 896 4937 930 4971
rect 964 4937 998 4971
rect 1032 4937 1066 4971
rect 1100 4937 1134 4971
rect 1168 4937 1202 4971
rect 1236 4937 1270 4971
rect 1304 4937 1338 4971
rect 1372 4937 1406 4971
rect 1440 4937 1474 4971
rect 1508 4937 1542 4971
rect 1576 4937 1610 4971
rect 1644 4937 1678 4971
rect 1712 4937 1746 4971
rect 1780 4937 1814 4971
rect 1848 4937 1882 4971
rect 1916 4937 1950 4971
rect 1984 4937 2018 4971
rect 2052 4937 2086 4971
rect 2120 4937 2154 4971
rect 2188 4937 2222 4971
rect 2256 4937 2290 4971
rect 2324 4937 2358 4971
rect 2392 4937 2426 4971
rect 2460 4937 2494 4971
rect 2528 4937 2562 4971
rect 2596 4937 2630 4971
rect 2664 4937 2698 4971
rect 2732 4937 2766 4971
rect 2800 4937 2834 4971
rect 2868 4937 2902 4971
rect 2936 4937 2970 4971
rect 3004 4937 3038 4971
rect 3072 4937 3106 4971
rect 3140 4937 3174 4971
rect 3208 4937 3242 4971
rect 3276 4937 3310 4971
rect 3344 4937 3378 4971
rect 3412 4937 3446 4971
rect 3480 4937 3514 4971
rect 3548 4937 3582 4971
rect 3616 4937 3650 4971
rect 3684 4937 3718 4971
rect 3752 4937 3786 4971
rect 3820 4937 3854 4971
rect 3888 4937 3922 4971
rect 3956 4937 3990 4971
rect 4024 4937 4058 4971
rect 4092 4937 4126 4971
rect 4160 4937 4194 4971
rect 4228 4937 4262 4971
rect 4296 4937 4330 4971
rect 4364 4937 4398 4971
rect 4432 4937 4466 4971
rect 4500 4937 4534 4971
rect 4568 4937 4602 4971
rect 4636 4937 4670 4971
rect 4704 4937 4738 4971
rect 4772 4937 4806 4971
rect 4840 4937 4874 4971
rect 4908 4937 4942 4971
rect 4976 4937 5010 4971
rect 5044 4937 5078 4971
rect 5112 4937 5146 4971
rect 5180 4937 5214 4971
rect 5248 4937 5282 4971
rect 5316 4937 5350 4971
rect 5384 4937 5418 4971
rect 5452 4937 5486 4971
rect 5520 4937 5554 4971
rect 5588 4937 5622 4971
rect 5656 4937 5690 4971
rect 5724 4937 5758 4971
rect 5792 4937 5826 4971
rect 5860 4937 5894 4971
rect 5928 4937 5962 4971
rect 5996 4937 6030 4971
rect 6064 4937 6098 4971
rect 6132 4937 6166 4971
rect 6200 4937 6234 4971
rect 6268 4937 6302 4971
rect 6336 4937 6370 4971
rect 6404 4937 6438 4971
rect 6472 4937 6506 4971
rect 6540 4937 6574 4971
rect 6608 4937 6642 4971
rect 6676 4937 6710 4971
rect 6744 4937 6778 4971
rect 6812 4937 6846 4971
rect 6880 4937 6914 4971
rect 6948 4937 6982 4971
rect 7016 4937 7050 4971
rect 7084 4937 7118 4971
rect 7152 4937 7186 4971
rect 7220 4937 7254 4971
rect 7288 4937 7322 4971
rect 7356 4937 7390 4971
rect 7424 4937 7458 4971
rect 7492 4937 7526 4971
rect 7560 4937 7594 4971
rect 7628 4937 7662 4971
rect 7696 4937 7730 4971
rect 7764 4937 7872 4971
rect 522 4896 713 4937
rect 556 4862 713 4896
rect 522 4861 713 4862
rect 522 4828 593 4861
rect 556 4827 593 4828
rect 627 4827 679 4861
rect 7838 4903 7872 4937
rect 556 4794 713 4827
rect 7838 4835 7872 4869
rect 522 4791 713 4794
rect 522 4760 593 4791
rect 556 4757 593 4760
rect 627 4757 679 4791
rect 556 4726 713 4757
rect 522 4721 713 4726
rect 522 4692 593 4721
rect 556 4687 593 4692
rect 627 4687 679 4721
rect 7838 4767 7872 4801
rect 556 4658 713 4687
rect 522 4651 713 4658
rect 522 4624 593 4651
rect 556 4617 593 4624
rect 627 4617 679 4651
rect 556 4590 713 4617
rect 7838 4699 7872 4733
rect 7838 4631 7872 4665
rect 522 4581 713 4590
rect 522 4556 593 4581
rect 556 4547 593 4556
rect 627 4547 679 4581
rect 556 4522 713 4547
rect 522 4511 713 4522
rect 522 4488 593 4511
rect 556 4477 593 4488
rect 627 4477 679 4511
rect 7838 4563 7872 4597
rect 556 4454 713 4477
rect 522 4441 713 4454
rect 522 4420 593 4441
rect 556 4407 593 4420
rect 627 4407 679 4441
rect 556 4386 713 4407
rect 7838 4495 7872 4529
rect 7838 4427 7872 4461
rect 522 4371 713 4386
rect 522 4352 593 4371
rect 556 4337 593 4352
rect 627 4337 679 4371
rect 556 4318 713 4337
rect 522 4301 713 4318
rect 522 4284 593 4301
rect 556 4267 593 4284
rect 627 4267 679 4301
rect 7838 4359 7872 4393
rect 7838 4291 7872 4325
rect 556 4250 713 4267
rect 522 4231 713 4250
rect 522 4216 593 4231
rect 556 4197 593 4216
rect 627 4197 679 4231
rect 556 4182 713 4197
rect 522 4161 713 4182
rect 522 4148 593 4161
rect 556 4127 593 4148
rect 627 4127 679 4161
rect 556 4114 713 4127
rect 522 4090 713 4114
rect 522 4080 593 4090
rect 556 4056 593 4080
rect 627 4056 679 4090
rect 556 4046 713 4056
rect 522 4019 713 4046
rect 522 4012 593 4019
rect 556 3985 593 4012
rect 627 3985 679 4019
rect 556 3978 713 3985
rect 522 3948 713 3978
rect 522 3944 593 3948
rect 556 3914 593 3944
rect 627 3914 679 3948
rect 556 3910 713 3914
rect 522 3877 713 3910
rect 522 3876 593 3877
rect 556 3843 593 3876
rect 627 3843 679 3877
rect 556 3842 713 3843
rect 522 3808 713 3842
rect 7838 4223 7872 4257
rect 7838 4155 7872 4189
rect 7838 4087 7872 4121
rect 7838 4019 7872 4053
rect 7838 3951 7872 3985
rect 7838 3883 7872 3917
rect 7838 3815 7872 3849
rect 556 3806 713 3808
rect 556 3774 593 3806
rect 522 3772 593 3774
rect 627 3772 679 3806
rect 522 3740 713 3772
rect 556 3735 713 3740
rect 556 3706 593 3735
rect 522 3701 593 3706
rect 627 3701 679 3735
rect 522 3672 713 3701
rect 556 3664 713 3672
rect 556 3638 593 3664
rect 522 3630 593 3638
rect 627 3630 679 3664
rect 522 3604 713 3630
rect 556 3593 713 3604
rect 7838 3674 7872 3781
rect 7838 3606 7872 3640
rect 556 3570 593 3593
rect 522 3559 593 3570
rect 627 3559 679 3593
rect 522 3536 713 3559
rect 556 3522 713 3536
rect 556 3502 593 3522
rect 522 3488 593 3502
rect 627 3488 679 3522
rect 7838 3538 7872 3572
rect 522 3468 713 3488
rect 556 3451 713 3468
rect 556 3434 593 3451
rect 522 3417 593 3434
rect 627 3417 679 3451
rect 522 3400 713 3417
rect 556 3380 713 3400
rect 7838 3470 7872 3504
rect 7838 3402 7872 3436
rect 556 3366 593 3380
rect 522 3346 593 3366
rect 627 3346 679 3380
rect 522 3332 713 3346
rect 556 3309 713 3332
rect 556 3298 593 3309
rect 522 3275 593 3298
rect 627 3275 679 3309
rect 7838 3334 7872 3368
rect 522 3264 713 3275
rect 556 3238 713 3264
rect 7838 3266 7872 3300
rect 556 3230 593 3238
rect 522 3204 593 3230
rect 627 3204 679 3238
rect 522 3196 713 3204
rect 556 3162 713 3196
rect 522 3128 713 3162
rect 7838 3198 7872 3232
rect 7838 3128 7872 3164
rect 522 3094 630 3128
rect 664 3094 698 3128
rect 732 3094 766 3128
rect 800 3094 834 3128
rect 868 3094 902 3128
rect 936 3094 970 3128
rect 1004 3094 1038 3128
rect 1072 3094 1106 3128
rect 1140 3094 1174 3128
rect 1208 3094 1242 3128
rect 1276 3094 1310 3128
rect 1344 3094 1378 3128
rect 1412 3094 1446 3128
rect 1480 3094 1514 3128
rect 1548 3094 1582 3128
rect 1616 3094 1650 3128
rect 1684 3094 1718 3128
rect 1752 3094 1786 3128
rect 1820 3094 1854 3128
rect 1888 3094 1922 3128
rect 1956 3094 1990 3128
rect 2024 3094 2058 3128
rect 2092 3094 2126 3128
rect 2160 3094 2194 3128
rect 2228 3094 2262 3128
rect 2296 3094 2330 3128
rect 2364 3094 2398 3128
rect 2432 3094 2466 3128
rect 2500 3094 2534 3128
rect 2568 3094 2602 3128
rect 2636 3094 2670 3128
rect 2704 3094 2738 3128
rect 2772 3094 2806 3128
rect 2840 3094 2874 3128
rect 2908 3094 2942 3128
rect 2976 3094 3010 3128
rect 3044 3094 3078 3128
rect 3112 3094 3146 3128
rect 3180 3094 3214 3128
rect 3248 3094 3282 3128
rect 3316 3094 3350 3128
rect 3384 3094 3418 3128
rect 3452 3094 3486 3128
rect 3520 3094 3554 3128
rect 3588 3094 3622 3128
rect 3656 3094 3690 3128
rect 3724 3094 3758 3128
rect 3792 3094 3826 3128
rect 3860 3094 3894 3128
rect 3928 3094 3962 3128
rect 3996 3094 4030 3128
rect 4064 3094 4098 3128
rect 4132 3094 4166 3128
rect 4200 3094 4234 3128
rect 4268 3094 4302 3128
rect 4336 3094 4370 3128
rect 4404 3094 4438 3128
rect 4472 3094 4506 3128
rect 4540 3094 4574 3128
rect 4608 3094 4642 3128
rect 4676 3094 4710 3128
rect 4744 3094 4778 3128
rect 4812 3094 4846 3128
rect 4880 3094 4914 3128
rect 4948 3094 4982 3128
rect 5016 3094 5050 3128
rect 5084 3094 5118 3128
rect 5152 3094 5186 3128
rect 5220 3094 5254 3128
rect 5288 3094 5322 3128
rect 5356 3094 5390 3128
rect 5424 3094 5458 3128
rect 5492 3094 5526 3128
rect 5560 3094 5594 3128
rect 5628 3094 5662 3128
rect 5696 3094 5730 3128
rect 5764 3094 5798 3128
rect 5832 3094 5866 3128
rect 5900 3094 5934 3128
rect 5968 3094 6002 3128
rect 6036 3094 6070 3128
rect 6104 3094 6138 3128
rect 6172 3094 6206 3128
rect 6240 3094 6274 3128
rect 6308 3094 6342 3128
rect 6376 3094 6410 3128
rect 6444 3094 6478 3128
rect 6512 3094 6546 3128
rect 6580 3094 6614 3128
rect 6648 3094 6682 3128
rect 6716 3094 6750 3128
rect 6784 3094 6818 3128
rect 6852 3094 6886 3128
rect 6920 3094 6954 3128
rect 6988 3094 7022 3128
rect 7056 3094 7090 3128
rect 7124 3094 7158 3128
rect 7192 3094 7226 3128
rect 7260 3094 7294 3128
rect 7328 3094 7362 3128
rect 7396 3094 7430 3128
rect 7464 3094 7498 3128
rect 7532 3094 7566 3128
rect 7600 3094 7634 3128
rect 7668 3094 7702 3128
rect 7736 3094 7770 3128
rect 7804 3094 7872 3128
<< mvpsubdiff >>
rect 11552 3598 11576 3632
rect 11610 3598 11645 3632
rect 11679 3598 11714 3632
rect 11748 3598 11783 3632
rect 11817 3598 11852 3632
rect 11886 3598 11921 3632
rect 11955 3598 11990 3632
rect 12024 3598 12059 3632
rect 12093 3598 12128 3632
rect 12162 3598 12197 3632
rect 12231 3598 12266 3632
rect 12300 3598 12335 3632
rect 12369 3598 12404 3632
rect 12438 3598 12473 3632
rect 12507 3598 12542 3632
rect 12576 3598 12611 3632
rect 12645 3598 12680 3632
rect 12714 3598 12749 3632
rect 12783 3598 12818 3632
rect 12852 3598 12887 3632
rect 12921 3598 12956 3632
rect 12990 3598 13025 3632
rect 13059 3598 13094 3632
rect 13128 3598 13163 3632
rect 13197 3598 13232 3632
rect 13266 3598 13301 3632
rect 13335 3598 13370 3632
rect 13404 3598 13439 3632
rect 13473 3598 13508 3632
rect 13542 3598 13577 3632
rect 13611 3598 13646 3632
rect 13680 3598 13715 3632
rect 13749 3598 13784 3632
rect 13818 3598 13853 3632
rect 13887 3598 13922 3632
rect 13956 3598 13991 3632
rect 14025 3598 14059 3632
rect 14093 3598 14127 3632
rect 14161 3598 14195 3632
rect 14229 3598 14263 3632
rect 14297 3598 14331 3632
rect 14365 3598 14399 3632
rect 14433 3598 14467 3632
rect 14501 3598 14535 3632
rect 14569 3598 14603 3632
rect 14637 3598 14671 3632
rect 14705 3598 14739 3632
rect 14773 3598 14807 3632
rect 14841 3598 14875 3632
rect 14909 3598 14943 3632
rect 14977 3598 15011 3632
rect 15045 3598 15079 3632
rect 15113 3598 15147 3632
rect 15181 3598 15215 3632
rect 15249 3598 15283 3632
rect 15317 3598 15351 3632
rect 15385 3598 15419 3632
rect 15453 3598 15487 3632
rect 15521 3598 15555 3632
rect 15589 3598 15623 3632
rect 15657 3598 15691 3632
rect 15725 3598 15759 3632
rect 15793 3598 15827 3632
rect 15861 3598 15895 3632
rect 15929 3598 15963 3632
rect 15997 3598 16031 3632
rect 16065 3598 16099 3632
rect 16133 3598 16167 3632
rect 16201 3598 16235 3632
rect 16269 3598 16303 3632
rect 16337 3598 16371 3632
rect 16405 3598 16439 3632
rect 16473 3598 16507 3632
rect 16541 3598 16575 3632
rect 16609 3598 16643 3632
rect 16677 3598 16711 3632
rect 16745 3598 16779 3632
rect 16813 3598 16847 3632
rect 16881 3598 16915 3632
rect 16949 3598 16983 3632
rect 17017 3598 17051 3632
rect 17085 3598 17119 3632
rect 17153 3598 17187 3632
rect 17221 3598 17255 3632
rect 17289 3598 17323 3632
rect 17357 3598 17391 3632
rect 17425 3598 17459 3632
rect 17493 3598 17527 3632
rect 17561 3598 17595 3632
rect 17629 3598 17663 3632
rect 17697 3598 17731 3632
rect 17765 3598 17799 3632
rect 17833 3598 17867 3632
rect 17901 3598 17935 3632
rect 17969 3598 18003 3632
rect 18037 3598 18071 3632
rect 18105 3598 18139 3632
rect 18173 3598 18207 3632
rect 18241 3598 18275 3632
rect 18309 3598 18343 3632
rect 18377 3598 18411 3632
rect 18445 3598 18479 3632
rect 18513 3598 18547 3632
rect 18581 3598 18615 3632
rect 18649 3598 18683 3632
rect 18717 3598 18751 3632
rect 18785 3598 18819 3632
rect 18853 3598 18887 3632
rect 18921 3598 18955 3632
rect 18989 3598 19023 3632
rect 19057 3598 19091 3632
rect 19125 3598 19159 3632
rect 19193 3598 19227 3632
rect 19261 3598 19295 3632
rect 19329 3598 19363 3632
rect 19397 3598 19431 3632
rect 19465 3598 19499 3632
rect 19533 3598 19567 3632
rect 19601 3598 19635 3632
rect 19669 3598 19703 3632
rect 19737 3598 19761 3632
rect 10488 2821 10562 2855
rect 10596 2821 10630 2855
rect 10664 2821 10698 2855
rect 10732 2821 10766 2855
rect 10800 2821 10834 2855
rect 10868 2821 10902 2855
rect 10936 2821 10970 2855
rect 11004 2821 11038 2855
rect 11072 2821 11106 2855
rect 11140 2821 11174 2855
rect 11208 2821 11242 2855
rect 11276 2821 11310 2855
rect 11344 2821 11378 2855
rect 11412 2821 11446 2855
rect 11480 2821 11514 2855
rect 11548 2821 11582 2855
rect 11616 2821 11650 2855
rect 11684 2821 11718 2855
rect 11752 2821 11786 2855
rect 11820 2821 11854 2855
rect 11888 2821 11922 2855
rect 11956 2821 11990 2855
rect 12024 2821 12058 2855
rect 12092 2821 12126 2855
rect 12160 2821 12194 2855
rect 12228 2821 12262 2855
rect 12296 2821 12330 2855
rect 12364 2821 12398 2855
rect 12432 2821 12466 2855
rect 12500 2821 12534 2855
rect 12568 2821 12602 2855
rect 12636 2821 12670 2855
rect 12704 2821 12738 2855
rect 12772 2821 12806 2855
rect 12840 2821 12874 2855
rect 12908 2821 12942 2855
rect 12976 2821 13010 2855
rect 13044 2821 13078 2855
rect 13112 2821 13146 2855
rect 13180 2821 13214 2855
rect 13248 2821 13282 2855
rect 13316 2821 13350 2855
rect 13384 2821 13418 2855
rect 13452 2821 13486 2855
rect 13520 2821 13554 2855
rect 13588 2821 13622 2855
rect 13656 2821 13690 2855
rect 13724 2821 13758 2855
rect 13792 2821 13826 2855
rect 13860 2821 13894 2855
rect 13928 2821 13962 2855
rect 13996 2821 14030 2855
rect 14064 2821 14098 2855
rect 14132 2821 14166 2855
rect 14200 2821 14234 2855
rect 14268 2821 14302 2855
rect 14336 2821 14370 2855
rect 14404 2821 14438 2855
rect 14472 2821 14506 2855
rect 14540 2821 14574 2855
rect 14608 2821 14642 2855
rect 14676 2821 14710 2855
rect 14744 2821 14778 2855
rect 14812 2821 14846 2855
rect 14880 2821 14914 2855
rect 14948 2821 14982 2855
rect 15016 2821 15050 2855
rect 15084 2821 15118 2855
rect 15152 2821 15186 2855
rect 15220 2821 15254 2855
rect 15288 2821 15322 2855
rect 15356 2821 15390 2855
rect 15424 2821 15458 2855
rect 15492 2821 15526 2855
rect 15560 2821 15594 2855
rect 15628 2821 15662 2855
rect 15696 2821 15730 2855
rect 15764 2821 15798 2855
rect 15832 2821 15866 2855
rect 15900 2821 15934 2855
rect 15968 2821 16002 2855
rect 16036 2821 16070 2855
rect 16104 2821 16138 2855
rect 16172 2821 16206 2855
rect 16240 2821 16274 2855
rect 16308 2821 16342 2855
rect 16376 2821 16444 2855
rect 9716 2778 10412 2812
rect 9716 2744 9723 2778
rect 9757 2744 9795 2778
rect 9829 2744 9867 2778
rect 9901 2744 9939 2778
rect 9973 2744 10011 2778
rect 10045 2744 10083 2778
rect 10117 2744 10155 2778
rect 10189 2744 10227 2778
rect 10261 2744 10299 2778
rect 10333 2744 10371 2778
rect 10405 2744 10412 2778
rect 9716 2705 10412 2744
rect 9716 2671 9723 2705
rect 9757 2671 9795 2705
rect 9829 2671 9867 2705
rect 9901 2671 9939 2705
rect 9973 2671 10011 2705
rect 10045 2671 10083 2705
rect 10117 2671 10155 2705
rect 10189 2671 10227 2705
rect 10261 2671 10299 2705
rect 10333 2671 10371 2705
rect 10405 2671 10412 2705
rect 9716 2632 10412 2671
rect 9716 2598 9723 2632
rect 9757 2598 9795 2632
rect 9829 2598 9867 2632
rect 9901 2598 9939 2632
rect 9973 2598 10011 2632
rect 10045 2598 10083 2632
rect 10117 2598 10155 2632
rect 10189 2598 10227 2632
rect 10261 2598 10299 2632
rect 10333 2598 10371 2632
rect 10405 2598 10412 2632
rect 9716 2558 10412 2598
rect 9716 2524 9723 2558
rect 9757 2524 9795 2558
rect 9829 2524 9867 2558
rect 9901 2524 9939 2558
rect 9973 2524 10011 2558
rect 10045 2524 10083 2558
rect 10117 2524 10155 2558
rect 10189 2524 10227 2558
rect 10261 2524 10299 2558
rect 10333 2524 10371 2558
rect 10405 2524 10412 2558
rect 2428 2219 2452 2253
rect 2486 2219 2521 2253
rect 2555 2219 2590 2253
rect 2624 2219 2659 2253
rect 2693 2219 2728 2253
rect 2762 2219 2797 2253
rect 2831 2219 2866 2253
rect 2900 2219 2935 2253
rect 2969 2219 3004 2253
rect 3038 2219 3073 2253
rect 3107 2219 3142 2253
rect 3176 2219 3211 2253
rect 3245 2219 3280 2253
rect 3314 2219 3349 2253
rect 3383 2219 3418 2253
rect 3452 2219 3487 2253
rect 3521 2219 3556 2253
rect 3590 2219 3625 2253
rect 3659 2219 3694 2253
rect 3728 2219 3762 2253
rect 3796 2219 3830 2253
rect 3864 2219 3898 2253
rect 3932 2219 3966 2253
rect 4000 2219 4034 2253
rect 4068 2219 4102 2253
rect 4136 2219 4170 2253
rect 4204 2219 4238 2253
rect 4272 2219 4306 2253
rect 4340 2219 4374 2253
rect 4408 2219 4442 2253
rect 4476 2219 4510 2253
rect 4544 2219 4578 2253
rect 4612 2219 4646 2253
rect 4680 2219 4714 2253
rect 4748 2219 4782 2253
rect 4816 2219 4850 2253
rect 4884 2219 4918 2253
rect 4952 2219 4986 2253
rect 5020 2219 5054 2253
rect 5088 2219 5122 2253
rect 5156 2219 5190 2253
rect 5224 2219 5258 2253
rect 5292 2219 5326 2253
rect 5360 2219 5394 2253
rect 5428 2219 5462 2253
rect 5496 2219 5530 2253
rect 5564 2219 5598 2253
rect 5632 2219 5666 2253
rect 5700 2219 5734 2253
rect 5768 2219 5802 2253
rect 5836 2219 5870 2253
rect 5904 2219 5938 2253
rect 5972 2219 6006 2253
rect 6040 2219 6074 2253
rect 6108 2219 6142 2253
rect 6176 2219 6210 2253
rect 6244 2219 6278 2253
rect 6312 2219 6346 2253
rect 6380 2219 6414 2253
rect 6448 2219 6482 2253
rect 6516 2219 6550 2253
rect 6584 2219 6618 2253
rect 6652 2219 6686 2253
rect 6720 2219 6754 2253
rect 6788 2219 6822 2253
rect 6856 2219 6890 2253
rect 6924 2219 6958 2253
rect 6992 2219 7016 2253
rect 9716 2484 10412 2524
rect 9716 2450 9723 2484
rect 9757 2450 9795 2484
rect 9829 2450 9867 2484
rect 9901 2450 9939 2484
rect 9973 2450 10011 2484
rect 10045 2450 10083 2484
rect 10117 2450 10155 2484
rect 10189 2450 10227 2484
rect 10261 2450 10299 2484
rect 10333 2450 10371 2484
rect 10405 2450 10412 2484
rect 9716 2410 10412 2450
rect 9716 2376 9723 2410
rect 9757 2376 9795 2410
rect 9829 2376 9867 2410
rect 9901 2376 9939 2410
rect 9973 2376 10011 2410
rect 10045 2376 10083 2410
rect 10117 2376 10155 2410
rect 10189 2376 10227 2410
rect 10261 2376 10299 2410
rect 10333 2376 10371 2410
rect 10405 2376 10412 2410
rect 9716 2336 10412 2376
rect 9716 2302 9723 2336
rect 9757 2302 9795 2336
rect 9829 2302 9867 2336
rect 9901 2302 9939 2336
rect 9973 2302 10011 2336
rect 10045 2302 10083 2336
rect 10117 2302 10155 2336
rect 10189 2302 10227 2336
rect 10261 2302 10299 2336
rect 10333 2302 10371 2336
rect 10405 2302 10412 2336
rect 9716 2262 10412 2302
rect 9716 2228 9723 2262
rect 9757 2228 9795 2262
rect 9829 2228 9867 2262
rect 9901 2228 9939 2262
rect 9973 2228 10011 2262
rect 10045 2228 10083 2262
rect 10117 2228 10155 2262
rect 10189 2228 10227 2262
rect 10261 2228 10299 2262
rect 10333 2228 10371 2262
rect 10405 2228 10412 2262
rect 9716 2188 10412 2228
rect 9716 2154 9723 2188
rect 9757 2154 9795 2188
rect 9829 2154 9867 2188
rect 9901 2154 9939 2188
rect 9973 2154 10011 2188
rect 10045 2154 10083 2188
rect 10117 2154 10155 2188
rect 10189 2154 10227 2188
rect 10261 2154 10299 2188
rect 10333 2154 10371 2188
rect 10405 2154 10412 2188
rect 9716 2114 10412 2154
rect 9716 2080 9723 2114
rect 9757 2080 9795 2114
rect 9829 2080 9867 2114
rect 9901 2080 9939 2114
rect 9973 2080 10011 2114
rect 10045 2080 10083 2114
rect 10117 2080 10155 2114
rect 10189 2080 10227 2114
rect 10261 2080 10299 2114
rect 10333 2080 10371 2114
rect 10405 2080 10412 2114
rect 9716 2040 10412 2080
rect 9716 2006 9723 2040
rect 9757 2006 9795 2040
rect 9829 2006 9867 2040
rect 9901 2006 9939 2040
rect 9973 2006 10011 2040
rect 10045 2006 10083 2040
rect 10117 2006 10155 2040
rect 10189 2006 10227 2040
rect 10261 2006 10299 2040
rect 10333 2006 10371 2040
rect 10405 2006 10412 2040
rect 10488 2787 10522 2821
rect 10488 2719 10522 2753
rect 10488 2651 10522 2685
rect 10488 2583 10522 2617
rect 10488 2515 10522 2549
rect 10488 2357 10522 2481
rect 10488 2289 10522 2323
rect 16410 2727 16444 2821
rect 16410 2659 16444 2693
rect 16410 2591 16444 2625
rect 16410 2523 16444 2557
rect 16410 2455 16444 2489
rect 10488 2221 10522 2255
rect 10488 2153 10522 2187
rect 16410 2387 16444 2421
rect 16410 2319 16444 2353
rect 16410 2251 16444 2285
rect 16410 2183 16444 2217
rect 10488 2047 10522 2119
rect 16410 2115 16444 2149
rect 16410 2047 16444 2081
rect 10488 2013 10556 2047
rect 10590 2013 10624 2047
rect 10658 2013 10692 2047
rect 10726 2013 10760 2047
rect 10794 2013 10828 2047
rect 10862 2013 10896 2047
rect 10930 2013 10964 2047
rect 10998 2013 11032 2047
rect 11066 2013 11100 2047
rect 11134 2013 11168 2047
rect 11202 2013 11236 2047
rect 11270 2013 11304 2047
rect 11338 2013 11372 2047
rect 11406 2013 11440 2047
rect 11474 2013 11508 2047
rect 11542 2013 11576 2047
rect 11610 2013 11644 2047
rect 11678 2013 11712 2047
rect 11746 2013 11780 2047
rect 11814 2013 11848 2047
rect 11882 2013 11916 2047
rect 11950 2013 11984 2047
rect 12018 2013 12052 2047
rect 12086 2013 12120 2047
rect 12154 2013 12188 2047
rect 12222 2013 12256 2047
rect 12290 2013 12324 2047
rect 12358 2013 12392 2047
rect 12426 2013 12460 2047
rect 12494 2013 12528 2047
rect 12562 2013 12596 2047
rect 12630 2013 12664 2047
rect 12698 2013 12732 2047
rect 12766 2013 12800 2047
rect 12834 2013 12868 2047
rect 12902 2013 12936 2047
rect 12970 2013 13004 2047
rect 13038 2013 13072 2047
rect 13106 2013 13140 2047
rect 13174 2013 13208 2047
rect 13242 2013 13276 2047
rect 13310 2013 13344 2047
rect 13378 2013 13412 2047
rect 13446 2013 13480 2047
rect 13514 2013 13548 2047
rect 13582 2013 13616 2047
rect 13650 2013 13684 2047
rect 13718 2013 13752 2047
rect 13786 2013 13820 2047
rect 13854 2013 13888 2047
rect 13922 2013 13956 2047
rect 13990 2013 14024 2047
rect 14058 2013 14092 2047
rect 14126 2013 14160 2047
rect 14194 2013 14228 2047
rect 14262 2013 14296 2047
rect 14330 2013 14364 2047
rect 14398 2013 14432 2047
rect 14466 2013 14500 2047
rect 14534 2013 14568 2047
rect 14602 2013 14636 2047
rect 14670 2013 14704 2047
rect 14738 2013 14772 2047
rect 14806 2013 14840 2047
rect 14874 2013 14908 2047
rect 14942 2013 14976 2047
rect 15010 2013 15044 2047
rect 15078 2013 15112 2047
rect 15146 2013 15180 2047
rect 15214 2013 15248 2047
rect 15282 2013 15316 2047
rect 15350 2013 15384 2047
rect 15418 2013 15452 2047
rect 15486 2013 15520 2047
rect 15554 2013 15588 2047
rect 15622 2013 15656 2047
rect 15690 2013 15724 2047
rect 15758 2013 15792 2047
rect 15826 2013 15860 2047
rect 15894 2013 15928 2047
rect 15962 2013 15996 2047
rect 16030 2013 16064 2047
rect 16098 2013 16132 2047
rect 16166 2013 16200 2047
rect 16234 2013 16268 2047
rect 16302 2013 16336 2047
rect 16370 2013 16444 2047
rect 16563 2376 19045 2410
rect 19045 2293 19585 2294
rect 19045 2259 19079 2293
rect 19113 2259 19152 2293
rect 19186 2259 19225 2293
rect 19259 2259 19298 2293
rect 19332 2259 19371 2293
rect 19405 2259 19444 2293
rect 19478 2259 19517 2293
rect 19551 2259 19585 2293
rect 19045 2219 19585 2259
rect 19045 2185 19079 2219
rect 19113 2185 19152 2219
rect 19186 2185 19225 2219
rect 19259 2185 19298 2219
rect 19332 2185 19371 2219
rect 19405 2185 19444 2219
rect 19478 2185 19517 2219
rect 19551 2185 19585 2219
rect 19045 2145 19585 2185
rect 19045 2111 19079 2145
rect 19113 2111 19152 2145
rect 19186 2111 19225 2145
rect 19259 2111 19298 2145
rect 19332 2111 19371 2145
rect 19405 2111 19444 2145
rect 19478 2111 19517 2145
rect 19551 2111 19585 2145
rect 19045 2071 19585 2111
rect 19045 2070 19079 2071
rect 16563 2037 19079 2070
rect 19113 2037 19152 2071
rect 19186 2037 19225 2071
rect 19259 2037 19298 2071
rect 19332 2037 19371 2071
rect 19405 2037 19444 2071
rect 19478 2037 19517 2071
rect 19551 2037 19585 2071
rect 16563 2035 19585 2037
rect 9716 1966 10412 2006
rect 9716 1932 9723 1966
rect 9757 1932 9795 1966
rect 9829 1932 9867 1966
rect 9901 1932 9939 1966
rect 9973 1932 10011 1966
rect 10045 1932 10083 1966
rect 10117 1932 10155 1966
rect 10189 1932 10227 1966
rect 10261 1932 10299 1966
rect 10333 1932 10371 1966
rect 10405 1932 10412 1966
rect 9716 1898 10412 1932
rect 16597 2001 16631 2035
rect 16665 2001 16699 2035
rect 16733 2001 16767 2035
rect 16801 2001 16835 2035
rect 16869 2001 16903 2035
rect 16937 2001 16971 2035
rect 17005 2001 17039 2035
rect 17073 2001 17107 2035
rect 17141 2001 17175 2035
rect 17209 2001 17243 2035
rect 17277 2001 17311 2035
rect 17345 2001 17379 2035
rect 17413 2001 17447 2035
rect 17481 2001 17515 2035
rect 17549 2001 17583 2035
rect 17617 2001 17651 2035
rect 17685 2001 17719 2035
rect 17753 2001 17787 2035
rect 17821 2001 17855 2035
rect 17889 2001 17923 2035
rect 17957 2001 17991 2035
rect 18025 2001 18059 2035
rect 18093 2001 18127 2035
rect 18161 2001 18195 2035
rect 18229 2001 18263 2035
rect 18297 2001 18331 2035
rect 18365 2001 18399 2035
rect 18433 2001 18467 2035
rect 18501 2001 18535 2035
rect 18569 2001 18603 2035
rect 18637 2001 18671 2035
rect 18705 2001 18739 2035
rect 18773 2001 18807 2035
rect 18841 2001 18875 2035
rect 18909 2001 18943 2035
rect 18977 2001 19011 2035
rect 19045 2001 19585 2035
rect 16563 1997 19585 2001
rect 16563 1966 19079 1997
rect 19045 1963 19079 1966
rect 19113 1963 19152 1997
rect 19186 1963 19225 1997
rect 19259 1963 19298 1997
rect 19332 1963 19371 1997
rect 19405 1963 19444 1997
rect 19478 1963 19517 1997
rect 19551 1963 19585 1997
rect 19045 1932 19585 1963
rect 19011 1923 19585 1932
rect 9716 1864 9750 1898
rect 9784 1864 9819 1898
rect 9853 1864 9888 1898
rect 9922 1864 9957 1898
rect 9991 1864 10026 1898
rect 10060 1864 10095 1898
rect 10129 1864 10164 1898
rect 10198 1864 10233 1898
rect 10267 1864 10302 1898
rect 10336 1864 10371 1898
rect 10405 1864 10440 1898
rect 10474 1864 10509 1898
rect 10543 1864 10578 1898
rect 10612 1864 10647 1898
rect 10681 1864 10716 1898
rect 10750 1864 10785 1898
rect 10819 1864 10854 1898
rect 10888 1864 10923 1898
rect 10957 1864 10992 1898
rect 11026 1864 11061 1898
rect 11095 1864 11130 1898
rect 11164 1864 11199 1898
rect 11233 1864 11268 1898
rect 11302 1864 11337 1898
rect 11371 1864 11406 1898
rect 11440 1864 11475 1898
rect 11509 1864 11544 1898
rect 11578 1864 11613 1898
rect 11647 1864 11682 1898
rect 11716 1864 11751 1898
rect 11785 1864 11820 1898
rect 11854 1864 11889 1898
rect 11923 1864 11958 1898
rect 11992 1864 12027 1898
rect 12061 1864 12096 1898
rect 12130 1864 12165 1898
rect 12199 1864 12234 1898
rect 12268 1864 12303 1898
rect 12337 1864 12372 1898
rect 12406 1864 12441 1898
rect 12475 1864 12510 1898
rect 12544 1864 12579 1898
rect 12613 1864 12648 1898
rect 12682 1864 12717 1898
rect 12751 1864 12786 1898
rect 12820 1864 12855 1898
rect 12889 1864 12924 1898
rect 12958 1864 12993 1898
rect 9716 1830 12993 1864
rect 9716 1796 9750 1830
rect 9784 1796 9819 1830
rect 9853 1796 9888 1830
rect 9922 1796 9957 1830
rect 9991 1796 10026 1830
rect 10060 1796 10095 1830
rect 10129 1796 10164 1830
rect 10198 1796 10233 1830
rect 10267 1796 10302 1830
rect 10336 1796 10371 1830
rect 10405 1796 10440 1830
rect 10474 1796 10509 1830
rect 10543 1796 10578 1830
rect 10612 1796 10647 1830
rect 10681 1796 10716 1830
rect 10750 1796 10785 1830
rect 10819 1796 10854 1830
rect 10888 1796 10923 1830
rect 10957 1796 10992 1830
rect 11026 1796 11061 1830
rect 11095 1796 11130 1830
rect 11164 1796 11199 1830
rect 11233 1796 11268 1830
rect 11302 1796 11337 1830
rect 11371 1796 11406 1830
rect 11440 1796 11475 1830
rect 11509 1796 11544 1830
rect 11578 1796 11613 1830
rect 11647 1796 11682 1830
rect 11716 1796 11751 1830
rect 11785 1796 11820 1830
rect 11854 1796 11889 1830
rect 11923 1796 11958 1830
rect 11992 1796 12027 1830
rect 12061 1796 12096 1830
rect 12130 1796 12165 1830
rect 12199 1796 12234 1830
rect 12268 1796 12303 1830
rect 12337 1796 12372 1830
rect 12406 1796 12441 1830
rect 12475 1796 12510 1830
rect 12544 1796 12579 1830
rect 12613 1796 12648 1830
rect 12682 1796 12717 1830
rect 12751 1796 12786 1830
rect 12820 1796 12855 1830
rect 12889 1796 12924 1830
rect 12958 1796 12993 1830
rect 9716 1762 12993 1796
rect 9716 1728 9750 1762
rect 9784 1728 9819 1762
rect 9853 1728 9888 1762
rect 9922 1728 9957 1762
rect 9991 1728 10026 1762
rect 10060 1728 10095 1762
rect 10129 1728 10164 1762
rect 10198 1728 10233 1762
rect 10267 1728 10302 1762
rect 10336 1728 10371 1762
rect 10405 1728 10440 1762
rect 10474 1728 10509 1762
rect 10543 1728 10578 1762
rect 10612 1728 10647 1762
rect 10681 1728 10716 1762
rect 10750 1728 10785 1762
rect 10819 1728 10854 1762
rect 10888 1728 10923 1762
rect 10957 1728 10992 1762
rect 11026 1728 11061 1762
rect 11095 1728 11130 1762
rect 11164 1728 11199 1762
rect 11233 1728 11268 1762
rect 11302 1728 11337 1762
rect 11371 1728 11406 1762
rect 11440 1728 11475 1762
rect 11509 1728 11544 1762
rect 11578 1728 11613 1762
rect 11647 1728 11682 1762
rect 11716 1728 11751 1762
rect 11785 1728 11820 1762
rect 11854 1728 11889 1762
rect 11923 1728 11958 1762
rect 11992 1728 12027 1762
rect 12061 1728 12096 1762
rect 12130 1728 12165 1762
rect 12199 1728 12234 1762
rect 12268 1728 12303 1762
rect 12337 1728 12372 1762
rect 12406 1728 12441 1762
rect 12475 1728 12510 1762
rect 12544 1728 12579 1762
rect 12613 1728 12648 1762
rect 12682 1728 12717 1762
rect 12751 1728 12786 1762
rect 12820 1728 12855 1762
rect 12889 1728 12924 1762
rect 12958 1728 12993 1762
rect 9716 1694 12993 1728
rect 9716 1660 9750 1694
rect 9784 1660 9819 1694
rect 9853 1660 9888 1694
rect 9922 1660 9957 1694
rect 9991 1660 10026 1694
rect 10060 1660 10095 1694
rect 10129 1660 10164 1694
rect 10198 1660 10233 1694
rect 10267 1660 10302 1694
rect 10336 1660 10371 1694
rect 10405 1660 10440 1694
rect 10474 1660 10509 1694
rect 10543 1660 10578 1694
rect 10612 1660 10647 1694
rect 10681 1660 10716 1694
rect 10750 1660 10785 1694
rect 10819 1660 10854 1694
rect 10888 1660 10923 1694
rect 10957 1660 10992 1694
rect 11026 1660 11061 1694
rect 11095 1660 11130 1694
rect 11164 1660 11199 1694
rect 11233 1660 11268 1694
rect 11302 1660 11337 1694
rect 11371 1660 11406 1694
rect 11440 1660 11475 1694
rect 11509 1660 11544 1694
rect 11578 1660 11613 1694
rect 11647 1660 11682 1694
rect 11716 1660 11751 1694
rect 11785 1660 11820 1694
rect 11854 1660 11889 1694
rect 11923 1660 11958 1694
rect 11992 1660 12027 1694
rect 12061 1660 12096 1694
rect 12130 1660 12165 1694
rect 12199 1660 12234 1694
rect 12268 1660 12303 1694
rect 12337 1660 12372 1694
rect 12406 1660 12441 1694
rect 12475 1660 12510 1694
rect 12544 1660 12579 1694
rect 12613 1660 12648 1694
rect 12682 1660 12717 1694
rect 12751 1660 12786 1694
rect 12820 1660 12855 1694
rect 12889 1660 12924 1694
rect 12958 1660 12993 1694
rect 9716 1626 12993 1660
rect 9716 1592 9750 1626
rect 9784 1592 9819 1626
rect 9853 1592 9888 1626
rect 9922 1592 9957 1626
rect 9991 1592 10026 1626
rect 10060 1592 10095 1626
rect 10129 1592 10164 1626
rect 10198 1592 10233 1626
rect 10267 1592 10302 1626
rect 10336 1592 10371 1626
rect 10405 1592 10440 1626
rect 10474 1592 10509 1626
rect 10543 1592 10578 1626
rect 10612 1592 10647 1626
rect 10681 1592 10716 1626
rect 10750 1592 10785 1626
rect 10819 1592 10854 1626
rect 10888 1592 10923 1626
rect 10957 1592 10992 1626
rect 11026 1592 11061 1626
rect 11095 1592 11130 1626
rect 11164 1592 11199 1626
rect 11233 1592 11268 1626
rect 11302 1592 11337 1626
rect 11371 1592 11406 1626
rect 11440 1592 11475 1626
rect 11509 1592 11544 1626
rect 11578 1592 11613 1626
rect 11647 1592 11682 1626
rect 11716 1592 11751 1626
rect 11785 1592 11820 1626
rect 11854 1592 11889 1626
rect 11923 1592 11958 1626
rect 11992 1592 12027 1626
rect 12061 1592 12096 1626
rect 12130 1592 12165 1626
rect 12199 1592 12234 1626
rect 12268 1592 12303 1626
rect 12337 1592 12372 1626
rect 12406 1592 12441 1626
rect 12475 1592 12510 1626
rect 12544 1592 12579 1626
rect 12613 1592 12648 1626
rect 12682 1592 12717 1626
rect 12751 1592 12786 1626
rect 12820 1592 12855 1626
rect 12889 1592 12924 1626
rect 12958 1592 12993 1626
rect 19011 1889 19079 1923
rect 19113 1889 19152 1923
rect 19186 1889 19225 1923
rect 19259 1889 19298 1923
rect 19332 1889 19371 1923
rect 19405 1889 19444 1923
rect 19478 1889 19517 1923
rect 19551 1889 19585 1923
rect 19011 1849 19585 1889
rect 19011 1815 19079 1849
rect 19113 1815 19152 1849
rect 19186 1815 19225 1849
rect 19259 1815 19298 1849
rect 19332 1815 19371 1849
rect 19405 1815 19444 1849
rect 19478 1815 19517 1849
rect 19551 1815 19585 1849
rect 19011 1775 19585 1815
rect 19011 1741 19079 1775
rect 19113 1741 19152 1775
rect 19186 1741 19225 1775
rect 19259 1741 19298 1775
rect 19332 1741 19371 1775
rect 19405 1741 19444 1775
rect 19478 1741 19517 1775
rect 19551 1741 19585 1775
rect 19011 1701 19585 1741
rect 19011 1667 19079 1701
rect 19113 1667 19152 1701
rect 19186 1667 19225 1701
rect 19259 1667 19298 1701
rect 19332 1667 19371 1701
rect 19405 1667 19444 1701
rect 19478 1667 19517 1701
rect 19551 1667 19585 1701
rect 19011 1627 19585 1667
rect 19011 1593 19079 1627
rect 19113 1593 19152 1627
rect 19186 1593 19225 1627
rect 19259 1593 19298 1627
rect 19332 1593 19371 1627
rect 19405 1593 19444 1627
rect 19478 1593 19517 1627
rect 19551 1593 19585 1627
rect 19011 1592 19585 1593
rect 25787 1761 25821 1785
rect 25787 1690 25821 1727
rect 25787 1619 25821 1656
rect 25787 1548 25821 1585
rect 25787 1476 25821 1514
rect 25787 1404 25821 1442
rect 25787 1332 25821 1370
rect 25787 1260 25821 1298
rect 25787 1202 25821 1226
rect 8168 942 8202 966
rect 16344 1061 16394 1085
rect 8168 870 8202 908
rect 8168 798 8202 836
rect 8168 726 8202 764
rect 8168 654 8202 692
rect 8168 582 8202 620
rect 8168 510 8202 548
rect 8168 438 8202 476
rect 8168 366 8202 404
rect 8168 294 8202 332
rect 8168 222 8202 260
rect 8168 150 8202 188
rect 8168 78 8202 116
rect 8168 6 8202 44
rect 8168 -52 8202 -28
rect 10604 924 10638 948
rect 10604 854 10638 890
rect 10604 784 10638 820
rect 10604 714 10638 750
rect 10604 644 10638 680
rect 10604 574 10638 610
rect 10604 503 10638 540
rect 10604 432 10638 469
rect 10604 361 10638 398
rect 10604 290 10638 327
rect 10604 219 10638 256
rect 10604 148 10638 185
rect 10604 77 10638 114
rect 10604 6 10638 43
rect 10604 -52 10638 -28
rect 16344 1027 16352 1061
rect 16386 1027 16394 1061
rect 16344 974 16394 1027
rect 16344 940 16352 974
rect 16386 940 16394 974
rect 16344 887 16394 940
rect 16344 853 16352 887
rect 16386 853 16394 887
rect 12678 620 12712 644
rect 16344 800 16394 853
rect 16344 766 16352 800
rect 16386 766 16394 800
rect 16344 713 16394 766
rect 16344 679 16352 713
rect 16386 679 16394 713
rect 12678 547 12712 586
rect 12678 474 12712 513
rect 12678 401 12712 440
rect 16344 626 16394 679
rect 16344 592 16352 626
rect 16386 592 16394 626
rect 16344 539 16394 592
rect 16344 505 16352 539
rect 16386 505 16394 539
rect 12678 328 12712 367
rect 12678 255 12712 294
rect 12678 182 12712 221
rect 12678 109 12712 148
rect 16344 452 16394 505
rect 16344 418 16352 452
rect 16386 418 16394 452
rect 16344 365 16394 418
rect 16344 331 16352 365
rect 16386 331 16394 365
rect 16344 278 16394 331
rect 16344 244 16352 278
rect 16386 244 16394 278
rect 16344 191 16394 244
rect 12678 36 12712 75
rect 12678 -37 12712 2
rect 2398 -92 2422 -58
rect 2456 -92 2491 -58
rect 2525 -92 2560 -58
rect 2594 -92 2629 -58
rect 2663 -92 2698 -58
rect 2732 -92 2767 -58
rect 2801 -92 2836 -58
rect 2870 -92 2905 -58
rect 2939 -92 2974 -58
rect 3008 -92 3043 -58
rect 3077 -92 3112 -58
rect 3146 -92 3181 -58
rect 3215 -92 3250 -58
rect 3284 -92 3319 -58
rect 3353 -92 3388 -58
rect 3422 -92 3457 -58
rect 3491 -92 3526 -58
rect 3560 -92 3595 -58
rect 3629 -92 3664 -58
rect 3698 -92 3733 -58
rect 3767 -92 3802 -58
rect 3836 -92 3871 -58
rect 3905 -92 3940 -58
rect 3974 -92 4008 -58
rect 4042 -92 4076 -58
rect 4110 -92 4144 -58
rect 4178 -92 4212 -58
rect 4246 -92 4280 -58
rect 4314 -92 4348 -58
rect 4382 -92 4416 -58
rect 4450 -92 4484 -58
rect 4518 -92 4552 -58
rect 4586 -92 4620 -58
rect 4654 -92 4688 -58
rect 4722 -92 4756 -58
rect 4790 -92 4824 -58
rect 4858 -92 4892 -58
rect 4926 -92 4960 -58
rect 4994 -92 5028 -58
rect 5062 -92 5096 -58
rect 5130 -92 5164 -58
rect 5198 -92 5232 -58
rect 5266 -92 5300 -58
rect 5334 -92 5368 -58
rect 5402 -92 5436 -58
rect 5470 -92 5504 -58
rect 5538 -92 5572 -58
rect 5606 -92 5640 -58
rect 5674 -92 5708 -58
rect 5742 -92 5776 -58
rect 5810 -92 5844 -58
rect 5878 -92 5912 -58
rect 5946 -92 5980 -58
rect 6014 -92 6048 -58
rect 6082 -92 6116 -58
rect 6150 -92 6184 -58
rect 6218 -92 6252 -58
rect 6286 -92 6320 -58
rect 6354 -92 6388 -58
rect 6422 -92 6456 -58
rect 6490 -92 6524 -58
rect 6558 -92 6592 -58
rect 6626 -92 6660 -58
rect 6694 -92 6728 -58
rect 6762 -92 6796 -58
rect 6830 -92 6864 -58
rect 6898 -92 6922 -58
rect 13118 -71 13142 -37
rect 13176 -71 13211 -37
rect 13245 -71 13280 -37
rect 13314 -71 13349 -37
rect 13383 -71 13418 -37
rect 13452 -71 13486 -37
rect 13520 -71 13554 -37
rect 13588 -71 13622 -37
rect 13656 -71 13690 -37
rect 13724 -71 13758 -37
rect 13792 -71 13826 -37
rect 13860 -71 13894 -37
rect 13928 -71 13962 -37
rect 13996 -71 14030 -37
rect 14064 -71 14098 -37
rect 14132 -71 14166 -37
rect 14200 -71 14234 -37
rect 14268 -71 14302 -37
rect 14336 -71 14370 -37
rect 14404 -71 14438 -37
rect 14472 -71 14506 -37
rect 14540 -71 14574 -37
rect 14608 -71 14642 -37
rect 14676 -71 14710 -37
rect 14744 -71 14778 -37
rect 14812 -71 14846 -37
rect 14880 -71 14914 -37
rect 14948 -71 14982 -37
rect 15016 -71 15050 -37
rect 15084 -71 15118 -37
rect 15152 -71 15186 -37
rect 15220 -71 15254 -37
rect 15288 -71 15322 -37
rect 15356 -71 15390 -37
rect 15424 -71 15458 -37
rect 15492 -71 15526 -37
rect 15560 -71 15594 -37
rect 15628 -71 15662 -37
rect 15696 -71 15730 -37
rect 15764 -71 15788 -37
rect 12678 -95 12712 -71
rect 16344 157 16352 191
rect 16386 157 16394 191
rect 16344 104 16394 157
rect 16344 70 16352 104
rect 16386 70 16394 104
rect 16344 17 16394 70
rect 16344 -17 16352 17
rect 16386 -17 16394 17
rect 16344 -70 16394 -17
rect 16344 -104 16352 -70
rect 16386 -104 16394 -70
rect 16344 -157 16394 -104
rect 16344 -191 16352 -157
rect 16386 -191 16394 -157
rect 16344 -245 16394 -191
rect 16344 -279 16352 -245
rect 16386 -279 16394 -245
rect 16344 -333 16394 -279
rect 16344 -367 16352 -333
rect 16386 -367 16394 -333
rect 16344 -421 16394 -367
rect 16344 -455 16352 -421
rect 16386 -455 16394 -421
rect 16344 -509 16394 -455
rect 16344 -543 16352 -509
rect 16386 -543 16394 -509
rect 16344 -597 16394 -543
rect 16344 -631 16352 -597
rect 16386 -631 16394 -597
rect 16344 -685 16394 -631
rect 16344 -719 16352 -685
rect 16386 -719 16394 -685
rect 16344 -773 16394 -719
rect 16344 -807 16352 -773
rect 16386 -807 16394 -773
rect 16344 -861 16394 -807
rect 16344 -895 16352 -861
rect 16386 -895 16394 -861
rect 16344 -929 16394 -895
rect 15874 -937 16394 -929
rect 15874 -971 15898 -937
rect 15932 -971 15991 -937
rect 16025 -971 16084 -937
rect 16118 -971 16176 -937
rect 16210 -971 16268 -937
rect 16302 -971 16394 -937
rect 15874 -979 16394 -971
rect 406 -3265 495 -3231
rect 529 -3265 563 -3231
rect 597 -3265 631 -3231
rect 665 -3265 699 -3231
rect 733 -3265 767 -3231
rect 801 -3265 835 -3231
rect 869 -3265 903 -3231
rect 937 -3265 971 -3231
rect 1005 -3265 1073 -3231
rect 406 -3299 440 -3265
rect 406 -3367 440 -3333
rect 1039 -3321 1073 -3265
rect 406 -3435 440 -3401
rect 406 -3503 440 -3469
rect 406 -3571 440 -3537
rect 406 -3639 440 -3605
rect 406 -3746 440 -3673
rect 406 -3814 440 -3780
rect 406 -3882 440 -3848
rect 406 -3950 440 -3916
rect 406 -4018 440 -3984
rect 406 -4086 440 -4052
rect 406 -4154 440 -4120
rect 406 -4222 440 -4188
rect 406 -4290 440 -4256
rect 406 -4358 440 -4324
rect 406 -4426 440 -4392
rect 406 -4494 440 -4460
rect 406 -4562 440 -4528
rect 406 -4630 440 -4596
rect 406 -4698 440 -4664
rect 406 -4766 440 -4732
rect 406 -4834 440 -4800
rect 406 -4902 440 -4868
rect 406 -4970 440 -4936
rect 406 -5038 440 -5004
rect 406 -5106 440 -5072
rect 406 -5174 440 -5140
rect 406 -5242 440 -5208
rect 406 -5310 440 -5276
rect 406 -5378 440 -5344
rect 406 -5446 440 -5412
rect 406 -5514 440 -5480
rect 406 -5582 440 -5548
rect 406 -5650 440 -5616
rect 406 -5718 440 -5684
rect 406 -5786 440 -5752
rect 406 -5854 440 -5820
rect 406 -5922 440 -5888
rect 406 -5990 440 -5956
rect 406 -6058 440 -6024
rect 406 -6126 440 -6092
rect 406 -6194 440 -6160
rect 406 -6262 440 -6228
rect 406 -6330 440 -6296
rect 406 -6398 440 -6364
rect 406 -6466 440 -6432
rect 406 -6534 440 -6500
rect 406 -6602 440 -6568
rect 406 -6670 440 -6636
rect 406 -6738 440 -6704
rect 406 -6806 440 -6772
rect 406 -6874 440 -6840
rect 406 -6942 440 -6908
rect 406 -7010 440 -6976
rect 406 -7078 440 -7044
rect 406 -7146 440 -7112
rect 406 -7214 440 -7180
rect 406 -7282 440 -7248
rect 406 -7350 440 -7316
rect 406 -7418 440 -7384
rect 406 -7486 440 -7452
rect 406 -7554 440 -7520
rect 406 -7622 440 -7588
rect 406 -7690 440 -7656
rect 406 -7758 440 -7724
rect 406 -7826 440 -7792
rect 406 -7894 440 -7860
rect 406 -7962 440 -7928
rect 406 -8030 440 -7996
rect 406 -8098 440 -8064
rect 406 -8166 440 -8132
rect 406 -8234 440 -8200
rect 406 -8302 440 -8268
rect 406 -8370 440 -8336
rect 406 -8438 440 -8404
rect 406 -8506 440 -8472
rect 406 -8574 440 -8540
rect 406 -8642 440 -8608
rect 406 -8710 440 -8676
rect 406 -8778 440 -8744
rect 406 -8846 440 -8812
rect 406 -8914 440 -8880
rect 406 -8982 440 -8948
rect 406 -9050 440 -9016
rect 406 -9118 440 -9084
rect 406 -9186 440 -9152
rect 406 -9254 440 -9220
rect 406 -9322 440 -9288
rect 406 -9390 440 -9356
rect 406 -9458 440 -9424
rect 406 -9526 440 -9492
rect 406 -9594 440 -9560
rect 406 -9662 440 -9628
rect 406 -9730 440 -9696
rect 406 -9798 440 -9764
rect 406 -9866 440 -9832
rect 406 -9934 440 -9900
rect 406 -10002 440 -9968
rect 406 -10070 440 -10036
rect 406 -10138 440 -10104
rect 406 -10206 440 -10172
rect 406 -10274 440 -10240
rect 406 -10342 440 -10308
rect 406 -10410 440 -10376
rect 406 -10478 440 -10444
rect 406 -10546 440 -10512
rect 406 -10614 440 -10580
rect 406 -10682 440 -10648
rect 406 -10750 440 -10716
rect 406 -10818 440 -10784
rect 406 -10886 440 -10852
rect 406 -10954 440 -10920
rect 1039 -3389 1073 -3355
rect 1039 -3457 1073 -3423
rect 1039 -3525 1073 -3491
rect 1039 -3593 1073 -3559
rect 1039 -3661 1073 -3627
rect 1039 -3729 1073 -3695
rect 1039 -3797 1073 -3763
rect 1039 -3865 1073 -3831
rect 1039 -3933 1073 -3899
rect 1039 -4001 1073 -3967
rect 1039 -4069 1073 -4035
rect 1039 -4137 1073 -4103
rect 1039 -4205 1073 -4171
rect 1039 -4273 1073 -4239
rect 1039 -4341 1073 -4307
rect 1039 -4409 1073 -4375
rect 1039 -4477 1073 -4443
rect 1039 -4545 1073 -4511
rect 1039 -4613 1073 -4579
rect 1039 -4681 1073 -4647
rect 1039 -4749 1073 -4715
rect 1039 -4817 1073 -4783
rect 1039 -4885 1073 -4851
rect 1039 -4953 1073 -4919
rect 1039 -5021 1073 -4987
rect 1039 -5089 1073 -5055
rect 1039 -5157 1073 -5123
rect 1039 -5225 1073 -5191
rect 1039 -5293 1073 -5259
rect 1039 -5361 1073 -5327
rect 1039 -5429 1073 -5395
rect 1039 -5497 1073 -5463
rect 1039 -5565 1073 -5531
rect 1039 -5633 1073 -5599
rect 1039 -5701 1073 -5667
rect 1039 -5769 1073 -5735
rect 1039 -5837 1073 -5803
rect 1039 -5905 1073 -5871
rect 1039 -5973 1073 -5939
rect 1039 -6041 1073 -6007
rect 1039 -6109 1073 -6075
rect 1039 -6177 1073 -6143
rect 1039 -6245 1073 -6211
rect 1039 -6313 1073 -6279
rect 1039 -6381 1073 -6347
rect 1039 -6449 1073 -6415
rect 1039 -6517 1073 -6483
rect 1039 -6585 1073 -6551
rect 1039 -6653 1073 -6619
rect 1039 -6721 1073 -6687
rect 1039 -6789 1073 -6755
rect 1039 -6857 1073 -6823
rect 1039 -6925 1073 -6891
rect 1039 -6993 1073 -6959
rect 1039 -7061 1073 -7027
rect 1039 -7129 1073 -7095
rect 1039 -7197 1073 -7163
rect 1039 -7265 1073 -7231
rect 1039 -7333 1073 -7299
rect 1039 -7401 1073 -7367
rect 1039 -7469 1073 -7435
rect 1039 -7537 1073 -7503
rect 1039 -7605 1073 -7571
rect 1039 -7673 1073 -7639
rect 1039 -7741 1073 -7707
rect 1039 -7809 1073 -7775
rect 1039 -7877 1073 -7843
rect 1039 -7945 1073 -7911
rect 1039 -8013 1073 -7979
rect 1039 -8081 1073 -8047
rect 1039 -8149 1073 -8115
rect 1039 -8217 1073 -8183
rect 1039 -8285 1073 -8251
rect 1039 -8353 1073 -8319
rect 1039 -8421 1073 -8387
rect 1039 -8489 1073 -8455
rect 1039 -8557 1073 -8523
rect 1039 -8625 1073 -8591
rect 1039 -8693 1073 -8659
rect 1039 -8761 1073 -8727
rect 1039 -8829 1073 -8795
rect 1039 -8897 1073 -8863
rect 1039 -8965 1073 -8931
rect 1039 -9033 1073 -8999
rect 1039 -9101 1073 -9067
rect 1039 -9169 1073 -9135
rect 1039 -9237 1073 -9203
rect 1039 -9305 1073 -9271
rect 1039 -9373 1073 -9339
rect 1039 -9441 1073 -9407
rect 1039 -9509 1073 -9475
rect 1039 -9577 1073 -9543
rect 1039 -9645 1073 -9611
rect 1039 -9713 1073 -9679
rect 1039 -9781 1073 -9747
rect 1039 -9849 1073 -9815
rect 1039 -9917 1073 -9883
rect 1039 -9985 1073 -9951
rect 1039 -10053 1073 -10019
rect 1039 -10121 1073 -10087
rect 1039 -10189 1073 -10155
rect 1039 -10257 1073 -10223
rect 1039 -10325 1073 -10291
rect 1039 -10393 1073 -10359
rect 1039 -10461 1073 -10427
rect 1039 -10529 1073 -10495
rect 1039 -10597 1073 -10563
rect 1039 -10665 1073 -10631
rect 1039 -10733 1073 -10699
rect 1039 -10801 1073 -10767
rect 1039 -10869 1073 -10835
rect 1039 -10937 1073 -10903
rect 406 -11073 440 -10988
rect 1039 -11005 1073 -10971
rect 1039 -11073 1073 -11039
rect 406 -11107 474 -11073
rect 508 -11107 542 -11073
rect 576 -11107 610 -11073
rect 644 -11107 678 -11073
rect 712 -11107 746 -11073
rect 780 -11107 814 -11073
rect 848 -11107 882 -11073
rect 916 -11107 950 -11073
rect 984 -11107 1073 -11073
<< mvnsubdiff >>
rect 8482 4883 8550 4917
rect 8584 4883 8620 4917
rect 8654 4883 8690 4917
rect 8724 4883 8760 4917
rect 8794 4883 8830 4917
rect 8864 4883 8900 4917
rect 8934 4883 8970 4917
rect 9004 4883 9040 4917
rect 9074 4883 9110 4917
rect 9144 4883 9180 4917
rect 9214 4883 9250 4917
rect 9284 4883 9320 4917
rect 9354 4883 9390 4917
rect 9424 4883 9460 4917
rect 9494 4883 9530 4917
rect 9564 4883 9599 4917
rect 9633 4883 9668 4917
rect 9702 4883 9737 4917
rect 9771 4883 9806 4917
rect 9840 4883 9875 4917
rect 9909 4883 9944 4917
rect 9978 4883 10013 4917
rect 10047 4883 10082 4917
rect 10116 4883 10151 4917
rect 10185 4883 10220 4917
rect 10254 4883 10289 4917
rect 10323 4883 10358 4917
rect 10392 4883 10427 4917
rect 10461 4883 10496 4917
rect 10530 4883 10565 4917
rect 10599 4883 10634 4917
rect 10668 4883 10703 4917
rect 10737 4883 10772 4917
rect 10806 4883 10841 4917
rect 10875 4883 10910 4917
rect 10944 4883 10979 4917
rect 11013 4883 11048 4917
rect 11082 4883 11117 4917
rect 11151 4883 11186 4917
rect 11220 4883 11322 4917
rect 11356 4883 11391 4917
rect 11425 4883 11460 4917
rect 11494 4883 11529 4917
rect 11563 4883 11598 4917
rect 11632 4883 11667 4917
rect 11701 4883 11736 4917
rect 11770 4883 11805 4917
rect 11839 4883 11874 4917
rect 11908 4883 11943 4917
rect 11977 4883 12012 4917
rect 12046 4883 12081 4917
rect 12115 4883 12150 4917
rect 12184 4883 12219 4917
rect 12253 4883 12288 4917
rect 12322 4883 12357 4917
rect 12391 4883 12426 4917
rect 12460 4883 12495 4917
rect 12529 4883 12563 4917
rect 12597 4883 12631 4917
rect 12665 4883 12699 4917
rect 12733 4883 12767 4917
rect 12801 4883 12835 4917
rect 12869 4883 12903 4917
rect 12937 4883 12971 4917
rect 13005 4883 13039 4917
rect 13073 4883 13107 4917
rect 13141 4883 13175 4917
rect 13209 4883 13243 4917
rect 13277 4883 13311 4917
rect 13345 4883 13379 4917
rect 13413 4883 13447 4917
rect 13481 4883 13515 4917
rect 13549 4883 13583 4917
rect 13617 4883 13651 4917
rect 13685 4883 13719 4917
rect 13753 4883 13787 4917
rect 13821 4883 13855 4917
rect 13889 4883 13923 4917
rect 13957 4883 13991 4917
rect 14025 4883 14059 4917
rect 14093 4883 14127 4917
rect 14161 4883 14195 4917
rect 14229 4883 14263 4917
rect 14297 4883 14331 4917
rect 14365 4883 14399 4917
rect 14433 4883 14467 4917
rect 14501 4883 14535 4917
rect 14569 4883 14603 4917
rect 14637 4883 14671 4917
rect 14705 4883 14739 4917
rect 14773 4883 14807 4917
rect 14841 4883 14875 4917
rect 14909 4883 14943 4917
rect 14977 4883 15011 4917
rect 15045 4883 15079 4917
rect 15113 4883 15147 4917
rect 15181 4883 15215 4917
rect 15249 4883 15283 4917
rect 15317 4883 15351 4917
rect 15385 4883 15419 4917
rect 15453 4883 15487 4917
rect 15521 4883 15555 4917
rect 15589 4883 15623 4917
rect 15657 4883 15691 4917
rect 15725 4883 15759 4917
rect 15793 4883 15827 4917
rect 15861 4883 15895 4917
rect 15929 4883 15963 4917
rect 15997 4883 16031 4917
rect 16065 4883 16099 4917
rect 16133 4883 16167 4917
rect 16201 4883 16235 4917
rect 16269 4883 16303 4917
rect 16337 4883 16371 4917
rect 16405 4883 16439 4917
rect 16473 4883 16507 4917
rect 16541 4883 16575 4917
rect 16609 4883 16643 4917
rect 16677 4883 16711 4917
rect 16745 4883 16779 4917
rect 16813 4883 16847 4917
rect 16881 4883 16915 4917
rect 16949 4883 16983 4917
rect 17017 4883 17051 4917
rect 17085 4883 17119 4917
rect 17153 4883 17187 4917
rect 17221 4883 17255 4917
rect 17289 4883 17323 4917
rect 17357 4883 17391 4917
rect 17425 4883 17459 4917
rect 17493 4883 17527 4917
rect 17561 4883 17595 4917
rect 17629 4883 17663 4917
rect 17697 4883 17731 4917
rect 17765 4883 17799 4917
rect 17833 4883 17867 4917
rect 17901 4883 17935 4917
rect 17969 4883 18003 4917
rect 18037 4883 18071 4917
rect 18105 4883 18139 4917
rect 18173 4883 18207 4917
rect 18241 4883 18275 4917
rect 18309 4883 18343 4917
rect 18377 4883 18411 4917
rect 18445 4883 18479 4917
rect 18513 4883 18547 4917
rect 18581 4883 18615 4917
rect 18649 4883 18683 4917
rect 18717 4883 18751 4917
rect 18785 4883 18819 4917
rect 18853 4883 18887 4917
rect 18921 4883 18955 4917
rect 18989 4883 19023 4917
rect 19057 4883 19091 4917
rect 19125 4883 19159 4917
rect 19193 4883 19227 4917
rect 19261 4883 19295 4917
rect 19329 4883 19363 4917
rect 19397 4883 19431 4917
rect 19465 4883 19499 4917
rect 19533 4883 19567 4917
rect 19601 4883 19635 4917
rect 19669 4883 19703 4917
rect 19737 4883 19771 4917
rect 19805 4883 19839 4917
rect 19873 4883 19907 4917
rect 19941 4883 20009 4917
rect 8482 4848 8516 4883
rect 8482 4779 8516 4814
rect 8482 4710 8516 4745
rect 8482 4641 8516 4676
rect 8482 4572 8516 4607
rect 8482 4503 8516 4538
rect 8482 4434 8516 4469
rect 8482 4365 8516 4400
rect 8482 4296 8516 4331
rect 8482 4226 8516 4262
rect 8482 4156 8516 4192
rect 8482 4086 8516 4122
rect 8482 4016 8516 4052
rect 8482 3946 8516 3982
rect 8482 3876 8516 3912
rect 8482 3806 8516 3842
rect 11254 4783 11288 4883
rect 11254 4715 11288 4749
rect 11254 4647 11288 4681
rect 11254 4579 11288 4613
rect 11254 4511 11288 4545
rect 11254 4443 11288 4477
rect 11254 4375 11288 4409
rect 11254 4307 11288 4341
rect 11254 4239 11288 4273
rect 11254 4171 11288 4205
rect 11254 4103 11288 4137
rect 11254 4035 11288 4069
rect 11254 3967 11288 4001
rect 11254 3899 11288 3933
rect 11254 3831 11288 3865
rect 8482 3736 8516 3772
rect 8482 3666 8516 3702
rect 8482 3596 8516 3632
rect 11254 3763 11288 3797
rect 11254 3695 11288 3729
rect 8482 3526 8516 3562
rect 11254 3627 11288 3661
rect 19975 4835 20009 4883
rect 19975 4674 20009 4801
rect 19975 4606 20009 4640
rect 19975 4538 20009 4572
rect 19975 4470 20009 4504
rect 19975 4402 20009 4436
rect 19975 4334 20009 4368
rect 19975 4266 20009 4300
rect 19975 4198 20009 4232
rect 19975 4130 20009 4164
rect 19975 4062 20009 4096
rect 19975 3994 20009 4028
rect 19975 3926 20009 3960
rect 19975 3858 20009 3892
rect 19975 3790 20009 3824
rect 19975 3722 20009 3756
rect 19975 3654 20009 3688
rect 8482 3456 8516 3492
rect 11254 3559 11288 3593
rect 11254 3491 11288 3525
rect 8482 3386 8516 3422
rect 11254 3382 11288 3457
rect 19975 3586 20009 3620
rect 19975 3518 20009 3552
rect 19975 3450 20009 3484
rect 19975 3382 20009 3416
rect 8482 3316 8516 3352
rect 8482 3246 8516 3282
rect 8482 3176 8516 3212
rect 11254 3348 11322 3382
rect 11356 3348 11390 3382
rect 11424 3348 11458 3382
rect 11492 3348 11526 3382
rect 11560 3348 11594 3382
rect 11628 3348 11662 3382
rect 11696 3348 11730 3382
rect 11764 3348 11798 3382
rect 11832 3348 11866 3382
rect 11900 3348 11934 3382
rect 11968 3348 12002 3382
rect 12036 3348 12070 3382
rect 12104 3348 12138 3382
rect 12172 3348 12206 3382
rect 12240 3348 12274 3382
rect 12308 3348 12342 3382
rect 12376 3348 12410 3382
rect 12444 3348 12478 3382
rect 12512 3348 12546 3382
rect 12580 3348 12614 3382
rect 12648 3348 12682 3382
rect 12716 3348 12750 3382
rect 12784 3348 12818 3382
rect 12852 3348 12886 3382
rect 12920 3348 12954 3382
rect 12988 3348 13022 3382
rect 13056 3348 13090 3382
rect 13124 3348 13158 3382
rect 13192 3348 13226 3382
rect 13260 3348 13294 3382
rect 13328 3348 13362 3382
rect 13396 3348 13430 3382
rect 13464 3348 13498 3382
rect 13532 3348 13566 3382
rect 13600 3348 13634 3382
rect 13668 3348 13702 3382
rect 13736 3348 13770 3382
rect 13804 3348 13838 3382
rect 13872 3348 13906 3382
rect 13940 3348 13974 3382
rect 14008 3348 14042 3382
rect 14076 3348 14110 3382
rect 14144 3348 14178 3382
rect 14212 3348 14246 3382
rect 14280 3348 14314 3382
rect 14348 3348 14382 3382
rect 14416 3348 14450 3382
rect 14484 3348 14518 3382
rect 14552 3348 14586 3382
rect 14620 3348 14654 3382
rect 14688 3348 14722 3382
rect 14756 3348 14790 3382
rect 14824 3348 14858 3382
rect 14892 3348 14926 3382
rect 14960 3348 14994 3382
rect 15028 3348 15062 3382
rect 15096 3348 15130 3382
rect 15164 3348 15198 3382
rect 15232 3348 15266 3382
rect 15300 3348 15334 3382
rect 15368 3348 15402 3382
rect 15436 3348 15470 3382
rect 15504 3348 15538 3382
rect 15572 3348 15606 3382
rect 15640 3348 15674 3382
rect 15708 3348 15742 3382
rect 15776 3348 15810 3382
rect 15844 3348 15878 3382
rect 15912 3348 15946 3382
rect 15980 3348 16014 3382
rect 16048 3348 16082 3382
rect 16116 3348 16150 3382
rect 16184 3348 16218 3382
rect 16252 3348 16286 3382
rect 16320 3348 16354 3382
rect 16388 3348 16422 3382
rect 16456 3348 16490 3382
rect 16524 3348 16558 3382
rect 16592 3348 16626 3382
rect 16660 3348 16694 3382
rect 16728 3348 16762 3382
rect 16796 3348 16830 3382
rect 16864 3348 16898 3382
rect 16932 3348 16966 3382
rect 17000 3348 17034 3382
rect 17068 3348 17102 3382
rect 17136 3348 17170 3382
rect 17204 3348 17238 3382
rect 17272 3348 17306 3382
rect 17340 3348 17374 3382
rect 17408 3348 17442 3382
rect 17476 3348 17510 3382
rect 17544 3348 17578 3382
rect 17612 3348 17646 3382
rect 17680 3348 17714 3382
rect 17748 3348 17782 3382
rect 17816 3348 17850 3382
rect 17884 3348 17918 3382
rect 17952 3348 17986 3382
rect 18020 3348 18054 3382
rect 18088 3348 18122 3382
rect 18156 3348 18190 3382
rect 18224 3348 18258 3382
rect 18292 3348 18326 3382
rect 18360 3348 18394 3382
rect 18428 3348 18462 3382
rect 18496 3348 18530 3382
rect 18564 3348 18598 3382
rect 18632 3348 18666 3382
rect 18700 3348 18734 3382
rect 18768 3348 18802 3382
rect 18836 3348 18870 3382
rect 18904 3348 18938 3382
rect 18972 3348 19006 3382
rect 19040 3348 19074 3382
rect 19108 3348 19142 3382
rect 19176 3348 19210 3382
rect 19244 3348 19278 3382
rect 19312 3348 19346 3382
rect 19380 3348 19414 3382
rect 19448 3348 19482 3382
rect 19516 3348 19550 3382
rect 19584 3348 19618 3382
rect 19652 3348 19686 3382
rect 19720 3348 19754 3382
rect 19788 3348 19822 3382
rect 19856 3348 19890 3382
rect 19924 3348 20009 3382
rect 11254 3314 11302 3348
rect 11254 3280 11261 3314
rect 11295 3280 11302 3314
rect 11254 3231 11302 3280
rect 11254 3197 11261 3231
rect 11295 3197 11302 3231
rect 8482 3106 8516 3142
rect 11254 3148 11302 3197
rect 11254 3114 11261 3148
rect 11295 3114 11302 3148
rect 11254 3094 11302 3114
rect 8482 3036 8516 3072
rect 10295 3087 11302 3094
rect 10295 3053 10401 3087
rect 10435 3053 10474 3087
rect 10508 3053 10547 3087
rect 10581 3053 10620 3087
rect 10654 3053 10692 3087
rect 10726 3053 10764 3087
rect 10798 3053 10836 3087
rect 10870 3053 10908 3087
rect 10942 3053 10980 3087
rect 11014 3053 11052 3087
rect 11086 3053 11124 3087
rect 11158 3053 11196 3087
rect 11230 3053 11302 3087
rect 10295 3046 11302 3053
rect 10295 3002 10337 3046
rect 8482 2968 8550 3002
rect 8584 2968 8619 3002
rect 8653 2968 8688 3002
rect 8722 2968 8757 3002
rect 8791 2968 8826 3002
rect 8860 2968 8895 3002
rect 8929 2968 8964 3002
rect 8998 2968 9033 3002
rect 9067 2968 9102 3002
rect 9136 2968 9171 3002
rect 9205 2968 9240 3002
rect 9274 2968 9309 3002
rect 9343 2968 9378 3002
rect 9412 2968 9447 3002
rect 9481 2968 9516 3002
rect 9550 2968 9585 3002
rect 9619 2968 9654 3002
rect 9688 2968 9723 3002
rect 9757 2968 9792 3002
rect 9826 2968 9861 3002
rect 9895 2968 9929 3002
rect 9963 2968 9997 3002
rect 10031 2968 10065 3002
rect 10099 2968 10133 3002
rect 10167 2968 10201 3002
rect 10235 2968 10269 3002
rect 10303 2968 10337 3002
rect 574 2518 598 2552
rect 632 2518 668 2552
rect 702 2518 738 2552
rect 772 2518 808 2552
rect 842 2518 878 2552
rect 912 2518 948 2552
rect 982 2518 1019 2552
rect 1053 2518 1090 2552
rect 1124 2518 1161 2552
rect 1195 2518 1232 2552
rect 1266 2518 1303 2552
rect 1337 2518 1374 2552
rect 1408 2518 1445 2552
rect 1479 2518 1516 2552
rect 1550 2518 1574 2552
rect 2151 2465 2271 2499
rect 2305 2465 2339 2499
rect 2373 2465 2407 2499
rect 2441 2465 2475 2499
rect 2509 2465 2543 2499
rect 2577 2465 2611 2499
rect 2645 2465 2679 2499
rect 2713 2465 2747 2499
rect 2781 2465 2815 2499
rect 2849 2465 2883 2499
rect 2917 2465 2951 2499
rect 2985 2465 3019 2499
rect 3053 2465 3087 2499
rect 3121 2465 3155 2499
rect 3189 2465 3223 2499
rect 3257 2465 3291 2499
rect 3325 2465 3359 2499
rect 3393 2465 3427 2499
rect 3461 2465 3495 2499
rect 3529 2465 3563 2499
rect 3597 2465 3631 2499
rect 3665 2465 3699 2499
rect 3733 2465 3767 2499
rect 3801 2465 3835 2499
rect 3869 2465 3903 2499
rect 3937 2465 3971 2499
rect 4005 2465 4039 2499
rect 4073 2465 4107 2499
rect 4141 2465 4175 2499
rect 4209 2465 4243 2499
rect 4277 2465 4311 2499
rect 4345 2465 4379 2499
rect 4413 2465 4447 2499
rect 4481 2465 4515 2499
rect 4549 2465 4583 2499
rect 4617 2465 4651 2499
rect 4685 2465 4719 2499
rect 4753 2465 4787 2499
rect 4821 2465 4855 2499
rect 4889 2465 4923 2499
rect 4957 2465 4991 2499
rect 5025 2465 5059 2499
rect 5093 2465 5127 2499
rect 5161 2465 5195 2499
rect 5229 2465 5263 2499
rect 5297 2465 5331 2499
rect 5365 2465 5399 2499
rect 5433 2465 5467 2499
rect 5501 2465 5535 2499
rect 5569 2465 5603 2499
rect 5637 2465 5671 2499
rect 5705 2465 5739 2499
rect 5773 2465 5807 2499
rect 5841 2465 5875 2499
rect 5909 2465 5943 2499
rect 5977 2465 6011 2499
rect 6045 2465 6079 2499
rect 6113 2465 6147 2499
rect 6181 2465 6215 2499
rect 6249 2465 6283 2499
rect 6317 2465 6351 2499
rect 6385 2465 6419 2499
rect 6453 2465 6487 2499
rect 6521 2465 6555 2499
rect 6589 2465 6623 2499
rect 6657 2465 6691 2499
rect 6725 2465 6759 2499
rect 6793 2465 6827 2499
rect 6861 2465 6895 2499
rect 6929 2465 6963 2499
rect 6997 2465 7031 2499
rect 7065 2465 7099 2499
rect 7133 2465 7167 2499
rect 7201 2465 7235 2499
rect 7269 2465 7303 2499
rect 7337 2465 7371 2499
rect 7405 2465 7439 2499
rect 7473 2465 7507 2499
rect 7541 2465 7575 2499
rect 7609 2465 7643 2499
rect 7677 2465 7711 2499
rect 7745 2465 7779 2499
rect 7813 2465 7847 2499
rect 7881 2465 7915 2499
rect 7949 2465 7983 2499
rect 8017 2465 8051 2499
rect 8085 2465 8119 2499
rect 8153 2465 8187 2499
rect 8221 2465 8255 2499
rect 8289 2465 8323 2499
rect 8357 2465 8391 2499
rect 8425 2465 8459 2499
rect 8493 2465 8527 2499
rect 8561 2465 8595 2499
rect 8629 2465 8663 2499
rect 8697 2465 8731 2499
rect 8765 2465 8799 2499
rect 8833 2465 8867 2499
rect 8901 2465 8935 2499
rect 8969 2465 9003 2499
rect 9037 2465 9071 2499
rect 9105 2465 9139 2499
rect 9173 2465 9207 2499
rect 9241 2465 9275 2499
rect 9309 2465 9343 2499
rect 9377 2465 9445 2499
rect 2151 2431 2185 2465
rect 2151 2363 2185 2397
rect 2151 2295 2185 2329
rect 2151 2227 2185 2261
rect 9411 2375 9445 2465
rect 9411 2307 9445 2341
rect 574 2130 598 2164
rect 632 2130 669 2164
rect 703 2130 740 2164
rect 774 2130 811 2164
rect 845 2130 882 2164
rect 916 2130 953 2164
rect 987 2130 1024 2164
rect 1058 2130 1095 2164
rect 1129 2130 1166 2164
rect 1200 2130 1236 2164
rect 1270 2130 1306 2164
rect 1340 2130 1376 2164
rect 1410 2130 1446 2164
rect 1480 2130 1516 2164
rect 1550 2130 1574 2164
rect 574 2096 1574 2130
rect 574 2062 598 2096
rect 632 2062 669 2096
rect 703 2062 740 2096
rect 774 2062 811 2096
rect 845 2062 882 2096
rect 916 2062 953 2096
rect 987 2062 1024 2096
rect 1058 2062 1095 2096
rect 1129 2062 1166 2096
rect 1200 2062 1236 2096
rect 1270 2062 1306 2096
rect 1340 2062 1376 2096
rect 1410 2062 1446 2096
rect 1480 2062 1516 2096
rect 1550 2062 1574 2096
rect 574 2028 1574 2062
rect 574 1994 598 2028
rect 632 1994 669 2028
rect 703 1994 740 2028
rect 774 1994 811 2028
rect 845 1994 882 2028
rect 916 1994 953 2028
rect 987 1994 1024 2028
rect 1058 1994 1095 2028
rect 1129 1994 1166 2028
rect 1200 1994 1236 2028
rect 1270 1994 1306 2028
rect 1340 1994 1376 2028
rect 1410 1994 1446 2028
rect 1480 1994 1516 2028
rect 1550 1994 1574 2028
rect 574 1960 1574 1994
rect 574 1926 598 1960
rect 632 1926 669 1960
rect 703 1926 740 1960
rect 774 1926 811 1960
rect 845 1926 882 1960
rect 916 1926 953 1960
rect 987 1926 1024 1960
rect 1058 1926 1095 1960
rect 1129 1926 1166 1960
rect 1200 1926 1236 1960
rect 1270 1926 1306 1960
rect 1340 1926 1376 1960
rect 1410 1926 1446 1960
rect 1480 1926 1516 1960
rect 1550 1926 1574 1960
rect 2151 2159 2185 2193
rect 9411 2239 9445 2273
rect 2151 2091 2185 2125
rect 9411 2171 9445 2205
rect 9411 2103 9445 2137
rect 2151 2023 2185 2057
rect 2151 1955 2185 1989
rect 2151 1887 2185 1921
rect 2151 1819 2185 1853
rect 2151 1751 2185 1785
rect 2151 1683 2185 1717
rect 9411 2035 9445 2069
rect 9411 1967 9445 2001
rect 9411 1899 9445 1933
rect 9411 1831 9445 1865
rect 9411 1763 9445 1797
rect 2151 1615 2185 1649
rect 9411 1695 9445 1729
rect 9411 1627 9445 1661
rect 2151 1547 2185 1581
rect 2151 1479 2185 1513
rect 2151 1411 2185 1445
rect 9411 1559 9445 1593
rect 17793 2572 17817 2606
rect 17851 2572 17889 2606
rect 17923 2572 17961 2606
rect 17995 2572 18033 2606
rect 18067 2572 18105 2606
rect 18139 2572 18176 2606
rect 18210 2572 18247 2606
rect 18281 2572 18318 2606
rect 18352 2572 18389 2606
rect 18423 2572 18460 2606
rect 18494 2572 18531 2606
rect 18565 2572 18602 2606
rect 18636 2572 18673 2606
rect 18707 2572 18744 2606
rect 18778 2572 18815 2606
rect 18849 2572 18886 2606
rect 18920 2572 18957 2606
rect 18991 2572 19028 2606
rect 19062 2572 19086 2606
rect 28031 1795 28065 1829
rect 9411 1491 9445 1525
rect 574 1367 598 1401
rect 632 1367 668 1401
rect 702 1367 738 1401
rect 772 1367 808 1401
rect 842 1367 878 1401
rect 912 1367 948 1401
rect 982 1367 1019 1401
rect 1053 1367 1090 1401
rect 1124 1367 1161 1401
rect 1195 1367 1232 1401
rect 1266 1367 1303 1401
rect 1337 1367 1374 1401
rect 1408 1367 1445 1401
rect 1479 1367 1516 1401
rect 1550 1367 1574 1401
rect 2151 1343 2185 1377
rect 2151 1275 2185 1309
rect 2151 1207 2185 1241
rect 9411 1423 9445 1457
rect 2151 1139 2185 1173
rect 2151 1071 2185 1105
rect 2151 1003 2185 1037
rect 2151 935 2185 969
rect 2151 867 2185 901
rect 2151 799 2185 833
rect 2151 731 2185 765
rect 2151 663 2185 697
rect 2151 595 2185 629
rect 2151 527 2185 561
rect 2151 459 2185 493
rect 2151 391 2185 425
rect 2151 323 2185 357
rect 2151 255 2185 289
rect 2151 187 2185 221
rect 2151 119 2185 153
rect 2151 51 2185 85
rect 2151 -17 2185 17
rect 9411 1355 9445 1389
rect 9411 1321 9479 1355
rect 9513 1321 9547 1355
rect 9581 1321 9615 1355
rect 9649 1321 9683 1355
rect 9717 1321 9751 1355
rect 9785 1321 9819 1355
rect 9853 1321 9887 1355
rect 9921 1321 9955 1355
rect 9989 1321 10023 1355
rect 10057 1321 10091 1355
rect 10125 1321 10159 1355
rect 10193 1321 10227 1355
rect 10261 1321 10295 1355
rect 10329 1321 10363 1355
rect 10397 1321 10431 1355
rect 10465 1321 10499 1355
rect 10533 1321 10567 1355
rect 10601 1321 10635 1355
rect 10669 1321 10703 1355
rect 10737 1321 10771 1355
rect 10805 1321 10839 1355
rect 10873 1321 10907 1355
rect 10941 1321 10975 1355
rect 11009 1321 11043 1355
rect 11077 1321 11111 1355
rect 11145 1321 11179 1355
rect 11213 1321 11247 1355
rect 11281 1321 11315 1355
rect 11349 1321 11383 1355
rect 11417 1321 11451 1355
rect 11485 1321 11519 1355
rect 11553 1321 11587 1355
rect 11621 1321 11655 1355
rect 11689 1321 11723 1355
rect 11757 1321 11791 1355
rect 11825 1321 11859 1355
rect 11893 1321 11927 1355
rect 11961 1321 11995 1355
rect 12029 1321 12063 1355
rect 12097 1321 12131 1355
rect 12165 1321 12199 1355
rect 12233 1321 12267 1355
rect 12301 1321 12335 1355
rect 12369 1321 12403 1355
rect 12437 1321 12471 1355
rect 12505 1321 12539 1355
rect 12573 1321 12607 1355
rect 12641 1321 12675 1355
rect 12709 1321 12743 1355
rect 12777 1321 12811 1355
rect 12845 1321 12879 1355
rect 12913 1321 12947 1355
rect 12981 1321 13015 1355
rect 13049 1321 13083 1355
rect 13117 1321 13151 1355
rect 13185 1321 13219 1355
rect 13253 1321 13287 1355
rect 13321 1321 13355 1355
rect 13389 1321 13423 1355
rect 13457 1321 13491 1355
rect 13525 1321 13559 1355
rect 13593 1321 13627 1355
rect 13661 1321 13695 1355
rect 13729 1321 13763 1355
rect 13797 1321 13831 1355
rect 13865 1321 13899 1355
rect 13933 1321 13967 1355
rect 14001 1321 14035 1355
rect 14069 1321 14103 1355
rect 14137 1321 14171 1355
rect 14205 1321 14239 1355
rect 14273 1321 14307 1355
rect 14341 1321 14375 1355
rect 14409 1321 14443 1355
rect 14477 1321 14511 1355
rect 14545 1321 14579 1355
rect 14613 1321 14647 1355
rect 14681 1321 14715 1355
rect 14749 1321 14783 1355
rect 14817 1321 14851 1355
rect 14885 1321 14919 1355
rect 14953 1321 14987 1355
rect 15021 1321 15055 1355
rect 15089 1321 15123 1355
rect 15157 1321 15191 1355
rect 15225 1321 15259 1355
rect 15293 1321 15327 1355
rect 15361 1321 15395 1355
rect 15429 1321 15463 1355
rect 15497 1321 15531 1355
rect 15565 1321 15599 1355
rect 15633 1321 15667 1355
rect 15701 1321 15735 1355
rect 15769 1321 15803 1355
rect 15837 1321 15871 1355
rect 15905 1321 15939 1355
rect 15973 1321 16007 1355
rect 16041 1321 16075 1355
rect 16109 1321 16143 1355
rect 16177 1321 16211 1355
rect 16245 1321 16279 1355
rect 16313 1321 16347 1355
rect 16381 1321 16415 1355
rect 16449 1321 16483 1355
rect 16517 1321 16551 1355
rect 16585 1321 16619 1355
rect 16653 1321 16687 1355
rect 16721 1321 16755 1355
rect 16789 1321 16823 1355
rect 16857 1321 16891 1355
rect 16925 1321 16959 1355
rect 16993 1321 17027 1355
rect 17061 1321 17095 1355
rect 17129 1321 17163 1355
rect 17197 1321 17231 1355
rect 17265 1321 17299 1355
rect 17333 1321 17367 1355
rect 17401 1321 17435 1355
rect 17469 1321 17503 1355
rect 17537 1321 17571 1355
rect 17605 1321 17639 1355
rect 17673 1321 17707 1355
rect 17741 1321 17775 1355
rect 17809 1321 17843 1355
rect 17877 1321 17911 1355
rect 17945 1321 17979 1355
rect 18013 1321 18047 1355
rect 18081 1321 18115 1355
rect 18149 1321 18183 1355
rect 18217 1321 18251 1355
rect 18285 1321 18319 1355
rect 18353 1321 18387 1355
rect 18421 1321 18455 1355
rect 18489 1321 18523 1355
rect 18557 1321 18591 1355
rect 18625 1321 18659 1355
rect 18693 1321 18727 1355
rect 18761 1321 18795 1355
rect 18829 1321 18897 1355
rect 18863 1248 18897 1321
rect 18863 1180 18897 1214
rect 28031 1727 28065 1761
rect 28031 1659 28065 1693
rect 28031 1591 28065 1625
rect 28031 1523 28065 1557
rect 28031 1455 28065 1489
rect 28031 1387 28065 1421
rect 28031 1319 28065 1353
rect 28031 1251 28065 1285
rect 18863 1112 18897 1146
rect 2151 -85 2185 -51
rect 18863 1044 18897 1078
rect 18863 976 18897 1010
rect 18863 908 18897 942
rect 18863 840 18897 874
rect 18863 772 18897 806
rect 18863 704 18897 738
rect 18863 636 18897 670
rect 18863 568 18897 602
rect 18863 500 18897 534
rect 18863 432 18897 466
rect 18863 364 18897 398
rect 18863 296 18897 330
rect 18863 228 18897 262
rect 2151 -234 2185 -119
rect 2151 -326 2185 -268
rect 2151 -360 2219 -326
rect 2253 -360 2287 -326
rect 2321 -360 2355 -326
rect 2389 -360 2423 -326
rect 2457 -360 2491 -326
rect 2525 -360 2559 -326
rect 2593 -360 2627 -326
rect 2661 -360 2695 -326
rect 2729 -360 2763 -326
rect 2797 -360 2831 -326
rect 2865 -360 2899 -326
rect 2933 -360 2967 -326
rect 3001 -360 3035 -326
rect 3069 -360 3103 -326
rect 3137 -360 3171 -326
rect 3205 -360 3239 -326
rect 3273 -360 3307 -326
rect 3341 -360 15632 -326
rect 574 -917 598 -883
rect 632 -917 668 -883
rect 702 -917 738 -883
rect 772 -917 808 -883
rect 842 -917 878 -883
rect 912 -917 948 -883
rect 982 -917 1019 -883
rect 1053 -917 1090 -883
rect 1124 -917 1161 -883
rect 1195 -917 1232 -883
rect 1266 -917 1303 -883
rect 1337 -917 1374 -883
rect 1408 -917 1445 -883
rect 1479 -917 1516 -883
rect 1550 -917 1574 -883
rect 15598 -1200 15632 -360
rect 18863 160 18897 194
rect 18863 92 18897 126
rect 18863 24 18897 58
rect 18863 -44 18897 -10
rect 18863 -112 18897 -78
rect 18863 -180 18897 -146
rect 18863 -248 18897 -214
rect 18863 -316 18897 -282
rect 18863 -384 18897 -350
rect 18863 -452 18897 -418
rect 18863 -520 18897 -486
rect 18863 -588 18897 -554
rect 18863 -656 18897 -622
rect 18863 -724 18897 -690
rect 18863 -792 18897 -758
rect 18863 -860 18897 -826
rect 18863 -928 18897 -894
rect 18863 -996 18897 -962
rect 18863 -1064 18897 -1030
rect 18863 -1132 18897 -1098
rect 18863 -1200 18897 -1166
rect 15598 -1234 18016 -1200
rect 18050 -1234 18096 -1200
rect 18130 -1234 18176 -1200
rect 18210 -1234 18255 -1200
rect 18289 -1234 18334 -1200
rect 18368 -1234 18413 -1200
rect 18447 -1234 18530 -1200
rect 18564 -1234 18598 -1200
rect 18632 -1234 18666 -1200
rect 18700 -1234 18734 -1200
rect 18768 -1234 18897 -1200
rect 28031 1183 28065 1217
rect 28031 1115 28065 1149
rect 28031 1047 28065 1081
rect 28031 979 28065 1013
rect 28031 911 28065 945
rect 28031 843 28065 877
rect 28031 775 28065 809
rect 28031 707 28065 741
rect 28031 639 28065 673
rect 28031 571 28065 605
rect 28031 503 28065 537
rect 28031 435 28065 469
rect 28031 367 28065 401
rect 28031 299 28065 333
rect 28031 231 28065 265
rect 28031 163 28065 197
rect 28031 95 28065 129
rect 28031 27 28065 61
rect 28031 -41 28065 -7
rect 28031 -109 28065 -75
rect 28031 -177 28065 -143
rect 28031 -245 28065 -211
rect 28031 -313 28065 -279
rect 28031 -381 28065 -347
rect 28031 -449 28065 -415
rect 28031 -517 28065 -483
rect 28031 -585 28065 -551
rect 28031 -653 28065 -619
rect 28031 -721 28065 -687
rect 28031 -789 28065 -755
rect 28031 -857 28065 -823
rect 28031 -925 28065 -891
rect 28031 -993 28065 -959
rect 28031 -1061 28065 -1027
rect 28031 -1129 28065 -1095
rect 28031 -1197 28065 -1163
rect 28031 -1265 28065 -1231
rect 28031 -1333 28065 -1299
rect 28031 -1401 28065 -1367
rect 28031 -1469 28065 -1435
rect 28031 -1537 28065 -1503
rect 28031 -1605 28065 -1571
rect 28031 -1673 28065 -1639
rect 28031 -1741 28065 -1707
rect 28031 -1809 28065 -1775
rect 28031 -1877 28065 -1843
rect 28031 -1945 28065 -1911
rect 28031 -2013 28065 -1979
rect 28031 -2081 28065 -2047
rect 28031 -2149 28065 -2115
rect 28031 -2217 28065 -2183
rect 28031 -2285 28065 -2251
rect 28031 -2353 28065 -2319
rect 574 -2432 598 -2398
rect 632 -2432 668 -2398
rect 702 -2432 738 -2398
rect 772 -2432 808 -2398
rect 842 -2432 878 -2398
rect 912 -2432 948 -2398
rect 982 -2432 1019 -2398
rect 1053 -2432 1090 -2398
rect 1124 -2432 1161 -2398
rect 1195 -2432 1232 -2398
rect 1266 -2432 1303 -2398
rect 1337 -2432 1374 -2398
rect 1408 -2432 1445 -2398
rect 1479 -2432 1516 -2398
rect 1550 -2432 1574 -2398
rect 28031 -2421 28065 -2387
rect 28031 -2489 28065 -2455
rect 28031 -2557 28065 -2523
rect 28031 -2625 28065 -2591
rect 28031 -2693 28065 -2659
rect 28031 -2761 28065 -2727
rect 28031 -2829 28065 -2795
rect 28031 -2897 28065 -2863
rect 28031 -2965 28065 -2931
rect 28031 -3033 28065 -2999
rect 28031 -3101 28065 -3067
rect 28031 -3169 28065 -3135
rect 28031 -3237 28065 -3203
rect 28031 -3305 28065 -3271
rect 28031 -3373 28065 -3339
rect 28031 -3441 28065 -3407
rect 28031 -3509 28065 -3475
rect 28031 -3577 28065 -3543
rect 28031 -3645 28065 -3611
rect 28031 -3713 28065 -3679
rect 28031 -3781 28065 -3747
rect 28031 -3849 28065 -3815
rect 28031 -3917 28065 -3883
rect 28031 -3985 28065 -3951
rect 28031 -4053 28065 -4019
rect 28031 -4121 28065 -4087
rect 28031 -4189 28065 -4155
rect 28031 -4257 28065 -4223
rect 28031 -4325 28065 -4291
rect 28031 -4393 28065 -4359
rect 28031 -4461 28065 -4427
rect 28031 -4529 28065 -4495
rect 28031 -4597 28065 -4563
rect 28031 -4665 28065 -4631
rect 28031 -4733 28065 -4699
rect 28031 -4801 28065 -4767
rect 28031 -4869 28065 -4835
rect 28031 -4937 28065 -4903
rect 28031 -5005 28065 -4971
rect 28031 -5073 28065 -5039
rect 28031 -5141 28065 -5107
rect 28031 -5209 28065 -5175
rect 28031 -5277 28065 -5243
rect 28031 -5345 28065 -5311
rect 28031 -5413 28065 -5379
rect 28031 -5481 28065 -5447
rect 28031 -5549 28065 -5515
rect 28031 -5617 28065 -5583
rect 28031 -5685 28065 -5651
rect 28031 -5753 28065 -5719
rect 28031 -5821 28065 -5787
rect 28031 -5889 28065 -5855
rect 28031 -5957 28065 -5923
rect 28031 -6025 28065 -5991
rect 28031 -6093 28065 -6059
rect 28031 -6161 28065 -6127
rect 28031 -6229 28065 -6195
rect 28031 -6297 28065 -6263
rect 28031 -6365 28065 -6331
rect 28031 -6433 28065 -6399
rect 28031 -6501 28065 -6467
rect 28031 -6569 28065 -6535
rect 28031 -6637 28065 -6603
rect 28031 -6705 28065 -6671
rect 28031 -6773 28065 -6739
rect 28031 -6841 28065 -6807
rect 28031 -6909 28065 -6875
rect 28031 -6977 28065 -6943
rect 28031 -7045 28065 -7011
rect 28031 -7113 28065 -7079
rect 28031 -7181 28065 -7147
rect 28031 -7249 28065 -7215
rect 28031 -7317 28065 -7283
rect 28031 -7385 28065 -7351
rect 28031 -7453 28065 -7419
rect 28031 -7521 28065 -7487
rect 28031 -7589 28065 -7555
rect 28031 -7657 28065 -7623
rect 28031 -7725 28065 -7691
rect 28031 -7793 28065 -7759
rect 28031 -7861 28065 -7827
rect 28031 -7929 28065 -7895
rect 28031 -7997 28065 -7963
rect 28031 -8065 28065 -8031
rect 28031 -8133 28065 -8099
rect 28031 -8201 28065 -8167
rect 28031 -8269 28065 -8235
rect 28031 -8337 28065 -8303
rect 28031 -8405 28065 -8371
rect 28031 -8473 28065 -8439
rect 28031 -8541 28065 -8507
rect 28031 -8609 28065 -8575
rect 28031 -8677 28065 -8643
rect 28031 -8745 28065 -8711
rect 28031 -8813 28065 -8779
rect 28031 -8881 28065 -8847
rect 28031 -8949 28065 -8915
rect 28031 -9017 28065 -8983
rect 28031 -9085 28065 -9051
rect 28031 -9153 28065 -9119
rect 28031 -9221 28065 -9187
rect 28031 -9289 28065 -9255
rect 28031 -9357 28065 -9323
rect 28031 -9425 28065 -9391
rect 28031 -9493 28065 -9459
rect 28031 -9561 28065 -9527
rect 28031 -9629 28065 -9595
rect 28031 -9697 28065 -9663
rect 28031 -9765 28065 -9731
rect 28031 -9833 28065 -9799
rect 28031 -9901 28065 -9867
rect 28031 -9969 28065 -9935
rect 28031 -10037 28065 -10003
rect 28031 -10105 28065 -10071
rect 28031 -10173 28065 -10139
rect 23953 -10608 24053 -10201
rect 28031 -10241 28065 -10207
rect 28031 -10309 28065 -10275
rect 28031 -10377 28065 -10343
rect 28031 -10445 28065 -10411
rect 28031 -10608 28065 -10479
rect 23953 -10642 23987 -10608
rect 24021 -10642 24055 -10608
rect 24089 -10642 24123 -10608
rect 24157 -10642 24191 -10608
rect 24225 -10642 24259 -10608
rect 24293 -10642 24327 -10608
rect 24361 -10642 24395 -10608
rect 24429 -10642 24463 -10608
rect 24497 -10642 24531 -10608
rect 24565 -10642 24599 -10608
rect 24633 -10642 24667 -10608
rect 24701 -10642 24735 -10608
rect 24769 -10642 24803 -10608
rect 24837 -10642 24871 -10608
rect 24905 -10642 24939 -10608
rect 24973 -10642 25007 -10608
rect 25041 -10642 25075 -10608
rect 25109 -10642 25143 -10608
rect 25177 -10642 25211 -10608
rect 25245 -10642 25279 -10608
rect 25313 -10642 25347 -10608
rect 25381 -10642 25415 -10608
rect 25449 -10642 25483 -10608
rect 25517 -10642 25551 -10608
rect 25585 -10642 25619 -10608
rect 25653 -10642 25687 -10608
rect 25721 -10642 25755 -10608
rect 25789 -10642 25823 -10608
rect 25857 -10642 25891 -10608
rect 25925 -10642 25959 -10608
rect 25993 -10642 26027 -10608
rect 26061 -10642 26095 -10608
rect 26129 -10642 26163 -10608
rect 26197 -10642 26231 -10608
rect 26265 -10642 26299 -10608
rect 26333 -10642 26367 -10608
rect 26401 -10642 26435 -10608
rect 26469 -10642 26503 -10608
rect 26537 -10642 26571 -10608
rect 26605 -10642 26639 -10608
rect 26673 -10642 26707 -10608
rect 26741 -10642 26775 -10608
rect 26809 -10642 26843 -10608
rect 26877 -10642 26911 -10608
rect 26945 -10642 26979 -10608
rect 27013 -10642 27047 -10608
rect 27081 -10642 27115 -10608
rect 27149 -10642 27183 -10608
rect 27217 -10642 27251 -10608
rect 27285 -10642 27319 -10608
rect 27353 -10642 27387 -10608
rect 27421 -10642 27455 -10608
rect 27489 -10642 27523 -10608
rect 27557 -10642 27591 -10608
rect 27625 -10642 27659 -10608
rect 27693 -10642 27727 -10608
rect 27761 -10642 27795 -10608
rect 27829 -10642 27863 -10608
rect 27897 -10642 27931 -10608
rect 27965 -10642 28065 -10608
<< psubdiffcont >>
rect 20252 1394 20286 1428
rect 20252 1276 20286 1310
<< nsubdiffcont >>
rect 590 4937 624 4971
rect 658 4937 692 4971
rect 726 4937 760 4971
rect 794 4937 828 4971
rect 862 4937 896 4971
rect 930 4937 964 4971
rect 998 4937 1032 4971
rect 1066 4937 1100 4971
rect 1134 4937 1168 4971
rect 1202 4937 1236 4971
rect 1270 4937 1304 4971
rect 1338 4937 1372 4971
rect 1406 4937 1440 4971
rect 1474 4937 1508 4971
rect 1542 4937 1576 4971
rect 1610 4937 1644 4971
rect 1678 4937 1712 4971
rect 1746 4937 1780 4971
rect 1814 4937 1848 4971
rect 1882 4937 1916 4971
rect 1950 4937 1984 4971
rect 2018 4937 2052 4971
rect 2086 4937 2120 4971
rect 2154 4937 2188 4971
rect 2222 4937 2256 4971
rect 2290 4937 2324 4971
rect 2358 4937 2392 4971
rect 2426 4937 2460 4971
rect 2494 4937 2528 4971
rect 2562 4937 2596 4971
rect 2630 4937 2664 4971
rect 2698 4937 2732 4971
rect 2766 4937 2800 4971
rect 2834 4937 2868 4971
rect 2902 4937 2936 4971
rect 2970 4937 3004 4971
rect 3038 4937 3072 4971
rect 3106 4937 3140 4971
rect 3174 4937 3208 4971
rect 3242 4937 3276 4971
rect 3310 4937 3344 4971
rect 3378 4937 3412 4971
rect 3446 4937 3480 4971
rect 3514 4937 3548 4971
rect 3582 4937 3616 4971
rect 3650 4937 3684 4971
rect 3718 4937 3752 4971
rect 3786 4937 3820 4971
rect 3854 4937 3888 4971
rect 3922 4937 3956 4971
rect 3990 4937 4024 4971
rect 4058 4937 4092 4971
rect 4126 4937 4160 4971
rect 4194 4937 4228 4971
rect 4262 4937 4296 4971
rect 4330 4937 4364 4971
rect 4398 4937 4432 4971
rect 4466 4937 4500 4971
rect 4534 4937 4568 4971
rect 4602 4937 4636 4971
rect 4670 4937 4704 4971
rect 4738 4937 4772 4971
rect 4806 4937 4840 4971
rect 4874 4937 4908 4971
rect 4942 4937 4976 4971
rect 5010 4937 5044 4971
rect 5078 4937 5112 4971
rect 5146 4937 5180 4971
rect 5214 4937 5248 4971
rect 5282 4937 5316 4971
rect 5350 4937 5384 4971
rect 5418 4937 5452 4971
rect 5486 4937 5520 4971
rect 5554 4937 5588 4971
rect 5622 4937 5656 4971
rect 5690 4937 5724 4971
rect 5758 4937 5792 4971
rect 5826 4937 5860 4971
rect 5894 4937 5928 4971
rect 5962 4937 5996 4971
rect 6030 4937 6064 4971
rect 6098 4937 6132 4971
rect 6166 4937 6200 4971
rect 6234 4937 6268 4971
rect 6302 4937 6336 4971
rect 6370 4937 6404 4971
rect 6438 4937 6472 4971
rect 6506 4937 6540 4971
rect 6574 4937 6608 4971
rect 6642 4937 6676 4971
rect 6710 4937 6744 4971
rect 6778 4937 6812 4971
rect 6846 4937 6880 4971
rect 6914 4937 6948 4971
rect 6982 4937 7016 4971
rect 7050 4937 7084 4971
rect 7118 4937 7152 4971
rect 7186 4937 7220 4971
rect 7254 4937 7288 4971
rect 7322 4937 7356 4971
rect 7390 4937 7424 4971
rect 7458 4937 7492 4971
rect 7526 4937 7560 4971
rect 7594 4937 7628 4971
rect 7662 4937 7696 4971
rect 7730 4937 7764 4971
rect 522 4862 556 4896
rect 522 4794 556 4828
rect 593 4827 627 4861
rect 679 4827 713 4861
rect 7838 4869 7872 4903
rect 522 4726 556 4760
rect 593 4757 627 4791
rect 679 4757 713 4791
rect 522 4658 556 4692
rect 593 4687 627 4721
rect 679 4687 713 4721
rect 7838 4801 7872 4835
rect 7838 4733 7872 4767
rect 522 4590 556 4624
rect 593 4617 627 4651
rect 679 4617 713 4651
rect 7838 4665 7872 4699
rect 522 4522 556 4556
rect 593 4547 627 4581
rect 679 4547 713 4581
rect 522 4454 556 4488
rect 593 4477 627 4511
rect 679 4477 713 4511
rect 7838 4597 7872 4631
rect 7838 4529 7872 4563
rect 522 4386 556 4420
rect 593 4407 627 4441
rect 679 4407 713 4441
rect 7838 4461 7872 4495
rect 522 4318 556 4352
rect 593 4337 627 4371
rect 679 4337 713 4371
rect 522 4250 556 4284
rect 593 4267 627 4301
rect 679 4267 713 4301
rect 7838 4393 7872 4427
rect 7838 4325 7872 4359
rect 522 4182 556 4216
rect 593 4197 627 4231
rect 679 4197 713 4231
rect 522 4114 556 4148
rect 593 4127 627 4161
rect 679 4127 713 4161
rect 522 4046 556 4080
rect 593 4056 627 4090
rect 679 4056 713 4090
rect 522 3978 556 4012
rect 593 3985 627 4019
rect 679 3985 713 4019
rect 522 3910 556 3944
rect 593 3914 627 3948
rect 679 3914 713 3948
rect 522 3842 556 3876
rect 593 3843 627 3877
rect 679 3843 713 3877
rect 7838 4257 7872 4291
rect 7838 4189 7872 4223
rect 7838 4121 7872 4155
rect 7838 4053 7872 4087
rect 7838 3985 7872 4019
rect 7838 3917 7872 3951
rect 7838 3849 7872 3883
rect 522 3774 556 3808
rect 593 3772 627 3806
rect 679 3772 713 3806
rect 522 3706 556 3740
rect 593 3701 627 3735
rect 679 3701 713 3735
rect 7838 3781 7872 3815
rect 522 3638 556 3672
rect 593 3630 627 3664
rect 679 3630 713 3664
rect 522 3570 556 3604
rect 7838 3640 7872 3674
rect 593 3559 627 3593
rect 679 3559 713 3593
rect 522 3502 556 3536
rect 593 3488 627 3522
rect 679 3488 713 3522
rect 7838 3572 7872 3606
rect 7838 3504 7872 3538
rect 522 3434 556 3468
rect 593 3417 627 3451
rect 679 3417 713 3451
rect 522 3366 556 3400
rect 7838 3436 7872 3470
rect 593 3346 627 3380
rect 679 3346 713 3380
rect 522 3298 556 3332
rect 593 3275 627 3309
rect 679 3275 713 3309
rect 7838 3368 7872 3402
rect 7838 3300 7872 3334
rect 522 3230 556 3264
rect 593 3204 627 3238
rect 679 3204 713 3238
rect 522 3162 556 3196
rect 7838 3232 7872 3266
rect 7838 3164 7872 3198
rect 630 3094 664 3128
rect 698 3094 732 3128
rect 766 3094 800 3128
rect 834 3094 868 3128
rect 902 3094 936 3128
rect 970 3094 1004 3128
rect 1038 3094 1072 3128
rect 1106 3094 1140 3128
rect 1174 3094 1208 3128
rect 1242 3094 1276 3128
rect 1310 3094 1344 3128
rect 1378 3094 1412 3128
rect 1446 3094 1480 3128
rect 1514 3094 1548 3128
rect 1582 3094 1616 3128
rect 1650 3094 1684 3128
rect 1718 3094 1752 3128
rect 1786 3094 1820 3128
rect 1854 3094 1888 3128
rect 1922 3094 1956 3128
rect 1990 3094 2024 3128
rect 2058 3094 2092 3128
rect 2126 3094 2160 3128
rect 2194 3094 2228 3128
rect 2262 3094 2296 3128
rect 2330 3094 2364 3128
rect 2398 3094 2432 3128
rect 2466 3094 2500 3128
rect 2534 3094 2568 3128
rect 2602 3094 2636 3128
rect 2670 3094 2704 3128
rect 2738 3094 2772 3128
rect 2806 3094 2840 3128
rect 2874 3094 2908 3128
rect 2942 3094 2976 3128
rect 3010 3094 3044 3128
rect 3078 3094 3112 3128
rect 3146 3094 3180 3128
rect 3214 3094 3248 3128
rect 3282 3094 3316 3128
rect 3350 3094 3384 3128
rect 3418 3094 3452 3128
rect 3486 3094 3520 3128
rect 3554 3094 3588 3128
rect 3622 3094 3656 3128
rect 3690 3094 3724 3128
rect 3758 3094 3792 3128
rect 3826 3094 3860 3128
rect 3894 3094 3928 3128
rect 3962 3094 3996 3128
rect 4030 3094 4064 3128
rect 4098 3094 4132 3128
rect 4166 3094 4200 3128
rect 4234 3094 4268 3128
rect 4302 3094 4336 3128
rect 4370 3094 4404 3128
rect 4438 3094 4472 3128
rect 4506 3094 4540 3128
rect 4574 3094 4608 3128
rect 4642 3094 4676 3128
rect 4710 3094 4744 3128
rect 4778 3094 4812 3128
rect 4846 3094 4880 3128
rect 4914 3094 4948 3128
rect 4982 3094 5016 3128
rect 5050 3094 5084 3128
rect 5118 3094 5152 3128
rect 5186 3094 5220 3128
rect 5254 3094 5288 3128
rect 5322 3094 5356 3128
rect 5390 3094 5424 3128
rect 5458 3094 5492 3128
rect 5526 3094 5560 3128
rect 5594 3094 5628 3128
rect 5662 3094 5696 3128
rect 5730 3094 5764 3128
rect 5798 3094 5832 3128
rect 5866 3094 5900 3128
rect 5934 3094 5968 3128
rect 6002 3094 6036 3128
rect 6070 3094 6104 3128
rect 6138 3094 6172 3128
rect 6206 3094 6240 3128
rect 6274 3094 6308 3128
rect 6342 3094 6376 3128
rect 6410 3094 6444 3128
rect 6478 3094 6512 3128
rect 6546 3094 6580 3128
rect 6614 3094 6648 3128
rect 6682 3094 6716 3128
rect 6750 3094 6784 3128
rect 6818 3094 6852 3128
rect 6886 3094 6920 3128
rect 6954 3094 6988 3128
rect 7022 3094 7056 3128
rect 7090 3094 7124 3128
rect 7158 3094 7192 3128
rect 7226 3094 7260 3128
rect 7294 3094 7328 3128
rect 7362 3094 7396 3128
rect 7430 3094 7464 3128
rect 7498 3094 7532 3128
rect 7566 3094 7600 3128
rect 7634 3094 7668 3128
rect 7702 3094 7736 3128
rect 7770 3094 7804 3128
<< mvpsubdiffcont >>
rect 11576 3598 11610 3632
rect 11645 3598 11679 3632
rect 11714 3598 11748 3632
rect 11783 3598 11817 3632
rect 11852 3598 11886 3632
rect 11921 3598 11955 3632
rect 11990 3598 12024 3632
rect 12059 3598 12093 3632
rect 12128 3598 12162 3632
rect 12197 3598 12231 3632
rect 12266 3598 12300 3632
rect 12335 3598 12369 3632
rect 12404 3598 12438 3632
rect 12473 3598 12507 3632
rect 12542 3598 12576 3632
rect 12611 3598 12645 3632
rect 12680 3598 12714 3632
rect 12749 3598 12783 3632
rect 12818 3598 12852 3632
rect 12887 3598 12921 3632
rect 12956 3598 12990 3632
rect 13025 3598 13059 3632
rect 13094 3598 13128 3632
rect 13163 3598 13197 3632
rect 13232 3598 13266 3632
rect 13301 3598 13335 3632
rect 13370 3598 13404 3632
rect 13439 3598 13473 3632
rect 13508 3598 13542 3632
rect 13577 3598 13611 3632
rect 13646 3598 13680 3632
rect 13715 3598 13749 3632
rect 13784 3598 13818 3632
rect 13853 3598 13887 3632
rect 13922 3598 13956 3632
rect 13991 3598 14025 3632
rect 14059 3598 14093 3632
rect 14127 3598 14161 3632
rect 14195 3598 14229 3632
rect 14263 3598 14297 3632
rect 14331 3598 14365 3632
rect 14399 3598 14433 3632
rect 14467 3598 14501 3632
rect 14535 3598 14569 3632
rect 14603 3598 14637 3632
rect 14671 3598 14705 3632
rect 14739 3598 14773 3632
rect 14807 3598 14841 3632
rect 14875 3598 14909 3632
rect 14943 3598 14977 3632
rect 15011 3598 15045 3632
rect 15079 3598 15113 3632
rect 15147 3598 15181 3632
rect 15215 3598 15249 3632
rect 15283 3598 15317 3632
rect 15351 3598 15385 3632
rect 15419 3598 15453 3632
rect 15487 3598 15521 3632
rect 15555 3598 15589 3632
rect 15623 3598 15657 3632
rect 15691 3598 15725 3632
rect 15759 3598 15793 3632
rect 15827 3598 15861 3632
rect 15895 3598 15929 3632
rect 15963 3598 15997 3632
rect 16031 3598 16065 3632
rect 16099 3598 16133 3632
rect 16167 3598 16201 3632
rect 16235 3598 16269 3632
rect 16303 3598 16337 3632
rect 16371 3598 16405 3632
rect 16439 3598 16473 3632
rect 16507 3598 16541 3632
rect 16575 3598 16609 3632
rect 16643 3598 16677 3632
rect 16711 3598 16745 3632
rect 16779 3598 16813 3632
rect 16847 3598 16881 3632
rect 16915 3598 16949 3632
rect 16983 3598 17017 3632
rect 17051 3598 17085 3632
rect 17119 3598 17153 3632
rect 17187 3598 17221 3632
rect 17255 3598 17289 3632
rect 17323 3598 17357 3632
rect 17391 3598 17425 3632
rect 17459 3598 17493 3632
rect 17527 3598 17561 3632
rect 17595 3598 17629 3632
rect 17663 3598 17697 3632
rect 17731 3598 17765 3632
rect 17799 3598 17833 3632
rect 17867 3598 17901 3632
rect 17935 3598 17969 3632
rect 18003 3598 18037 3632
rect 18071 3598 18105 3632
rect 18139 3598 18173 3632
rect 18207 3598 18241 3632
rect 18275 3598 18309 3632
rect 18343 3598 18377 3632
rect 18411 3598 18445 3632
rect 18479 3598 18513 3632
rect 18547 3598 18581 3632
rect 18615 3598 18649 3632
rect 18683 3598 18717 3632
rect 18751 3598 18785 3632
rect 18819 3598 18853 3632
rect 18887 3598 18921 3632
rect 18955 3598 18989 3632
rect 19023 3598 19057 3632
rect 19091 3598 19125 3632
rect 19159 3598 19193 3632
rect 19227 3598 19261 3632
rect 19295 3598 19329 3632
rect 19363 3598 19397 3632
rect 19431 3598 19465 3632
rect 19499 3598 19533 3632
rect 19567 3598 19601 3632
rect 19635 3598 19669 3632
rect 19703 3598 19737 3632
rect 10562 2821 10596 2855
rect 10630 2821 10664 2855
rect 10698 2821 10732 2855
rect 10766 2821 10800 2855
rect 10834 2821 10868 2855
rect 10902 2821 10936 2855
rect 10970 2821 11004 2855
rect 11038 2821 11072 2855
rect 11106 2821 11140 2855
rect 11174 2821 11208 2855
rect 11242 2821 11276 2855
rect 11310 2821 11344 2855
rect 11378 2821 11412 2855
rect 11446 2821 11480 2855
rect 11514 2821 11548 2855
rect 11582 2821 11616 2855
rect 11650 2821 11684 2855
rect 11718 2821 11752 2855
rect 11786 2821 11820 2855
rect 11854 2821 11888 2855
rect 11922 2821 11956 2855
rect 11990 2821 12024 2855
rect 12058 2821 12092 2855
rect 12126 2821 12160 2855
rect 12194 2821 12228 2855
rect 12262 2821 12296 2855
rect 12330 2821 12364 2855
rect 12398 2821 12432 2855
rect 12466 2821 12500 2855
rect 12534 2821 12568 2855
rect 12602 2821 12636 2855
rect 12670 2821 12704 2855
rect 12738 2821 12772 2855
rect 12806 2821 12840 2855
rect 12874 2821 12908 2855
rect 12942 2821 12976 2855
rect 13010 2821 13044 2855
rect 13078 2821 13112 2855
rect 13146 2821 13180 2855
rect 13214 2821 13248 2855
rect 13282 2821 13316 2855
rect 13350 2821 13384 2855
rect 13418 2821 13452 2855
rect 13486 2821 13520 2855
rect 13554 2821 13588 2855
rect 13622 2821 13656 2855
rect 13690 2821 13724 2855
rect 13758 2821 13792 2855
rect 13826 2821 13860 2855
rect 13894 2821 13928 2855
rect 13962 2821 13996 2855
rect 14030 2821 14064 2855
rect 14098 2821 14132 2855
rect 14166 2821 14200 2855
rect 14234 2821 14268 2855
rect 14302 2821 14336 2855
rect 14370 2821 14404 2855
rect 14438 2821 14472 2855
rect 14506 2821 14540 2855
rect 14574 2821 14608 2855
rect 14642 2821 14676 2855
rect 14710 2821 14744 2855
rect 14778 2821 14812 2855
rect 14846 2821 14880 2855
rect 14914 2821 14948 2855
rect 14982 2821 15016 2855
rect 15050 2821 15084 2855
rect 15118 2821 15152 2855
rect 15186 2821 15220 2855
rect 15254 2821 15288 2855
rect 15322 2821 15356 2855
rect 15390 2821 15424 2855
rect 15458 2821 15492 2855
rect 15526 2821 15560 2855
rect 15594 2821 15628 2855
rect 15662 2821 15696 2855
rect 15730 2821 15764 2855
rect 15798 2821 15832 2855
rect 15866 2821 15900 2855
rect 15934 2821 15968 2855
rect 16002 2821 16036 2855
rect 16070 2821 16104 2855
rect 16138 2821 16172 2855
rect 16206 2821 16240 2855
rect 16274 2821 16308 2855
rect 16342 2821 16376 2855
rect 9723 2744 9757 2778
rect 9795 2744 9829 2778
rect 9867 2744 9901 2778
rect 9939 2744 9973 2778
rect 10011 2744 10045 2778
rect 10083 2744 10117 2778
rect 10155 2744 10189 2778
rect 10227 2744 10261 2778
rect 10299 2744 10333 2778
rect 10371 2744 10405 2778
rect 9723 2671 9757 2705
rect 9795 2671 9829 2705
rect 9867 2671 9901 2705
rect 9939 2671 9973 2705
rect 10011 2671 10045 2705
rect 10083 2671 10117 2705
rect 10155 2671 10189 2705
rect 10227 2671 10261 2705
rect 10299 2671 10333 2705
rect 10371 2671 10405 2705
rect 9723 2598 9757 2632
rect 9795 2598 9829 2632
rect 9867 2598 9901 2632
rect 9939 2598 9973 2632
rect 10011 2598 10045 2632
rect 10083 2598 10117 2632
rect 10155 2598 10189 2632
rect 10227 2598 10261 2632
rect 10299 2598 10333 2632
rect 10371 2598 10405 2632
rect 9723 2524 9757 2558
rect 9795 2524 9829 2558
rect 9867 2524 9901 2558
rect 9939 2524 9973 2558
rect 10011 2524 10045 2558
rect 10083 2524 10117 2558
rect 10155 2524 10189 2558
rect 10227 2524 10261 2558
rect 10299 2524 10333 2558
rect 10371 2524 10405 2558
rect 2452 2219 2486 2253
rect 2521 2219 2555 2253
rect 2590 2219 2624 2253
rect 2659 2219 2693 2253
rect 2728 2219 2762 2253
rect 2797 2219 2831 2253
rect 2866 2219 2900 2253
rect 2935 2219 2969 2253
rect 3004 2219 3038 2253
rect 3073 2219 3107 2253
rect 3142 2219 3176 2253
rect 3211 2219 3245 2253
rect 3280 2219 3314 2253
rect 3349 2219 3383 2253
rect 3418 2219 3452 2253
rect 3487 2219 3521 2253
rect 3556 2219 3590 2253
rect 3625 2219 3659 2253
rect 3694 2219 3728 2253
rect 3762 2219 3796 2253
rect 3830 2219 3864 2253
rect 3898 2219 3932 2253
rect 3966 2219 4000 2253
rect 4034 2219 4068 2253
rect 4102 2219 4136 2253
rect 4170 2219 4204 2253
rect 4238 2219 4272 2253
rect 4306 2219 4340 2253
rect 4374 2219 4408 2253
rect 4442 2219 4476 2253
rect 4510 2219 4544 2253
rect 4578 2219 4612 2253
rect 4646 2219 4680 2253
rect 4714 2219 4748 2253
rect 4782 2219 4816 2253
rect 4850 2219 4884 2253
rect 4918 2219 4952 2253
rect 4986 2219 5020 2253
rect 5054 2219 5088 2253
rect 5122 2219 5156 2253
rect 5190 2219 5224 2253
rect 5258 2219 5292 2253
rect 5326 2219 5360 2253
rect 5394 2219 5428 2253
rect 5462 2219 5496 2253
rect 5530 2219 5564 2253
rect 5598 2219 5632 2253
rect 5666 2219 5700 2253
rect 5734 2219 5768 2253
rect 5802 2219 5836 2253
rect 5870 2219 5904 2253
rect 5938 2219 5972 2253
rect 6006 2219 6040 2253
rect 6074 2219 6108 2253
rect 6142 2219 6176 2253
rect 6210 2219 6244 2253
rect 6278 2219 6312 2253
rect 6346 2219 6380 2253
rect 6414 2219 6448 2253
rect 6482 2219 6516 2253
rect 6550 2219 6584 2253
rect 6618 2219 6652 2253
rect 6686 2219 6720 2253
rect 6754 2219 6788 2253
rect 6822 2219 6856 2253
rect 6890 2219 6924 2253
rect 6958 2219 6992 2253
rect 9723 2450 9757 2484
rect 9795 2450 9829 2484
rect 9867 2450 9901 2484
rect 9939 2450 9973 2484
rect 10011 2450 10045 2484
rect 10083 2450 10117 2484
rect 10155 2450 10189 2484
rect 10227 2450 10261 2484
rect 10299 2450 10333 2484
rect 10371 2450 10405 2484
rect 9723 2376 9757 2410
rect 9795 2376 9829 2410
rect 9867 2376 9901 2410
rect 9939 2376 9973 2410
rect 10011 2376 10045 2410
rect 10083 2376 10117 2410
rect 10155 2376 10189 2410
rect 10227 2376 10261 2410
rect 10299 2376 10333 2410
rect 10371 2376 10405 2410
rect 9723 2302 9757 2336
rect 9795 2302 9829 2336
rect 9867 2302 9901 2336
rect 9939 2302 9973 2336
rect 10011 2302 10045 2336
rect 10083 2302 10117 2336
rect 10155 2302 10189 2336
rect 10227 2302 10261 2336
rect 10299 2302 10333 2336
rect 10371 2302 10405 2336
rect 9723 2228 9757 2262
rect 9795 2228 9829 2262
rect 9867 2228 9901 2262
rect 9939 2228 9973 2262
rect 10011 2228 10045 2262
rect 10083 2228 10117 2262
rect 10155 2228 10189 2262
rect 10227 2228 10261 2262
rect 10299 2228 10333 2262
rect 10371 2228 10405 2262
rect 9723 2154 9757 2188
rect 9795 2154 9829 2188
rect 9867 2154 9901 2188
rect 9939 2154 9973 2188
rect 10011 2154 10045 2188
rect 10083 2154 10117 2188
rect 10155 2154 10189 2188
rect 10227 2154 10261 2188
rect 10299 2154 10333 2188
rect 10371 2154 10405 2188
rect 9723 2080 9757 2114
rect 9795 2080 9829 2114
rect 9867 2080 9901 2114
rect 9939 2080 9973 2114
rect 10011 2080 10045 2114
rect 10083 2080 10117 2114
rect 10155 2080 10189 2114
rect 10227 2080 10261 2114
rect 10299 2080 10333 2114
rect 10371 2080 10405 2114
rect 9723 2006 9757 2040
rect 9795 2006 9829 2040
rect 9867 2006 9901 2040
rect 9939 2006 9973 2040
rect 10011 2006 10045 2040
rect 10083 2006 10117 2040
rect 10155 2006 10189 2040
rect 10227 2006 10261 2040
rect 10299 2006 10333 2040
rect 10371 2006 10405 2040
rect 10488 2753 10522 2787
rect 10488 2685 10522 2719
rect 10488 2617 10522 2651
rect 10488 2549 10522 2583
rect 10488 2481 10522 2515
rect 10488 2323 10522 2357
rect 16410 2693 16444 2727
rect 16410 2625 16444 2659
rect 16410 2557 16444 2591
rect 16410 2489 16444 2523
rect 16410 2421 16444 2455
rect 10488 2255 10522 2289
rect 10488 2187 10522 2221
rect 10488 2119 10522 2153
rect 16410 2353 16444 2387
rect 16410 2285 16444 2319
rect 16410 2217 16444 2251
rect 16410 2149 16444 2183
rect 16410 2081 16444 2115
rect 10556 2013 10590 2047
rect 10624 2013 10658 2047
rect 10692 2013 10726 2047
rect 10760 2013 10794 2047
rect 10828 2013 10862 2047
rect 10896 2013 10930 2047
rect 10964 2013 10998 2047
rect 11032 2013 11066 2047
rect 11100 2013 11134 2047
rect 11168 2013 11202 2047
rect 11236 2013 11270 2047
rect 11304 2013 11338 2047
rect 11372 2013 11406 2047
rect 11440 2013 11474 2047
rect 11508 2013 11542 2047
rect 11576 2013 11610 2047
rect 11644 2013 11678 2047
rect 11712 2013 11746 2047
rect 11780 2013 11814 2047
rect 11848 2013 11882 2047
rect 11916 2013 11950 2047
rect 11984 2013 12018 2047
rect 12052 2013 12086 2047
rect 12120 2013 12154 2047
rect 12188 2013 12222 2047
rect 12256 2013 12290 2047
rect 12324 2013 12358 2047
rect 12392 2013 12426 2047
rect 12460 2013 12494 2047
rect 12528 2013 12562 2047
rect 12596 2013 12630 2047
rect 12664 2013 12698 2047
rect 12732 2013 12766 2047
rect 12800 2013 12834 2047
rect 12868 2013 12902 2047
rect 12936 2013 12970 2047
rect 13004 2013 13038 2047
rect 13072 2013 13106 2047
rect 13140 2013 13174 2047
rect 13208 2013 13242 2047
rect 13276 2013 13310 2047
rect 13344 2013 13378 2047
rect 13412 2013 13446 2047
rect 13480 2013 13514 2047
rect 13548 2013 13582 2047
rect 13616 2013 13650 2047
rect 13684 2013 13718 2047
rect 13752 2013 13786 2047
rect 13820 2013 13854 2047
rect 13888 2013 13922 2047
rect 13956 2013 13990 2047
rect 14024 2013 14058 2047
rect 14092 2013 14126 2047
rect 14160 2013 14194 2047
rect 14228 2013 14262 2047
rect 14296 2013 14330 2047
rect 14364 2013 14398 2047
rect 14432 2013 14466 2047
rect 14500 2013 14534 2047
rect 14568 2013 14602 2047
rect 14636 2013 14670 2047
rect 14704 2013 14738 2047
rect 14772 2013 14806 2047
rect 14840 2013 14874 2047
rect 14908 2013 14942 2047
rect 14976 2013 15010 2047
rect 15044 2013 15078 2047
rect 15112 2013 15146 2047
rect 15180 2013 15214 2047
rect 15248 2013 15282 2047
rect 15316 2013 15350 2047
rect 15384 2013 15418 2047
rect 15452 2013 15486 2047
rect 15520 2013 15554 2047
rect 15588 2013 15622 2047
rect 15656 2013 15690 2047
rect 15724 2013 15758 2047
rect 15792 2013 15826 2047
rect 15860 2013 15894 2047
rect 15928 2013 15962 2047
rect 15996 2013 16030 2047
rect 16064 2013 16098 2047
rect 16132 2013 16166 2047
rect 16200 2013 16234 2047
rect 16268 2013 16302 2047
rect 16336 2013 16370 2047
rect 16563 2070 19045 2376
rect 19079 2259 19113 2293
rect 19152 2259 19186 2293
rect 19225 2259 19259 2293
rect 19298 2259 19332 2293
rect 19371 2259 19405 2293
rect 19444 2259 19478 2293
rect 19517 2259 19551 2293
rect 19079 2185 19113 2219
rect 19152 2185 19186 2219
rect 19225 2185 19259 2219
rect 19298 2185 19332 2219
rect 19371 2185 19405 2219
rect 19444 2185 19478 2219
rect 19517 2185 19551 2219
rect 19079 2111 19113 2145
rect 19152 2111 19186 2145
rect 19225 2111 19259 2145
rect 19298 2111 19332 2145
rect 19371 2111 19405 2145
rect 19444 2111 19478 2145
rect 19517 2111 19551 2145
rect 19079 2037 19113 2071
rect 19152 2037 19186 2071
rect 19225 2037 19259 2071
rect 19298 2037 19332 2071
rect 19371 2037 19405 2071
rect 19444 2037 19478 2071
rect 19517 2037 19551 2071
rect 9723 1932 9757 1966
rect 9795 1932 9829 1966
rect 9867 1932 9901 1966
rect 9939 1932 9973 1966
rect 10011 1932 10045 1966
rect 10083 1932 10117 1966
rect 10155 1932 10189 1966
rect 10227 1932 10261 1966
rect 10299 1932 10333 1966
rect 10371 1932 10405 1966
rect 16563 2001 16597 2035
rect 16631 2001 16665 2035
rect 16699 2001 16733 2035
rect 16767 2001 16801 2035
rect 16835 2001 16869 2035
rect 16903 2001 16937 2035
rect 16971 2001 17005 2035
rect 17039 2001 17073 2035
rect 17107 2001 17141 2035
rect 17175 2001 17209 2035
rect 17243 2001 17277 2035
rect 17311 2001 17345 2035
rect 17379 2001 17413 2035
rect 17447 2001 17481 2035
rect 17515 2001 17549 2035
rect 17583 2001 17617 2035
rect 17651 2001 17685 2035
rect 17719 2001 17753 2035
rect 17787 2001 17821 2035
rect 17855 2001 17889 2035
rect 17923 2001 17957 2035
rect 17991 2001 18025 2035
rect 18059 2001 18093 2035
rect 18127 2001 18161 2035
rect 18195 2001 18229 2035
rect 18263 2001 18297 2035
rect 18331 2001 18365 2035
rect 18399 2001 18433 2035
rect 18467 2001 18501 2035
rect 18535 2001 18569 2035
rect 18603 2001 18637 2035
rect 18671 2001 18705 2035
rect 18739 2001 18773 2035
rect 18807 2001 18841 2035
rect 18875 2001 18909 2035
rect 18943 2001 18977 2035
rect 19011 2001 19045 2035
rect 16563 1932 19045 1966
rect 19079 1963 19113 1997
rect 19152 1963 19186 1997
rect 19225 1963 19259 1997
rect 19298 1963 19332 1997
rect 19371 1963 19405 1997
rect 19444 1963 19478 1997
rect 19517 1963 19551 1997
rect 16563 1898 19011 1932
rect 9750 1864 9784 1898
rect 9819 1864 9853 1898
rect 9888 1864 9922 1898
rect 9957 1864 9991 1898
rect 10026 1864 10060 1898
rect 10095 1864 10129 1898
rect 10164 1864 10198 1898
rect 10233 1864 10267 1898
rect 10302 1864 10336 1898
rect 10371 1864 10405 1898
rect 10440 1864 10474 1898
rect 10509 1864 10543 1898
rect 10578 1864 10612 1898
rect 10647 1864 10681 1898
rect 10716 1864 10750 1898
rect 10785 1864 10819 1898
rect 10854 1864 10888 1898
rect 10923 1864 10957 1898
rect 10992 1864 11026 1898
rect 11061 1864 11095 1898
rect 11130 1864 11164 1898
rect 11199 1864 11233 1898
rect 11268 1864 11302 1898
rect 11337 1864 11371 1898
rect 11406 1864 11440 1898
rect 11475 1864 11509 1898
rect 11544 1864 11578 1898
rect 11613 1864 11647 1898
rect 11682 1864 11716 1898
rect 11751 1864 11785 1898
rect 11820 1864 11854 1898
rect 11889 1864 11923 1898
rect 11958 1864 11992 1898
rect 12027 1864 12061 1898
rect 12096 1864 12130 1898
rect 12165 1864 12199 1898
rect 12234 1864 12268 1898
rect 12303 1864 12337 1898
rect 12372 1864 12406 1898
rect 12441 1864 12475 1898
rect 12510 1864 12544 1898
rect 12579 1864 12613 1898
rect 12648 1864 12682 1898
rect 12717 1864 12751 1898
rect 12786 1864 12820 1898
rect 12855 1864 12889 1898
rect 12924 1864 12958 1898
rect 9750 1796 9784 1830
rect 9819 1796 9853 1830
rect 9888 1796 9922 1830
rect 9957 1796 9991 1830
rect 10026 1796 10060 1830
rect 10095 1796 10129 1830
rect 10164 1796 10198 1830
rect 10233 1796 10267 1830
rect 10302 1796 10336 1830
rect 10371 1796 10405 1830
rect 10440 1796 10474 1830
rect 10509 1796 10543 1830
rect 10578 1796 10612 1830
rect 10647 1796 10681 1830
rect 10716 1796 10750 1830
rect 10785 1796 10819 1830
rect 10854 1796 10888 1830
rect 10923 1796 10957 1830
rect 10992 1796 11026 1830
rect 11061 1796 11095 1830
rect 11130 1796 11164 1830
rect 11199 1796 11233 1830
rect 11268 1796 11302 1830
rect 11337 1796 11371 1830
rect 11406 1796 11440 1830
rect 11475 1796 11509 1830
rect 11544 1796 11578 1830
rect 11613 1796 11647 1830
rect 11682 1796 11716 1830
rect 11751 1796 11785 1830
rect 11820 1796 11854 1830
rect 11889 1796 11923 1830
rect 11958 1796 11992 1830
rect 12027 1796 12061 1830
rect 12096 1796 12130 1830
rect 12165 1796 12199 1830
rect 12234 1796 12268 1830
rect 12303 1796 12337 1830
rect 12372 1796 12406 1830
rect 12441 1796 12475 1830
rect 12510 1796 12544 1830
rect 12579 1796 12613 1830
rect 12648 1796 12682 1830
rect 12717 1796 12751 1830
rect 12786 1796 12820 1830
rect 12855 1796 12889 1830
rect 12924 1796 12958 1830
rect 9750 1728 9784 1762
rect 9819 1728 9853 1762
rect 9888 1728 9922 1762
rect 9957 1728 9991 1762
rect 10026 1728 10060 1762
rect 10095 1728 10129 1762
rect 10164 1728 10198 1762
rect 10233 1728 10267 1762
rect 10302 1728 10336 1762
rect 10371 1728 10405 1762
rect 10440 1728 10474 1762
rect 10509 1728 10543 1762
rect 10578 1728 10612 1762
rect 10647 1728 10681 1762
rect 10716 1728 10750 1762
rect 10785 1728 10819 1762
rect 10854 1728 10888 1762
rect 10923 1728 10957 1762
rect 10992 1728 11026 1762
rect 11061 1728 11095 1762
rect 11130 1728 11164 1762
rect 11199 1728 11233 1762
rect 11268 1728 11302 1762
rect 11337 1728 11371 1762
rect 11406 1728 11440 1762
rect 11475 1728 11509 1762
rect 11544 1728 11578 1762
rect 11613 1728 11647 1762
rect 11682 1728 11716 1762
rect 11751 1728 11785 1762
rect 11820 1728 11854 1762
rect 11889 1728 11923 1762
rect 11958 1728 11992 1762
rect 12027 1728 12061 1762
rect 12096 1728 12130 1762
rect 12165 1728 12199 1762
rect 12234 1728 12268 1762
rect 12303 1728 12337 1762
rect 12372 1728 12406 1762
rect 12441 1728 12475 1762
rect 12510 1728 12544 1762
rect 12579 1728 12613 1762
rect 12648 1728 12682 1762
rect 12717 1728 12751 1762
rect 12786 1728 12820 1762
rect 12855 1728 12889 1762
rect 12924 1728 12958 1762
rect 9750 1660 9784 1694
rect 9819 1660 9853 1694
rect 9888 1660 9922 1694
rect 9957 1660 9991 1694
rect 10026 1660 10060 1694
rect 10095 1660 10129 1694
rect 10164 1660 10198 1694
rect 10233 1660 10267 1694
rect 10302 1660 10336 1694
rect 10371 1660 10405 1694
rect 10440 1660 10474 1694
rect 10509 1660 10543 1694
rect 10578 1660 10612 1694
rect 10647 1660 10681 1694
rect 10716 1660 10750 1694
rect 10785 1660 10819 1694
rect 10854 1660 10888 1694
rect 10923 1660 10957 1694
rect 10992 1660 11026 1694
rect 11061 1660 11095 1694
rect 11130 1660 11164 1694
rect 11199 1660 11233 1694
rect 11268 1660 11302 1694
rect 11337 1660 11371 1694
rect 11406 1660 11440 1694
rect 11475 1660 11509 1694
rect 11544 1660 11578 1694
rect 11613 1660 11647 1694
rect 11682 1660 11716 1694
rect 11751 1660 11785 1694
rect 11820 1660 11854 1694
rect 11889 1660 11923 1694
rect 11958 1660 11992 1694
rect 12027 1660 12061 1694
rect 12096 1660 12130 1694
rect 12165 1660 12199 1694
rect 12234 1660 12268 1694
rect 12303 1660 12337 1694
rect 12372 1660 12406 1694
rect 12441 1660 12475 1694
rect 12510 1660 12544 1694
rect 12579 1660 12613 1694
rect 12648 1660 12682 1694
rect 12717 1660 12751 1694
rect 12786 1660 12820 1694
rect 12855 1660 12889 1694
rect 12924 1660 12958 1694
rect 9750 1592 9784 1626
rect 9819 1592 9853 1626
rect 9888 1592 9922 1626
rect 9957 1592 9991 1626
rect 10026 1592 10060 1626
rect 10095 1592 10129 1626
rect 10164 1592 10198 1626
rect 10233 1592 10267 1626
rect 10302 1592 10336 1626
rect 10371 1592 10405 1626
rect 10440 1592 10474 1626
rect 10509 1592 10543 1626
rect 10578 1592 10612 1626
rect 10647 1592 10681 1626
rect 10716 1592 10750 1626
rect 10785 1592 10819 1626
rect 10854 1592 10888 1626
rect 10923 1592 10957 1626
rect 10992 1592 11026 1626
rect 11061 1592 11095 1626
rect 11130 1592 11164 1626
rect 11199 1592 11233 1626
rect 11268 1592 11302 1626
rect 11337 1592 11371 1626
rect 11406 1592 11440 1626
rect 11475 1592 11509 1626
rect 11544 1592 11578 1626
rect 11613 1592 11647 1626
rect 11682 1592 11716 1626
rect 11751 1592 11785 1626
rect 11820 1592 11854 1626
rect 11889 1592 11923 1626
rect 11958 1592 11992 1626
rect 12027 1592 12061 1626
rect 12096 1592 12130 1626
rect 12165 1592 12199 1626
rect 12234 1592 12268 1626
rect 12303 1592 12337 1626
rect 12372 1592 12406 1626
rect 12441 1592 12475 1626
rect 12510 1592 12544 1626
rect 12579 1592 12613 1626
rect 12648 1592 12682 1626
rect 12717 1592 12751 1626
rect 12786 1592 12820 1626
rect 12855 1592 12889 1626
rect 12924 1592 12958 1626
rect 12993 1592 19011 1898
rect 19079 1889 19113 1923
rect 19152 1889 19186 1923
rect 19225 1889 19259 1923
rect 19298 1889 19332 1923
rect 19371 1889 19405 1923
rect 19444 1889 19478 1923
rect 19517 1889 19551 1923
rect 19079 1815 19113 1849
rect 19152 1815 19186 1849
rect 19225 1815 19259 1849
rect 19298 1815 19332 1849
rect 19371 1815 19405 1849
rect 19444 1815 19478 1849
rect 19517 1815 19551 1849
rect 19079 1741 19113 1775
rect 19152 1741 19186 1775
rect 19225 1741 19259 1775
rect 19298 1741 19332 1775
rect 19371 1741 19405 1775
rect 19444 1741 19478 1775
rect 19517 1741 19551 1775
rect 19079 1667 19113 1701
rect 19152 1667 19186 1701
rect 19225 1667 19259 1701
rect 19298 1667 19332 1701
rect 19371 1667 19405 1701
rect 19444 1667 19478 1701
rect 19517 1667 19551 1701
rect 19079 1593 19113 1627
rect 19152 1593 19186 1627
rect 19225 1593 19259 1627
rect 19298 1593 19332 1627
rect 19371 1593 19405 1627
rect 19444 1593 19478 1627
rect 19517 1593 19551 1627
rect 25787 1727 25821 1761
rect 25787 1656 25821 1690
rect 25787 1585 25821 1619
rect 25787 1514 25821 1548
rect 25787 1442 25821 1476
rect 25787 1370 25821 1404
rect 25787 1298 25821 1332
rect 25787 1226 25821 1260
rect 8168 908 8202 942
rect 8168 836 8202 870
rect 8168 764 8202 798
rect 8168 692 8202 726
rect 8168 620 8202 654
rect 8168 548 8202 582
rect 8168 476 8202 510
rect 8168 404 8202 438
rect 8168 332 8202 366
rect 8168 260 8202 294
rect 8168 188 8202 222
rect 8168 116 8202 150
rect 8168 44 8202 78
rect 8168 -28 8202 6
rect 10604 890 10638 924
rect 10604 820 10638 854
rect 10604 750 10638 784
rect 10604 680 10638 714
rect 10604 610 10638 644
rect 10604 540 10638 574
rect 10604 469 10638 503
rect 10604 398 10638 432
rect 10604 327 10638 361
rect 10604 256 10638 290
rect 10604 185 10638 219
rect 10604 114 10638 148
rect 10604 43 10638 77
rect 10604 -28 10638 6
rect 16352 1027 16386 1061
rect 16352 940 16386 974
rect 16352 853 16386 887
rect 12678 586 12712 620
rect 16352 766 16386 800
rect 16352 679 16386 713
rect 12678 513 12712 547
rect 12678 440 12712 474
rect 12678 367 12712 401
rect 16352 592 16386 626
rect 16352 505 16386 539
rect 12678 294 12712 328
rect 12678 221 12712 255
rect 12678 148 12712 182
rect 16352 418 16386 452
rect 16352 331 16386 365
rect 12678 75 12712 109
rect 16352 244 16386 278
rect 12678 2 12712 36
rect 2422 -92 2456 -58
rect 2491 -92 2525 -58
rect 2560 -92 2594 -58
rect 2629 -92 2663 -58
rect 2698 -92 2732 -58
rect 2767 -92 2801 -58
rect 2836 -92 2870 -58
rect 2905 -92 2939 -58
rect 2974 -92 3008 -58
rect 3043 -92 3077 -58
rect 3112 -92 3146 -58
rect 3181 -92 3215 -58
rect 3250 -92 3284 -58
rect 3319 -92 3353 -58
rect 3388 -92 3422 -58
rect 3457 -92 3491 -58
rect 3526 -92 3560 -58
rect 3595 -92 3629 -58
rect 3664 -92 3698 -58
rect 3733 -92 3767 -58
rect 3802 -92 3836 -58
rect 3871 -92 3905 -58
rect 3940 -92 3974 -58
rect 4008 -92 4042 -58
rect 4076 -92 4110 -58
rect 4144 -92 4178 -58
rect 4212 -92 4246 -58
rect 4280 -92 4314 -58
rect 4348 -92 4382 -58
rect 4416 -92 4450 -58
rect 4484 -92 4518 -58
rect 4552 -92 4586 -58
rect 4620 -92 4654 -58
rect 4688 -92 4722 -58
rect 4756 -92 4790 -58
rect 4824 -92 4858 -58
rect 4892 -92 4926 -58
rect 4960 -92 4994 -58
rect 5028 -92 5062 -58
rect 5096 -92 5130 -58
rect 5164 -92 5198 -58
rect 5232 -92 5266 -58
rect 5300 -92 5334 -58
rect 5368 -92 5402 -58
rect 5436 -92 5470 -58
rect 5504 -92 5538 -58
rect 5572 -92 5606 -58
rect 5640 -92 5674 -58
rect 5708 -92 5742 -58
rect 5776 -92 5810 -58
rect 5844 -92 5878 -58
rect 5912 -92 5946 -58
rect 5980 -92 6014 -58
rect 6048 -92 6082 -58
rect 6116 -92 6150 -58
rect 6184 -92 6218 -58
rect 6252 -92 6286 -58
rect 6320 -92 6354 -58
rect 6388 -92 6422 -58
rect 6456 -92 6490 -58
rect 6524 -92 6558 -58
rect 6592 -92 6626 -58
rect 6660 -92 6694 -58
rect 6728 -92 6762 -58
rect 6796 -92 6830 -58
rect 6864 -92 6898 -58
rect 12678 -71 12712 -37
rect 13142 -71 13176 -37
rect 13211 -71 13245 -37
rect 13280 -71 13314 -37
rect 13349 -71 13383 -37
rect 13418 -71 13452 -37
rect 13486 -71 13520 -37
rect 13554 -71 13588 -37
rect 13622 -71 13656 -37
rect 13690 -71 13724 -37
rect 13758 -71 13792 -37
rect 13826 -71 13860 -37
rect 13894 -71 13928 -37
rect 13962 -71 13996 -37
rect 14030 -71 14064 -37
rect 14098 -71 14132 -37
rect 14166 -71 14200 -37
rect 14234 -71 14268 -37
rect 14302 -71 14336 -37
rect 14370 -71 14404 -37
rect 14438 -71 14472 -37
rect 14506 -71 14540 -37
rect 14574 -71 14608 -37
rect 14642 -71 14676 -37
rect 14710 -71 14744 -37
rect 14778 -71 14812 -37
rect 14846 -71 14880 -37
rect 14914 -71 14948 -37
rect 14982 -71 15016 -37
rect 15050 -71 15084 -37
rect 15118 -71 15152 -37
rect 15186 -71 15220 -37
rect 15254 -71 15288 -37
rect 15322 -71 15356 -37
rect 15390 -71 15424 -37
rect 15458 -71 15492 -37
rect 15526 -71 15560 -37
rect 15594 -71 15628 -37
rect 15662 -71 15696 -37
rect 15730 -71 15764 -37
rect 16352 157 16386 191
rect 16352 70 16386 104
rect 16352 -17 16386 17
rect 16352 -104 16386 -70
rect 16352 -191 16386 -157
rect 16352 -279 16386 -245
rect 16352 -367 16386 -333
rect 16352 -455 16386 -421
rect 16352 -543 16386 -509
rect 16352 -631 16386 -597
rect 16352 -719 16386 -685
rect 16352 -807 16386 -773
rect 16352 -895 16386 -861
rect 15898 -971 15932 -937
rect 15991 -971 16025 -937
rect 16084 -971 16118 -937
rect 16176 -971 16210 -937
rect 16268 -971 16302 -937
rect 495 -3265 529 -3231
rect 563 -3265 597 -3231
rect 631 -3265 665 -3231
rect 699 -3265 733 -3231
rect 767 -3265 801 -3231
rect 835 -3265 869 -3231
rect 903 -3265 937 -3231
rect 971 -3265 1005 -3231
rect 406 -3333 440 -3299
rect 1039 -3355 1073 -3321
rect 406 -3401 440 -3367
rect 406 -3469 440 -3435
rect 406 -3537 440 -3503
rect 406 -3605 440 -3571
rect 406 -3673 440 -3639
rect 406 -3780 440 -3746
rect 406 -3848 440 -3814
rect 406 -3916 440 -3882
rect 406 -3984 440 -3950
rect 406 -4052 440 -4018
rect 406 -4120 440 -4086
rect 406 -4188 440 -4154
rect 406 -4256 440 -4222
rect 406 -4324 440 -4290
rect 406 -4392 440 -4358
rect 406 -4460 440 -4426
rect 406 -4528 440 -4494
rect 406 -4596 440 -4562
rect 406 -4664 440 -4630
rect 406 -4732 440 -4698
rect 406 -4800 440 -4766
rect 406 -4868 440 -4834
rect 406 -4936 440 -4902
rect 406 -5004 440 -4970
rect 406 -5072 440 -5038
rect 406 -5140 440 -5106
rect 406 -5208 440 -5174
rect 406 -5276 440 -5242
rect 406 -5344 440 -5310
rect 406 -5412 440 -5378
rect 406 -5480 440 -5446
rect 406 -5548 440 -5514
rect 406 -5616 440 -5582
rect 406 -5684 440 -5650
rect 406 -5752 440 -5718
rect 406 -5820 440 -5786
rect 406 -5888 440 -5854
rect 406 -5956 440 -5922
rect 406 -6024 440 -5990
rect 406 -6092 440 -6058
rect 406 -6160 440 -6126
rect 406 -6228 440 -6194
rect 406 -6296 440 -6262
rect 406 -6364 440 -6330
rect 406 -6432 440 -6398
rect 406 -6500 440 -6466
rect 406 -6568 440 -6534
rect 406 -6636 440 -6602
rect 406 -6704 440 -6670
rect 406 -6772 440 -6738
rect 406 -6840 440 -6806
rect 406 -6908 440 -6874
rect 406 -6976 440 -6942
rect 406 -7044 440 -7010
rect 406 -7112 440 -7078
rect 406 -7180 440 -7146
rect 406 -7248 440 -7214
rect 406 -7316 440 -7282
rect 406 -7384 440 -7350
rect 406 -7452 440 -7418
rect 406 -7520 440 -7486
rect 406 -7588 440 -7554
rect 406 -7656 440 -7622
rect 406 -7724 440 -7690
rect 406 -7792 440 -7758
rect 406 -7860 440 -7826
rect 406 -7928 440 -7894
rect 406 -7996 440 -7962
rect 406 -8064 440 -8030
rect 406 -8132 440 -8098
rect 406 -8200 440 -8166
rect 406 -8268 440 -8234
rect 406 -8336 440 -8302
rect 406 -8404 440 -8370
rect 406 -8472 440 -8438
rect 406 -8540 440 -8506
rect 406 -8608 440 -8574
rect 406 -8676 440 -8642
rect 406 -8744 440 -8710
rect 406 -8812 440 -8778
rect 406 -8880 440 -8846
rect 406 -8948 440 -8914
rect 406 -9016 440 -8982
rect 406 -9084 440 -9050
rect 406 -9152 440 -9118
rect 406 -9220 440 -9186
rect 406 -9288 440 -9254
rect 406 -9356 440 -9322
rect 406 -9424 440 -9390
rect 406 -9492 440 -9458
rect 406 -9560 440 -9526
rect 406 -9628 440 -9594
rect 406 -9696 440 -9662
rect 406 -9764 440 -9730
rect 406 -9832 440 -9798
rect 406 -9900 440 -9866
rect 406 -9968 440 -9934
rect 406 -10036 440 -10002
rect 406 -10104 440 -10070
rect 406 -10172 440 -10138
rect 406 -10240 440 -10206
rect 406 -10308 440 -10274
rect 406 -10376 440 -10342
rect 406 -10444 440 -10410
rect 406 -10512 440 -10478
rect 406 -10580 440 -10546
rect 406 -10648 440 -10614
rect 406 -10716 440 -10682
rect 406 -10784 440 -10750
rect 406 -10852 440 -10818
rect 406 -10920 440 -10886
rect 406 -10988 440 -10954
rect 1039 -3423 1073 -3389
rect 1039 -3491 1073 -3457
rect 1039 -3559 1073 -3525
rect 1039 -3627 1073 -3593
rect 1039 -3695 1073 -3661
rect 1039 -3763 1073 -3729
rect 1039 -3831 1073 -3797
rect 1039 -3899 1073 -3865
rect 1039 -3967 1073 -3933
rect 1039 -4035 1073 -4001
rect 1039 -4103 1073 -4069
rect 1039 -4171 1073 -4137
rect 1039 -4239 1073 -4205
rect 1039 -4307 1073 -4273
rect 1039 -4375 1073 -4341
rect 1039 -4443 1073 -4409
rect 1039 -4511 1073 -4477
rect 1039 -4579 1073 -4545
rect 1039 -4647 1073 -4613
rect 1039 -4715 1073 -4681
rect 1039 -4783 1073 -4749
rect 1039 -4851 1073 -4817
rect 1039 -4919 1073 -4885
rect 1039 -4987 1073 -4953
rect 1039 -5055 1073 -5021
rect 1039 -5123 1073 -5089
rect 1039 -5191 1073 -5157
rect 1039 -5259 1073 -5225
rect 1039 -5327 1073 -5293
rect 1039 -5395 1073 -5361
rect 1039 -5463 1073 -5429
rect 1039 -5531 1073 -5497
rect 1039 -5599 1073 -5565
rect 1039 -5667 1073 -5633
rect 1039 -5735 1073 -5701
rect 1039 -5803 1073 -5769
rect 1039 -5871 1073 -5837
rect 1039 -5939 1073 -5905
rect 1039 -6007 1073 -5973
rect 1039 -6075 1073 -6041
rect 1039 -6143 1073 -6109
rect 1039 -6211 1073 -6177
rect 1039 -6279 1073 -6245
rect 1039 -6347 1073 -6313
rect 1039 -6415 1073 -6381
rect 1039 -6483 1073 -6449
rect 1039 -6551 1073 -6517
rect 1039 -6619 1073 -6585
rect 1039 -6687 1073 -6653
rect 1039 -6755 1073 -6721
rect 1039 -6823 1073 -6789
rect 1039 -6891 1073 -6857
rect 1039 -6959 1073 -6925
rect 1039 -7027 1073 -6993
rect 1039 -7095 1073 -7061
rect 1039 -7163 1073 -7129
rect 1039 -7231 1073 -7197
rect 1039 -7299 1073 -7265
rect 1039 -7367 1073 -7333
rect 1039 -7435 1073 -7401
rect 1039 -7503 1073 -7469
rect 1039 -7571 1073 -7537
rect 1039 -7639 1073 -7605
rect 1039 -7707 1073 -7673
rect 1039 -7775 1073 -7741
rect 1039 -7843 1073 -7809
rect 1039 -7911 1073 -7877
rect 1039 -7979 1073 -7945
rect 1039 -8047 1073 -8013
rect 1039 -8115 1073 -8081
rect 1039 -8183 1073 -8149
rect 1039 -8251 1073 -8217
rect 1039 -8319 1073 -8285
rect 1039 -8387 1073 -8353
rect 1039 -8455 1073 -8421
rect 1039 -8523 1073 -8489
rect 1039 -8591 1073 -8557
rect 1039 -8659 1073 -8625
rect 1039 -8727 1073 -8693
rect 1039 -8795 1073 -8761
rect 1039 -8863 1073 -8829
rect 1039 -8931 1073 -8897
rect 1039 -8999 1073 -8965
rect 1039 -9067 1073 -9033
rect 1039 -9135 1073 -9101
rect 1039 -9203 1073 -9169
rect 1039 -9271 1073 -9237
rect 1039 -9339 1073 -9305
rect 1039 -9407 1073 -9373
rect 1039 -9475 1073 -9441
rect 1039 -9543 1073 -9509
rect 1039 -9611 1073 -9577
rect 1039 -9679 1073 -9645
rect 1039 -9747 1073 -9713
rect 1039 -9815 1073 -9781
rect 1039 -9883 1073 -9849
rect 1039 -9951 1073 -9917
rect 1039 -10019 1073 -9985
rect 1039 -10087 1073 -10053
rect 1039 -10155 1073 -10121
rect 1039 -10223 1073 -10189
rect 1039 -10291 1073 -10257
rect 1039 -10359 1073 -10325
rect 1039 -10427 1073 -10393
rect 1039 -10495 1073 -10461
rect 1039 -10563 1073 -10529
rect 1039 -10631 1073 -10597
rect 1039 -10699 1073 -10665
rect 1039 -10767 1073 -10733
rect 1039 -10835 1073 -10801
rect 1039 -10903 1073 -10869
rect 1039 -10971 1073 -10937
rect 1039 -11039 1073 -11005
rect 474 -11107 508 -11073
rect 542 -11107 576 -11073
rect 610 -11107 644 -11073
rect 678 -11107 712 -11073
rect 746 -11107 780 -11073
rect 814 -11107 848 -11073
rect 882 -11107 916 -11073
rect 950 -11107 984 -11073
<< mvnsubdiffcont >>
rect 8550 4883 8584 4917
rect 8620 4883 8654 4917
rect 8690 4883 8724 4917
rect 8760 4883 8794 4917
rect 8830 4883 8864 4917
rect 8900 4883 8934 4917
rect 8970 4883 9004 4917
rect 9040 4883 9074 4917
rect 9110 4883 9144 4917
rect 9180 4883 9214 4917
rect 9250 4883 9284 4917
rect 9320 4883 9354 4917
rect 9390 4883 9424 4917
rect 9460 4883 9494 4917
rect 9530 4883 9564 4917
rect 9599 4883 9633 4917
rect 9668 4883 9702 4917
rect 9737 4883 9771 4917
rect 9806 4883 9840 4917
rect 9875 4883 9909 4917
rect 9944 4883 9978 4917
rect 10013 4883 10047 4917
rect 10082 4883 10116 4917
rect 10151 4883 10185 4917
rect 10220 4883 10254 4917
rect 10289 4883 10323 4917
rect 10358 4883 10392 4917
rect 10427 4883 10461 4917
rect 10496 4883 10530 4917
rect 10565 4883 10599 4917
rect 10634 4883 10668 4917
rect 10703 4883 10737 4917
rect 10772 4883 10806 4917
rect 10841 4883 10875 4917
rect 10910 4883 10944 4917
rect 10979 4883 11013 4917
rect 11048 4883 11082 4917
rect 11117 4883 11151 4917
rect 11186 4883 11220 4917
rect 11322 4883 11356 4917
rect 11391 4883 11425 4917
rect 11460 4883 11494 4917
rect 11529 4883 11563 4917
rect 11598 4883 11632 4917
rect 11667 4883 11701 4917
rect 11736 4883 11770 4917
rect 11805 4883 11839 4917
rect 11874 4883 11908 4917
rect 11943 4883 11977 4917
rect 12012 4883 12046 4917
rect 12081 4883 12115 4917
rect 12150 4883 12184 4917
rect 12219 4883 12253 4917
rect 12288 4883 12322 4917
rect 12357 4883 12391 4917
rect 12426 4883 12460 4917
rect 12495 4883 12529 4917
rect 12563 4883 12597 4917
rect 12631 4883 12665 4917
rect 12699 4883 12733 4917
rect 12767 4883 12801 4917
rect 12835 4883 12869 4917
rect 12903 4883 12937 4917
rect 12971 4883 13005 4917
rect 13039 4883 13073 4917
rect 13107 4883 13141 4917
rect 13175 4883 13209 4917
rect 13243 4883 13277 4917
rect 13311 4883 13345 4917
rect 13379 4883 13413 4917
rect 13447 4883 13481 4917
rect 13515 4883 13549 4917
rect 13583 4883 13617 4917
rect 13651 4883 13685 4917
rect 13719 4883 13753 4917
rect 13787 4883 13821 4917
rect 13855 4883 13889 4917
rect 13923 4883 13957 4917
rect 13991 4883 14025 4917
rect 14059 4883 14093 4917
rect 14127 4883 14161 4917
rect 14195 4883 14229 4917
rect 14263 4883 14297 4917
rect 14331 4883 14365 4917
rect 14399 4883 14433 4917
rect 14467 4883 14501 4917
rect 14535 4883 14569 4917
rect 14603 4883 14637 4917
rect 14671 4883 14705 4917
rect 14739 4883 14773 4917
rect 14807 4883 14841 4917
rect 14875 4883 14909 4917
rect 14943 4883 14977 4917
rect 15011 4883 15045 4917
rect 15079 4883 15113 4917
rect 15147 4883 15181 4917
rect 15215 4883 15249 4917
rect 15283 4883 15317 4917
rect 15351 4883 15385 4917
rect 15419 4883 15453 4917
rect 15487 4883 15521 4917
rect 15555 4883 15589 4917
rect 15623 4883 15657 4917
rect 15691 4883 15725 4917
rect 15759 4883 15793 4917
rect 15827 4883 15861 4917
rect 15895 4883 15929 4917
rect 15963 4883 15997 4917
rect 16031 4883 16065 4917
rect 16099 4883 16133 4917
rect 16167 4883 16201 4917
rect 16235 4883 16269 4917
rect 16303 4883 16337 4917
rect 16371 4883 16405 4917
rect 16439 4883 16473 4917
rect 16507 4883 16541 4917
rect 16575 4883 16609 4917
rect 16643 4883 16677 4917
rect 16711 4883 16745 4917
rect 16779 4883 16813 4917
rect 16847 4883 16881 4917
rect 16915 4883 16949 4917
rect 16983 4883 17017 4917
rect 17051 4883 17085 4917
rect 17119 4883 17153 4917
rect 17187 4883 17221 4917
rect 17255 4883 17289 4917
rect 17323 4883 17357 4917
rect 17391 4883 17425 4917
rect 17459 4883 17493 4917
rect 17527 4883 17561 4917
rect 17595 4883 17629 4917
rect 17663 4883 17697 4917
rect 17731 4883 17765 4917
rect 17799 4883 17833 4917
rect 17867 4883 17901 4917
rect 17935 4883 17969 4917
rect 18003 4883 18037 4917
rect 18071 4883 18105 4917
rect 18139 4883 18173 4917
rect 18207 4883 18241 4917
rect 18275 4883 18309 4917
rect 18343 4883 18377 4917
rect 18411 4883 18445 4917
rect 18479 4883 18513 4917
rect 18547 4883 18581 4917
rect 18615 4883 18649 4917
rect 18683 4883 18717 4917
rect 18751 4883 18785 4917
rect 18819 4883 18853 4917
rect 18887 4883 18921 4917
rect 18955 4883 18989 4917
rect 19023 4883 19057 4917
rect 19091 4883 19125 4917
rect 19159 4883 19193 4917
rect 19227 4883 19261 4917
rect 19295 4883 19329 4917
rect 19363 4883 19397 4917
rect 19431 4883 19465 4917
rect 19499 4883 19533 4917
rect 19567 4883 19601 4917
rect 19635 4883 19669 4917
rect 19703 4883 19737 4917
rect 19771 4883 19805 4917
rect 19839 4883 19873 4917
rect 19907 4883 19941 4917
rect 8482 4814 8516 4848
rect 8482 4745 8516 4779
rect 8482 4676 8516 4710
rect 8482 4607 8516 4641
rect 8482 4538 8516 4572
rect 8482 4469 8516 4503
rect 8482 4400 8516 4434
rect 8482 4331 8516 4365
rect 8482 4262 8516 4296
rect 8482 4192 8516 4226
rect 8482 4122 8516 4156
rect 8482 4052 8516 4086
rect 8482 3982 8516 4016
rect 8482 3912 8516 3946
rect 8482 3842 8516 3876
rect 8482 3772 8516 3806
rect 11254 4749 11288 4783
rect 11254 4681 11288 4715
rect 11254 4613 11288 4647
rect 11254 4545 11288 4579
rect 11254 4477 11288 4511
rect 11254 4409 11288 4443
rect 11254 4341 11288 4375
rect 11254 4273 11288 4307
rect 11254 4205 11288 4239
rect 11254 4137 11288 4171
rect 11254 4069 11288 4103
rect 11254 4001 11288 4035
rect 11254 3933 11288 3967
rect 11254 3865 11288 3899
rect 8482 3702 8516 3736
rect 8482 3632 8516 3666
rect 11254 3797 11288 3831
rect 11254 3729 11288 3763
rect 11254 3661 11288 3695
rect 8482 3562 8516 3596
rect 19975 4801 20009 4835
rect 19975 4640 20009 4674
rect 19975 4572 20009 4606
rect 19975 4504 20009 4538
rect 19975 4436 20009 4470
rect 19975 4368 20009 4402
rect 19975 4300 20009 4334
rect 19975 4232 20009 4266
rect 19975 4164 20009 4198
rect 19975 4096 20009 4130
rect 19975 4028 20009 4062
rect 19975 3960 20009 3994
rect 19975 3892 20009 3926
rect 19975 3824 20009 3858
rect 19975 3756 20009 3790
rect 19975 3688 20009 3722
rect 11254 3593 11288 3627
rect 19975 3620 20009 3654
rect 8482 3492 8516 3526
rect 11254 3525 11288 3559
rect 8482 3422 8516 3456
rect 8482 3352 8516 3386
rect 11254 3457 11288 3491
rect 19975 3552 20009 3586
rect 19975 3484 20009 3518
rect 19975 3416 20009 3450
rect 8482 3282 8516 3316
rect 8482 3212 8516 3246
rect 11322 3348 11356 3382
rect 11390 3348 11424 3382
rect 11458 3348 11492 3382
rect 11526 3348 11560 3382
rect 11594 3348 11628 3382
rect 11662 3348 11696 3382
rect 11730 3348 11764 3382
rect 11798 3348 11832 3382
rect 11866 3348 11900 3382
rect 11934 3348 11968 3382
rect 12002 3348 12036 3382
rect 12070 3348 12104 3382
rect 12138 3348 12172 3382
rect 12206 3348 12240 3382
rect 12274 3348 12308 3382
rect 12342 3348 12376 3382
rect 12410 3348 12444 3382
rect 12478 3348 12512 3382
rect 12546 3348 12580 3382
rect 12614 3348 12648 3382
rect 12682 3348 12716 3382
rect 12750 3348 12784 3382
rect 12818 3348 12852 3382
rect 12886 3348 12920 3382
rect 12954 3348 12988 3382
rect 13022 3348 13056 3382
rect 13090 3348 13124 3382
rect 13158 3348 13192 3382
rect 13226 3348 13260 3382
rect 13294 3348 13328 3382
rect 13362 3348 13396 3382
rect 13430 3348 13464 3382
rect 13498 3348 13532 3382
rect 13566 3348 13600 3382
rect 13634 3348 13668 3382
rect 13702 3348 13736 3382
rect 13770 3348 13804 3382
rect 13838 3348 13872 3382
rect 13906 3348 13940 3382
rect 13974 3348 14008 3382
rect 14042 3348 14076 3382
rect 14110 3348 14144 3382
rect 14178 3348 14212 3382
rect 14246 3348 14280 3382
rect 14314 3348 14348 3382
rect 14382 3348 14416 3382
rect 14450 3348 14484 3382
rect 14518 3348 14552 3382
rect 14586 3348 14620 3382
rect 14654 3348 14688 3382
rect 14722 3348 14756 3382
rect 14790 3348 14824 3382
rect 14858 3348 14892 3382
rect 14926 3348 14960 3382
rect 14994 3348 15028 3382
rect 15062 3348 15096 3382
rect 15130 3348 15164 3382
rect 15198 3348 15232 3382
rect 15266 3348 15300 3382
rect 15334 3348 15368 3382
rect 15402 3348 15436 3382
rect 15470 3348 15504 3382
rect 15538 3348 15572 3382
rect 15606 3348 15640 3382
rect 15674 3348 15708 3382
rect 15742 3348 15776 3382
rect 15810 3348 15844 3382
rect 15878 3348 15912 3382
rect 15946 3348 15980 3382
rect 16014 3348 16048 3382
rect 16082 3348 16116 3382
rect 16150 3348 16184 3382
rect 16218 3348 16252 3382
rect 16286 3348 16320 3382
rect 16354 3348 16388 3382
rect 16422 3348 16456 3382
rect 16490 3348 16524 3382
rect 16558 3348 16592 3382
rect 16626 3348 16660 3382
rect 16694 3348 16728 3382
rect 16762 3348 16796 3382
rect 16830 3348 16864 3382
rect 16898 3348 16932 3382
rect 16966 3348 17000 3382
rect 17034 3348 17068 3382
rect 17102 3348 17136 3382
rect 17170 3348 17204 3382
rect 17238 3348 17272 3382
rect 17306 3348 17340 3382
rect 17374 3348 17408 3382
rect 17442 3348 17476 3382
rect 17510 3348 17544 3382
rect 17578 3348 17612 3382
rect 17646 3348 17680 3382
rect 17714 3348 17748 3382
rect 17782 3348 17816 3382
rect 17850 3348 17884 3382
rect 17918 3348 17952 3382
rect 17986 3348 18020 3382
rect 18054 3348 18088 3382
rect 18122 3348 18156 3382
rect 18190 3348 18224 3382
rect 18258 3348 18292 3382
rect 18326 3348 18360 3382
rect 18394 3348 18428 3382
rect 18462 3348 18496 3382
rect 18530 3348 18564 3382
rect 18598 3348 18632 3382
rect 18666 3348 18700 3382
rect 18734 3348 18768 3382
rect 18802 3348 18836 3382
rect 18870 3348 18904 3382
rect 18938 3348 18972 3382
rect 19006 3348 19040 3382
rect 19074 3348 19108 3382
rect 19142 3348 19176 3382
rect 19210 3348 19244 3382
rect 19278 3348 19312 3382
rect 19346 3348 19380 3382
rect 19414 3348 19448 3382
rect 19482 3348 19516 3382
rect 19550 3348 19584 3382
rect 19618 3348 19652 3382
rect 19686 3348 19720 3382
rect 19754 3348 19788 3382
rect 19822 3348 19856 3382
rect 19890 3348 19924 3382
rect 11261 3280 11295 3314
rect 8482 3142 8516 3176
rect 11261 3197 11295 3231
rect 8482 3072 8516 3106
rect 11261 3114 11295 3148
rect 8482 3002 8516 3036
rect 10401 3053 10435 3087
rect 10474 3053 10508 3087
rect 10547 3053 10581 3087
rect 10620 3053 10654 3087
rect 10692 3053 10726 3087
rect 10764 3053 10798 3087
rect 10836 3053 10870 3087
rect 10908 3053 10942 3087
rect 10980 3053 11014 3087
rect 11052 3053 11086 3087
rect 11124 3053 11158 3087
rect 11196 3053 11230 3087
rect 8550 2968 8584 3002
rect 8619 2968 8653 3002
rect 8688 2968 8722 3002
rect 8757 2968 8791 3002
rect 8826 2968 8860 3002
rect 8895 2968 8929 3002
rect 8964 2968 8998 3002
rect 9033 2968 9067 3002
rect 9102 2968 9136 3002
rect 9171 2968 9205 3002
rect 9240 2968 9274 3002
rect 9309 2968 9343 3002
rect 9378 2968 9412 3002
rect 9447 2968 9481 3002
rect 9516 2968 9550 3002
rect 9585 2968 9619 3002
rect 9654 2968 9688 3002
rect 9723 2968 9757 3002
rect 9792 2968 9826 3002
rect 9861 2968 9895 3002
rect 9929 2968 9963 3002
rect 9997 2968 10031 3002
rect 10065 2968 10099 3002
rect 10133 2968 10167 3002
rect 10201 2968 10235 3002
rect 10269 2968 10303 3002
rect 598 2518 632 2552
rect 668 2518 702 2552
rect 738 2518 772 2552
rect 808 2518 842 2552
rect 878 2518 912 2552
rect 948 2518 982 2552
rect 1019 2518 1053 2552
rect 1090 2518 1124 2552
rect 1161 2518 1195 2552
rect 1232 2518 1266 2552
rect 1303 2518 1337 2552
rect 1374 2518 1408 2552
rect 1445 2518 1479 2552
rect 1516 2518 1550 2552
rect 2271 2465 2305 2499
rect 2339 2465 2373 2499
rect 2407 2465 2441 2499
rect 2475 2465 2509 2499
rect 2543 2465 2577 2499
rect 2611 2465 2645 2499
rect 2679 2465 2713 2499
rect 2747 2465 2781 2499
rect 2815 2465 2849 2499
rect 2883 2465 2917 2499
rect 2951 2465 2985 2499
rect 3019 2465 3053 2499
rect 3087 2465 3121 2499
rect 3155 2465 3189 2499
rect 3223 2465 3257 2499
rect 3291 2465 3325 2499
rect 3359 2465 3393 2499
rect 3427 2465 3461 2499
rect 3495 2465 3529 2499
rect 3563 2465 3597 2499
rect 3631 2465 3665 2499
rect 3699 2465 3733 2499
rect 3767 2465 3801 2499
rect 3835 2465 3869 2499
rect 3903 2465 3937 2499
rect 3971 2465 4005 2499
rect 4039 2465 4073 2499
rect 4107 2465 4141 2499
rect 4175 2465 4209 2499
rect 4243 2465 4277 2499
rect 4311 2465 4345 2499
rect 4379 2465 4413 2499
rect 4447 2465 4481 2499
rect 4515 2465 4549 2499
rect 4583 2465 4617 2499
rect 4651 2465 4685 2499
rect 4719 2465 4753 2499
rect 4787 2465 4821 2499
rect 4855 2465 4889 2499
rect 4923 2465 4957 2499
rect 4991 2465 5025 2499
rect 5059 2465 5093 2499
rect 5127 2465 5161 2499
rect 5195 2465 5229 2499
rect 5263 2465 5297 2499
rect 5331 2465 5365 2499
rect 5399 2465 5433 2499
rect 5467 2465 5501 2499
rect 5535 2465 5569 2499
rect 5603 2465 5637 2499
rect 5671 2465 5705 2499
rect 5739 2465 5773 2499
rect 5807 2465 5841 2499
rect 5875 2465 5909 2499
rect 5943 2465 5977 2499
rect 6011 2465 6045 2499
rect 6079 2465 6113 2499
rect 6147 2465 6181 2499
rect 6215 2465 6249 2499
rect 6283 2465 6317 2499
rect 6351 2465 6385 2499
rect 6419 2465 6453 2499
rect 6487 2465 6521 2499
rect 6555 2465 6589 2499
rect 6623 2465 6657 2499
rect 6691 2465 6725 2499
rect 6759 2465 6793 2499
rect 6827 2465 6861 2499
rect 6895 2465 6929 2499
rect 6963 2465 6997 2499
rect 7031 2465 7065 2499
rect 7099 2465 7133 2499
rect 7167 2465 7201 2499
rect 7235 2465 7269 2499
rect 7303 2465 7337 2499
rect 7371 2465 7405 2499
rect 7439 2465 7473 2499
rect 7507 2465 7541 2499
rect 7575 2465 7609 2499
rect 7643 2465 7677 2499
rect 7711 2465 7745 2499
rect 7779 2465 7813 2499
rect 7847 2465 7881 2499
rect 7915 2465 7949 2499
rect 7983 2465 8017 2499
rect 8051 2465 8085 2499
rect 8119 2465 8153 2499
rect 8187 2465 8221 2499
rect 8255 2465 8289 2499
rect 8323 2465 8357 2499
rect 8391 2465 8425 2499
rect 8459 2465 8493 2499
rect 8527 2465 8561 2499
rect 8595 2465 8629 2499
rect 8663 2465 8697 2499
rect 8731 2465 8765 2499
rect 8799 2465 8833 2499
rect 8867 2465 8901 2499
rect 8935 2465 8969 2499
rect 9003 2465 9037 2499
rect 9071 2465 9105 2499
rect 9139 2465 9173 2499
rect 9207 2465 9241 2499
rect 9275 2465 9309 2499
rect 9343 2465 9377 2499
rect 2151 2397 2185 2431
rect 2151 2329 2185 2363
rect 2151 2261 2185 2295
rect 9411 2341 9445 2375
rect 9411 2273 9445 2307
rect 2151 2193 2185 2227
rect 598 2130 632 2164
rect 669 2130 703 2164
rect 740 2130 774 2164
rect 811 2130 845 2164
rect 882 2130 916 2164
rect 953 2130 987 2164
rect 1024 2130 1058 2164
rect 1095 2130 1129 2164
rect 1166 2130 1200 2164
rect 1236 2130 1270 2164
rect 1306 2130 1340 2164
rect 1376 2130 1410 2164
rect 1446 2130 1480 2164
rect 1516 2130 1550 2164
rect 598 2062 632 2096
rect 669 2062 703 2096
rect 740 2062 774 2096
rect 811 2062 845 2096
rect 882 2062 916 2096
rect 953 2062 987 2096
rect 1024 2062 1058 2096
rect 1095 2062 1129 2096
rect 1166 2062 1200 2096
rect 1236 2062 1270 2096
rect 1306 2062 1340 2096
rect 1376 2062 1410 2096
rect 1446 2062 1480 2096
rect 1516 2062 1550 2096
rect 598 1994 632 2028
rect 669 1994 703 2028
rect 740 1994 774 2028
rect 811 1994 845 2028
rect 882 1994 916 2028
rect 953 1994 987 2028
rect 1024 1994 1058 2028
rect 1095 1994 1129 2028
rect 1166 1994 1200 2028
rect 1236 1994 1270 2028
rect 1306 1994 1340 2028
rect 1376 1994 1410 2028
rect 1446 1994 1480 2028
rect 1516 1994 1550 2028
rect 598 1926 632 1960
rect 669 1926 703 1960
rect 740 1926 774 1960
rect 811 1926 845 1960
rect 882 1926 916 1960
rect 953 1926 987 1960
rect 1024 1926 1058 1960
rect 1095 1926 1129 1960
rect 1166 1926 1200 1960
rect 1236 1926 1270 1960
rect 1306 1926 1340 1960
rect 1376 1926 1410 1960
rect 1446 1926 1480 1960
rect 1516 1926 1550 1960
rect 9411 2205 9445 2239
rect 2151 2125 2185 2159
rect 9411 2137 9445 2171
rect 2151 2057 2185 2091
rect 2151 1989 2185 2023
rect 2151 1921 2185 1955
rect 2151 1853 2185 1887
rect 2151 1785 2185 1819
rect 2151 1717 2185 1751
rect 2151 1649 2185 1683
rect 9411 2069 9445 2103
rect 9411 2001 9445 2035
rect 9411 1933 9445 1967
rect 9411 1865 9445 1899
rect 9411 1797 9445 1831
rect 9411 1729 9445 1763
rect 9411 1661 9445 1695
rect 2151 1581 2185 1615
rect 2151 1513 2185 1547
rect 2151 1445 2185 1479
rect 9411 1593 9445 1627
rect 17817 2572 17851 2606
rect 17889 2572 17923 2606
rect 17961 2572 17995 2606
rect 18033 2572 18067 2606
rect 18105 2572 18139 2606
rect 18176 2572 18210 2606
rect 18247 2572 18281 2606
rect 18318 2572 18352 2606
rect 18389 2572 18423 2606
rect 18460 2572 18494 2606
rect 18531 2572 18565 2606
rect 18602 2572 18636 2606
rect 18673 2572 18707 2606
rect 18744 2572 18778 2606
rect 18815 2572 18849 2606
rect 18886 2572 18920 2606
rect 18957 2572 18991 2606
rect 19028 2572 19062 2606
rect 9411 1525 9445 1559
rect 598 1367 632 1401
rect 668 1367 702 1401
rect 738 1367 772 1401
rect 808 1367 842 1401
rect 878 1367 912 1401
rect 948 1367 982 1401
rect 1019 1367 1053 1401
rect 1090 1367 1124 1401
rect 1161 1367 1195 1401
rect 1232 1367 1266 1401
rect 1303 1367 1337 1401
rect 1374 1367 1408 1401
rect 1445 1367 1479 1401
rect 1516 1367 1550 1401
rect 2151 1377 2185 1411
rect 2151 1309 2185 1343
rect 2151 1241 2185 1275
rect 2151 1173 2185 1207
rect 9411 1457 9445 1491
rect 2151 1105 2185 1139
rect 2151 1037 2185 1071
rect 2151 969 2185 1003
rect 2151 901 2185 935
rect 2151 833 2185 867
rect 2151 765 2185 799
rect 2151 697 2185 731
rect 2151 629 2185 663
rect 2151 561 2185 595
rect 2151 493 2185 527
rect 2151 425 2185 459
rect 2151 357 2185 391
rect 2151 289 2185 323
rect 2151 221 2185 255
rect 2151 153 2185 187
rect 2151 85 2185 119
rect 2151 17 2185 51
rect 9411 1389 9445 1423
rect 9479 1321 9513 1355
rect 9547 1321 9581 1355
rect 9615 1321 9649 1355
rect 9683 1321 9717 1355
rect 9751 1321 9785 1355
rect 9819 1321 9853 1355
rect 9887 1321 9921 1355
rect 9955 1321 9989 1355
rect 10023 1321 10057 1355
rect 10091 1321 10125 1355
rect 10159 1321 10193 1355
rect 10227 1321 10261 1355
rect 10295 1321 10329 1355
rect 10363 1321 10397 1355
rect 10431 1321 10465 1355
rect 10499 1321 10533 1355
rect 10567 1321 10601 1355
rect 10635 1321 10669 1355
rect 10703 1321 10737 1355
rect 10771 1321 10805 1355
rect 10839 1321 10873 1355
rect 10907 1321 10941 1355
rect 10975 1321 11009 1355
rect 11043 1321 11077 1355
rect 11111 1321 11145 1355
rect 11179 1321 11213 1355
rect 11247 1321 11281 1355
rect 11315 1321 11349 1355
rect 11383 1321 11417 1355
rect 11451 1321 11485 1355
rect 11519 1321 11553 1355
rect 11587 1321 11621 1355
rect 11655 1321 11689 1355
rect 11723 1321 11757 1355
rect 11791 1321 11825 1355
rect 11859 1321 11893 1355
rect 11927 1321 11961 1355
rect 11995 1321 12029 1355
rect 12063 1321 12097 1355
rect 12131 1321 12165 1355
rect 12199 1321 12233 1355
rect 12267 1321 12301 1355
rect 12335 1321 12369 1355
rect 12403 1321 12437 1355
rect 12471 1321 12505 1355
rect 12539 1321 12573 1355
rect 12607 1321 12641 1355
rect 12675 1321 12709 1355
rect 12743 1321 12777 1355
rect 12811 1321 12845 1355
rect 12879 1321 12913 1355
rect 12947 1321 12981 1355
rect 13015 1321 13049 1355
rect 13083 1321 13117 1355
rect 13151 1321 13185 1355
rect 13219 1321 13253 1355
rect 13287 1321 13321 1355
rect 13355 1321 13389 1355
rect 13423 1321 13457 1355
rect 13491 1321 13525 1355
rect 13559 1321 13593 1355
rect 13627 1321 13661 1355
rect 13695 1321 13729 1355
rect 13763 1321 13797 1355
rect 13831 1321 13865 1355
rect 13899 1321 13933 1355
rect 13967 1321 14001 1355
rect 14035 1321 14069 1355
rect 14103 1321 14137 1355
rect 14171 1321 14205 1355
rect 14239 1321 14273 1355
rect 14307 1321 14341 1355
rect 14375 1321 14409 1355
rect 14443 1321 14477 1355
rect 14511 1321 14545 1355
rect 14579 1321 14613 1355
rect 14647 1321 14681 1355
rect 14715 1321 14749 1355
rect 14783 1321 14817 1355
rect 14851 1321 14885 1355
rect 14919 1321 14953 1355
rect 14987 1321 15021 1355
rect 15055 1321 15089 1355
rect 15123 1321 15157 1355
rect 15191 1321 15225 1355
rect 15259 1321 15293 1355
rect 15327 1321 15361 1355
rect 15395 1321 15429 1355
rect 15463 1321 15497 1355
rect 15531 1321 15565 1355
rect 15599 1321 15633 1355
rect 15667 1321 15701 1355
rect 15735 1321 15769 1355
rect 15803 1321 15837 1355
rect 15871 1321 15905 1355
rect 15939 1321 15973 1355
rect 16007 1321 16041 1355
rect 16075 1321 16109 1355
rect 16143 1321 16177 1355
rect 16211 1321 16245 1355
rect 16279 1321 16313 1355
rect 16347 1321 16381 1355
rect 16415 1321 16449 1355
rect 16483 1321 16517 1355
rect 16551 1321 16585 1355
rect 16619 1321 16653 1355
rect 16687 1321 16721 1355
rect 16755 1321 16789 1355
rect 16823 1321 16857 1355
rect 16891 1321 16925 1355
rect 16959 1321 16993 1355
rect 17027 1321 17061 1355
rect 17095 1321 17129 1355
rect 17163 1321 17197 1355
rect 17231 1321 17265 1355
rect 17299 1321 17333 1355
rect 17367 1321 17401 1355
rect 17435 1321 17469 1355
rect 17503 1321 17537 1355
rect 17571 1321 17605 1355
rect 17639 1321 17673 1355
rect 17707 1321 17741 1355
rect 17775 1321 17809 1355
rect 17843 1321 17877 1355
rect 17911 1321 17945 1355
rect 17979 1321 18013 1355
rect 18047 1321 18081 1355
rect 18115 1321 18149 1355
rect 18183 1321 18217 1355
rect 18251 1321 18285 1355
rect 18319 1321 18353 1355
rect 18387 1321 18421 1355
rect 18455 1321 18489 1355
rect 18523 1321 18557 1355
rect 18591 1321 18625 1355
rect 18659 1321 18693 1355
rect 18727 1321 18761 1355
rect 18795 1321 18829 1355
rect 18863 1214 18897 1248
rect 28031 1761 28065 1795
rect 28031 1693 28065 1727
rect 28031 1625 28065 1659
rect 28031 1557 28065 1591
rect 28031 1489 28065 1523
rect 28031 1421 28065 1455
rect 28031 1353 28065 1387
rect 28031 1285 28065 1319
rect 28031 1217 28065 1251
rect 18863 1146 18897 1180
rect 2151 -51 2185 -17
rect 18863 1078 18897 1112
rect 18863 1010 18897 1044
rect 18863 942 18897 976
rect 18863 874 18897 908
rect 18863 806 18897 840
rect 18863 738 18897 772
rect 18863 670 18897 704
rect 18863 602 18897 636
rect 18863 534 18897 568
rect 18863 466 18897 500
rect 18863 398 18897 432
rect 18863 330 18897 364
rect 18863 262 18897 296
rect 18863 194 18897 228
rect 2151 -119 2185 -85
rect 2151 -268 2185 -234
rect 2219 -360 2253 -326
rect 2287 -360 2321 -326
rect 2355 -360 2389 -326
rect 2423 -360 2457 -326
rect 2491 -360 2525 -326
rect 2559 -360 2593 -326
rect 2627 -360 2661 -326
rect 2695 -360 2729 -326
rect 2763 -360 2797 -326
rect 2831 -360 2865 -326
rect 2899 -360 2933 -326
rect 2967 -360 3001 -326
rect 3035 -360 3069 -326
rect 3103 -360 3137 -326
rect 3171 -360 3205 -326
rect 3239 -360 3273 -326
rect 3307 -360 3341 -326
rect 598 -917 632 -883
rect 668 -917 702 -883
rect 738 -917 772 -883
rect 808 -917 842 -883
rect 878 -917 912 -883
rect 948 -917 982 -883
rect 1019 -917 1053 -883
rect 1090 -917 1124 -883
rect 1161 -917 1195 -883
rect 1232 -917 1266 -883
rect 1303 -917 1337 -883
rect 1374 -917 1408 -883
rect 1445 -917 1479 -883
rect 1516 -917 1550 -883
rect 18863 126 18897 160
rect 18863 58 18897 92
rect 18863 -10 18897 24
rect 18863 -78 18897 -44
rect 18863 -146 18897 -112
rect 18863 -214 18897 -180
rect 18863 -282 18897 -248
rect 18863 -350 18897 -316
rect 18863 -418 18897 -384
rect 18863 -486 18897 -452
rect 18863 -554 18897 -520
rect 18863 -622 18897 -588
rect 18863 -690 18897 -656
rect 18863 -758 18897 -724
rect 18863 -826 18897 -792
rect 18863 -894 18897 -860
rect 18863 -962 18897 -928
rect 18863 -1030 18897 -996
rect 18863 -1098 18897 -1064
rect 18863 -1166 18897 -1132
rect 18016 -1234 18050 -1200
rect 18096 -1234 18130 -1200
rect 18176 -1234 18210 -1200
rect 18255 -1234 18289 -1200
rect 18334 -1234 18368 -1200
rect 18413 -1234 18447 -1200
rect 18530 -1234 18564 -1200
rect 18598 -1234 18632 -1200
rect 18666 -1234 18700 -1200
rect 18734 -1234 18768 -1200
rect 28031 1149 28065 1183
rect 28031 1081 28065 1115
rect 28031 1013 28065 1047
rect 28031 945 28065 979
rect 28031 877 28065 911
rect 28031 809 28065 843
rect 28031 741 28065 775
rect 28031 673 28065 707
rect 28031 605 28065 639
rect 28031 537 28065 571
rect 28031 469 28065 503
rect 28031 401 28065 435
rect 28031 333 28065 367
rect 28031 265 28065 299
rect 28031 197 28065 231
rect 28031 129 28065 163
rect 28031 61 28065 95
rect 28031 -7 28065 27
rect 28031 -75 28065 -41
rect 28031 -143 28065 -109
rect 28031 -211 28065 -177
rect 28031 -279 28065 -245
rect 28031 -347 28065 -313
rect 28031 -415 28065 -381
rect 28031 -483 28065 -449
rect 28031 -551 28065 -517
rect 28031 -619 28065 -585
rect 28031 -687 28065 -653
rect 28031 -755 28065 -721
rect 28031 -823 28065 -789
rect 28031 -891 28065 -857
rect 28031 -959 28065 -925
rect 28031 -1027 28065 -993
rect 28031 -1095 28065 -1061
rect 28031 -1163 28065 -1129
rect 28031 -1231 28065 -1197
rect 28031 -1299 28065 -1265
rect 28031 -1367 28065 -1333
rect 28031 -1435 28065 -1401
rect 28031 -1503 28065 -1469
rect 28031 -1571 28065 -1537
rect 28031 -1639 28065 -1605
rect 28031 -1707 28065 -1673
rect 28031 -1775 28065 -1741
rect 28031 -1843 28065 -1809
rect 28031 -1911 28065 -1877
rect 28031 -1979 28065 -1945
rect 28031 -2047 28065 -2013
rect 28031 -2115 28065 -2081
rect 28031 -2183 28065 -2149
rect 28031 -2251 28065 -2217
rect 28031 -2319 28065 -2285
rect 28031 -2387 28065 -2353
rect 598 -2432 632 -2398
rect 668 -2432 702 -2398
rect 738 -2432 772 -2398
rect 808 -2432 842 -2398
rect 878 -2432 912 -2398
rect 948 -2432 982 -2398
rect 1019 -2432 1053 -2398
rect 1090 -2432 1124 -2398
rect 1161 -2432 1195 -2398
rect 1232 -2432 1266 -2398
rect 1303 -2432 1337 -2398
rect 1374 -2432 1408 -2398
rect 1445 -2432 1479 -2398
rect 1516 -2432 1550 -2398
rect 28031 -2455 28065 -2421
rect 28031 -2523 28065 -2489
rect 28031 -2591 28065 -2557
rect 28031 -2659 28065 -2625
rect 28031 -2727 28065 -2693
rect 28031 -2795 28065 -2761
rect 28031 -2863 28065 -2829
rect 28031 -2931 28065 -2897
rect 28031 -2999 28065 -2965
rect 28031 -3067 28065 -3033
rect 28031 -3135 28065 -3101
rect 28031 -3203 28065 -3169
rect 28031 -3271 28065 -3237
rect 28031 -3339 28065 -3305
rect 28031 -3407 28065 -3373
rect 28031 -3475 28065 -3441
rect 28031 -3543 28065 -3509
rect 28031 -3611 28065 -3577
rect 28031 -3679 28065 -3645
rect 28031 -3747 28065 -3713
rect 28031 -3815 28065 -3781
rect 28031 -3883 28065 -3849
rect 28031 -3951 28065 -3917
rect 28031 -4019 28065 -3985
rect 28031 -4087 28065 -4053
rect 28031 -4155 28065 -4121
rect 28031 -4223 28065 -4189
rect 28031 -4291 28065 -4257
rect 28031 -4359 28065 -4325
rect 28031 -4427 28065 -4393
rect 28031 -4495 28065 -4461
rect 28031 -4563 28065 -4529
rect 28031 -4631 28065 -4597
rect 28031 -4699 28065 -4665
rect 28031 -4767 28065 -4733
rect 28031 -4835 28065 -4801
rect 28031 -4903 28065 -4869
rect 28031 -4971 28065 -4937
rect 28031 -5039 28065 -5005
rect 28031 -5107 28065 -5073
rect 28031 -5175 28065 -5141
rect 28031 -5243 28065 -5209
rect 28031 -5311 28065 -5277
rect 28031 -5379 28065 -5345
rect 28031 -5447 28065 -5413
rect 28031 -5515 28065 -5481
rect 28031 -5583 28065 -5549
rect 28031 -5651 28065 -5617
rect 28031 -5719 28065 -5685
rect 28031 -5787 28065 -5753
rect 28031 -5855 28065 -5821
rect 28031 -5923 28065 -5889
rect 28031 -5991 28065 -5957
rect 28031 -6059 28065 -6025
rect 28031 -6127 28065 -6093
rect 28031 -6195 28065 -6161
rect 28031 -6263 28065 -6229
rect 28031 -6331 28065 -6297
rect 28031 -6399 28065 -6365
rect 28031 -6467 28065 -6433
rect 28031 -6535 28065 -6501
rect 28031 -6603 28065 -6569
rect 28031 -6671 28065 -6637
rect 28031 -6739 28065 -6705
rect 28031 -6807 28065 -6773
rect 28031 -6875 28065 -6841
rect 28031 -6943 28065 -6909
rect 28031 -7011 28065 -6977
rect 28031 -7079 28065 -7045
rect 28031 -7147 28065 -7113
rect 28031 -7215 28065 -7181
rect 28031 -7283 28065 -7249
rect 28031 -7351 28065 -7317
rect 28031 -7419 28065 -7385
rect 28031 -7487 28065 -7453
rect 28031 -7555 28065 -7521
rect 28031 -7623 28065 -7589
rect 28031 -7691 28065 -7657
rect 28031 -7759 28065 -7725
rect 28031 -7827 28065 -7793
rect 28031 -7895 28065 -7861
rect 28031 -7963 28065 -7929
rect 28031 -8031 28065 -7997
rect 28031 -8099 28065 -8065
rect 28031 -8167 28065 -8133
rect 28031 -8235 28065 -8201
rect 28031 -8303 28065 -8269
rect 28031 -8371 28065 -8337
rect 28031 -8439 28065 -8405
rect 28031 -8507 28065 -8473
rect 28031 -8575 28065 -8541
rect 28031 -8643 28065 -8609
rect 28031 -8711 28065 -8677
rect 28031 -8779 28065 -8745
rect 28031 -8847 28065 -8813
rect 28031 -8915 28065 -8881
rect 28031 -8983 28065 -8949
rect 28031 -9051 28065 -9017
rect 28031 -9119 28065 -9085
rect 28031 -9187 28065 -9153
rect 28031 -9255 28065 -9221
rect 28031 -9323 28065 -9289
rect 28031 -9391 28065 -9357
rect 28031 -9459 28065 -9425
rect 28031 -9527 28065 -9493
rect 28031 -9595 28065 -9561
rect 28031 -9663 28065 -9629
rect 28031 -9731 28065 -9697
rect 28031 -9799 28065 -9765
rect 28031 -9867 28065 -9833
rect 28031 -9935 28065 -9901
rect 28031 -10003 28065 -9969
rect 28031 -10071 28065 -10037
rect 28031 -10139 28065 -10105
rect 28031 -10207 28065 -10173
rect 28031 -10275 28065 -10241
rect 28031 -10343 28065 -10309
rect 28031 -10411 28065 -10377
rect 28031 -10479 28065 -10445
rect 23987 -10642 24021 -10608
rect 24055 -10642 24089 -10608
rect 24123 -10642 24157 -10608
rect 24191 -10642 24225 -10608
rect 24259 -10642 24293 -10608
rect 24327 -10642 24361 -10608
rect 24395 -10642 24429 -10608
rect 24463 -10642 24497 -10608
rect 24531 -10642 24565 -10608
rect 24599 -10642 24633 -10608
rect 24667 -10642 24701 -10608
rect 24735 -10642 24769 -10608
rect 24803 -10642 24837 -10608
rect 24871 -10642 24905 -10608
rect 24939 -10642 24973 -10608
rect 25007 -10642 25041 -10608
rect 25075 -10642 25109 -10608
rect 25143 -10642 25177 -10608
rect 25211 -10642 25245 -10608
rect 25279 -10642 25313 -10608
rect 25347 -10642 25381 -10608
rect 25415 -10642 25449 -10608
rect 25483 -10642 25517 -10608
rect 25551 -10642 25585 -10608
rect 25619 -10642 25653 -10608
rect 25687 -10642 25721 -10608
rect 25755 -10642 25789 -10608
rect 25823 -10642 25857 -10608
rect 25891 -10642 25925 -10608
rect 25959 -10642 25993 -10608
rect 26027 -10642 26061 -10608
rect 26095 -10642 26129 -10608
rect 26163 -10642 26197 -10608
rect 26231 -10642 26265 -10608
rect 26299 -10642 26333 -10608
rect 26367 -10642 26401 -10608
rect 26435 -10642 26469 -10608
rect 26503 -10642 26537 -10608
rect 26571 -10642 26605 -10608
rect 26639 -10642 26673 -10608
rect 26707 -10642 26741 -10608
rect 26775 -10642 26809 -10608
rect 26843 -10642 26877 -10608
rect 26911 -10642 26945 -10608
rect 26979 -10642 27013 -10608
rect 27047 -10642 27081 -10608
rect 27115 -10642 27149 -10608
rect 27183 -10642 27217 -10608
rect 27251 -10642 27285 -10608
rect 27319 -10642 27353 -10608
rect 27387 -10642 27421 -10608
rect 27455 -10642 27489 -10608
rect 27523 -10642 27557 -10608
rect 27591 -10642 27625 -10608
rect 27659 -10642 27693 -10608
rect 27727 -10642 27761 -10608
rect 27795 -10642 27829 -10608
rect 27863 -10642 27897 -10608
rect 27931 -10642 27965 -10608
<< poly >>
rect 916 4819 1716 4851
rect 1772 4819 1972 4851
rect 2028 4819 2228 4851
rect 2284 4819 2484 4851
rect 2540 4819 2740 4851
rect 2796 4819 2996 4851
rect 3052 4819 3252 4851
rect 3308 4819 3508 4851
rect 3564 4819 3764 4851
rect 3820 4819 4020 4851
rect 4076 4819 4276 4851
rect 4332 4819 4532 4851
rect 4588 4819 4788 4851
rect 4844 4819 5044 4851
rect 5100 4819 5300 4851
rect 5356 4819 5556 4851
rect 5612 4819 5812 4851
rect 5868 4819 6068 4851
rect 6124 4819 6324 4851
rect 6380 4819 6580 4851
rect 6636 4819 6836 4851
rect 6892 4819 7692 4851
rect 916 4677 1716 4709
rect 1772 4677 1972 4709
rect 916 4661 1972 4677
rect 916 4627 932 4661
rect 966 4627 1003 4661
rect 1037 4627 1074 4661
rect 1108 4627 1145 4661
rect 1179 4627 1216 4661
rect 1250 4627 1287 4661
rect 1321 4627 1358 4661
rect 1392 4627 1429 4661
rect 1463 4627 1500 4661
rect 1534 4627 1571 4661
rect 1605 4627 1642 4661
rect 1676 4627 1712 4661
rect 1746 4627 1782 4661
rect 1816 4627 1852 4661
rect 1886 4627 1922 4661
rect 1956 4627 1972 4661
rect 916 4611 1972 4627
rect 2028 4677 2228 4709
rect 2284 4677 2484 4709
rect 2540 4677 2740 4709
rect 2796 4677 2996 4709
rect 3052 4677 3252 4709
rect 2028 4661 3252 4677
rect 2028 4627 2044 4661
rect 2078 4627 2112 4661
rect 2146 4627 2180 4661
rect 2214 4627 2248 4661
rect 2282 4627 2316 4661
rect 2350 4627 2384 4661
rect 2418 4627 2452 4661
rect 2486 4627 2520 4661
rect 2554 4627 2588 4661
rect 2622 4627 2656 4661
rect 2690 4627 2724 4661
rect 2758 4627 2792 4661
rect 2826 4627 2860 4661
rect 2894 4627 2928 4661
rect 2962 4627 2996 4661
rect 3030 4627 3064 4661
rect 3098 4627 3133 4661
rect 3167 4627 3202 4661
rect 3236 4627 3252 4661
rect 2028 4611 3252 4627
rect 3308 4661 3508 4709
rect 3308 4627 3324 4661
rect 3358 4627 3458 4661
rect 3492 4627 3508 4661
rect 3308 4611 3508 4627
rect 3564 4677 3764 4709
rect 3820 4677 4020 4709
rect 4076 4677 4276 4709
rect 4332 4677 4532 4709
rect 4588 4677 4788 4709
rect 4844 4677 5044 4709
rect 5100 4677 5300 4709
rect 5356 4677 5556 4709
rect 5612 4677 5812 4709
rect 5868 4677 6068 4709
rect 6124 4677 6324 4709
rect 6380 4677 6580 4709
rect 6636 4677 6836 4709
rect 3564 4661 6836 4677
rect 3564 4627 3580 4661
rect 3614 4627 3648 4661
rect 3682 4627 3716 4661
rect 3750 4627 3784 4661
rect 3818 4627 3852 4661
rect 3886 4627 3920 4661
rect 3954 4627 3988 4661
rect 4022 4627 4056 4661
rect 4090 4627 4124 4661
rect 4158 4627 4192 4661
rect 4226 4627 4260 4661
rect 4294 4627 4328 4661
rect 4362 4627 4396 4661
rect 4430 4627 4464 4661
rect 4498 4627 4532 4661
rect 4566 4627 4600 4661
rect 4634 4627 4668 4661
rect 4702 4627 4736 4661
rect 4770 4627 4804 4661
rect 4838 4627 4872 4661
rect 4906 4627 4940 4661
rect 4974 4627 5008 4661
rect 5042 4627 5076 4661
rect 5110 4627 5144 4661
rect 5178 4627 5212 4661
rect 5246 4627 5280 4661
rect 5314 4627 5348 4661
rect 5382 4627 5416 4661
rect 5450 4627 5484 4661
rect 5518 4627 5552 4661
rect 5586 4627 5620 4661
rect 5654 4627 5688 4661
rect 5722 4627 5756 4661
rect 5790 4627 5824 4661
rect 5858 4627 5892 4661
rect 5926 4627 5960 4661
rect 5994 4627 6028 4661
rect 6062 4627 6096 4661
rect 6130 4627 6165 4661
rect 6199 4627 6234 4661
rect 6268 4627 6303 4661
rect 6337 4627 6372 4661
rect 6406 4627 6441 4661
rect 6475 4627 6510 4661
rect 6544 4627 6579 4661
rect 6613 4627 6648 4661
rect 6682 4627 6717 4661
rect 6751 4627 6786 4661
rect 6820 4627 6836 4661
rect 3564 4611 6836 4627
rect 6892 4661 7692 4709
rect 6892 4627 7010 4661
rect 7044 4627 7080 4661
rect 7114 4627 7150 4661
rect 7184 4627 7220 4661
rect 7254 4627 7290 4661
rect 7324 4627 7360 4661
rect 7394 4627 7430 4661
rect 7464 4627 7500 4661
rect 7534 4627 7571 4661
rect 7605 4627 7642 4661
rect 7676 4627 7692 4661
rect 6892 4611 7692 4627
rect 916 4483 1716 4499
rect 916 4449 932 4483
rect 966 4449 1006 4483
rect 1040 4449 1080 4483
rect 1114 4449 1154 4483
rect 1188 4449 1228 4483
rect 1262 4449 1301 4483
rect 1335 4449 1374 4483
rect 1408 4449 1447 4483
rect 1481 4449 1520 4483
rect 1554 4449 1593 4483
rect 1627 4449 1666 4483
rect 1700 4449 1716 4483
rect 916 4401 1716 4449
rect 1772 4483 3764 4499
rect 1772 4449 1788 4483
rect 1822 4449 1856 4483
rect 1890 4449 1924 4483
rect 1958 4449 1992 4483
rect 2026 4449 2060 4483
rect 2094 4449 2128 4483
rect 2162 4449 2196 4483
rect 2230 4449 2265 4483
rect 2299 4449 2334 4483
rect 2368 4449 2403 4483
rect 2437 4449 2472 4483
rect 2506 4449 2541 4483
rect 2575 4449 2610 4483
rect 2644 4449 2679 4483
rect 2713 4449 2748 4483
rect 2782 4449 2817 4483
rect 2851 4449 2886 4483
rect 2920 4449 2955 4483
rect 2989 4449 3024 4483
rect 3058 4449 3093 4483
rect 3127 4449 3162 4483
rect 3196 4449 3231 4483
rect 3265 4449 3300 4483
rect 3334 4449 3369 4483
rect 3403 4449 3438 4483
rect 3472 4449 3507 4483
rect 3541 4449 3576 4483
rect 3610 4449 3645 4483
rect 3679 4449 3714 4483
rect 3748 4449 3764 4483
rect 1772 4433 3764 4449
rect 1772 4401 1972 4433
rect 2028 4401 2228 4433
rect 2284 4401 2484 4433
rect 2540 4401 2740 4433
rect 2796 4401 2996 4433
rect 3052 4401 3252 4433
rect 3308 4401 3508 4433
rect 3564 4401 3764 4433
rect 3820 4483 4020 4499
rect 3820 4449 3836 4483
rect 3870 4449 3970 4483
rect 4004 4449 4020 4483
rect 3820 4401 4020 4449
rect 4076 4483 4276 4499
rect 4076 4449 4092 4483
rect 4126 4449 4226 4483
rect 4260 4449 4276 4483
rect 4076 4401 4276 4449
rect 4332 4483 4532 4499
rect 4332 4449 4348 4483
rect 4382 4449 4482 4483
rect 4516 4449 4532 4483
rect 4332 4401 4532 4449
rect 4588 4483 6581 4499
rect 4588 4449 4604 4483
rect 4638 4449 4672 4483
rect 4706 4449 4740 4483
rect 4774 4449 4808 4483
rect 4842 4449 4876 4483
rect 4910 4449 4944 4483
rect 4978 4449 5013 4483
rect 5047 4449 5082 4483
rect 5116 4449 5151 4483
rect 5185 4449 5220 4483
rect 5254 4449 5289 4483
rect 5323 4449 5358 4483
rect 5392 4449 5427 4483
rect 5461 4449 5496 4483
rect 5530 4449 5565 4483
rect 5599 4449 5634 4483
rect 5668 4449 5703 4483
rect 5737 4449 5772 4483
rect 5806 4449 5841 4483
rect 5875 4449 5910 4483
rect 5944 4449 5979 4483
rect 6013 4449 6048 4483
rect 6082 4449 6117 4483
rect 6151 4449 6186 4483
rect 6220 4449 6255 4483
rect 6289 4449 6324 4483
rect 6358 4449 6393 4483
rect 6427 4449 6462 4483
rect 6496 4449 6531 4483
rect 6565 4449 6581 4483
rect 4588 4433 6581 4449
rect 6636 4483 7692 4499
rect 6636 4449 6652 4483
rect 6686 4449 6722 4483
rect 6756 4449 6792 4483
rect 6826 4449 6862 4483
rect 6896 4449 6932 4483
rect 6966 4449 7003 4483
rect 7037 4449 7074 4483
rect 7108 4449 7145 4483
rect 7179 4449 7216 4483
rect 7250 4449 7287 4483
rect 7321 4449 7358 4483
rect 7392 4449 7429 4483
rect 7463 4449 7500 4483
rect 7534 4449 7571 4483
rect 7605 4449 7642 4483
rect 7676 4449 7692 4483
rect 6636 4433 7692 4449
rect 4588 4401 4788 4433
rect 4844 4401 5044 4433
rect 5100 4401 5300 4433
rect 5356 4401 5556 4433
rect 5612 4401 5812 4433
rect 5868 4401 6068 4433
rect 6124 4401 6324 4433
rect 6380 4401 6580 4433
rect 6636 4401 6836 4433
rect 6892 4401 7692 4433
rect 916 4259 1716 4291
rect 1772 4259 1972 4291
rect 2028 4259 2228 4291
rect 2284 4259 2484 4291
rect 2540 4259 2740 4291
rect 2796 4259 2996 4291
rect 3052 4259 3252 4291
rect 3308 4259 3508 4291
rect 3564 4259 3764 4291
rect 3820 4259 4020 4291
rect 4076 4259 4276 4291
rect 4332 4259 4532 4291
rect 4588 4259 4788 4291
rect 4844 4259 5044 4291
rect 5100 4259 5300 4291
rect 5356 4259 5556 4291
rect 5612 4259 5812 4291
rect 5868 4259 6068 4291
rect 6124 4259 6324 4291
rect 6380 4259 6580 4291
rect 6636 4259 6836 4291
rect 6892 4259 7692 4291
rect 916 3809 1716 3841
rect 1772 3809 1972 3841
rect 2028 3809 2228 3841
rect 2284 3809 2484 3841
rect 2540 3809 2740 3841
rect 2796 3809 2996 3841
rect 3052 3809 3252 3841
rect 3308 3809 3508 3841
rect 3564 3809 3764 3841
rect 3820 3809 4020 3841
rect 4076 3809 4276 3841
rect 4332 3809 4532 3841
rect 4588 3809 4788 3841
rect 4844 3809 5044 3841
rect 5100 3809 5300 3841
rect 5356 3809 5556 3841
rect 5612 3809 5812 3841
rect 5868 3809 6068 3841
rect 6124 3809 6324 3841
rect 6380 3809 6580 3841
rect 6636 3809 6836 3841
rect 6892 3809 7692 3841
rect 916 3667 1716 3699
rect 1772 3667 1972 3699
rect 916 3651 1972 3667
rect 916 3617 932 3651
rect 966 3617 1003 3651
rect 1037 3617 1074 3651
rect 1108 3617 1145 3651
rect 1179 3617 1216 3651
rect 1250 3617 1287 3651
rect 1321 3617 1358 3651
rect 1392 3617 1429 3651
rect 1463 3617 1500 3651
rect 1534 3617 1571 3651
rect 1605 3617 1642 3651
rect 1676 3617 1712 3651
rect 1746 3617 1782 3651
rect 1816 3617 1852 3651
rect 1886 3617 1922 3651
rect 1956 3617 1972 3651
rect 916 3601 1972 3617
rect 2028 3667 2228 3699
rect 2284 3667 2484 3699
rect 2540 3667 2740 3699
rect 2796 3667 2996 3699
rect 3052 3667 3252 3699
rect 3308 3667 3508 3699
rect 3564 3667 3764 3699
rect 3820 3667 4020 3699
rect 2028 3651 4020 3667
rect 2028 3617 2044 3651
rect 2078 3617 2112 3651
rect 2146 3617 2180 3651
rect 2214 3617 2248 3651
rect 2282 3617 2316 3651
rect 2350 3617 2384 3651
rect 2418 3617 2452 3651
rect 2486 3617 2521 3651
rect 2555 3617 2590 3651
rect 2624 3617 2659 3651
rect 2693 3617 2728 3651
rect 2762 3617 2797 3651
rect 2831 3617 2866 3651
rect 2900 3617 2935 3651
rect 2969 3617 3004 3651
rect 3038 3617 3073 3651
rect 3107 3617 3142 3651
rect 3176 3617 3211 3651
rect 3245 3617 3280 3651
rect 3314 3617 3349 3651
rect 3383 3617 3418 3651
rect 3452 3617 3487 3651
rect 3521 3617 3556 3651
rect 3590 3617 3625 3651
rect 3659 3617 3694 3651
rect 3728 3617 3763 3651
rect 3797 3617 3832 3651
rect 3866 3617 3901 3651
rect 3935 3617 3970 3651
rect 4004 3617 4020 3651
rect 2028 3601 4020 3617
rect 4076 3651 4276 3699
rect 4076 3617 4092 3651
rect 4126 3617 4226 3651
rect 4260 3617 4276 3651
rect 4076 3601 4276 3617
rect 4332 3651 4532 3699
rect 4332 3617 4348 3651
rect 4382 3617 4482 3651
rect 4516 3617 4532 3651
rect 4332 3601 4532 3617
rect 4588 3651 4788 3699
rect 4588 3617 4604 3651
rect 4638 3617 4738 3651
rect 4772 3617 4788 3651
rect 4588 3601 4788 3617
rect 4844 3667 5044 3699
rect 5100 3667 5300 3699
rect 5356 3667 5556 3699
rect 5612 3667 5812 3699
rect 5868 3667 6068 3699
rect 6124 3667 6324 3699
rect 6380 3667 6580 3699
rect 4844 3651 6580 3667
rect 4844 3617 4860 3651
rect 4894 3617 4929 3651
rect 4963 3617 4998 3651
rect 5032 3617 5067 3651
rect 5101 3617 5136 3651
rect 5170 3617 5205 3651
rect 5239 3617 5274 3651
rect 5308 3617 5343 3651
rect 5377 3617 5412 3651
rect 5446 3617 5481 3651
rect 5515 3617 5550 3651
rect 5584 3617 5620 3651
rect 5654 3617 5690 3651
rect 5724 3617 5760 3651
rect 5794 3617 5830 3651
rect 5864 3617 5900 3651
rect 5934 3617 5970 3651
rect 6004 3617 6040 3651
rect 6074 3617 6110 3651
rect 6144 3617 6180 3651
rect 6214 3617 6250 3651
rect 6284 3617 6320 3651
rect 6354 3617 6390 3651
rect 6424 3617 6460 3651
rect 6494 3617 6530 3651
rect 6564 3617 6580 3651
rect 4844 3601 6580 3617
rect 6636 3667 6836 3699
rect 6892 3667 7692 3699
rect 6636 3651 7692 3667
rect 6636 3617 6652 3651
rect 6686 3617 6722 3651
rect 6756 3617 6792 3651
rect 6826 3617 6862 3651
rect 6896 3617 6932 3651
rect 6966 3617 7003 3651
rect 7037 3617 7074 3651
rect 7108 3617 7145 3651
rect 7179 3617 7216 3651
rect 7250 3617 7287 3651
rect 7321 3617 7358 3651
rect 7392 3617 7429 3651
rect 7463 3617 7500 3651
rect 7534 3617 7571 3651
rect 7605 3617 7642 3651
rect 7676 3617 7692 3651
rect 6636 3601 7692 3617
rect 916 3473 1716 3489
rect 916 3439 932 3473
rect 966 3439 1006 3473
rect 1040 3439 1080 3473
rect 1114 3439 1154 3473
rect 1188 3439 1228 3473
rect 1262 3439 1301 3473
rect 1335 3439 1374 3473
rect 1408 3439 1447 3473
rect 1481 3439 1520 3473
rect 1554 3439 1593 3473
rect 1627 3439 1666 3473
rect 1700 3439 1716 3473
rect 916 3391 1716 3439
rect 1772 3473 5044 3489
rect 1772 3439 1788 3473
rect 1822 3439 1856 3473
rect 1890 3439 1924 3473
rect 1958 3439 1992 3473
rect 2026 3439 2060 3473
rect 2094 3439 2128 3473
rect 2162 3439 2196 3473
rect 2230 3439 2264 3473
rect 2298 3439 2332 3473
rect 2366 3439 2400 3473
rect 2434 3439 2468 3473
rect 2502 3439 2536 3473
rect 2570 3439 2604 3473
rect 2638 3439 2672 3473
rect 2706 3439 2740 3473
rect 2774 3439 2808 3473
rect 2842 3439 2876 3473
rect 2910 3439 2944 3473
rect 2978 3439 3012 3473
rect 3046 3439 3080 3473
rect 3114 3439 3148 3473
rect 3182 3439 3216 3473
rect 3250 3439 3284 3473
rect 3318 3439 3352 3473
rect 3386 3439 3420 3473
rect 3454 3439 3488 3473
rect 3522 3439 3556 3473
rect 3590 3439 3624 3473
rect 3658 3439 3692 3473
rect 3726 3439 3760 3473
rect 3794 3439 3828 3473
rect 3862 3439 3896 3473
rect 3930 3439 3964 3473
rect 3998 3439 4032 3473
rect 4066 3439 4100 3473
rect 4134 3439 4168 3473
rect 4202 3439 4236 3473
rect 4270 3439 4304 3473
rect 4338 3439 4373 3473
rect 4407 3439 4442 3473
rect 4476 3439 4511 3473
rect 4545 3439 4580 3473
rect 4614 3439 4649 3473
rect 4683 3439 4718 3473
rect 4752 3439 4787 3473
rect 4821 3439 4856 3473
rect 4890 3439 4925 3473
rect 4959 3439 4994 3473
rect 5028 3439 5044 3473
rect 1772 3423 5044 3439
rect 1772 3391 1972 3423
rect 2028 3391 2228 3423
rect 2284 3391 2484 3423
rect 2540 3391 2740 3423
rect 2796 3391 2996 3423
rect 3052 3391 3252 3423
rect 3308 3391 3508 3423
rect 3564 3391 3764 3423
rect 3820 3391 4020 3423
rect 4076 3391 4276 3423
rect 4332 3391 4532 3423
rect 4588 3391 4788 3423
rect 4844 3391 5044 3423
rect 5100 3473 5556 3489
rect 5100 3439 5116 3473
rect 5150 3439 5194 3473
rect 5228 3439 5272 3473
rect 5306 3439 5350 3473
rect 5384 3439 5428 3473
rect 5462 3439 5506 3473
rect 5540 3439 5556 3473
rect 5100 3423 5556 3439
rect 5100 3391 5300 3423
rect 5356 3391 5556 3423
rect 5612 3473 6580 3489
rect 5612 3439 5628 3473
rect 5662 3439 5697 3473
rect 5731 3439 5766 3473
rect 5800 3439 5835 3473
rect 5869 3439 5904 3473
rect 5938 3439 5973 3473
rect 6007 3439 6042 3473
rect 6076 3439 6111 3473
rect 6145 3439 6180 3473
rect 6214 3439 6250 3473
rect 6284 3439 6320 3473
rect 6354 3439 6390 3473
rect 6424 3439 6460 3473
rect 6494 3439 6530 3473
rect 6564 3439 6580 3473
rect 5612 3423 6580 3439
rect 5612 3391 5812 3423
rect 5868 3391 6068 3423
rect 6124 3391 6324 3423
rect 6380 3391 6580 3423
rect 6636 3473 7692 3489
rect 6636 3439 6652 3473
rect 6686 3439 6722 3473
rect 6756 3439 6792 3473
rect 6826 3439 6862 3473
rect 6896 3439 6932 3473
rect 6966 3439 7003 3473
rect 7037 3439 7074 3473
rect 7108 3439 7145 3473
rect 7179 3439 7216 3473
rect 7250 3439 7287 3473
rect 7321 3439 7358 3473
rect 7392 3439 7429 3473
rect 7463 3439 7500 3473
rect 7534 3439 7571 3473
rect 7605 3439 7642 3473
rect 7676 3439 7692 3473
rect 6636 3423 7692 3439
rect 6636 3391 6836 3423
rect 6892 3391 7692 3423
rect 916 3249 1716 3281
rect 1772 3249 1972 3281
rect 2028 3249 2228 3281
rect 2284 3249 2484 3281
rect 2540 3249 2740 3281
rect 2796 3249 2996 3281
rect 3052 3249 3252 3281
rect 3308 3249 3508 3281
rect 3564 3249 3764 3281
rect 3820 3249 4020 3281
rect 4076 3249 4276 3281
rect 4332 3249 4532 3281
rect 4588 3249 4788 3281
rect 4844 3249 5044 3281
rect 5100 3249 5300 3281
rect 5356 3249 5556 3281
rect 5612 3249 5812 3281
rect 5868 3249 6068 3281
rect 6124 3249 6324 3281
rect 6380 3249 6580 3281
rect 6636 3249 6836 3281
rect 6892 3249 7692 3281
rect 8759 4804 8859 4836
rect 8915 4804 9015 4836
rect 9071 4804 9171 4836
rect 9227 4804 9327 4836
rect 9507 4804 9607 4836
rect 9787 4804 9887 4836
rect 9943 4804 10043 4836
rect 10376 4804 10476 4836
rect 10532 4804 10632 4836
rect 10688 4804 10788 4836
rect 10844 4804 10944 4836
rect 11000 4804 11100 4836
rect 8759 3772 8859 3804
rect 8915 3772 9015 3804
rect 8759 3756 9015 3772
rect 8759 3722 8775 3756
rect 8809 3722 8870 3756
rect 8904 3722 8965 3756
rect 8999 3722 9015 3756
rect 8759 3706 9015 3722
rect 9071 3772 9171 3804
rect 9227 3772 9327 3804
rect 9071 3756 9327 3772
rect 9071 3722 9087 3756
rect 9121 3722 9182 3756
rect 9216 3722 9277 3756
rect 9311 3722 9327 3756
rect 9071 3706 9327 3722
rect 9507 3736 9607 3804
rect 9507 3702 9541 3736
rect 9575 3702 9607 3736
rect 9787 3772 9887 3804
rect 9943 3772 10043 3804
rect 9787 3756 10043 3772
rect 9787 3722 9803 3756
rect 9837 3722 9898 3756
rect 9932 3722 9993 3756
rect 10027 3722 10043 3756
rect 9787 3706 10043 3722
rect 10376 3772 10476 3804
rect 10532 3772 10632 3804
rect 10688 3772 10788 3804
rect 10844 3772 10944 3804
rect 11000 3772 11100 3804
rect 10376 3756 11100 3772
rect 10376 3722 10392 3756
rect 10426 3722 10466 3756
rect 10500 3722 10539 3756
rect 10573 3722 10612 3756
rect 10646 3722 10685 3756
rect 10719 3722 10758 3756
rect 10792 3722 10831 3756
rect 10865 3722 10904 3756
rect 10938 3722 10977 3756
rect 11011 3722 11050 3756
rect 11084 3722 11100 3756
rect 10376 3706 11100 3722
rect 9507 3668 9607 3702
rect 9507 3634 9541 3668
rect 9575 3634 9607 3668
rect 9507 3618 9607 3634
rect 10624 3643 10824 3659
rect 10624 3609 10640 3643
rect 10674 3609 10774 3643
rect 10808 3609 10824 3643
rect 10624 3561 10824 3609
rect 8861 3364 8893 3464
rect 9893 3448 9991 3464
rect 9893 3414 9941 3448
rect 9975 3414 9991 3448
rect 10624 3445 10824 3477
rect 9893 3364 9991 3414
rect 9925 3353 9991 3364
rect 9925 3319 9941 3353
rect 9975 3319 9991 3353
rect 9925 3308 9991 3319
rect 8861 3208 8893 3308
rect 9893 3258 9991 3308
rect 9893 3224 9941 3258
rect 9975 3224 9991 3258
rect 9893 3208 9991 3224
rect 10054 3335 10120 3351
rect 10054 3301 10070 3335
rect 10104 3325 10120 3335
rect 10104 3301 10152 3325
rect 10054 3267 10152 3301
rect 10054 3233 10070 3267
rect 10104 3233 10152 3267
rect 10054 3225 10152 3233
rect 11152 3225 11184 3325
rect 10054 3217 10120 3225
rect 17843 3234 17943 3266
rect 17999 3234 18099 3266
rect 18327 3234 18427 3266
rect 18483 3234 18583 3266
rect 18789 3234 18889 3266
rect 18945 3234 19045 3266
rect 16939 3064 16971 3184
rect 17571 3168 17669 3184
rect 17571 3134 17619 3168
rect 17653 3134 17669 3168
rect 17571 3100 17669 3134
rect 17571 3066 17619 3100
rect 17653 3066 17669 3100
rect 17571 3064 17669 3066
rect 17603 3050 17669 3064
rect 17843 3002 17943 3034
rect 17999 3002 18099 3034
rect 18327 3002 18427 3034
rect 18483 3002 18583 3034
rect 18789 3002 18889 3034
rect 18945 3002 19045 3034
rect 1606 2388 1672 2397
rect 542 2288 574 2388
rect 1574 2381 1672 2388
rect 1574 2347 1622 2381
rect 1656 2347 1672 2381
rect 1574 2313 1672 2347
rect 1574 2288 1622 2313
rect 1606 2279 1622 2288
rect 1656 2279 1672 2313
rect 1606 2263 1672 2279
rect 7471 2092 7503 2192
rect 8503 2158 8689 2192
rect 8503 2124 8571 2158
rect 8605 2124 8639 2158
rect 8673 2124 8689 2158
rect 8503 2092 8689 2124
rect 2392 1912 2424 2092
rect 4424 2076 4522 2092
rect 4424 2042 4472 2076
rect 4506 2042 4522 2076
rect 4424 2008 4522 2042
rect 4424 1974 4472 2008
rect 4506 1974 4522 2008
rect 4424 1940 4522 1974
rect 4424 1912 4472 1940
rect 4456 1906 4472 1912
rect 4506 1906 4522 1940
rect 4456 1872 4522 1906
rect 4456 1856 4472 1872
rect 542 1696 574 1796
rect 1574 1780 1672 1796
rect 1574 1746 1622 1780
rect 1656 1746 1672 1780
rect 1574 1696 1672 1746
rect 1606 1685 1672 1696
rect 1606 1651 1622 1685
rect 1656 1651 1672 1685
rect 1606 1640 1672 1651
rect 542 1540 574 1640
rect 1574 1590 1672 1640
rect 1574 1556 1622 1590
rect 1656 1556 1672 1590
rect 1574 1540 1672 1556
rect 2392 1676 2424 1856
rect 4424 1838 4472 1856
rect 4506 1838 4522 1872
rect 4424 1804 4522 1838
rect 4424 1770 4472 1804
rect 4506 1770 4522 1804
rect 4424 1736 4522 1770
rect 4424 1702 4472 1736
rect 4506 1702 4522 1736
rect 4424 1676 4522 1702
rect 4564 2076 4662 2092
rect 4564 2042 4580 2076
rect 4614 2042 4662 2076
rect 4564 2006 4662 2042
rect 4564 1972 4580 2006
rect 4614 1972 4662 2006
rect 4564 1936 4662 1972
rect 4564 1902 4580 1936
rect 4614 1912 4662 1936
rect 6662 1912 6694 2092
rect 6874 1954 8474 1986
rect 4614 1902 4630 1912
rect 4564 1866 4630 1902
rect 4564 1832 4580 1866
rect 4614 1856 4630 1866
rect 4614 1832 4662 1856
rect 4564 1796 4662 1832
rect 4564 1762 4580 1796
rect 4614 1762 4662 1796
rect 4564 1726 4662 1762
rect 4564 1692 4580 1726
rect 4614 1692 4662 1726
rect 4564 1676 4662 1692
rect 6662 1676 6694 1856
rect 6874 1822 8474 1870
rect 6874 1788 6909 1822
rect 6943 1788 6977 1822
rect 7011 1788 7045 1822
rect 7079 1788 7113 1822
rect 7147 1788 7181 1822
rect 7215 1788 7249 1822
rect 7283 1788 7317 1822
rect 7351 1788 7385 1822
rect 7419 1788 7453 1822
rect 7487 1788 7521 1822
rect 7555 1788 7589 1822
rect 7623 1788 7657 1822
rect 7691 1788 7725 1822
rect 7759 1788 7793 1822
rect 7827 1788 7862 1822
rect 7896 1788 7931 1822
rect 7965 1788 8000 1822
rect 8034 1788 8069 1822
rect 8103 1788 8138 1822
rect 8172 1788 8207 1822
rect 8241 1788 8276 1822
rect 8310 1788 8345 1822
rect 8379 1788 8414 1822
rect 8448 1788 8474 1822
rect 6874 1740 8474 1788
rect 4456 1668 4522 1676
rect 4456 1634 4472 1668
rect 4506 1634 4522 1668
rect 4456 1620 4522 1634
rect 6874 1624 8474 1656
rect 2392 1440 2424 1620
rect 4424 1599 4522 1620
rect 4424 1565 4472 1599
rect 4506 1565 4522 1599
rect 4424 1530 4522 1565
rect 4424 1496 4472 1530
rect 4506 1496 4522 1530
rect 4424 1461 4522 1496
rect 17910 2802 18086 2838
rect 17910 2768 17932 2802
rect 17966 2768 18000 2802
rect 18034 2768 18086 2802
rect 17910 2738 18086 2768
rect 19086 2738 19118 2838
rect 4424 1440 4472 1461
rect 4456 1427 4472 1440
rect 4506 1427 4522 1461
rect 7469 1473 7843 1489
rect 7469 1439 7485 1473
rect 7519 1439 7562 1473
rect 7596 1439 7639 1473
rect 7673 1439 7716 1473
rect 7750 1439 7793 1473
rect 7827 1439 7843 1473
rect 4456 1392 4522 1427
rect 4456 1384 4472 1392
rect 542 1134 574 1234
rect 1574 1218 1672 1234
rect 1574 1184 1622 1218
rect 1656 1184 1672 1218
rect 1574 1134 1672 1184
rect 1606 1123 1672 1134
rect 1606 1089 1622 1123
rect 1656 1089 1672 1123
rect 1606 1078 1672 1089
rect 542 978 574 1078
rect 1574 1028 1672 1078
rect 1574 994 1622 1028
rect 1656 994 1672 1028
rect 1574 978 1672 994
rect 2392 1204 2424 1384
rect 4424 1358 4472 1384
rect 4506 1358 4522 1392
rect 7469 1423 7843 1439
rect 7469 1391 7499 1423
rect 7555 1391 7585 1423
rect 7641 1391 7671 1423
rect 7727 1391 7757 1423
rect 7813 1391 7843 1423
rect 4424 1323 4522 1358
rect 4424 1289 4472 1323
rect 4506 1289 4522 1323
rect 4424 1254 4522 1289
rect 4424 1220 4472 1254
rect 4506 1220 4522 1254
rect 4424 1204 4522 1220
rect 4564 1368 4662 1384
rect 4564 1334 4580 1368
rect 4614 1334 4662 1368
rect 4564 1254 4662 1334
rect 4564 1220 4580 1254
rect 4614 1220 4662 1254
rect 4564 1204 4662 1220
rect 6662 1204 6694 1384
rect 2451 1098 3019 1114
rect 2451 1064 2467 1098
rect 2501 1064 2539 1098
rect 2573 1064 2611 1098
rect 2645 1064 2683 1098
rect 2717 1064 2755 1098
rect 2789 1064 2827 1098
rect 2861 1064 2898 1098
rect 2932 1064 2969 1098
rect 3003 1064 3019 1098
rect 2451 1048 3019 1064
rect 2451 1016 2551 1048
rect 2607 1016 2707 1048
rect 2763 1016 2863 1048
rect 2919 1016 3019 1048
rect 3075 1098 3643 1114
rect 3075 1064 3091 1098
rect 3125 1064 3162 1098
rect 3196 1064 3233 1098
rect 3267 1064 3305 1098
rect 3339 1064 3377 1098
rect 3411 1064 3449 1098
rect 3483 1064 3521 1098
rect 3555 1064 3593 1098
rect 3627 1064 3643 1098
rect 3075 1048 3643 1064
rect 3075 1016 3175 1048
rect 3231 1016 3331 1048
rect 3387 1016 3487 1048
rect 3543 1016 3643 1048
rect 3823 1098 4079 1114
rect 3823 1064 3839 1098
rect 3873 1064 3934 1098
rect 3968 1064 4029 1098
rect 4063 1064 4079 1098
rect 3823 1048 4079 1064
rect 3823 1016 3923 1048
rect 3979 1016 4079 1048
rect 4135 1098 4391 1114
rect 4135 1064 4151 1098
rect 4185 1064 4246 1098
rect 4280 1064 4341 1098
rect 4375 1064 4391 1098
rect 4135 1048 4391 1064
rect 4135 1016 4235 1048
rect 4291 1016 4391 1048
rect 4447 1098 4547 1114
rect 4447 1064 4463 1098
rect 4497 1064 4547 1098
rect 4447 1016 4547 1064
rect 4603 1098 4859 1114
rect 4603 1064 4619 1098
rect 4653 1064 4714 1098
rect 4748 1064 4809 1098
rect 4843 1064 4859 1098
rect 4603 1048 4859 1064
rect 4603 1016 4703 1048
rect 4759 1016 4859 1048
rect 4915 1098 5015 1114
rect 4915 1064 4931 1098
rect 4965 1064 5015 1098
rect 4915 1016 5015 1064
rect 5071 1098 5483 1114
rect 5071 1064 5087 1098
rect 5121 1064 5157 1098
rect 5191 1064 5226 1098
rect 5260 1064 5295 1098
rect 5329 1064 5364 1098
rect 5398 1064 5433 1098
rect 5467 1064 5483 1098
rect 5071 1048 5483 1064
rect 5071 1016 5171 1048
rect 5227 1016 5327 1048
rect 5383 1016 5483 1048
rect 5713 1098 5969 1114
rect 5713 1064 5729 1098
rect 5763 1064 5824 1098
rect 5858 1064 5919 1098
rect 5953 1064 5969 1098
rect 5713 1048 5969 1064
rect 5713 1016 5813 1048
rect 5869 1016 5969 1048
rect 6025 1098 6281 1114
rect 6025 1064 6041 1098
rect 6075 1064 6136 1098
rect 6170 1064 6231 1098
rect 6265 1064 6281 1098
rect 6025 1048 6281 1064
rect 6445 1098 6841 1114
rect 6445 1064 6461 1098
rect 6495 1064 6544 1098
rect 6578 1064 6627 1098
rect 6661 1064 6709 1098
rect 6743 1064 6791 1098
rect 6825 1064 6841 1098
rect 6445 1048 6841 1064
rect 6025 1016 6125 1048
rect 6181 1016 6281 1048
rect 6461 1016 6561 1048
rect 6741 1016 6841 1048
rect 6897 1098 7033 1114
rect 6897 1064 6913 1098
rect 6947 1064 6983 1098
rect 7017 1064 7033 1098
rect 6897 1048 7033 1064
rect 6897 1016 6997 1048
rect 542 822 574 922
rect 1574 872 1740 922
rect 1574 838 1622 872
rect 1656 838 1690 872
rect 1724 838 1740 872
rect 1574 822 1740 838
rect 542 666 574 766
rect 1574 750 1672 766
rect 1574 716 1622 750
rect 1656 716 1672 750
rect 1574 666 1672 716
rect 1606 655 1672 666
rect 1606 621 1622 655
rect 1656 621 1672 655
rect 1606 610 1672 621
rect 542 510 574 610
rect 1574 560 1672 610
rect 1574 526 1622 560
rect 1656 526 1672 560
rect 1574 510 1672 526
rect 542 354 574 454
rect 1574 404 1740 454
rect 1574 370 1622 404
rect 1656 370 1690 404
rect 1724 370 1740 404
rect 1574 354 1740 370
rect 542 198 574 298
rect 1574 282 1672 298
rect 1574 248 1622 282
rect 1656 248 1672 282
rect 1574 198 1672 248
rect 1606 187 1672 198
rect 1606 153 1622 187
rect 1656 153 1672 187
rect 1606 142 1672 153
rect 542 42 574 142
rect 1574 92 1672 142
rect 1574 58 1622 92
rect 1656 58 1672 92
rect 1574 42 1672 58
rect 542 -114 574 -14
rect 1574 -64 1740 -14
rect 1574 -98 1622 -64
rect 1656 -98 1690 -64
rect 1724 -98 1740 -64
rect 1574 -114 1740 -98
rect 2451 -16 2551 16
rect 2607 -16 2707 16
rect 2763 -16 2863 16
rect 2919 -16 3019 16
rect 3075 -16 3175 16
rect 3231 -16 3331 16
rect 3387 -16 3487 16
rect 3543 -16 3643 16
rect 3823 -16 3923 16
rect 3979 -16 4079 16
rect 4135 -16 4235 16
rect 4291 -16 4391 16
rect 4447 -16 4547 16
rect 4603 -16 4703 16
rect 4759 -16 4859 16
rect 4915 -16 5015 16
rect 5071 -16 5171 16
rect 5227 -16 5327 16
rect 5383 -16 5483 16
rect 5713 -16 5813 16
rect 5869 -16 5969 16
rect 6025 -16 6125 16
rect 6181 -16 6281 16
rect 6461 -16 6561 16
rect 6741 -16 6841 16
rect 6897 -16 6997 16
rect 8329 1030 8897 1046
rect 8329 996 8345 1030
rect 8379 996 8416 1030
rect 8450 996 8487 1030
rect 8521 996 8559 1030
rect 8593 996 8631 1030
rect 8665 996 8703 1030
rect 8737 996 8775 1030
rect 8809 996 8847 1030
rect 8881 996 8897 1030
rect 8329 980 8897 996
rect 8329 948 8429 980
rect 8485 948 8585 980
rect 8641 948 8741 980
rect 8797 948 8897 980
rect 8953 1030 9677 1046
rect 8953 996 8969 1030
rect 9003 996 9043 1030
rect 9077 996 9116 1030
rect 9150 996 9189 1030
rect 9223 996 9262 1030
rect 9296 996 9335 1030
rect 9369 996 9408 1030
rect 9442 996 9481 1030
rect 9515 996 9554 1030
rect 9588 996 9627 1030
rect 9661 996 9677 1030
rect 8953 980 9677 996
rect 8953 948 9053 980
rect 9109 948 9209 980
rect 9265 948 9365 980
rect 9421 948 9521 980
rect 9577 948 9677 980
rect 9733 1030 10457 1046
rect 9733 996 9749 1030
rect 9783 996 9822 1030
rect 9856 996 9895 1030
rect 9929 996 9968 1030
rect 10002 996 10041 1030
rect 10075 996 10114 1030
rect 10148 996 10187 1030
rect 10221 996 10260 1030
rect 10294 996 10333 1030
rect 10367 996 10407 1030
rect 10441 996 10457 1030
rect 9733 980 10457 996
rect 10788 1030 12550 1046
rect 10788 996 10804 1030
rect 10838 996 10875 1030
rect 10909 996 10946 1030
rect 10980 996 11017 1030
rect 11051 996 11088 1030
rect 11122 996 11159 1030
rect 11193 996 11230 1030
rect 11264 996 11301 1030
rect 11335 996 11372 1030
rect 11406 996 11443 1030
rect 11477 996 11514 1030
rect 11548 996 11585 1030
rect 11619 996 11656 1030
rect 11690 996 11727 1030
rect 11761 996 11798 1030
rect 11832 996 11869 1030
rect 11903 996 11940 1030
rect 11974 996 12010 1030
rect 12044 996 12080 1030
rect 12114 996 12150 1030
rect 12184 996 12220 1030
rect 12254 996 12290 1030
rect 12324 996 12360 1030
rect 12394 996 12430 1030
rect 12464 996 12500 1030
rect 12534 996 12550 1030
rect 10788 980 12550 996
rect 9733 948 9833 980
rect 9889 948 9989 980
rect 10045 948 10145 980
rect 10201 948 10301 980
rect 10357 948 10457 980
rect 10782 948 11182 980
rect 11238 948 11638 980
rect 11694 948 12094 980
rect 12150 948 12550 980
rect 12828 1030 12962 1046
rect 12828 996 12844 1030
rect 12878 996 12912 1030
rect 12946 996 12962 1030
rect 15268 1034 15448 1066
rect 15504 1034 15684 1066
rect 15740 1034 15920 1066
rect 15976 1034 16156 1066
rect 12828 980 12962 996
rect 12828 948 12948 980
rect 7469 -41 7499 -9
rect 7555 -41 7585 -9
rect 7641 -41 7671 -9
rect 7727 -41 7757 -9
rect 7813 -41 7843 -9
rect 13044 844 13076 1024
rect 15076 1008 15174 1024
rect 15076 974 15124 1008
rect 15158 974 15174 1008
rect 15076 940 15174 974
rect 15076 906 15124 940
rect 15158 906 15174 940
rect 15076 872 15174 906
rect 15076 844 15124 872
rect 15108 838 15124 844
rect 15158 838 15174 872
rect 15108 804 15174 838
rect 15108 788 15124 804
rect 12828 716 12948 748
rect 13044 608 13076 788
rect 15076 770 15124 788
rect 15158 770 15174 804
rect 15076 736 15174 770
rect 15076 702 15124 736
rect 15158 702 15174 736
rect 15076 668 15174 702
rect 15268 802 15448 834
rect 15504 802 15684 834
rect 15740 802 15920 834
rect 15976 802 16156 834
rect 15268 778 16156 802
rect 15268 744 15284 778
rect 15318 744 15353 778
rect 15387 744 15422 778
rect 15456 744 15491 778
rect 15525 744 15560 778
rect 15594 744 15629 778
rect 15663 744 15698 778
rect 15732 744 15766 778
rect 15800 744 15834 778
rect 15868 744 15902 778
rect 15936 744 15970 778
rect 16004 744 16038 778
rect 16072 744 16106 778
rect 16140 744 16156 778
rect 15268 711 16156 744
rect 15268 679 15448 711
rect 15504 679 15684 711
rect 15740 679 15920 711
rect 15976 679 16156 711
rect 15076 634 15124 668
rect 15158 634 15174 668
rect 15076 608 15174 634
rect 15108 599 15174 608
rect 15108 565 15124 599
rect 15158 565 15174 599
rect 15108 552 15174 565
rect 13044 372 13076 552
rect 15076 530 15174 552
rect 15076 496 15124 530
rect 15158 496 15174 530
rect 15076 461 15174 496
rect 15076 427 15124 461
rect 15158 427 15174 461
rect 15076 392 15174 427
rect 15076 372 15124 392
rect 15108 358 15124 372
rect 15158 358 15174 392
rect 15108 323 15174 358
rect 15108 316 15124 323
rect 13044 136 13076 316
rect 15076 289 15124 316
rect 15158 289 15174 323
rect 15268 447 15448 479
rect 15504 447 15684 479
rect 15740 447 15920 479
rect 15976 447 16156 479
rect 15268 398 16156 447
rect 15268 364 15284 398
rect 15318 364 15353 398
rect 15387 364 15422 398
rect 15456 364 15491 398
rect 15525 364 15560 398
rect 15594 364 15629 398
rect 15663 364 15698 398
rect 15732 364 15766 398
rect 15800 364 15834 398
rect 15868 364 15902 398
rect 15936 364 15970 398
rect 16004 364 16038 398
rect 16072 364 16106 398
rect 16140 364 16156 398
rect 15268 326 16156 364
rect 15268 294 15448 326
rect 15504 294 15684 326
rect 15076 254 15174 289
rect 15076 220 15124 254
rect 15158 220 15174 254
rect 15076 185 15174 220
rect 15076 151 15124 185
rect 15158 151 15174 185
rect 15076 136 15174 151
rect 15108 135 15174 136
rect 15895 259 16029 275
rect 15895 225 15911 259
rect 15945 225 15979 259
rect 16013 225 16029 259
rect 15895 209 16029 225
rect 15929 177 16029 209
rect 16085 259 16219 275
rect 16085 225 16101 259
rect 16135 225 16169 259
rect 16203 225 16219 259
rect 16085 209 16219 225
rect 16085 177 16185 209
rect 18370 193 18396 293
rect 18596 257 18766 293
rect 18596 223 18644 257
rect 18678 223 18712 257
rect 18746 223 18766 257
rect 18596 193 18766 223
rect 15268 62 15448 94
rect 15504 62 15684 94
rect 8329 -84 8429 -52
rect 8485 -84 8585 -52
rect 8641 -84 8741 -52
rect 8797 -84 8897 -52
rect 8953 -84 9053 -52
rect 9109 -84 9209 -52
rect 9265 -84 9365 -52
rect 9421 -84 9521 -52
rect 9577 -84 9677 -52
rect 9733 -84 9833 -52
rect 9889 -84 9989 -52
rect 10045 -84 10145 -52
rect 10201 -84 10301 -52
rect 10357 -84 10457 -52
rect 10782 -84 11182 -52
rect 11238 -84 11638 -52
rect 11694 -84 12094 -52
rect 12150 -84 12550 -52
rect 542 -270 574 -170
rect 1574 -186 1672 -170
rect 1574 -220 1622 -186
rect 1656 -220 1672 -186
rect 1574 -270 1672 -220
rect 1606 -281 1672 -270
rect 1606 -315 1622 -281
rect 1656 -315 1672 -281
rect 1606 -326 1672 -315
rect 542 -426 574 -326
rect 1574 -376 1672 -326
rect 1574 -410 1622 -376
rect 1656 -410 1672 -376
rect 1574 -426 1672 -410
rect 542 -582 574 -482
rect 1574 -532 1740 -482
rect 1574 -566 1622 -532
rect 1656 -566 1690 -532
rect 1724 -566 1740 -532
rect 1574 -582 1740 -566
rect 542 -738 574 -638
rect 1574 -688 1740 -638
rect 1574 -722 1622 -688
rect 1656 -722 1690 -688
rect 1724 -722 1740 -688
rect 1574 -738 1740 -722
rect 542 -1179 574 -1079
rect 1574 -1095 1672 -1079
rect 1574 -1129 1622 -1095
rect 1656 -1129 1672 -1095
rect 1574 -1179 1672 -1129
rect 1606 -1190 1672 -1179
rect 1606 -1224 1622 -1190
rect 1656 -1224 1672 -1190
rect 1606 -1235 1672 -1224
rect 18370 37 18396 137
rect 18596 105 18766 137
rect 18596 71 18644 105
rect 18678 71 18712 105
rect 18746 71 18766 105
rect 18596 37 18766 71
rect 15929 -855 16029 -823
rect 16085 -855 16185 -823
rect 542 -1335 574 -1235
rect 1574 -1285 1672 -1235
rect 1574 -1319 1622 -1285
rect 1656 -1319 1672 -1285
rect 1574 -1335 1672 -1319
rect 542 -1491 574 -1391
rect 1574 -1407 1672 -1391
rect 1574 -1441 1622 -1407
rect 1656 -1441 1672 -1407
rect 1574 -1491 1672 -1441
rect 1606 -1502 1672 -1491
rect 1606 -1536 1622 -1502
rect 1656 -1536 1672 -1502
rect 1606 -1547 1672 -1536
rect 542 -1647 574 -1547
rect 1574 -1597 1672 -1547
rect 1574 -1631 1622 -1597
rect 1656 -1631 1672 -1597
rect 1574 -1647 1672 -1631
rect 542 -1803 574 -1703
rect 1574 -1719 1672 -1703
rect 1574 -1753 1622 -1719
rect 1656 -1753 1672 -1719
rect 1574 -1803 1672 -1753
rect 1606 -1814 1672 -1803
rect 1606 -1848 1622 -1814
rect 1656 -1848 1672 -1814
rect 1606 -1859 1672 -1848
rect 542 -1959 574 -1859
rect 1574 -1909 1672 -1859
rect 1574 -1943 1622 -1909
rect 1656 -1943 1672 -1909
rect 1574 -1959 1672 -1943
rect 542 -2115 574 -2015
rect 1574 -2031 1672 -2015
rect 1574 -2065 1622 -2031
rect 1656 -2065 1672 -2031
rect 1574 -2115 1672 -2065
rect 1606 -2126 1672 -2115
rect 1606 -2160 1622 -2126
rect 1656 -2160 1672 -2126
rect 1606 -2171 1672 -2160
rect 542 -2271 574 -2171
rect 1574 -2221 1672 -2171
rect 1574 -2255 1622 -2221
rect 1656 -2255 1672 -2221
rect 1574 -2271 1672 -2255
rect 2669 -9584 2769 -9552
rect 2825 -9584 2925 -9552
rect 2669 -10216 2769 -10184
rect 2825 -10216 2925 -10184
rect 2669 -10232 2925 -10216
rect 2669 -10266 2685 -10232
rect 2719 -10266 2780 -10232
rect 2814 -10266 2875 -10232
rect 2909 -10266 2925 -10232
rect 2669 -10282 2925 -10266
rect 18870 -11617 18924 -11593
rect 18904 -11651 18924 -11617
rect 18870 -11685 18924 -11651
rect 18904 -11719 18924 -11685
rect 18870 -11743 18924 -11719
rect 18874 -12867 18924 -12843
rect 18908 -12901 18924 -12867
rect 18874 -12935 18924 -12901
rect 18908 -12969 18924 -12935
rect 18874 -12993 18924 -12969
rect 3068 -17018 3324 -17002
rect 3068 -17052 3084 -17018
rect 3118 -17052 3179 -17018
rect 3213 -17052 3274 -17018
rect 3308 -17052 3324 -17018
rect 3068 -17068 3324 -17052
rect 3068 -17100 3168 -17068
rect 3224 -17100 3324 -17068
rect 3068 -17732 3168 -17700
rect 3224 -17732 3324 -17700
rect 2625 -17833 2881 -17817
rect 2625 -17867 2641 -17833
rect 2675 -17867 2736 -17833
rect 2770 -17867 2831 -17833
rect 2865 -17867 2881 -17833
rect 2625 -17883 2881 -17867
rect 2625 -17915 2725 -17883
rect 2781 -17915 2881 -17883
rect 2625 -18947 2725 -18915
rect 2781 -18947 2881 -18915
<< polycont >>
rect 932 4627 966 4661
rect 1003 4627 1037 4661
rect 1074 4627 1108 4661
rect 1145 4627 1179 4661
rect 1216 4627 1250 4661
rect 1287 4627 1321 4661
rect 1358 4627 1392 4661
rect 1429 4627 1463 4661
rect 1500 4627 1534 4661
rect 1571 4627 1605 4661
rect 1642 4627 1676 4661
rect 1712 4627 1746 4661
rect 1782 4627 1816 4661
rect 1852 4627 1886 4661
rect 1922 4627 1956 4661
rect 2044 4627 2078 4661
rect 2112 4627 2146 4661
rect 2180 4627 2214 4661
rect 2248 4627 2282 4661
rect 2316 4627 2350 4661
rect 2384 4627 2418 4661
rect 2452 4627 2486 4661
rect 2520 4627 2554 4661
rect 2588 4627 2622 4661
rect 2656 4627 2690 4661
rect 2724 4627 2758 4661
rect 2792 4627 2826 4661
rect 2860 4627 2894 4661
rect 2928 4627 2962 4661
rect 2996 4627 3030 4661
rect 3064 4627 3098 4661
rect 3133 4627 3167 4661
rect 3202 4627 3236 4661
rect 3324 4627 3358 4661
rect 3458 4627 3492 4661
rect 3580 4627 3614 4661
rect 3648 4627 3682 4661
rect 3716 4627 3750 4661
rect 3784 4627 3818 4661
rect 3852 4627 3886 4661
rect 3920 4627 3954 4661
rect 3988 4627 4022 4661
rect 4056 4627 4090 4661
rect 4124 4627 4158 4661
rect 4192 4627 4226 4661
rect 4260 4627 4294 4661
rect 4328 4627 4362 4661
rect 4396 4627 4430 4661
rect 4464 4627 4498 4661
rect 4532 4627 4566 4661
rect 4600 4627 4634 4661
rect 4668 4627 4702 4661
rect 4736 4627 4770 4661
rect 4804 4627 4838 4661
rect 4872 4627 4906 4661
rect 4940 4627 4974 4661
rect 5008 4627 5042 4661
rect 5076 4627 5110 4661
rect 5144 4627 5178 4661
rect 5212 4627 5246 4661
rect 5280 4627 5314 4661
rect 5348 4627 5382 4661
rect 5416 4627 5450 4661
rect 5484 4627 5518 4661
rect 5552 4627 5586 4661
rect 5620 4627 5654 4661
rect 5688 4627 5722 4661
rect 5756 4627 5790 4661
rect 5824 4627 5858 4661
rect 5892 4627 5926 4661
rect 5960 4627 5994 4661
rect 6028 4627 6062 4661
rect 6096 4627 6130 4661
rect 6165 4627 6199 4661
rect 6234 4627 6268 4661
rect 6303 4627 6337 4661
rect 6372 4627 6406 4661
rect 6441 4627 6475 4661
rect 6510 4627 6544 4661
rect 6579 4627 6613 4661
rect 6648 4627 6682 4661
rect 6717 4627 6751 4661
rect 6786 4627 6820 4661
rect 7010 4627 7044 4661
rect 7080 4627 7114 4661
rect 7150 4627 7184 4661
rect 7220 4627 7254 4661
rect 7290 4627 7324 4661
rect 7360 4627 7394 4661
rect 7430 4627 7464 4661
rect 7500 4627 7534 4661
rect 7571 4627 7605 4661
rect 7642 4627 7676 4661
rect 932 4449 966 4483
rect 1006 4449 1040 4483
rect 1080 4449 1114 4483
rect 1154 4449 1188 4483
rect 1228 4449 1262 4483
rect 1301 4449 1335 4483
rect 1374 4449 1408 4483
rect 1447 4449 1481 4483
rect 1520 4449 1554 4483
rect 1593 4449 1627 4483
rect 1666 4449 1700 4483
rect 1788 4449 1822 4483
rect 1856 4449 1890 4483
rect 1924 4449 1958 4483
rect 1992 4449 2026 4483
rect 2060 4449 2094 4483
rect 2128 4449 2162 4483
rect 2196 4449 2230 4483
rect 2265 4449 2299 4483
rect 2334 4449 2368 4483
rect 2403 4449 2437 4483
rect 2472 4449 2506 4483
rect 2541 4449 2575 4483
rect 2610 4449 2644 4483
rect 2679 4449 2713 4483
rect 2748 4449 2782 4483
rect 2817 4449 2851 4483
rect 2886 4449 2920 4483
rect 2955 4449 2989 4483
rect 3024 4449 3058 4483
rect 3093 4449 3127 4483
rect 3162 4449 3196 4483
rect 3231 4449 3265 4483
rect 3300 4449 3334 4483
rect 3369 4449 3403 4483
rect 3438 4449 3472 4483
rect 3507 4449 3541 4483
rect 3576 4449 3610 4483
rect 3645 4449 3679 4483
rect 3714 4449 3748 4483
rect 3836 4449 3870 4483
rect 3970 4449 4004 4483
rect 4092 4449 4126 4483
rect 4226 4449 4260 4483
rect 4348 4449 4382 4483
rect 4482 4449 4516 4483
rect 4604 4449 4638 4483
rect 4672 4449 4706 4483
rect 4740 4449 4774 4483
rect 4808 4449 4842 4483
rect 4876 4449 4910 4483
rect 4944 4449 4978 4483
rect 5013 4449 5047 4483
rect 5082 4449 5116 4483
rect 5151 4449 5185 4483
rect 5220 4449 5254 4483
rect 5289 4449 5323 4483
rect 5358 4449 5392 4483
rect 5427 4449 5461 4483
rect 5496 4449 5530 4483
rect 5565 4449 5599 4483
rect 5634 4449 5668 4483
rect 5703 4449 5737 4483
rect 5772 4449 5806 4483
rect 5841 4449 5875 4483
rect 5910 4449 5944 4483
rect 5979 4449 6013 4483
rect 6048 4449 6082 4483
rect 6117 4449 6151 4483
rect 6186 4449 6220 4483
rect 6255 4449 6289 4483
rect 6324 4449 6358 4483
rect 6393 4449 6427 4483
rect 6462 4449 6496 4483
rect 6531 4449 6565 4483
rect 6652 4449 6686 4483
rect 6722 4449 6756 4483
rect 6792 4449 6826 4483
rect 6862 4449 6896 4483
rect 6932 4449 6966 4483
rect 7003 4449 7037 4483
rect 7074 4449 7108 4483
rect 7145 4449 7179 4483
rect 7216 4449 7250 4483
rect 7287 4449 7321 4483
rect 7358 4449 7392 4483
rect 7429 4449 7463 4483
rect 7500 4449 7534 4483
rect 7571 4449 7605 4483
rect 7642 4449 7676 4483
rect 932 3617 966 3651
rect 1003 3617 1037 3651
rect 1074 3617 1108 3651
rect 1145 3617 1179 3651
rect 1216 3617 1250 3651
rect 1287 3617 1321 3651
rect 1358 3617 1392 3651
rect 1429 3617 1463 3651
rect 1500 3617 1534 3651
rect 1571 3617 1605 3651
rect 1642 3617 1676 3651
rect 1712 3617 1746 3651
rect 1782 3617 1816 3651
rect 1852 3617 1886 3651
rect 1922 3617 1956 3651
rect 2044 3617 2078 3651
rect 2112 3617 2146 3651
rect 2180 3617 2214 3651
rect 2248 3617 2282 3651
rect 2316 3617 2350 3651
rect 2384 3617 2418 3651
rect 2452 3617 2486 3651
rect 2521 3617 2555 3651
rect 2590 3617 2624 3651
rect 2659 3617 2693 3651
rect 2728 3617 2762 3651
rect 2797 3617 2831 3651
rect 2866 3617 2900 3651
rect 2935 3617 2969 3651
rect 3004 3617 3038 3651
rect 3073 3617 3107 3651
rect 3142 3617 3176 3651
rect 3211 3617 3245 3651
rect 3280 3617 3314 3651
rect 3349 3617 3383 3651
rect 3418 3617 3452 3651
rect 3487 3617 3521 3651
rect 3556 3617 3590 3651
rect 3625 3617 3659 3651
rect 3694 3617 3728 3651
rect 3763 3617 3797 3651
rect 3832 3617 3866 3651
rect 3901 3617 3935 3651
rect 3970 3617 4004 3651
rect 4092 3617 4126 3651
rect 4226 3617 4260 3651
rect 4348 3617 4382 3651
rect 4482 3617 4516 3651
rect 4604 3617 4638 3651
rect 4738 3617 4772 3651
rect 4860 3617 4894 3651
rect 4929 3617 4963 3651
rect 4998 3617 5032 3651
rect 5067 3617 5101 3651
rect 5136 3617 5170 3651
rect 5205 3617 5239 3651
rect 5274 3617 5308 3651
rect 5343 3617 5377 3651
rect 5412 3617 5446 3651
rect 5481 3617 5515 3651
rect 5550 3617 5584 3651
rect 5620 3617 5654 3651
rect 5690 3617 5724 3651
rect 5760 3617 5794 3651
rect 5830 3617 5864 3651
rect 5900 3617 5934 3651
rect 5970 3617 6004 3651
rect 6040 3617 6074 3651
rect 6110 3617 6144 3651
rect 6180 3617 6214 3651
rect 6250 3617 6284 3651
rect 6320 3617 6354 3651
rect 6390 3617 6424 3651
rect 6460 3617 6494 3651
rect 6530 3617 6564 3651
rect 6652 3617 6686 3651
rect 6722 3617 6756 3651
rect 6792 3617 6826 3651
rect 6862 3617 6896 3651
rect 6932 3617 6966 3651
rect 7003 3617 7037 3651
rect 7074 3617 7108 3651
rect 7145 3617 7179 3651
rect 7216 3617 7250 3651
rect 7287 3617 7321 3651
rect 7358 3617 7392 3651
rect 7429 3617 7463 3651
rect 7500 3617 7534 3651
rect 7571 3617 7605 3651
rect 7642 3617 7676 3651
rect 932 3439 966 3473
rect 1006 3439 1040 3473
rect 1080 3439 1114 3473
rect 1154 3439 1188 3473
rect 1228 3439 1262 3473
rect 1301 3439 1335 3473
rect 1374 3439 1408 3473
rect 1447 3439 1481 3473
rect 1520 3439 1554 3473
rect 1593 3439 1627 3473
rect 1666 3439 1700 3473
rect 1788 3439 1822 3473
rect 1856 3439 1890 3473
rect 1924 3439 1958 3473
rect 1992 3439 2026 3473
rect 2060 3439 2094 3473
rect 2128 3439 2162 3473
rect 2196 3439 2230 3473
rect 2264 3439 2298 3473
rect 2332 3439 2366 3473
rect 2400 3439 2434 3473
rect 2468 3439 2502 3473
rect 2536 3439 2570 3473
rect 2604 3439 2638 3473
rect 2672 3439 2706 3473
rect 2740 3439 2774 3473
rect 2808 3439 2842 3473
rect 2876 3439 2910 3473
rect 2944 3439 2978 3473
rect 3012 3439 3046 3473
rect 3080 3439 3114 3473
rect 3148 3439 3182 3473
rect 3216 3439 3250 3473
rect 3284 3439 3318 3473
rect 3352 3439 3386 3473
rect 3420 3439 3454 3473
rect 3488 3439 3522 3473
rect 3556 3439 3590 3473
rect 3624 3439 3658 3473
rect 3692 3439 3726 3473
rect 3760 3439 3794 3473
rect 3828 3439 3862 3473
rect 3896 3439 3930 3473
rect 3964 3439 3998 3473
rect 4032 3439 4066 3473
rect 4100 3439 4134 3473
rect 4168 3439 4202 3473
rect 4236 3439 4270 3473
rect 4304 3439 4338 3473
rect 4373 3439 4407 3473
rect 4442 3439 4476 3473
rect 4511 3439 4545 3473
rect 4580 3439 4614 3473
rect 4649 3439 4683 3473
rect 4718 3439 4752 3473
rect 4787 3439 4821 3473
rect 4856 3439 4890 3473
rect 4925 3439 4959 3473
rect 4994 3439 5028 3473
rect 5116 3439 5150 3473
rect 5194 3439 5228 3473
rect 5272 3439 5306 3473
rect 5350 3439 5384 3473
rect 5428 3439 5462 3473
rect 5506 3439 5540 3473
rect 5628 3439 5662 3473
rect 5697 3439 5731 3473
rect 5766 3439 5800 3473
rect 5835 3439 5869 3473
rect 5904 3439 5938 3473
rect 5973 3439 6007 3473
rect 6042 3439 6076 3473
rect 6111 3439 6145 3473
rect 6180 3439 6214 3473
rect 6250 3439 6284 3473
rect 6320 3439 6354 3473
rect 6390 3439 6424 3473
rect 6460 3439 6494 3473
rect 6530 3439 6564 3473
rect 6652 3439 6686 3473
rect 6722 3439 6756 3473
rect 6792 3439 6826 3473
rect 6862 3439 6896 3473
rect 6932 3439 6966 3473
rect 7003 3439 7037 3473
rect 7074 3439 7108 3473
rect 7145 3439 7179 3473
rect 7216 3439 7250 3473
rect 7287 3439 7321 3473
rect 7358 3439 7392 3473
rect 7429 3439 7463 3473
rect 7500 3439 7534 3473
rect 7571 3439 7605 3473
rect 7642 3439 7676 3473
rect 8775 3722 8809 3756
rect 8870 3722 8904 3756
rect 8965 3722 8999 3756
rect 9087 3722 9121 3756
rect 9182 3722 9216 3756
rect 9277 3722 9311 3756
rect 9541 3702 9575 3736
rect 9803 3722 9837 3756
rect 9898 3722 9932 3756
rect 9993 3722 10027 3756
rect 10392 3722 10426 3756
rect 10466 3722 10500 3756
rect 10539 3722 10573 3756
rect 10612 3722 10646 3756
rect 10685 3722 10719 3756
rect 10758 3722 10792 3756
rect 10831 3722 10865 3756
rect 10904 3722 10938 3756
rect 10977 3722 11011 3756
rect 11050 3722 11084 3756
rect 9541 3634 9575 3668
rect 10640 3609 10674 3643
rect 10774 3609 10808 3643
rect 9941 3414 9975 3448
rect 9941 3319 9975 3353
rect 9941 3224 9975 3258
rect 10070 3301 10104 3335
rect 10070 3233 10104 3267
rect 17619 3134 17653 3168
rect 17619 3066 17653 3100
rect 1622 2347 1656 2381
rect 1622 2279 1656 2313
rect 8571 2124 8605 2158
rect 8639 2124 8673 2158
rect 4472 2042 4506 2076
rect 4472 1974 4506 2008
rect 4472 1906 4506 1940
rect 1622 1746 1656 1780
rect 1622 1651 1656 1685
rect 1622 1556 1656 1590
rect 4472 1838 4506 1872
rect 4472 1770 4506 1804
rect 4472 1702 4506 1736
rect 4580 2042 4614 2076
rect 4580 1972 4614 2006
rect 4580 1902 4614 1936
rect 4580 1832 4614 1866
rect 4580 1762 4614 1796
rect 4580 1692 4614 1726
rect 6909 1788 6943 1822
rect 6977 1788 7011 1822
rect 7045 1788 7079 1822
rect 7113 1788 7147 1822
rect 7181 1788 7215 1822
rect 7249 1788 7283 1822
rect 7317 1788 7351 1822
rect 7385 1788 7419 1822
rect 7453 1788 7487 1822
rect 7521 1788 7555 1822
rect 7589 1788 7623 1822
rect 7657 1788 7691 1822
rect 7725 1788 7759 1822
rect 7793 1788 7827 1822
rect 7862 1788 7896 1822
rect 7931 1788 7965 1822
rect 8000 1788 8034 1822
rect 8069 1788 8103 1822
rect 8138 1788 8172 1822
rect 8207 1788 8241 1822
rect 8276 1788 8310 1822
rect 8345 1788 8379 1822
rect 8414 1788 8448 1822
rect 4472 1634 4506 1668
rect 4472 1565 4506 1599
rect 4472 1496 4506 1530
rect 17932 2768 17966 2802
rect 18000 2768 18034 2802
rect 4472 1427 4506 1461
rect 7485 1439 7519 1473
rect 7562 1439 7596 1473
rect 7639 1439 7673 1473
rect 7716 1439 7750 1473
rect 7793 1439 7827 1473
rect 1622 1184 1656 1218
rect 1622 1089 1656 1123
rect 1622 994 1656 1028
rect 4472 1358 4506 1392
rect 4472 1289 4506 1323
rect 4472 1220 4506 1254
rect 4580 1334 4614 1368
rect 4580 1220 4614 1254
rect 2467 1064 2501 1098
rect 2539 1064 2573 1098
rect 2611 1064 2645 1098
rect 2683 1064 2717 1098
rect 2755 1064 2789 1098
rect 2827 1064 2861 1098
rect 2898 1064 2932 1098
rect 2969 1064 3003 1098
rect 3091 1064 3125 1098
rect 3162 1064 3196 1098
rect 3233 1064 3267 1098
rect 3305 1064 3339 1098
rect 3377 1064 3411 1098
rect 3449 1064 3483 1098
rect 3521 1064 3555 1098
rect 3593 1064 3627 1098
rect 3839 1064 3873 1098
rect 3934 1064 3968 1098
rect 4029 1064 4063 1098
rect 4151 1064 4185 1098
rect 4246 1064 4280 1098
rect 4341 1064 4375 1098
rect 4463 1064 4497 1098
rect 4619 1064 4653 1098
rect 4714 1064 4748 1098
rect 4809 1064 4843 1098
rect 4931 1064 4965 1098
rect 5087 1064 5121 1098
rect 5157 1064 5191 1098
rect 5226 1064 5260 1098
rect 5295 1064 5329 1098
rect 5364 1064 5398 1098
rect 5433 1064 5467 1098
rect 5729 1064 5763 1098
rect 5824 1064 5858 1098
rect 5919 1064 5953 1098
rect 6041 1064 6075 1098
rect 6136 1064 6170 1098
rect 6231 1064 6265 1098
rect 6461 1064 6495 1098
rect 6544 1064 6578 1098
rect 6627 1064 6661 1098
rect 6709 1064 6743 1098
rect 6791 1064 6825 1098
rect 6913 1064 6947 1098
rect 6983 1064 7017 1098
rect 1622 838 1656 872
rect 1690 838 1724 872
rect 1622 716 1656 750
rect 1622 621 1656 655
rect 1622 526 1656 560
rect 1622 370 1656 404
rect 1690 370 1724 404
rect 1622 248 1656 282
rect 1622 153 1656 187
rect 1622 58 1656 92
rect 1622 -98 1656 -64
rect 1690 -98 1724 -64
rect 8345 996 8379 1030
rect 8416 996 8450 1030
rect 8487 996 8521 1030
rect 8559 996 8593 1030
rect 8631 996 8665 1030
rect 8703 996 8737 1030
rect 8775 996 8809 1030
rect 8847 996 8881 1030
rect 8969 996 9003 1030
rect 9043 996 9077 1030
rect 9116 996 9150 1030
rect 9189 996 9223 1030
rect 9262 996 9296 1030
rect 9335 996 9369 1030
rect 9408 996 9442 1030
rect 9481 996 9515 1030
rect 9554 996 9588 1030
rect 9627 996 9661 1030
rect 9749 996 9783 1030
rect 9822 996 9856 1030
rect 9895 996 9929 1030
rect 9968 996 10002 1030
rect 10041 996 10075 1030
rect 10114 996 10148 1030
rect 10187 996 10221 1030
rect 10260 996 10294 1030
rect 10333 996 10367 1030
rect 10407 996 10441 1030
rect 10804 996 10838 1030
rect 10875 996 10909 1030
rect 10946 996 10980 1030
rect 11017 996 11051 1030
rect 11088 996 11122 1030
rect 11159 996 11193 1030
rect 11230 996 11264 1030
rect 11301 996 11335 1030
rect 11372 996 11406 1030
rect 11443 996 11477 1030
rect 11514 996 11548 1030
rect 11585 996 11619 1030
rect 11656 996 11690 1030
rect 11727 996 11761 1030
rect 11798 996 11832 1030
rect 11869 996 11903 1030
rect 11940 996 11974 1030
rect 12010 996 12044 1030
rect 12080 996 12114 1030
rect 12150 996 12184 1030
rect 12220 996 12254 1030
rect 12290 996 12324 1030
rect 12360 996 12394 1030
rect 12430 996 12464 1030
rect 12500 996 12534 1030
rect 12844 996 12878 1030
rect 12912 996 12946 1030
rect 15124 974 15158 1008
rect 15124 906 15158 940
rect 15124 838 15158 872
rect 15124 770 15158 804
rect 15124 702 15158 736
rect 15284 744 15318 778
rect 15353 744 15387 778
rect 15422 744 15456 778
rect 15491 744 15525 778
rect 15560 744 15594 778
rect 15629 744 15663 778
rect 15698 744 15732 778
rect 15766 744 15800 778
rect 15834 744 15868 778
rect 15902 744 15936 778
rect 15970 744 16004 778
rect 16038 744 16072 778
rect 16106 744 16140 778
rect 15124 634 15158 668
rect 15124 565 15158 599
rect 15124 496 15158 530
rect 15124 427 15158 461
rect 15124 358 15158 392
rect 15124 289 15158 323
rect 15284 364 15318 398
rect 15353 364 15387 398
rect 15422 364 15456 398
rect 15491 364 15525 398
rect 15560 364 15594 398
rect 15629 364 15663 398
rect 15698 364 15732 398
rect 15766 364 15800 398
rect 15834 364 15868 398
rect 15902 364 15936 398
rect 15970 364 16004 398
rect 16038 364 16072 398
rect 16106 364 16140 398
rect 15124 220 15158 254
rect 15124 151 15158 185
rect 15911 225 15945 259
rect 15979 225 16013 259
rect 16101 225 16135 259
rect 16169 225 16203 259
rect 18644 223 18678 257
rect 18712 223 18746 257
rect 1622 -220 1656 -186
rect 1622 -315 1656 -281
rect 1622 -410 1656 -376
rect 1622 -566 1656 -532
rect 1690 -566 1724 -532
rect 1622 -722 1656 -688
rect 1690 -722 1724 -688
rect 1622 -1129 1656 -1095
rect 1622 -1224 1656 -1190
rect 18644 71 18678 105
rect 18712 71 18746 105
rect 1622 -1319 1656 -1285
rect 1622 -1441 1656 -1407
rect 1622 -1536 1656 -1502
rect 1622 -1631 1656 -1597
rect 1622 -1753 1656 -1719
rect 1622 -1848 1656 -1814
rect 1622 -1943 1656 -1909
rect 1622 -2065 1656 -2031
rect 1622 -2160 1656 -2126
rect 1622 -2255 1656 -2221
rect 2685 -10266 2719 -10232
rect 2780 -10266 2814 -10232
rect 2875 -10266 2909 -10232
rect 18870 -11651 18904 -11617
rect 18870 -11719 18904 -11685
rect 18874 -12901 18908 -12867
rect 18874 -12969 18908 -12935
rect 3084 -17052 3118 -17018
rect 3179 -17052 3213 -17018
rect 3274 -17052 3308 -17018
rect 2641 -17867 2675 -17833
rect 2736 -17867 2770 -17833
rect 2831 -17867 2865 -17833
<< npolyres >>
rect 1765 -11743 18870 -11593
rect 1765 -11843 1915 -11743
rect 1765 -11993 18924 -11843
rect 18774 -12093 18924 -11993
rect 1765 -12243 18924 -12093
rect 1765 -12343 1915 -12243
rect 1765 -12493 18924 -12343
rect 18774 -12593 18924 -12493
rect 1765 -12743 18924 -12593
rect 1765 -12843 1915 -12743
rect 1765 -12993 18874 -12843
<< mvndiffres >>
rect 10671 2643 16336 2743
rect 16236 2569 16336 2643
rect 10626 2469 16336 2569
rect 10626 2395 10726 2469
rect 10626 2295 16336 2395
rect 16236 2221 16336 2295
rect 10668 2121 16336 2221
rect 515 -3460 789 -3360
rect 515 -10922 615 -3460
rect 689 -10864 789 -3460
rect 863 -10864 963 -3403
rect 689 -10964 963 -10864
<< locali >>
rect 467 4960 539 4994
rect 573 4971 611 4994
rect 645 4971 683 4994
rect 717 4971 755 4994
rect 789 4971 827 4994
rect 861 4971 899 4994
rect 933 4971 971 4994
rect 1005 4971 1043 4994
rect 1077 4971 1115 4994
rect 1149 4971 1187 4994
rect 1221 4971 1259 4994
rect 1293 4971 1331 4994
rect 1365 4971 1403 4994
rect 1437 4971 1475 4994
rect 1509 4971 1547 4994
rect 1581 4971 1619 4994
rect 1653 4971 1691 4994
rect 1725 4971 1763 4994
rect 1797 4971 1835 4994
rect 1869 4971 1907 4994
rect 1941 4971 1979 4994
rect 2013 4971 2051 4994
rect 2085 4971 2123 4994
rect 2157 4971 2195 4994
rect 2229 4971 2267 4994
rect 2301 4971 2339 4994
rect 2373 4971 2411 4994
rect 2445 4971 2483 4994
rect 2517 4971 2555 4994
rect 2589 4971 2627 4994
rect 2661 4971 2699 4994
rect 2733 4971 2771 4994
rect 2805 4971 2843 4994
rect 2877 4971 2915 4994
rect 2949 4971 2987 4994
rect 3021 4971 3059 4994
rect 3093 4971 3131 4994
rect 3165 4971 3203 4994
rect 3237 4971 3275 4994
rect 3309 4971 3347 4994
rect 3381 4971 3419 4994
rect 3453 4971 3491 4994
rect 3525 4971 3563 4994
rect 3597 4971 3635 4994
rect 3669 4971 3707 4994
rect 3741 4971 3779 4994
rect 3813 4971 3851 4994
rect 3885 4971 3923 4994
rect 3957 4971 3995 4994
rect 4029 4971 4067 4994
rect 4101 4971 4139 4994
rect 4173 4971 4211 4994
rect 4245 4971 4283 4994
rect 4317 4971 4355 4994
rect 4389 4971 4427 4994
rect 4461 4971 4499 4994
rect 4533 4971 4571 4994
rect 4605 4971 4643 4994
rect 4677 4971 4715 4994
rect 4749 4971 4787 4994
rect 4821 4971 4859 4994
rect 4893 4971 4931 4994
rect 4965 4971 5003 4994
rect 5037 4971 5075 4994
rect 5109 4971 5147 4994
rect 5181 4971 5219 4994
rect 5253 4971 5291 4994
rect 5325 4971 5363 4994
rect 5397 4971 5435 4994
rect 5469 4971 5507 4994
rect 5541 4971 5579 4994
rect 5613 4971 5651 4994
rect 5685 4971 5723 4994
rect 5757 4971 5795 4994
rect 5829 4971 5868 4994
rect 5902 4971 5941 4994
rect 5975 4971 6014 4994
rect 6048 4971 6087 4994
rect 6121 4971 6160 4994
rect 6194 4971 6233 4994
rect 6267 4971 6306 4994
rect 6340 4971 6379 4994
rect 6413 4971 6452 4994
rect 6486 4971 6525 4994
rect 6559 4971 6598 4994
rect 6632 4971 6671 4994
rect 6705 4971 6744 4994
rect 573 4960 590 4971
rect 645 4960 658 4971
rect 717 4960 726 4971
rect 789 4960 794 4971
rect 861 4960 862 4971
rect 467 4937 590 4960
rect 624 4937 658 4960
rect 692 4937 726 4960
rect 760 4937 794 4960
rect 828 4937 862 4960
rect 896 4960 899 4971
rect 964 4960 971 4971
rect 1032 4960 1043 4971
rect 1100 4960 1115 4971
rect 1168 4960 1187 4971
rect 1236 4960 1259 4971
rect 1304 4960 1331 4971
rect 1372 4960 1403 4971
rect 896 4937 930 4960
rect 964 4937 998 4960
rect 1032 4937 1066 4960
rect 1100 4937 1134 4960
rect 1168 4937 1202 4960
rect 1236 4937 1270 4960
rect 1304 4937 1338 4960
rect 1372 4937 1406 4960
rect 1440 4937 1474 4971
rect 1509 4960 1542 4971
rect 1581 4960 1610 4971
rect 1653 4960 1678 4971
rect 1725 4960 1746 4971
rect 1797 4960 1814 4971
rect 1869 4960 1882 4971
rect 1941 4960 1950 4971
rect 2013 4960 2018 4971
rect 2085 4960 2086 4971
rect 1508 4937 1542 4960
rect 1576 4937 1610 4960
rect 1644 4937 1678 4960
rect 1712 4937 1746 4960
rect 1780 4937 1814 4960
rect 1848 4937 1882 4960
rect 1916 4937 1950 4960
rect 1984 4937 2018 4960
rect 2052 4937 2086 4960
rect 2120 4960 2123 4971
rect 2188 4960 2195 4971
rect 2256 4960 2267 4971
rect 2324 4960 2339 4971
rect 2392 4960 2411 4971
rect 2460 4960 2483 4971
rect 2528 4960 2555 4971
rect 2596 4960 2627 4971
rect 2120 4937 2154 4960
rect 2188 4937 2222 4960
rect 2256 4937 2290 4960
rect 2324 4937 2358 4960
rect 2392 4937 2426 4960
rect 2460 4937 2494 4960
rect 2528 4937 2562 4960
rect 2596 4937 2630 4960
rect 2664 4937 2698 4971
rect 2733 4960 2766 4971
rect 2805 4960 2834 4971
rect 2877 4960 2902 4971
rect 2949 4960 2970 4971
rect 3021 4960 3038 4971
rect 3093 4960 3106 4971
rect 3165 4960 3174 4971
rect 3237 4960 3242 4971
rect 3309 4960 3310 4971
rect 2732 4937 2766 4960
rect 2800 4937 2834 4960
rect 2868 4937 2902 4960
rect 2936 4937 2970 4960
rect 3004 4937 3038 4960
rect 3072 4937 3106 4960
rect 3140 4937 3174 4960
rect 3208 4937 3242 4960
rect 3276 4937 3310 4960
rect 3344 4960 3347 4971
rect 3412 4960 3419 4971
rect 3480 4960 3491 4971
rect 3548 4960 3563 4971
rect 3616 4960 3635 4971
rect 3684 4960 3707 4971
rect 3752 4960 3779 4971
rect 3820 4960 3851 4971
rect 3344 4937 3378 4960
rect 3412 4937 3446 4960
rect 3480 4937 3514 4960
rect 3548 4937 3582 4960
rect 3616 4937 3650 4960
rect 3684 4937 3718 4960
rect 3752 4937 3786 4960
rect 3820 4937 3854 4960
rect 3888 4937 3922 4971
rect 3957 4960 3990 4971
rect 4029 4960 4058 4971
rect 4101 4960 4126 4971
rect 4173 4960 4194 4971
rect 4245 4960 4262 4971
rect 4317 4960 4330 4971
rect 4389 4960 4398 4971
rect 4461 4960 4466 4971
rect 4533 4960 4534 4971
rect 3956 4937 3990 4960
rect 4024 4937 4058 4960
rect 4092 4937 4126 4960
rect 4160 4937 4194 4960
rect 4228 4937 4262 4960
rect 4296 4937 4330 4960
rect 4364 4937 4398 4960
rect 4432 4937 4466 4960
rect 4500 4937 4534 4960
rect 4568 4960 4571 4971
rect 4636 4960 4643 4971
rect 4704 4960 4715 4971
rect 4772 4960 4787 4971
rect 4840 4960 4859 4971
rect 4908 4960 4931 4971
rect 4976 4960 5003 4971
rect 5044 4960 5075 4971
rect 4568 4937 4602 4960
rect 4636 4937 4670 4960
rect 4704 4937 4738 4960
rect 4772 4937 4806 4960
rect 4840 4937 4874 4960
rect 4908 4937 4942 4960
rect 4976 4937 5010 4960
rect 5044 4937 5078 4960
rect 5112 4937 5146 4971
rect 5181 4960 5214 4971
rect 5253 4960 5282 4971
rect 5325 4960 5350 4971
rect 5397 4960 5418 4971
rect 5469 4960 5486 4971
rect 5541 4960 5554 4971
rect 5613 4960 5622 4971
rect 5685 4960 5690 4971
rect 5757 4960 5758 4971
rect 5180 4937 5214 4960
rect 5248 4937 5282 4960
rect 5316 4937 5350 4960
rect 5384 4937 5418 4960
rect 5452 4937 5486 4960
rect 5520 4937 5554 4960
rect 5588 4937 5622 4960
rect 5656 4937 5690 4960
rect 5724 4937 5758 4960
rect 5792 4960 5795 4971
rect 5860 4960 5868 4971
rect 5928 4960 5941 4971
rect 5996 4960 6014 4971
rect 6064 4960 6087 4971
rect 6132 4960 6160 4971
rect 6200 4960 6233 4971
rect 5792 4937 5826 4960
rect 5860 4937 5894 4960
rect 5928 4937 5962 4960
rect 5996 4937 6030 4960
rect 6064 4937 6098 4960
rect 6132 4937 6166 4960
rect 6200 4937 6234 4960
rect 6268 4937 6302 4971
rect 6340 4960 6370 4971
rect 6413 4960 6438 4971
rect 6486 4960 6506 4971
rect 6559 4960 6574 4971
rect 6632 4960 6642 4971
rect 6705 4960 6710 4971
rect 6336 4937 6370 4960
rect 6404 4937 6438 4960
rect 6472 4937 6506 4960
rect 6540 4937 6574 4960
rect 6608 4937 6642 4960
rect 6676 4937 6710 4960
rect 6778 4971 6817 4994
rect 6851 4971 6890 4994
rect 6924 4971 6963 4994
rect 6997 4971 7036 4994
rect 7070 4971 7109 4994
rect 7143 4971 7182 4994
rect 7216 4971 7255 4994
rect 7289 4971 7328 4994
rect 7362 4971 7401 4994
rect 7435 4971 7474 4994
rect 7508 4971 7547 4994
rect 7581 4971 7620 4994
rect 7654 4971 7693 4994
rect 7727 4971 7766 4994
rect 6744 4937 6778 4960
rect 6812 4960 6817 4971
rect 6880 4960 6890 4971
rect 6948 4960 6963 4971
rect 7016 4960 7036 4971
rect 7084 4960 7109 4971
rect 7152 4960 7182 4971
rect 6812 4937 6846 4960
rect 6880 4937 6914 4960
rect 6948 4937 6982 4960
rect 7016 4937 7050 4960
rect 7084 4937 7118 4960
rect 7152 4937 7186 4960
rect 7220 4937 7254 4971
rect 7289 4960 7322 4971
rect 7362 4960 7390 4971
rect 7435 4960 7458 4971
rect 7508 4960 7526 4971
rect 7581 4960 7594 4971
rect 7654 4960 7662 4971
rect 7727 4960 7730 4971
rect 7288 4937 7322 4960
rect 7356 4937 7390 4960
rect 7424 4937 7458 4960
rect 7492 4937 7526 4960
rect 7560 4937 7594 4960
rect 7628 4937 7662 4960
rect 7696 4937 7730 4960
rect 7764 4960 7766 4971
rect 7800 4960 7872 4994
rect 7764 4937 7872 4960
rect 467 4922 713 4937
rect 501 4896 713 4922
rect 501 4888 522 4896
rect 467 4862 522 4888
rect 556 4862 713 4896
rect 467 4861 713 4862
rect 467 4847 593 4861
rect 501 4828 593 4847
rect 501 4813 522 4828
rect 467 4794 522 4813
rect 556 4827 593 4828
rect 627 4827 679 4861
rect 556 4823 713 4827
rect 7838 4920 7872 4937
rect 7838 4846 7872 4869
rect 556 4794 663 4823
rect 467 4791 663 4794
rect 697 4791 713 4823
rect 467 4772 593 4791
rect 501 4760 593 4772
rect 501 4738 522 4760
rect 467 4726 522 4738
rect 556 4757 593 4760
rect 627 4789 663 4791
rect 627 4757 679 4789
rect 556 4740 713 4757
rect 556 4726 663 4740
rect 467 4721 663 4726
rect 697 4721 713 4740
rect 467 4697 593 4721
rect 501 4692 593 4697
rect 501 4663 522 4692
rect 467 4658 522 4663
rect 556 4687 593 4692
rect 627 4706 663 4721
rect 871 4751 905 4773
rect 1727 4751 1761 4773
rect 1983 4751 2017 4773
rect 2239 4751 2273 4773
rect 2495 4751 2529 4773
rect 2751 4751 2785 4773
rect 3007 4751 3041 4773
rect 3263 4751 3297 4773
rect 3519 4751 3553 4773
rect 3775 4751 3809 4773
rect 4031 4751 4065 4773
rect 4287 4751 4321 4773
rect 4543 4751 4577 4773
rect 4799 4751 4833 4773
rect 5055 4751 5089 4773
rect 5311 4751 5345 4773
rect 5567 4751 5601 4773
rect 5823 4751 5857 4773
rect 6079 4751 6113 4773
rect 6335 4751 6369 4773
rect 6591 4751 6625 4773
rect 6847 4751 6881 4773
rect 7703 4751 7737 4773
rect 7838 4772 7872 4801
rect 627 4687 679 4706
rect 556 4658 713 4687
rect 7838 4699 7872 4733
rect 467 4657 713 4658
rect 467 4651 663 4657
rect 697 4651 713 4657
rect 467 4624 593 4651
rect 467 4622 522 4624
rect 501 4590 522 4622
rect 556 4617 593 4624
rect 627 4623 663 4651
rect 916 4652 932 4661
rect 916 4627 928 4652
rect 966 4627 1003 4661
rect 1037 4652 1074 4661
rect 1108 4652 1145 4661
rect 1179 4652 1216 4661
rect 1250 4652 1287 4661
rect 1321 4652 1358 4661
rect 1040 4627 1074 4652
rect 1118 4627 1145 4652
rect 1196 4627 1216 4652
rect 1273 4627 1287 4652
rect 1350 4627 1358 4652
rect 1392 4652 1429 4661
rect 1392 4627 1393 4652
rect 627 4617 679 4623
rect 962 4618 1006 4627
rect 1040 4618 1084 4627
rect 1118 4618 1162 4627
rect 1196 4618 1239 4627
rect 1273 4618 1316 4627
rect 1350 4618 1393 4627
rect 1427 4627 1429 4652
rect 1463 4652 1500 4661
rect 1534 4652 1571 4661
rect 1605 4652 1642 4661
rect 1463 4627 1470 4652
rect 1534 4627 1547 4652
rect 1605 4627 1624 4652
rect 1676 4627 1712 4661
rect 1746 4627 1782 4661
rect 1816 4627 1852 4661
rect 1886 4627 1922 4661
rect 1956 4627 1972 4661
rect 2028 4627 2044 4661
rect 2085 4627 2112 4661
rect 2164 4627 2180 4661
rect 2214 4627 2248 4661
rect 2282 4627 2316 4661
rect 2376 4627 2384 4661
rect 2418 4627 2421 4661
rect 2486 4627 2500 4661
rect 2554 4627 2578 4661
rect 2622 4627 2656 4661
rect 2690 4627 2724 4661
rect 2758 4627 2792 4661
rect 2826 4627 2837 4661
rect 2894 4627 2922 4661
rect 2962 4627 2996 4661
rect 3041 4627 3064 4661
rect 3125 4627 3133 4661
rect 3167 4627 3175 4661
rect 3236 4627 3252 4661
rect 3308 4627 3324 4661
rect 3358 4627 3385 4661
rect 3419 4627 3458 4661
rect 3496 4627 3508 4661
rect 3564 4627 3576 4661
rect 3614 4627 3648 4661
rect 3682 4627 3691 4661
rect 3750 4627 3784 4661
rect 3818 4627 3852 4661
rect 3892 4627 3920 4661
rect 3979 4627 3988 4661
rect 4022 4627 4032 4661
rect 4090 4627 4119 4661
rect 4158 4627 4192 4661
rect 4240 4627 4260 4661
rect 4294 4627 4328 4661
rect 4362 4627 4371 4661
rect 4430 4627 4457 4661
rect 4498 4627 4532 4661
rect 4577 4627 4600 4661
rect 4663 4627 4668 4661
rect 4702 4627 4715 4661
rect 4770 4627 4804 4661
rect 4838 4627 4872 4661
rect 4915 4627 4940 4661
rect 4989 4627 5008 4661
rect 5063 4627 5076 4661
rect 5136 4627 5144 4661
rect 5209 4627 5212 4661
rect 5246 4627 5248 4661
rect 5314 4627 5321 4661
rect 5382 4627 5394 4661
rect 5450 4627 5467 4661
rect 5518 4627 5540 4661
rect 5586 4627 5613 4661
rect 5654 4627 5686 4661
rect 5722 4627 5756 4661
rect 5793 4627 5824 4661
rect 5866 4627 5892 4661
rect 5939 4627 5960 4661
rect 6012 4627 6028 4661
rect 6085 4627 6096 4661
rect 6158 4627 6165 4661
rect 6231 4627 6234 4661
rect 6268 4627 6270 4661
rect 6337 4627 6343 4661
rect 6406 4627 6416 4661
rect 6475 4627 6489 4661
rect 6544 4627 6579 4661
rect 6613 4627 6648 4661
rect 6682 4627 6717 4661
rect 6751 4627 6786 4661
rect 6820 4627 6836 4661
rect 6994 4627 7010 4661
rect 7044 4652 7080 4661
rect 7044 4627 7066 4652
rect 7114 4627 7150 4661
rect 7184 4627 7220 4661
rect 7254 4652 7290 4661
rect 7324 4652 7360 4661
rect 7269 4627 7290 4652
rect 7354 4627 7360 4652
rect 7394 4652 7430 4661
rect 7464 4652 7500 4661
rect 7394 4627 7405 4652
rect 7464 4627 7490 4652
rect 7534 4627 7571 4661
rect 7605 4627 7642 4661
rect 7676 4627 7692 4661
rect 7838 4631 7872 4664
rect 1427 4618 1470 4627
rect 1504 4618 1547 4627
rect 1581 4618 1624 4627
rect 7100 4618 7150 4627
rect 7184 4618 7235 4627
rect 7269 4618 7320 4627
rect 7354 4618 7405 4627
rect 7439 4618 7490 4627
rect 556 4590 713 4617
rect 501 4588 713 4590
rect 467 4581 713 4588
rect 467 4556 593 4581
rect 467 4547 522 4556
rect 501 4522 522 4547
rect 556 4547 593 4556
rect 627 4547 679 4581
rect 556 4522 713 4547
rect 501 4513 713 4522
rect 467 4511 713 4513
rect 467 4488 593 4511
rect 467 4472 522 4488
rect 501 4454 522 4472
rect 556 4477 593 4488
rect 627 4486 679 4511
rect 7838 4563 7872 4590
rect 7838 4495 7872 4516
rect 627 4477 660 4486
rect 962 4483 1006 4492
rect 1040 4483 1084 4492
rect 1118 4483 1162 4492
rect 1196 4483 1239 4492
rect 1273 4483 1316 4492
rect 1350 4483 1393 4492
rect 1427 4483 1470 4492
rect 1504 4483 1547 4492
rect 1581 4483 1624 4492
rect 1823 4483 1865 4486
rect 1899 4483 1941 4486
rect 1975 4483 2017 4486
rect 2051 4483 2093 4486
rect 2127 4483 2169 4486
rect 2203 4483 2244 4486
rect 2278 4483 2319 4486
rect 2353 4483 2394 4486
rect 2428 4483 2469 4486
rect 2503 4483 2544 4486
rect 2578 4483 2619 4486
rect 2653 4483 2694 4486
rect 2728 4483 2769 4486
rect 2803 4483 2844 4486
rect 2878 4483 2919 4486
rect 3129 4483 3173 4486
rect 3207 4483 3251 4486
rect 3285 4483 3329 4486
rect 3363 4483 3407 4486
rect 3441 4483 3485 4486
rect 3519 4483 3563 4486
rect 3597 4483 3641 4486
rect 3675 4483 3718 4486
rect 3866 4483 3929 4486
rect 556 4454 660 4477
rect 501 4452 660 4454
rect 694 4452 713 4477
rect 501 4441 713 4452
rect 916 4458 928 4483
rect 916 4449 932 4458
rect 966 4449 1006 4483
rect 1040 4449 1080 4483
rect 1118 4458 1154 4483
rect 1196 4458 1228 4483
rect 1273 4458 1301 4483
rect 1350 4458 1374 4483
rect 1427 4458 1447 4483
rect 1504 4458 1520 4483
rect 1581 4458 1593 4483
rect 1658 4458 1666 4483
rect 1114 4449 1154 4458
rect 1188 4449 1228 4458
rect 1262 4449 1301 4458
rect 1335 4449 1374 4458
rect 1408 4449 1447 4458
rect 1481 4449 1520 4458
rect 1554 4449 1593 4458
rect 1627 4449 1666 4458
rect 1700 4449 1716 4483
rect 1772 4449 1788 4483
rect 1823 4452 1856 4483
rect 1899 4452 1924 4483
rect 1975 4452 1992 4483
rect 2051 4452 2060 4483
rect 2127 4452 2128 4483
rect 1822 4449 1856 4452
rect 1890 4449 1924 4452
rect 1958 4449 1992 4452
rect 2026 4449 2060 4452
rect 2094 4449 2128 4452
rect 2162 4452 2169 4483
rect 2230 4452 2244 4483
rect 2299 4452 2319 4483
rect 2368 4452 2394 4483
rect 2437 4452 2469 4483
rect 2162 4449 2196 4452
rect 2230 4449 2265 4452
rect 2299 4449 2334 4452
rect 2368 4449 2403 4452
rect 2437 4449 2472 4452
rect 2506 4449 2541 4483
rect 2578 4452 2610 4483
rect 2653 4452 2679 4483
rect 2728 4452 2748 4483
rect 2803 4452 2817 4483
rect 2878 4452 2886 4483
rect 2953 4452 2955 4483
rect 2575 4449 2610 4452
rect 2644 4449 2679 4452
rect 2713 4449 2748 4452
rect 2782 4449 2817 4452
rect 2851 4449 2886 4452
rect 2920 4449 2955 4452
rect 2989 4449 3024 4483
rect 3058 4449 3093 4483
rect 3129 4452 3162 4483
rect 3207 4452 3231 4483
rect 3285 4452 3300 4483
rect 3363 4452 3369 4483
rect 3127 4449 3162 4452
rect 3196 4449 3231 4452
rect 3265 4449 3300 4452
rect 3334 4449 3369 4452
rect 3403 4452 3407 4483
rect 3472 4452 3485 4483
rect 3541 4452 3563 4483
rect 3610 4452 3641 4483
rect 3403 4449 3438 4452
rect 3472 4449 3507 4452
rect 3541 4449 3576 4452
rect 3610 4449 3645 4452
rect 3679 4449 3714 4483
rect 3752 4452 3764 4483
rect 3748 4449 3764 4452
rect 3820 4452 3832 4483
rect 3870 4452 3929 4483
rect 3963 4452 3970 4483
rect 3820 4449 3836 4452
rect 3870 4449 3970 4452
rect 4004 4449 4020 4483
rect 4076 4449 4092 4483
rect 4126 4452 4133 4483
rect 4167 4483 4230 4486
rect 4378 4483 4451 4486
rect 4634 4483 4675 4486
rect 4709 4483 4750 4486
rect 4784 4483 4825 4486
rect 4859 4483 4900 4486
rect 4934 4483 4975 4486
rect 5009 4483 5050 4486
rect 5084 4483 5125 4486
rect 5159 4483 5199 4486
rect 5233 4483 5273 4486
rect 5307 4483 5347 4486
rect 5381 4483 5421 4486
rect 5455 4483 5495 4486
rect 5529 4483 5569 4486
rect 5603 4483 5643 4486
rect 5677 4483 5717 4486
rect 5751 4483 5791 4486
rect 5825 4483 5865 4486
rect 5899 4483 5939 4486
rect 5973 4483 6013 4486
rect 4167 4452 4226 4483
rect 4264 4452 4276 4483
rect 4126 4449 4226 4452
rect 4260 4449 4276 4452
rect 4332 4452 4344 4483
rect 4382 4452 4451 4483
rect 4332 4449 4348 4452
rect 4382 4449 4482 4452
rect 4516 4449 4532 4483
rect 4588 4452 4600 4483
rect 4588 4449 4604 4452
rect 4638 4449 4672 4483
rect 4709 4452 4740 4483
rect 4784 4452 4808 4483
rect 4859 4452 4876 4483
rect 4934 4452 4944 4483
rect 5009 4452 5013 4483
rect 4706 4449 4740 4452
rect 4774 4449 4808 4452
rect 4842 4449 4876 4452
rect 4910 4449 4944 4452
rect 4978 4449 5013 4452
rect 5047 4452 5050 4483
rect 5116 4452 5125 4483
rect 5185 4452 5199 4483
rect 5254 4452 5273 4483
rect 5323 4452 5347 4483
rect 5392 4452 5421 4483
rect 5461 4452 5495 4483
rect 5047 4449 5082 4452
rect 5116 4449 5151 4452
rect 5185 4449 5220 4452
rect 5254 4449 5289 4452
rect 5323 4449 5358 4452
rect 5392 4449 5427 4452
rect 5461 4449 5496 4452
rect 5530 4449 5565 4483
rect 5603 4452 5634 4483
rect 5677 4452 5703 4483
rect 5751 4452 5772 4483
rect 5825 4452 5841 4483
rect 5899 4452 5910 4483
rect 5973 4452 5979 4483
rect 5599 4449 5634 4452
rect 5668 4449 5703 4452
rect 5737 4449 5772 4452
rect 5806 4449 5841 4452
rect 5875 4449 5910 4452
rect 5944 4449 5979 4452
rect 6047 4483 6087 4486
rect 6121 4483 6161 4486
rect 6195 4483 6235 4486
rect 6269 4483 6309 4486
rect 6343 4483 6383 4486
rect 6417 4483 6457 4486
rect 6491 4483 6531 4486
rect 7100 4483 7138 4492
rect 7172 4483 7210 4492
rect 7244 4483 7282 4492
rect 7316 4483 7355 4492
rect 7389 4483 7428 4492
rect 7462 4483 7501 4492
rect 7535 4483 7574 4492
rect 7608 4483 7647 4492
rect 6047 4452 6048 4483
rect 6013 4449 6048 4452
rect 6082 4452 6087 4483
rect 6151 4452 6161 4483
rect 6220 4452 6235 4483
rect 6289 4452 6309 4483
rect 6358 4452 6383 4483
rect 6427 4452 6457 4483
rect 6082 4449 6117 4452
rect 6151 4449 6186 4452
rect 6220 4449 6255 4452
rect 6289 4449 6324 4452
rect 6358 4449 6393 4452
rect 6427 4449 6462 4452
rect 6496 4449 6531 4483
rect 6565 4449 6581 4483
rect 6636 4449 6652 4483
rect 6686 4449 6722 4483
rect 6756 4449 6792 4483
rect 6826 4449 6862 4483
rect 6896 4449 6932 4483
rect 6966 4449 7003 4483
rect 7037 4458 7066 4483
rect 7108 4458 7138 4483
rect 7179 4458 7210 4483
rect 7250 4458 7282 4483
rect 7321 4458 7355 4483
rect 7392 4458 7428 4483
rect 7037 4449 7074 4458
rect 7108 4449 7145 4458
rect 7179 4449 7216 4458
rect 7250 4449 7287 4458
rect 7321 4449 7358 4458
rect 7392 4449 7429 4458
rect 7463 4449 7500 4483
rect 7535 4458 7571 4483
rect 7608 4458 7642 4483
rect 7681 4458 7692 4483
rect 7534 4449 7571 4458
rect 7605 4449 7642 4458
rect 7676 4449 7692 4458
rect 501 4438 593 4441
rect 467 4420 593 4438
rect 467 4397 522 4420
rect 501 4386 522 4397
rect 556 4407 593 4420
rect 627 4407 679 4441
rect 556 4404 713 4407
rect 556 4386 660 4404
rect 501 4371 660 4386
rect 694 4371 713 4404
rect 7838 4427 7872 4441
rect 501 4363 593 4371
rect 467 4352 593 4363
rect 467 4322 522 4352
rect 501 4318 522 4322
rect 556 4337 593 4352
rect 627 4370 660 4371
rect 627 4337 679 4370
rect 556 4321 713 4337
rect 556 4318 660 4321
rect 501 4301 660 4318
rect 694 4301 713 4321
rect 501 4288 593 4301
rect 467 4284 593 4288
rect 467 4250 522 4284
rect 556 4267 593 4284
rect 627 4287 660 4301
rect 871 4337 905 4359
rect 1727 4337 1761 4359
rect 1983 4337 2017 4359
rect 2239 4337 2273 4359
rect 2495 4337 2529 4359
rect 2751 4337 2785 4359
rect 3007 4337 3041 4359
rect 3263 4337 3297 4359
rect 3519 4337 3553 4359
rect 3775 4337 3809 4359
rect 4031 4337 4065 4359
rect 4287 4337 4321 4359
rect 4543 4337 4577 4359
rect 4799 4337 4833 4359
rect 5055 4337 5089 4359
rect 5311 4337 5345 4359
rect 5567 4337 5601 4359
rect 5823 4337 5857 4359
rect 6079 4337 6113 4359
rect 6335 4337 6369 4359
rect 6591 4337 6625 4359
rect 6847 4337 6881 4359
rect 7703 4337 7737 4359
rect 7838 4359 7872 4366
rect 627 4267 679 4287
rect 556 4250 713 4267
rect 467 4247 713 4250
rect 501 4231 713 4247
rect 501 4216 593 4231
rect 501 4213 522 4216
rect 467 4182 522 4213
rect 556 4197 593 4216
rect 627 4197 679 4231
rect 556 4182 713 4197
rect 467 4172 713 4182
rect 501 4161 713 4172
rect 501 4148 593 4161
rect 501 4138 522 4148
rect 467 4114 522 4138
rect 556 4127 593 4148
rect 627 4127 679 4161
rect 556 4114 713 4127
rect 467 4097 713 4114
rect 501 4090 713 4097
rect 501 4080 593 4090
rect 501 4063 522 4080
rect 467 4046 522 4063
rect 556 4056 593 4080
rect 627 4056 679 4090
rect 556 4046 713 4056
rect 467 4022 713 4046
rect 501 4019 713 4022
rect 501 4012 593 4019
rect 501 3988 522 4012
rect 467 3978 522 3988
rect 556 3985 593 4012
rect 627 3985 679 4019
rect 556 3978 713 3985
rect 467 3948 713 3978
rect 467 3947 593 3948
rect 501 3944 593 3947
rect 501 3913 522 3944
rect 467 3910 522 3913
rect 556 3914 593 3944
rect 627 3914 679 3948
rect 556 3910 713 3914
rect 467 3877 713 3910
rect 467 3876 593 3877
rect 467 3872 522 3876
rect 501 3842 522 3872
rect 556 3843 593 3876
rect 627 3843 679 3877
rect 556 3842 713 3843
rect 501 3838 713 3842
rect 467 3813 713 3838
rect 7838 4250 7872 4257
rect 7838 4175 7872 4189
rect 7838 4100 7872 4121
rect 7838 4025 7872 4053
rect 7838 3951 7872 3985
rect 7838 3883 7872 3916
rect 7838 3815 7872 3841
rect 467 3808 660 3813
rect 467 3797 522 3808
rect 501 3774 522 3797
rect 556 3806 660 3808
rect 694 3806 713 3813
rect 556 3774 593 3806
rect 501 3772 593 3774
rect 627 3779 660 3806
rect 627 3772 679 3779
rect 501 3763 713 3772
rect 467 3740 713 3763
rect 467 3722 522 3740
rect 501 3706 522 3722
rect 556 3735 713 3740
rect 556 3706 593 3735
rect 501 3701 593 3706
rect 627 3731 679 3735
rect 627 3701 660 3731
rect 871 3741 905 3763
rect 1727 3741 1761 3763
rect 1983 3741 2017 3763
rect 2239 3741 2273 3763
rect 2495 3741 2529 3763
rect 2751 3741 2785 3763
rect 3007 3741 3041 3763
rect 3263 3741 3297 3763
rect 3519 3741 3553 3763
rect 3775 3741 3809 3763
rect 4031 3741 4065 3763
rect 4287 3741 4321 3763
rect 4543 3741 4577 3763
rect 4799 3741 4833 3763
rect 5055 3741 5089 3763
rect 5311 3741 5345 3763
rect 5567 3741 5601 3763
rect 5823 3741 5857 3763
rect 6079 3741 6113 3763
rect 6335 3741 6369 3763
rect 6591 3741 6625 3763
rect 6847 3741 6881 3763
rect 7703 3741 7737 3763
rect 7838 3725 7872 3766
rect 501 3697 660 3701
rect 694 3697 713 3701
rect 501 3688 713 3697
rect 467 3672 713 3688
rect 467 3647 522 3672
rect 501 3638 522 3647
rect 556 3664 713 3672
rect 556 3638 593 3664
rect 501 3630 593 3638
rect 627 3648 679 3664
rect 7838 3674 7872 3691
rect 627 3630 660 3648
rect 501 3614 660 3630
rect 694 3614 713 3630
rect 916 3642 932 3651
rect 916 3617 928 3642
rect 966 3617 1003 3651
rect 1037 3642 1074 3651
rect 1108 3642 1145 3651
rect 1179 3642 1216 3651
rect 1250 3642 1287 3651
rect 1321 3642 1358 3651
rect 1040 3617 1074 3642
rect 1118 3617 1145 3642
rect 1196 3617 1216 3642
rect 1273 3617 1287 3642
rect 1350 3617 1358 3642
rect 1392 3642 1429 3651
rect 1392 3617 1393 3642
rect 501 3613 713 3614
rect 467 3604 713 3613
rect 962 3608 1006 3617
rect 1040 3608 1084 3617
rect 1118 3608 1162 3617
rect 1196 3608 1239 3617
rect 1273 3608 1316 3617
rect 1350 3608 1393 3617
rect 1427 3617 1429 3642
rect 1463 3642 1500 3651
rect 1534 3642 1571 3651
rect 1605 3642 1642 3651
rect 1463 3617 1470 3642
rect 1534 3617 1547 3642
rect 1605 3617 1624 3642
rect 1676 3617 1712 3651
rect 1746 3617 1782 3651
rect 1816 3617 1852 3651
rect 1886 3617 1922 3651
rect 1956 3617 1972 3651
rect 2028 3617 2044 3651
rect 2078 3617 2112 3651
rect 2146 3617 2180 3651
rect 2214 3617 2248 3651
rect 2282 3617 2316 3651
rect 2350 3617 2384 3651
rect 2418 3617 2452 3651
rect 2486 3617 2521 3651
rect 2555 3645 2590 3651
rect 2624 3645 2659 3651
rect 2693 3645 2728 3651
rect 2762 3645 2797 3651
rect 2831 3645 2866 3651
rect 2555 3617 2557 3645
rect 2624 3617 2633 3645
rect 2693 3617 2709 3645
rect 2762 3617 2785 3645
rect 2831 3617 2861 3645
rect 2900 3617 2935 3651
rect 2969 3645 3004 3651
rect 3038 3645 3073 3651
rect 3107 3645 3142 3651
rect 3176 3645 3211 3651
rect 3245 3645 3280 3651
rect 3314 3645 3349 3651
rect 2970 3617 3004 3645
rect 3045 3617 3073 3645
rect 3120 3617 3142 3645
rect 3195 3617 3211 3645
rect 3270 3617 3280 3645
rect 3345 3617 3349 3645
rect 3383 3645 3418 3651
rect 3452 3645 3487 3651
rect 3521 3645 3556 3651
rect 3590 3645 3625 3651
rect 3659 3645 3694 3651
rect 3728 3645 3763 3651
rect 3383 3617 3386 3645
rect 3452 3617 3461 3645
rect 3521 3617 3536 3645
rect 3590 3617 3611 3645
rect 3659 3617 3686 3645
rect 3728 3617 3761 3645
rect 3797 3617 3832 3651
rect 3866 3645 3901 3651
rect 3935 3645 3970 3651
rect 4004 3645 4020 3651
rect 3870 3617 3901 3645
rect 3945 3617 3970 3645
rect 4076 3648 4092 3651
rect 4126 3648 4226 3651
rect 4076 3617 4088 3648
rect 4126 3617 4195 3648
rect 4260 3617 4276 3651
rect 4332 3645 4348 3651
rect 4382 3645 4482 3651
rect 4382 3617 4445 3645
rect 1427 3608 1470 3617
rect 1504 3608 1547 3617
rect 1581 3608 1624 3617
rect 2591 3611 2633 3617
rect 2667 3611 2709 3617
rect 2743 3611 2785 3617
rect 2819 3611 2861 3617
rect 2895 3611 2936 3617
rect 2970 3611 3011 3617
rect 3045 3611 3086 3617
rect 3120 3611 3161 3617
rect 3195 3611 3236 3617
rect 3270 3611 3311 3617
rect 3345 3611 3386 3617
rect 3420 3611 3461 3617
rect 3495 3611 3536 3617
rect 3570 3611 3611 3617
rect 3645 3611 3686 3617
rect 3720 3611 3761 3617
rect 3795 3611 3836 3617
rect 3870 3611 3911 3617
rect 3945 3611 3986 3617
rect 4122 3614 4195 3617
rect 4366 3611 4445 3617
rect 4479 3617 4482 3645
rect 4516 3617 4532 3651
rect 4588 3617 4604 3651
rect 4638 3648 4738 3651
rect 4772 3648 4788 3651
rect 4638 3617 4641 3648
rect 4675 3617 4738 3648
rect 4776 3617 4788 3648
rect 4844 3645 4860 3651
rect 4894 3645 4929 3651
rect 4963 3645 4998 3651
rect 5032 3645 5067 3651
rect 5101 3645 5136 3651
rect 5170 3645 5205 3651
rect 4894 3617 4916 3645
rect 4963 3617 4988 3645
rect 5032 3617 5060 3645
rect 5101 3617 5132 3645
rect 5170 3617 5204 3645
rect 5239 3617 5274 3651
rect 5308 3645 5343 3651
rect 5377 3645 5412 3651
rect 5446 3645 5481 3651
rect 5515 3645 5550 3651
rect 5584 3645 5620 3651
rect 5310 3617 5343 3645
rect 5382 3617 5412 3645
rect 5454 3617 5481 3645
rect 5526 3617 5550 3645
rect 5598 3617 5620 3645
rect 5654 3645 5690 3651
rect 5654 3617 5655 3645
rect 4675 3614 4742 3617
rect 4878 3611 4916 3617
rect 4950 3611 4988 3617
rect 5022 3611 5060 3617
rect 5094 3611 5132 3617
rect 5166 3611 5204 3617
rect 5238 3611 5276 3617
rect 5310 3611 5348 3617
rect 5382 3611 5420 3617
rect 5454 3611 5492 3617
rect 5526 3611 5564 3617
rect 5598 3611 5655 3617
rect 5689 3617 5690 3645
rect 5724 3645 5760 3651
rect 5794 3645 5830 3651
rect 5864 3645 5900 3651
rect 5934 3645 5970 3651
rect 6004 3645 6040 3651
rect 6074 3645 6110 3651
rect 6144 3645 6180 3651
rect 6214 3645 6250 3651
rect 5724 3617 5729 3645
rect 5794 3617 5803 3645
rect 5864 3617 5877 3645
rect 5934 3617 5951 3645
rect 6004 3617 6025 3645
rect 6074 3617 6099 3645
rect 6144 3617 6173 3645
rect 6214 3617 6247 3645
rect 6284 3617 6320 3651
rect 6354 3617 6390 3651
rect 6424 3645 6460 3651
rect 6450 3617 6460 3645
rect 6494 3617 6530 3651
rect 6564 3645 6580 3651
rect 6569 3617 6580 3645
rect 6636 3617 6652 3651
rect 6686 3617 6722 3651
rect 6756 3617 6792 3651
rect 6826 3617 6862 3651
rect 6896 3617 6932 3651
rect 6966 3642 7003 3651
rect 7037 3642 7074 3651
rect 7108 3642 7145 3651
rect 7179 3642 7216 3651
rect 7250 3642 7287 3651
rect 7321 3642 7358 3651
rect 7392 3642 7429 3651
rect 7463 3642 7500 3651
rect 6966 3617 6992 3642
rect 7037 3617 7064 3642
rect 7108 3617 7136 3642
rect 7179 3617 7208 3642
rect 7250 3617 7280 3642
rect 7321 3617 7353 3642
rect 7392 3617 7426 3642
rect 7463 3617 7499 3642
rect 7534 3617 7571 3651
rect 7605 3617 7642 3651
rect 7676 3617 7692 3651
rect 5689 3611 5729 3617
rect 5763 3611 5803 3617
rect 5837 3611 5877 3617
rect 5911 3611 5951 3617
rect 5985 3611 6025 3617
rect 6059 3611 6099 3617
rect 6133 3611 6173 3617
rect 6207 3611 6247 3617
rect 6450 3611 6535 3617
rect 7026 3608 7064 3617
rect 7098 3608 7136 3617
rect 7170 3608 7208 3617
rect 7242 3608 7280 3617
rect 7314 3608 7353 3617
rect 7387 3608 7426 3617
rect 7460 3608 7499 3617
rect 467 3572 522 3604
rect 501 3570 522 3572
rect 556 3593 713 3604
rect 556 3570 593 3593
rect 501 3559 593 3570
rect 627 3559 679 3593
rect 501 3538 713 3559
rect 467 3536 713 3538
rect 467 3502 522 3536
rect 556 3522 713 3536
rect 556 3502 593 3522
rect 467 3498 593 3502
rect 501 3488 593 3498
rect 627 3488 679 3522
rect 501 3476 713 3488
rect 7838 3606 7872 3616
rect 7838 3538 7872 3541
rect 7838 3500 7872 3504
rect 501 3468 660 3476
rect 501 3464 522 3468
rect 467 3434 522 3464
rect 556 3451 660 3468
rect 694 3451 713 3476
rect 962 3473 1006 3482
rect 1040 3473 1084 3482
rect 1118 3473 1162 3482
rect 1196 3473 1239 3482
rect 1273 3473 1316 3482
rect 1350 3473 1393 3482
rect 1427 3473 1470 3482
rect 1504 3473 1547 3482
rect 1581 3473 1624 3482
rect 1819 3473 1859 3476
rect 1893 3473 1932 3476
rect 1966 3473 2005 3476
rect 2039 3473 2078 3476
rect 2112 3473 2151 3476
rect 2185 3473 2224 3476
rect 2258 3473 2297 3476
rect 2331 3473 2370 3476
rect 2404 3473 2443 3476
rect 2477 3473 2516 3476
rect 2550 3473 2589 3476
rect 2623 3473 2662 3476
rect 2696 3473 2735 3476
rect 2769 3473 2808 3476
rect 2842 3473 2881 3476
rect 2915 3473 2954 3476
rect 2988 3473 3027 3476
rect 3061 3473 3100 3476
rect 3134 3473 3173 3476
rect 3207 3473 3246 3476
rect 3280 3473 3319 3476
rect 3353 3473 3392 3476
rect 3426 3473 3465 3476
rect 3499 3473 3538 3476
rect 3572 3473 3611 3476
rect 3645 3473 3684 3476
rect 3895 3473 3946 3476
rect 3980 3473 4031 3476
rect 4065 3473 4116 3476
rect 4150 3473 4201 3476
rect 4407 3473 4458 3476
rect 4492 3473 4543 3476
rect 4577 3473 4628 3476
rect 4662 3473 4713 3476
rect 4919 3473 4998 3476
rect 5146 3473 5192 3476
rect 5226 3473 5272 3476
rect 5306 3473 5352 3476
rect 5386 3473 5431 3476
rect 5465 3473 5510 3476
rect 5658 3473 5700 3476
rect 5734 3473 5776 3476
rect 5810 3473 5852 3476
rect 5886 3473 5928 3476
rect 5962 3473 6004 3476
rect 6038 3473 6080 3476
rect 6114 3473 6156 3476
rect 6190 3473 6232 3476
rect 6266 3473 6308 3476
rect 6342 3473 6384 3476
rect 6418 3473 6459 3476
rect 6493 3473 6534 3476
rect 7026 3473 7064 3482
rect 7098 3473 7136 3482
rect 7170 3473 7208 3482
rect 7242 3473 7280 3482
rect 7314 3473 7353 3482
rect 7387 3473 7426 3482
rect 7460 3473 7499 3482
rect 556 3434 593 3451
rect 467 3424 593 3434
rect 501 3417 593 3424
rect 627 3442 660 3451
rect 627 3417 679 3442
rect 916 3448 928 3473
rect 916 3439 932 3448
rect 966 3439 1006 3473
rect 1040 3439 1080 3473
rect 1118 3448 1154 3473
rect 1196 3448 1228 3473
rect 1273 3448 1301 3473
rect 1350 3448 1374 3473
rect 1427 3448 1447 3473
rect 1504 3448 1520 3473
rect 1581 3448 1593 3473
rect 1658 3448 1666 3473
rect 1114 3439 1154 3448
rect 1188 3439 1228 3448
rect 1262 3439 1301 3448
rect 1335 3439 1374 3448
rect 1408 3439 1447 3448
rect 1481 3439 1520 3448
rect 1554 3439 1593 3448
rect 1627 3439 1666 3448
rect 1700 3439 1716 3473
rect 1772 3442 1785 3473
rect 1772 3439 1788 3442
rect 1822 3439 1856 3473
rect 1893 3442 1924 3473
rect 1966 3442 1992 3473
rect 2039 3442 2060 3473
rect 2112 3442 2128 3473
rect 2185 3442 2196 3473
rect 2258 3442 2264 3473
rect 2331 3442 2332 3473
rect 1890 3439 1924 3442
rect 1958 3439 1992 3442
rect 2026 3439 2060 3442
rect 2094 3439 2128 3442
rect 2162 3439 2196 3442
rect 2230 3439 2264 3442
rect 2298 3439 2332 3442
rect 2366 3442 2370 3473
rect 2434 3442 2443 3473
rect 2502 3442 2516 3473
rect 2570 3442 2589 3473
rect 2638 3442 2662 3473
rect 2706 3442 2735 3473
rect 2366 3439 2400 3442
rect 2434 3439 2468 3442
rect 2502 3439 2536 3442
rect 2570 3439 2604 3442
rect 2638 3439 2672 3442
rect 2706 3439 2740 3442
rect 2774 3439 2808 3473
rect 2842 3439 2876 3473
rect 2915 3442 2944 3473
rect 2988 3442 3012 3473
rect 3061 3442 3080 3473
rect 3134 3442 3148 3473
rect 3207 3442 3216 3473
rect 3280 3442 3284 3473
rect 2910 3439 2944 3442
rect 2978 3439 3012 3442
rect 3046 3439 3080 3442
rect 3114 3439 3148 3442
rect 3182 3439 3216 3442
rect 3250 3439 3284 3442
rect 3318 3442 3319 3473
rect 3386 3442 3392 3473
rect 3454 3442 3465 3473
rect 3522 3442 3538 3473
rect 3590 3442 3611 3473
rect 3658 3442 3684 3473
rect 3318 3439 3352 3442
rect 3386 3439 3420 3442
rect 3454 3439 3488 3442
rect 3522 3439 3556 3442
rect 3590 3439 3624 3442
rect 3658 3439 3692 3442
rect 3726 3439 3760 3473
rect 3794 3439 3828 3473
rect 3895 3442 3896 3473
rect 3862 3439 3896 3442
rect 3930 3442 3946 3473
rect 3998 3442 4031 3473
rect 3930 3439 3964 3442
rect 3998 3439 4032 3442
rect 4066 3439 4100 3473
rect 4150 3442 4168 3473
rect 4235 3442 4236 3473
rect 4134 3439 4168 3442
rect 4202 3439 4236 3442
rect 4270 3439 4304 3473
rect 4338 3439 4373 3473
rect 4407 3439 4442 3473
rect 4492 3442 4511 3473
rect 4577 3442 4580 3473
rect 4476 3439 4511 3442
rect 4545 3439 4580 3442
rect 4614 3442 4628 3473
rect 4683 3442 4713 3473
rect 4614 3439 4649 3442
rect 4683 3439 4718 3442
rect 4752 3439 4787 3473
rect 4821 3439 4856 3473
rect 4919 3442 4925 3473
rect 4890 3439 4925 3442
rect 4959 3439 4994 3473
rect 5032 3442 5044 3473
rect 5028 3439 5044 3442
rect 5100 3442 5112 3473
rect 5150 3442 5192 3473
rect 5100 3439 5116 3442
rect 5150 3439 5194 3442
rect 5228 3439 5272 3473
rect 5306 3439 5350 3473
rect 5386 3442 5428 3473
rect 5465 3442 5506 3473
rect 5544 3442 5556 3473
rect 5384 3439 5428 3442
rect 5462 3439 5506 3442
rect 5540 3439 5556 3442
rect 5612 3442 5624 3473
rect 5612 3439 5628 3442
rect 5662 3439 5697 3473
rect 5734 3442 5766 3473
rect 5810 3442 5835 3473
rect 5886 3442 5904 3473
rect 5962 3442 5973 3473
rect 6038 3442 6042 3473
rect 5731 3439 5766 3442
rect 5800 3439 5835 3442
rect 5869 3439 5904 3442
rect 5938 3439 5973 3442
rect 6007 3439 6042 3442
rect 6076 3442 6080 3473
rect 6145 3442 6156 3473
rect 6214 3442 6232 3473
rect 6284 3442 6308 3473
rect 6354 3442 6384 3473
rect 6424 3442 6459 3473
rect 6076 3439 6111 3442
rect 6145 3439 6180 3442
rect 6214 3439 6250 3442
rect 6284 3439 6320 3442
rect 6354 3439 6390 3442
rect 6424 3439 6460 3442
rect 6494 3439 6530 3473
rect 6568 3442 6580 3473
rect 6564 3439 6580 3442
rect 6636 3439 6652 3473
rect 6686 3439 6722 3473
rect 6756 3439 6792 3473
rect 6826 3439 6862 3473
rect 6896 3439 6932 3473
rect 6966 3448 6992 3473
rect 7037 3448 7064 3473
rect 7108 3448 7136 3473
rect 7179 3448 7208 3473
rect 7250 3448 7280 3473
rect 7321 3448 7353 3473
rect 7392 3448 7426 3473
rect 7463 3448 7499 3473
rect 6966 3439 7003 3448
rect 7037 3439 7074 3448
rect 7108 3439 7145 3448
rect 7179 3439 7216 3448
rect 7250 3439 7287 3448
rect 7321 3439 7358 3448
rect 7392 3439 7429 3448
rect 7463 3439 7500 3448
rect 7534 3439 7571 3473
rect 7605 3439 7642 3473
rect 7676 3439 7692 3473
rect 501 3400 713 3417
rect 501 3390 522 3400
rect 467 3366 522 3390
rect 556 3394 713 3400
rect 556 3380 660 3394
rect 694 3380 713 3394
rect 7838 3425 7872 3436
rect 556 3366 593 3380
rect 467 3350 593 3366
rect 501 3346 593 3350
rect 627 3360 660 3380
rect 627 3346 679 3360
rect 501 3332 713 3346
rect 501 3316 522 3332
rect 467 3298 522 3316
rect 556 3311 713 3332
rect 556 3309 660 3311
rect 694 3309 713 3311
rect 556 3298 593 3309
rect 467 3276 593 3298
rect 501 3275 593 3276
rect 627 3277 660 3309
rect 871 3327 905 3349
rect 1727 3327 1761 3349
rect 1983 3327 2017 3349
rect 2239 3327 2273 3349
rect 2495 3327 2529 3349
rect 2751 3327 2785 3349
rect 3007 3327 3041 3349
rect 3263 3327 3297 3349
rect 3519 3327 3553 3349
rect 3775 3327 3809 3349
rect 4031 3327 4065 3349
rect 4287 3327 4321 3349
rect 4543 3327 4577 3349
rect 4799 3327 4833 3349
rect 5055 3327 5089 3349
rect 5311 3327 5345 3349
rect 5567 3327 5601 3349
rect 5823 3327 5857 3349
rect 6079 3327 6113 3349
rect 6335 3327 6369 3349
rect 6591 3327 6625 3349
rect 6847 3327 6881 3349
rect 7703 3327 7737 3349
rect 7838 3350 7872 3368
rect 627 3275 679 3277
rect 501 3264 713 3275
rect 501 3242 522 3264
rect 467 3230 522 3242
rect 556 3238 713 3264
rect 556 3230 593 3238
rect 467 3204 593 3230
rect 627 3204 679 3238
rect 467 3202 713 3204
rect 501 3196 713 3202
rect 501 3168 522 3196
rect 467 3162 522 3168
rect 556 3162 713 3196
rect 467 3128 713 3162
rect 7838 3275 7872 3300
rect 7838 3200 7872 3232
rect 7838 3128 7872 3164
rect 467 3094 482 3128
rect 516 3094 630 3128
rect 664 3094 698 3128
rect 732 3094 766 3128
rect 800 3094 834 3128
rect 868 3094 902 3128
rect 936 3094 970 3128
rect 1004 3094 1038 3128
rect 1072 3111 1106 3128
rect 1140 3111 1174 3128
rect 1208 3111 1242 3128
rect 1276 3111 1310 3128
rect 1344 3111 1378 3128
rect 1412 3111 1446 3128
rect 1480 3111 1514 3128
rect 1072 3094 1077 3111
rect 1140 3094 1150 3111
rect 1208 3094 1223 3111
rect 1276 3094 1296 3111
rect 1344 3094 1368 3111
rect 1412 3094 1440 3111
rect 1480 3094 1512 3111
rect 1548 3094 1582 3128
rect 1616 3111 1650 3128
rect 1684 3111 1718 3128
rect 1752 3111 1786 3128
rect 1820 3111 1854 3128
rect 1888 3111 1922 3128
rect 1956 3111 1990 3128
rect 2024 3111 2058 3128
rect 2092 3111 2126 3128
rect 1618 3094 1650 3111
rect 1690 3094 1718 3111
rect 1762 3094 1786 3111
rect 1834 3094 1854 3111
rect 1906 3094 1922 3111
rect 1978 3094 1990 3111
rect 2050 3094 2058 3111
rect 2122 3094 2126 3111
rect 2160 3111 2194 3128
rect 1111 3077 1150 3094
rect 1184 3077 1223 3094
rect 1257 3077 1296 3094
rect 1330 3077 1368 3094
rect 1402 3077 1440 3094
rect 1474 3077 1512 3094
rect 1546 3077 1584 3094
rect 1618 3077 1656 3094
rect 1690 3077 1728 3094
rect 1762 3077 1800 3094
rect 1834 3077 1872 3094
rect 1906 3077 1944 3094
rect 1978 3077 2016 3094
rect 2050 3077 2088 3094
rect 2122 3077 2160 3094
rect 2228 3111 2262 3128
rect 2296 3111 2330 3128
rect 2364 3111 2398 3128
rect 2432 3111 2466 3128
rect 2500 3111 2534 3128
rect 2568 3111 2602 3128
rect 2636 3111 2670 3128
rect 2704 3111 2738 3128
rect 2228 3094 2232 3111
rect 2296 3094 2304 3111
rect 2364 3094 2376 3111
rect 2432 3094 2448 3111
rect 2500 3094 2520 3111
rect 2568 3094 2592 3111
rect 2636 3094 2664 3111
rect 2704 3094 2736 3111
rect 2772 3094 2806 3128
rect 2840 3111 2874 3128
rect 2908 3111 2942 3128
rect 2976 3111 3010 3128
rect 3044 3111 3078 3128
rect 3112 3111 3146 3128
rect 3180 3111 3214 3128
rect 3248 3111 3282 3128
rect 3316 3111 3350 3128
rect 2842 3094 2874 3111
rect 2914 3094 2942 3111
rect 2986 3094 3010 3111
rect 3058 3094 3078 3111
rect 3130 3094 3146 3111
rect 3202 3094 3214 3111
rect 3274 3094 3282 3111
rect 3346 3094 3350 3111
rect 3384 3111 3418 3128
rect 2194 3077 2232 3094
rect 2266 3077 2304 3094
rect 2338 3077 2376 3094
rect 2410 3077 2448 3094
rect 2482 3077 2520 3094
rect 2554 3077 2592 3094
rect 2626 3077 2664 3094
rect 2698 3077 2736 3094
rect 2770 3077 2808 3094
rect 2842 3077 2880 3094
rect 2914 3077 2952 3094
rect 2986 3077 3024 3094
rect 3058 3077 3096 3094
rect 3130 3077 3168 3094
rect 3202 3077 3240 3094
rect 3274 3077 3312 3094
rect 3346 3077 3384 3094
rect 3452 3111 3486 3128
rect 3520 3111 3554 3128
rect 3588 3111 3622 3128
rect 3656 3111 3690 3128
rect 3724 3111 3758 3128
rect 3452 3094 3456 3111
rect 3520 3094 3528 3111
rect 3588 3094 3600 3111
rect 3656 3094 3672 3111
rect 3724 3094 3744 3111
rect 3792 3094 3826 3128
rect 3860 3094 3888 3128
rect 3928 3094 3962 3128
rect 3996 3094 4030 3128
rect 4070 3094 4098 3128
rect 4144 3094 4166 3128
rect 4218 3094 4234 3128
rect 4292 3094 4302 3128
rect 4366 3094 4370 3128
rect 4404 3094 4406 3128
rect 4472 3094 4480 3128
rect 4540 3094 4553 3128
rect 4608 3094 4626 3128
rect 4676 3094 4699 3128
rect 4744 3094 4772 3128
rect 4812 3094 4845 3128
rect 4880 3094 4914 3128
rect 4952 3094 4982 3128
rect 5025 3094 5050 3128
rect 5098 3094 5118 3128
rect 5171 3094 5186 3128
rect 5244 3094 5254 3128
rect 5317 3094 5322 3128
rect 5424 3094 5429 3128
rect 5492 3094 5502 3128
rect 5560 3094 5575 3128
rect 5628 3094 5648 3128
rect 5696 3094 5721 3128
rect 5764 3094 5794 3128
rect 5832 3094 5866 3128
rect 5901 3094 5934 3128
rect 5974 3094 6002 3128
rect 6047 3094 6070 3128
rect 6120 3094 6138 3128
rect 6193 3094 6206 3128
rect 6266 3094 6274 3128
rect 6339 3094 6342 3128
rect 6376 3094 6378 3128
rect 6444 3094 6451 3128
rect 6512 3094 6524 3128
rect 6580 3094 6597 3128
rect 6648 3094 6670 3128
rect 6716 3094 6743 3128
rect 6784 3094 6816 3128
rect 6852 3094 6886 3128
rect 6923 3094 6954 3128
rect 6996 3094 7022 3128
rect 7069 3094 7090 3128
rect 7142 3094 7158 3128
rect 7215 3094 7226 3128
rect 7288 3094 7294 3128
rect 7361 3094 7362 3128
rect 7396 3094 7400 3128
rect 7464 3094 7473 3128
rect 7532 3094 7546 3128
rect 7600 3094 7619 3128
rect 7668 3094 7692 3128
rect 7736 3094 7765 3128
rect 7804 3094 7872 3128
rect 8476 4917 20013 4918
rect 8476 4883 8550 4917
rect 8584 4912 8620 4917
rect 8654 4912 8690 4917
rect 8724 4912 8760 4917
rect 8794 4912 8830 4917
rect 8864 4912 8900 4917
rect 8934 4912 8970 4917
rect 9004 4912 9040 4917
rect 9074 4912 9110 4917
rect 9144 4912 9180 4917
rect 9214 4912 9250 4917
rect 8588 4883 8620 4912
rect 8661 4883 8690 4912
rect 8734 4883 8760 4912
rect 8807 4883 8830 4912
rect 8880 4883 8900 4912
rect 8953 4883 8970 4912
rect 9026 4883 9040 4912
rect 9099 4883 9110 4912
rect 9172 4883 9180 4912
rect 9245 4883 9250 4912
rect 9284 4912 9320 4917
rect 8476 4878 8554 4883
rect 8588 4878 8627 4883
rect 8661 4878 8700 4883
rect 8734 4878 8773 4883
rect 8807 4878 8846 4883
rect 8880 4878 8919 4883
rect 8953 4878 8992 4883
rect 9026 4878 9065 4883
rect 9099 4878 9138 4883
rect 9172 4878 9211 4883
rect 9245 4878 9284 4883
rect 9318 4883 9320 4912
rect 9354 4912 9390 4917
rect 9424 4912 9460 4917
rect 9494 4912 9530 4917
rect 9564 4912 9599 4917
rect 9633 4912 9668 4917
rect 9702 4912 9737 4917
rect 9771 4912 9806 4917
rect 9840 4912 9875 4917
rect 9909 4912 9944 4917
rect 9354 4883 9357 4912
rect 9424 4883 9430 4912
rect 9494 4883 9503 4912
rect 9564 4883 9576 4912
rect 9633 4883 9649 4912
rect 9702 4883 9722 4912
rect 9771 4883 9795 4912
rect 9840 4883 9868 4912
rect 9909 4883 9941 4912
rect 9978 4883 10013 4917
rect 10047 4912 10082 4917
rect 10116 4912 10151 4917
rect 10185 4912 10220 4917
rect 10254 4912 10289 4917
rect 10323 4912 10358 4917
rect 10392 4912 10427 4917
rect 10461 4912 10496 4917
rect 10530 4912 10565 4917
rect 10599 4912 10634 4917
rect 10048 4883 10082 4912
rect 10121 4883 10151 4912
rect 10194 4883 10220 4912
rect 10267 4883 10289 4912
rect 10340 4883 10358 4912
rect 10413 4883 10427 4912
rect 10486 4883 10496 4912
rect 10559 4883 10565 4912
rect 10632 4883 10634 4912
rect 10668 4912 10703 4917
rect 10737 4912 10772 4917
rect 10806 4912 10841 4917
rect 10875 4912 10910 4917
rect 10944 4912 10979 4917
rect 11013 4912 11048 4917
rect 11082 4912 11117 4917
rect 11151 4912 11186 4917
rect 11220 4912 11322 4917
rect 11356 4912 11391 4917
rect 11425 4912 11460 4917
rect 11494 4912 11529 4917
rect 11563 4912 11598 4917
rect 11632 4912 11667 4917
rect 11701 4912 11736 4917
rect 11770 4912 11805 4917
rect 11839 4912 11874 4917
rect 10668 4883 10671 4912
rect 10737 4883 10744 4912
rect 10806 4883 10817 4912
rect 10875 4883 10890 4912
rect 10944 4883 10963 4912
rect 11013 4883 11036 4912
rect 11082 4883 11109 4912
rect 11151 4883 11182 4912
rect 11220 4883 11255 4912
rect 9318 4878 9357 4883
rect 9391 4878 9430 4883
rect 9464 4878 9503 4883
rect 9537 4878 9576 4883
rect 9610 4878 9649 4883
rect 9683 4878 9722 4883
rect 9756 4878 9795 4883
rect 9829 4878 9868 4883
rect 9902 4878 9941 4883
rect 9975 4878 10014 4883
rect 10048 4878 10087 4883
rect 10121 4878 10160 4883
rect 10194 4878 10233 4883
rect 10267 4878 10306 4883
rect 10340 4878 10379 4883
rect 10413 4878 10452 4883
rect 10486 4878 10525 4883
rect 10559 4878 10598 4883
rect 10632 4878 10671 4883
rect 10705 4878 10744 4883
rect 10778 4878 10817 4883
rect 10851 4878 10890 4883
rect 10924 4878 10963 4883
rect 10997 4878 11036 4883
rect 11070 4878 11109 4883
rect 11143 4878 11182 4883
rect 11216 4878 11255 4883
rect 11289 4883 11322 4912
rect 11362 4883 11391 4912
rect 11435 4883 11460 4912
rect 11508 4883 11529 4912
rect 11581 4883 11598 4912
rect 11654 4883 11667 4912
rect 11727 4883 11736 4912
rect 11799 4883 11805 4912
rect 11871 4883 11874 4912
rect 11908 4912 11943 4917
rect 11908 4883 11909 4912
rect 11289 4878 11328 4883
rect 11362 4878 11401 4883
rect 11435 4878 11474 4883
rect 11508 4878 11547 4883
rect 11581 4878 11620 4883
rect 11654 4878 11693 4883
rect 11727 4878 11765 4883
rect 11799 4878 11837 4883
rect 11871 4878 11909 4883
rect 11977 4912 12012 4917
rect 12046 4912 12081 4917
rect 12115 4912 12150 4917
rect 12184 4912 12219 4917
rect 12253 4912 12288 4917
rect 12322 4912 12357 4917
rect 12391 4912 12426 4917
rect 12460 4912 12495 4917
rect 12529 4912 12563 4917
rect 12597 4912 12631 4917
rect 11977 4883 11981 4912
rect 12046 4883 12053 4912
rect 12115 4883 12125 4912
rect 12184 4883 12197 4912
rect 12253 4883 12269 4912
rect 12322 4883 12341 4912
rect 12391 4883 12413 4912
rect 12460 4883 12485 4912
rect 12529 4883 12557 4912
rect 12597 4883 12629 4912
rect 12665 4883 12699 4917
rect 12733 4912 12767 4917
rect 12801 4912 12835 4917
rect 12869 4912 12903 4917
rect 12937 4912 12971 4917
rect 13005 4912 13039 4917
rect 13073 4912 13107 4917
rect 13141 4912 13175 4917
rect 13209 4912 13243 4917
rect 12735 4883 12767 4912
rect 12807 4883 12835 4912
rect 12879 4883 12903 4912
rect 12951 4883 12971 4912
rect 13023 4883 13039 4912
rect 13095 4883 13107 4912
rect 13167 4883 13175 4912
rect 13239 4883 13243 4912
rect 13277 4912 13311 4917
rect 11943 4878 11981 4883
rect 12015 4878 12053 4883
rect 12087 4878 12125 4883
rect 12159 4878 12197 4883
rect 12231 4878 12269 4883
rect 12303 4878 12341 4883
rect 12375 4878 12413 4883
rect 12447 4878 12485 4883
rect 12519 4878 12557 4883
rect 12591 4878 12629 4883
rect 12663 4878 12701 4883
rect 12735 4878 12773 4883
rect 12807 4878 12845 4883
rect 12879 4878 12917 4883
rect 12951 4878 12989 4883
rect 13023 4878 13061 4883
rect 13095 4878 13133 4883
rect 13167 4878 13205 4883
rect 13239 4878 13277 4883
rect 13345 4912 13379 4917
rect 13413 4912 13447 4917
rect 13481 4912 13515 4917
rect 13549 4912 13583 4917
rect 13617 4912 13651 4917
rect 13685 4912 13719 4917
rect 13753 4912 13787 4917
rect 13821 4912 13855 4917
rect 13345 4883 13349 4912
rect 13413 4883 13421 4912
rect 13481 4883 13493 4912
rect 13549 4883 13565 4912
rect 13617 4883 13637 4912
rect 13685 4883 13709 4912
rect 13753 4883 13781 4912
rect 13821 4883 13853 4912
rect 13889 4883 13923 4917
rect 13957 4912 13991 4917
rect 14025 4912 14059 4917
rect 14093 4912 14127 4917
rect 14161 4912 14195 4917
rect 14229 4912 14263 4917
rect 14297 4912 14331 4917
rect 14365 4912 14399 4917
rect 14433 4912 14467 4917
rect 13959 4883 13991 4912
rect 14031 4883 14059 4912
rect 14103 4883 14127 4912
rect 14175 4883 14195 4912
rect 14247 4883 14263 4912
rect 14319 4883 14331 4912
rect 14391 4883 14399 4912
rect 14463 4883 14467 4912
rect 14501 4912 14535 4917
rect 13311 4878 13349 4883
rect 13383 4878 13421 4883
rect 13455 4878 13493 4883
rect 13527 4878 13565 4883
rect 13599 4878 13637 4883
rect 13671 4878 13709 4883
rect 13743 4878 13781 4883
rect 13815 4878 13853 4883
rect 13887 4878 13925 4883
rect 13959 4878 13997 4883
rect 14031 4878 14069 4883
rect 14103 4878 14141 4883
rect 14175 4878 14213 4883
rect 14247 4878 14285 4883
rect 14319 4878 14357 4883
rect 14391 4878 14429 4883
rect 14463 4878 14501 4883
rect 14569 4912 14603 4917
rect 14637 4912 14671 4917
rect 14705 4912 14739 4917
rect 14773 4912 14807 4917
rect 14841 4912 14875 4917
rect 14909 4912 14943 4917
rect 14977 4912 15011 4917
rect 15045 4912 15079 4917
rect 14569 4883 14573 4912
rect 14637 4883 14645 4912
rect 14705 4883 14717 4912
rect 14773 4883 14789 4912
rect 14841 4883 14861 4912
rect 14909 4883 14933 4912
rect 14977 4883 15005 4912
rect 15045 4883 15077 4912
rect 15113 4883 15147 4917
rect 15181 4912 15215 4917
rect 15249 4912 15283 4917
rect 15317 4912 15351 4917
rect 15385 4912 15419 4917
rect 15453 4912 15487 4917
rect 15521 4912 15555 4917
rect 15589 4912 15623 4917
rect 15657 4912 15691 4917
rect 15183 4883 15215 4912
rect 15255 4883 15283 4912
rect 15327 4883 15351 4912
rect 15399 4883 15419 4912
rect 15471 4883 15487 4912
rect 15543 4883 15555 4912
rect 15615 4883 15623 4912
rect 15687 4883 15691 4912
rect 15725 4912 15759 4917
rect 14535 4878 14573 4883
rect 14607 4878 14645 4883
rect 14679 4878 14717 4883
rect 14751 4878 14789 4883
rect 14823 4878 14861 4883
rect 14895 4878 14933 4883
rect 14967 4878 15005 4883
rect 15039 4878 15077 4883
rect 15111 4878 15149 4883
rect 15183 4878 15221 4883
rect 15255 4878 15293 4883
rect 15327 4878 15365 4883
rect 15399 4878 15437 4883
rect 15471 4878 15509 4883
rect 15543 4878 15581 4883
rect 15615 4878 15653 4883
rect 15687 4878 15725 4883
rect 15793 4912 15827 4917
rect 15861 4912 15895 4917
rect 15929 4912 15963 4917
rect 15997 4912 16031 4917
rect 16065 4912 16099 4917
rect 16133 4912 16167 4917
rect 16201 4912 16235 4917
rect 16269 4912 16303 4917
rect 15793 4883 15797 4912
rect 15861 4883 15869 4912
rect 15929 4883 15941 4912
rect 15997 4883 16013 4912
rect 16065 4883 16085 4912
rect 16133 4883 16157 4912
rect 16201 4883 16229 4912
rect 16269 4883 16301 4912
rect 16337 4883 16371 4917
rect 16405 4912 16439 4917
rect 16473 4912 16507 4917
rect 16541 4912 16575 4917
rect 16609 4912 16643 4917
rect 16677 4912 16711 4917
rect 16745 4912 16779 4917
rect 16813 4912 16847 4917
rect 16881 4912 16915 4917
rect 16407 4883 16439 4912
rect 16479 4883 16507 4912
rect 16551 4883 16575 4912
rect 16623 4883 16643 4912
rect 16695 4883 16711 4912
rect 16767 4883 16779 4912
rect 16839 4883 16847 4912
rect 16911 4883 16915 4912
rect 16949 4912 16983 4917
rect 15759 4878 15797 4883
rect 15831 4878 15869 4883
rect 15903 4878 15941 4883
rect 15975 4878 16013 4883
rect 16047 4878 16085 4883
rect 16119 4878 16157 4883
rect 16191 4878 16229 4883
rect 16263 4878 16301 4883
rect 16335 4878 16373 4883
rect 16407 4878 16445 4883
rect 16479 4878 16517 4883
rect 16551 4878 16589 4883
rect 16623 4878 16661 4883
rect 16695 4878 16733 4883
rect 16767 4878 16805 4883
rect 16839 4878 16877 4883
rect 16911 4878 16949 4883
rect 17017 4912 17051 4917
rect 17085 4912 17119 4917
rect 17153 4912 17187 4917
rect 17221 4912 17255 4917
rect 17289 4912 17323 4917
rect 17357 4912 17391 4917
rect 17425 4912 17459 4917
rect 17493 4912 17527 4917
rect 17017 4883 17021 4912
rect 17085 4883 17093 4912
rect 17153 4883 17165 4912
rect 17221 4883 17237 4912
rect 17289 4883 17309 4912
rect 17357 4883 17381 4912
rect 17425 4883 17453 4912
rect 17493 4883 17525 4912
rect 17561 4883 17595 4917
rect 17629 4912 17663 4917
rect 17697 4912 17731 4917
rect 17765 4912 17799 4917
rect 17833 4912 17867 4917
rect 17901 4912 17935 4917
rect 17969 4912 18003 4917
rect 18037 4912 18071 4917
rect 18105 4912 18139 4917
rect 17631 4883 17663 4912
rect 17703 4883 17731 4912
rect 17775 4883 17799 4912
rect 17847 4883 17867 4912
rect 17919 4883 17935 4912
rect 17991 4883 18003 4912
rect 18063 4883 18071 4912
rect 18135 4883 18139 4912
rect 18173 4912 18207 4917
rect 16983 4878 17021 4883
rect 17055 4878 17093 4883
rect 17127 4878 17165 4883
rect 17199 4878 17237 4883
rect 17271 4878 17309 4883
rect 17343 4878 17381 4883
rect 17415 4878 17453 4883
rect 17487 4878 17525 4883
rect 17559 4878 17597 4883
rect 17631 4878 17669 4883
rect 17703 4878 17741 4883
rect 17775 4878 17813 4883
rect 17847 4878 17885 4883
rect 17919 4878 17957 4883
rect 17991 4878 18029 4883
rect 18063 4878 18101 4883
rect 18135 4878 18173 4883
rect 18241 4912 18275 4917
rect 18309 4912 18343 4917
rect 18377 4912 18411 4917
rect 18445 4912 18479 4917
rect 18513 4912 18547 4917
rect 18581 4912 18615 4917
rect 18649 4912 18683 4917
rect 18717 4912 18751 4917
rect 18241 4883 18245 4912
rect 18309 4883 18317 4912
rect 18377 4883 18389 4912
rect 18445 4883 18461 4912
rect 18513 4883 18533 4912
rect 18581 4883 18605 4912
rect 18649 4883 18677 4912
rect 18717 4883 18749 4912
rect 18785 4883 18819 4917
rect 18853 4912 18887 4917
rect 18921 4912 18955 4917
rect 18989 4912 19023 4917
rect 19057 4912 19091 4917
rect 19125 4912 19159 4917
rect 19193 4912 19227 4917
rect 19261 4912 19295 4917
rect 19329 4912 19363 4917
rect 18855 4883 18887 4912
rect 18927 4883 18955 4912
rect 18999 4883 19023 4912
rect 19071 4883 19091 4912
rect 19143 4883 19159 4912
rect 19215 4883 19227 4912
rect 19287 4883 19295 4912
rect 19359 4883 19363 4912
rect 19397 4912 19431 4917
rect 18207 4878 18245 4883
rect 18279 4878 18317 4883
rect 18351 4878 18389 4883
rect 18423 4878 18461 4883
rect 18495 4878 18533 4883
rect 18567 4878 18605 4883
rect 18639 4878 18677 4883
rect 18711 4878 18749 4883
rect 18783 4878 18821 4883
rect 18855 4878 18893 4883
rect 18927 4878 18965 4883
rect 18999 4878 19037 4883
rect 19071 4878 19109 4883
rect 19143 4878 19181 4883
rect 19215 4878 19253 4883
rect 19287 4878 19325 4883
rect 19359 4878 19397 4883
rect 19465 4912 19499 4917
rect 19533 4912 19567 4917
rect 19601 4912 19635 4917
rect 19669 4912 19703 4917
rect 19737 4912 19771 4917
rect 19805 4912 19839 4917
rect 19873 4912 19907 4917
rect 19465 4883 19469 4912
rect 19533 4883 19541 4912
rect 19601 4883 19613 4912
rect 19669 4883 19685 4912
rect 19737 4883 19757 4912
rect 19805 4883 19829 4912
rect 19873 4883 19901 4912
rect 19941 4883 20013 4917
rect 19431 4878 19469 4883
rect 19503 4878 19541 4883
rect 19575 4878 19613 4883
rect 19647 4878 19685 4883
rect 19719 4878 19757 4883
rect 19791 4878 19829 4883
rect 19863 4878 19901 4883
rect 19935 4878 20013 4883
rect 8476 4872 20013 4878
rect 8476 4848 8522 4872
rect 8476 4804 8482 4848
rect 8516 4804 8522 4848
rect 11254 4840 11338 4872
rect 8476 4779 8522 4804
rect 8476 4730 8482 4779
rect 8516 4730 8522 4779
rect 8476 4710 8522 4730
rect 8476 4656 8482 4710
rect 8516 4656 8522 4710
rect 8476 4641 8522 4656
rect 8476 4582 8482 4641
rect 8516 4582 8522 4641
rect 8476 4572 8522 4582
rect 8476 4508 8482 4572
rect 8516 4508 8522 4572
rect 8476 4503 8522 4508
rect 8476 4469 8482 4503
rect 8516 4469 8522 4503
rect 8476 4468 8522 4469
rect 8476 4400 8482 4468
rect 8516 4400 8522 4468
rect 8476 4394 8522 4400
rect 8476 4331 8482 4394
rect 8516 4331 8522 4394
rect 8476 4320 8522 4331
rect 8476 4262 8482 4320
rect 8516 4262 8522 4320
rect 8476 4246 8522 4262
rect 8476 4192 8482 4246
rect 8516 4192 8522 4246
rect 8476 4172 8522 4192
rect 8476 4122 8482 4172
rect 8516 4122 8522 4172
rect 8476 4098 8522 4122
rect 8476 4052 8482 4098
rect 8516 4052 8522 4098
rect 8476 4024 8522 4052
rect 8476 3982 8482 4024
rect 8516 3982 8522 4024
rect 8476 3950 8522 3982
rect 8476 3912 8482 3950
rect 8516 3912 8522 3950
rect 8476 3876 8522 3912
rect 8476 3842 8482 3876
rect 8516 3842 8522 3876
rect 8476 3806 8522 3842
rect 8714 4736 8748 4758
rect 8714 4664 8748 4690
rect 8714 4592 8748 4622
rect 8714 4520 8748 4554
rect 8714 4452 8748 4486
rect 8714 4384 8748 4414
rect 8714 4316 8748 4342
rect 8714 4248 8748 4270
rect 8714 4180 8748 4198
rect 8714 4112 8748 4126
rect 8714 4044 8748 4054
rect 8714 3976 8748 3982
rect 8714 3908 8748 3910
rect 8714 3872 8748 3874
rect 8870 4736 8904 4758
rect 8870 4664 8904 4690
rect 8870 4592 8904 4622
rect 8870 4520 8904 4554
rect 8870 4452 8904 4486
rect 8870 4384 8904 4414
rect 8870 4316 8904 4342
rect 8870 4248 8904 4270
rect 8870 4180 8904 4198
rect 8870 4112 8904 4126
rect 8870 4044 8904 4054
rect 8870 3976 8904 3982
rect 8870 3908 8904 3910
rect 8870 3872 8904 3874
rect 9026 4736 9060 4758
rect 9026 4664 9060 4690
rect 9026 4592 9060 4622
rect 9026 4520 9060 4554
rect 9026 4452 9060 4486
rect 9026 4384 9060 4414
rect 9026 4316 9060 4342
rect 9026 4248 9060 4270
rect 9026 4180 9060 4198
rect 9026 4112 9060 4126
rect 9026 4044 9060 4054
rect 9026 3976 9060 3982
rect 9026 3908 9060 3910
rect 9026 3872 9060 3874
rect 9182 4736 9216 4758
rect 9182 4664 9216 4690
rect 9182 4592 9216 4622
rect 9182 4520 9216 4554
rect 9182 4452 9216 4486
rect 9182 4384 9216 4414
rect 9182 4316 9216 4342
rect 9182 4248 9216 4270
rect 9182 4180 9216 4198
rect 9182 4112 9216 4126
rect 9182 4044 9216 4054
rect 9182 3976 9216 3982
rect 9182 3908 9216 3910
rect 9182 3872 9216 3874
rect 9338 4736 9372 4758
rect 9338 4664 9372 4690
rect 9338 4592 9372 4622
rect 9338 4520 9372 4554
rect 9338 4452 9372 4486
rect 9338 4384 9372 4414
rect 9338 4316 9372 4342
rect 9338 4248 9372 4270
rect 9338 4180 9372 4198
rect 9338 4112 9372 4126
rect 9338 4044 9372 4054
rect 9338 3976 9372 3982
rect 9338 3908 9372 3910
rect 9338 3872 9372 3874
rect 9462 4736 9496 4758
rect 9462 4664 9496 4690
rect 9462 4592 9496 4622
rect 9462 4520 9496 4554
rect 9462 4452 9496 4486
rect 9462 4384 9496 4414
rect 9462 4316 9496 4342
rect 9462 4248 9496 4270
rect 9462 4180 9496 4198
rect 9462 4112 9496 4126
rect 9462 4044 9496 4054
rect 9462 3976 9496 3982
rect 9462 3908 9496 3910
rect 9462 3872 9496 3874
rect 9618 4736 9652 4758
rect 9618 4664 9652 4690
rect 9618 4592 9652 4622
rect 9618 4520 9652 4554
rect 9618 4452 9652 4486
rect 9618 4384 9652 4414
rect 9618 4316 9652 4342
rect 9618 4248 9652 4270
rect 9618 4180 9652 4198
rect 9618 4112 9652 4126
rect 9618 4044 9652 4054
rect 9618 3976 9652 3982
rect 9618 3908 9652 3910
rect 9618 3872 9652 3874
rect 9742 4736 9776 4758
rect 9742 4664 9776 4690
rect 9742 4592 9776 4622
rect 9742 4520 9776 4554
rect 9742 4452 9776 4486
rect 9742 4384 9776 4414
rect 9742 4316 9776 4342
rect 9742 4248 9776 4270
rect 9742 4180 9776 4198
rect 9742 4112 9776 4126
rect 9742 4044 9776 4054
rect 9742 3976 9776 3982
rect 9742 3908 9776 3910
rect 9742 3872 9776 3874
rect 9898 4736 9932 4758
rect 9898 4664 9932 4690
rect 9898 4592 9932 4622
rect 9898 4520 9932 4554
rect 9898 4452 9932 4486
rect 9898 4384 9932 4414
rect 9898 4316 9932 4342
rect 9898 4248 9932 4270
rect 9898 4180 9932 4198
rect 9898 4112 9932 4126
rect 9898 4044 9932 4054
rect 9898 3976 9932 3982
rect 9898 3908 9932 3910
rect 9898 3872 9932 3874
rect 10054 4736 10088 4758
rect 10054 4664 10088 4690
rect 10054 4592 10088 4622
rect 10054 4520 10088 4554
rect 10054 4452 10088 4486
rect 10054 4384 10088 4414
rect 10054 4316 10088 4342
rect 10054 4248 10088 4270
rect 10054 4180 10088 4198
rect 10054 4112 10088 4126
rect 10054 4044 10088 4054
rect 10054 3976 10088 3982
rect 10054 3908 10088 3910
rect 10054 3872 10088 3874
rect 10331 4736 10365 4758
rect 10331 4664 10365 4690
rect 10331 4592 10365 4622
rect 10331 4520 10365 4554
rect 10331 4452 10365 4486
rect 10331 4384 10365 4414
rect 10331 4316 10365 4342
rect 10331 4248 10365 4270
rect 10331 4180 10365 4198
rect 10331 4112 10365 4126
rect 10331 4044 10365 4054
rect 10331 3976 10365 3982
rect 10331 3908 10365 3910
rect 10331 3872 10365 3874
rect 10487 4736 10521 4758
rect 10487 4664 10521 4690
rect 10487 4592 10521 4622
rect 10487 4520 10521 4554
rect 10487 4452 10521 4486
rect 10487 4384 10521 4414
rect 10487 4316 10521 4342
rect 10487 4248 10521 4270
rect 10487 4180 10521 4198
rect 10487 4112 10521 4126
rect 10487 4044 10521 4054
rect 10487 3976 10521 3982
rect 10487 3908 10521 3910
rect 10487 3872 10521 3874
rect 10643 4736 10677 4758
rect 10643 4664 10677 4690
rect 10643 4592 10677 4622
rect 10643 4520 10677 4554
rect 10643 4452 10677 4486
rect 10643 4384 10677 4414
rect 10643 4316 10677 4342
rect 10643 4248 10677 4270
rect 10643 4180 10677 4198
rect 10643 4112 10677 4126
rect 10643 4044 10677 4054
rect 10643 3976 10677 3982
rect 10643 3908 10677 3910
rect 10643 3872 10677 3874
rect 10799 4736 10833 4758
rect 10799 4664 10833 4690
rect 10799 4592 10833 4622
rect 10799 4520 10833 4554
rect 10799 4452 10833 4486
rect 10799 4384 10833 4414
rect 10799 4316 10833 4342
rect 10799 4248 10833 4270
rect 10799 4180 10833 4198
rect 10799 4112 10833 4126
rect 10799 4044 10833 4054
rect 10799 3976 10833 3982
rect 10799 3908 10833 3910
rect 10799 3872 10833 3874
rect 10955 4736 10989 4758
rect 10955 4664 10989 4690
rect 10955 4592 10989 4622
rect 10955 4520 10989 4554
rect 10955 4452 10989 4486
rect 10955 4384 10989 4414
rect 10955 4316 10989 4342
rect 10955 4248 10989 4270
rect 10955 4180 10989 4198
rect 10955 4112 10989 4126
rect 10955 4044 10989 4054
rect 10955 3976 10989 3982
rect 10955 3908 10989 3910
rect 10955 3872 10989 3874
rect 11111 4736 11145 4758
rect 11111 4664 11145 4690
rect 11111 4592 11145 4622
rect 11111 4520 11145 4554
rect 11111 4452 11145 4486
rect 11111 4384 11145 4414
rect 11111 4316 11145 4342
rect 11111 4248 11145 4270
rect 11111 4180 11145 4198
rect 11111 4112 11145 4126
rect 11111 4044 11145 4054
rect 11111 3976 11145 3982
rect 11111 3908 11145 3910
rect 11111 3872 11145 3874
rect 11254 4806 11298 4840
rect 11332 4806 11338 4840
rect 11254 4783 11338 4806
rect 11288 4766 11338 4783
rect 11288 4749 11298 4766
rect 11254 4732 11298 4749
rect 11332 4732 11338 4766
rect 11254 4715 11338 4732
rect 11288 4692 11338 4715
rect 11288 4681 11298 4692
rect 11254 4658 11298 4681
rect 11332 4658 11338 4692
rect 19967 4840 20013 4872
rect 19967 4806 19973 4840
rect 20007 4835 20013 4840
rect 19967 4801 19975 4806
rect 20009 4801 20013 4835
rect 19967 4767 20013 4801
rect 19967 4733 19973 4767
rect 20007 4733 20013 4767
rect 19967 4694 20013 4733
rect 19967 4660 19973 4694
rect 20007 4674 20013 4694
rect 11254 4647 11338 4658
rect 11288 4618 11338 4647
rect 11288 4613 11298 4618
rect 11254 4584 11298 4613
rect 11332 4584 11338 4618
rect 13527 4599 13584 4633
rect 11254 4579 11338 4584
rect 11288 4545 11338 4579
rect 17403 4588 17437 4626
rect 11254 4544 11338 4545
rect 11254 4511 11298 4544
rect 11288 4510 11298 4511
rect 11332 4510 11338 4544
rect 16755 4525 16793 4559
rect 17996 4588 18030 4626
rect 19967 4640 19975 4660
rect 20009 4640 20013 4674
rect 19967 4621 20013 4640
rect 19967 4587 19973 4621
rect 20007 4606 20013 4621
rect 19967 4572 19975 4587
rect 20009 4572 20013 4606
rect 11288 4477 11338 4510
rect 11254 4470 11338 4477
rect 11254 4443 11298 4470
rect 11288 4436 11298 4443
rect 11332 4436 11338 4470
rect 17684 4491 17718 4529
rect 19365 4492 19399 4530
rect 19609 4530 19627 4564
rect 19661 4530 19675 4564
rect 19609 4492 19675 4530
rect 19609 4458 19627 4492
rect 19661 4458 19675 4492
rect 11288 4409 11338 4436
rect 11254 4396 11338 4409
rect 11254 4375 11298 4396
rect 11288 4362 11298 4375
rect 11332 4362 11338 4396
rect 11288 4341 11338 4362
rect 14759 4377 14797 4411
rect 18503 4377 18541 4411
rect 19438 4405 19504 4423
rect 11254 4322 11338 4341
rect 13921 4337 13987 4353
rect 11254 4307 11298 4322
rect 11288 4288 11298 4307
rect 11332 4288 11338 4322
rect 11288 4273 11338 4288
rect 11254 4248 11338 4273
rect 11254 4239 11298 4248
rect 11288 4214 11298 4239
rect 11332 4214 11338 4248
rect 11288 4205 11338 4214
rect 11254 4174 11338 4205
rect 11254 4171 11298 4174
rect 11288 4140 11298 4171
rect 11332 4140 11338 4174
rect 11784 4311 11850 4324
rect 11784 4277 11801 4311
rect 11835 4277 11850 4311
rect 11784 4239 11850 4277
rect 13921 4303 13933 4337
rect 13967 4303 14005 4337
rect 11784 4205 11801 4239
rect 11835 4205 11850 4239
rect 13284 4220 13322 4254
rect 13356 4220 13358 4254
rect 11288 4137 11338 4140
rect 11254 4103 11338 4137
rect 11288 4100 11338 4103
rect 11288 4069 11298 4100
rect 11254 4066 11298 4069
rect 11332 4066 11338 4100
rect 11254 4035 11338 4066
rect 11784 4156 11850 4205
rect 12412 4157 12688 4196
rect 11580 4088 11614 4126
rect 12434 4123 12472 4157
rect 12506 4123 12688 4157
rect 13292 4156 13358 4220
rect 13921 4156 13987 4303
rect 14725 4156 14791 4377
rect 15144 4229 15182 4263
rect 16502 4231 16540 4265
rect 16574 4231 16575 4265
rect 17706 4231 17744 4265
rect 15529 4189 15595 4203
rect 15563 4155 15601 4189
rect 16509 4156 16575 4231
rect 18469 4156 18535 4377
rect 19438 4371 19450 4405
rect 19484 4371 19504 4405
rect 19077 4303 19115 4337
rect 19438 4333 19504 4371
rect 19438 4299 19450 4333
rect 19484 4299 19504 4333
rect 11972 4081 12003 4119
rect 12412 4117 12688 4123
rect 12622 4104 12688 4117
rect 15771 4114 15919 4156
rect 11288 4026 11338 4035
rect 11288 4001 11298 4026
rect 11254 3992 11298 4001
rect 11332 3992 11338 4026
rect 12068 4000 12267 4090
rect 13123 4080 13161 4114
rect 12482 4024 12520 4058
rect 11254 3967 11338 3992
rect 11288 3952 11338 3967
rect 11288 3933 11298 3952
rect 11254 3918 11298 3933
rect 11332 3918 11338 3952
rect 11932 3988 12267 4000
rect 11932 3944 12171 3988
rect 12739 3984 12773 4022
rect 12996 4002 13254 4020
rect 13677 4002 13820 4104
rect 14123 4080 14161 4114
rect 14481 4002 14673 4104
rect 14924 4080 14962 4114
rect 15285 4002 15428 4104
rect 15755 4080 15794 4114
rect 15828 4080 15866 4114
rect 15900 4080 15938 4114
rect 15771 4054 15919 4080
rect 16089 4002 16232 4104
rect 16351 4087 16389 4121
rect 16977 4085 17015 4119
rect 16843 4068 16877 4081
rect 16843 4043 16880 4068
rect 16877 4024 16880 4043
rect 17014 4031 17045 4071
rect 12930 3944 13254 4002
rect 17165 3981 17298 4083
rect 17482 3965 17675 4099
rect 17779 4073 17988 4120
rect 18105 4088 18135 4117
rect 18283 4076 18318 4111
rect 17813 4039 17855 4073
rect 17889 4039 17931 4073
rect 17965 4039 17988 4073
rect 18469 4070 18505 4106
rect 18639 4065 18677 4099
rect 17779 3986 17988 4039
rect 18469 4003 18535 4054
rect 18463 3969 18501 4003
rect 18812 4002 18955 4104
rect 19260 4056 19268 4061
rect 19438 4083 19504 4299
rect 19609 4104 19675 4458
rect 19967 4548 20013 4572
rect 19967 4514 19973 4548
rect 20007 4538 20013 4548
rect 19967 4504 19975 4514
rect 20009 4504 20013 4538
rect 19967 4475 20013 4504
rect 19967 4441 19973 4475
rect 20007 4470 20013 4475
rect 19967 4436 19975 4441
rect 20009 4436 20013 4470
rect 19967 4402 20013 4436
rect 19967 4368 19973 4402
rect 20009 4368 20013 4402
rect 19967 4334 20013 4368
rect 19967 4329 19975 4334
rect 19967 4295 19973 4329
rect 20009 4300 20013 4334
rect 20007 4295 20013 4300
rect 19967 4266 20013 4295
rect 19967 4256 19975 4266
rect 19967 4222 19973 4256
rect 20009 4232 20013 4266
rect 20007 4222 20013 4232
rect 19967 4198 20013 4222
rect 19967 4183 19975 4198
rect 19729 4111 19763 4149
rect 19967 4149 19973 4183
rect 20009 4164 20013 4198
rect 20007 4149 20013 4164
rect 19967 4130 20013 4149
rect 19967 4110 19975 4130
rect 19967 4076 19973 4110
rect 20009 4096 20013 4130
rect 20007 4076 20013 4096
rect 19967 4062 20013 4076
rect 19302 4056 19316 4061
rect 19260 4018 19316 4056
rect 19260 4017 19268 4018
rect 19302 4017 19316 4018
rect 19967 4037 19975 4062
rect 19967 4003 19973 4037
rect 20009 4028 20013 4062
rect 20007 4003 20013 4028
rect 19967 3994 20013 4003
rect 18469 3966 18535 3969
rect 19967 3964 19975 3994
rect 19967 3930 19973 3964
rect 20009 3960 20013 3994
rect 20007 3930 20013 3960
rect 19967 3926 20013 3930
rect 11254 3899 11338 3918
rect 11288 3878 11338 3899
rect 11288 3865 11298 3878
rect 11254 3844 11298 3865
rect 11332 3844 11338 3878
rect 14332 3864 14370 3898
rect 8476 3768 8482 3806
rect 8516 3768 8522 3806
rect 8476 3736 8522 3768
rect 11254 3831 11338 3844
rect 11288 3804 11338 3831
rect 17116 3854 17150 3892
rect 19967 3892 19975 3926
rect 20009 3892 20013 3926
rect 19967 3891 20013 3892
rect 19967 3857 19973 3891
rect 20007 3858 20013 3891
rect 19967 3824 19975 3857
rect 20009 3824 20013 3858
rect 11288 3797 11298 3804
rect 11254 3770 11298 3797
rect 11332 3770 11338 3804
rect 11254 3763 11338 3770
rect 8476 3694 8482 3736
rect 8516 3694 8522 3736
rect 8476 3666 8522 3694
rect 8476 3620 8482 3666
rect 8516 3620 8522 3666
rect 8691 3722 8775 3756
rect 8809 3722 8870 3756
rect 8904 3722 8965 3756
rect 8999 3722 9015 3756
rect 9071 3722 9087 3756
rect 9121 3722 9182 3756
rect 9216 3751 9277 3756
rect 9311 3751 9327 3756
rect 9216 3722 9223 3751
rect 8657 3704 9015 3722
rect 9257 3722 9277 3751
rect 9257 3717 9295 3722
rect 9454 3736 9575 3752
rect 8657 3684 8691 3704
rect 9454 3702 9541 3736
rect 9787 3722 9803 3756
rect 9846 3723 9895 3757
rect 9929 3756 9977 3757
rect 9932 3723 9977 3756
rect 9837 3722 9898 3723
rect 9932 3722 9993 3723
rect 10027 3722 10043 3756
rect 10376 3722 10392 3756
rect 10433 3722 10466 3756
rect 10507 3722 10539 3756
rect 10580 3722 10612 3756
rect 10653 3722 10685 3756
rect 10726 3722 10758 3756
rect 10799 3722 10831 3756
rect 10872 3722 10904 3756
rect 10945 3722 10977 3756
rect 11018 3722 11050 3756
rect 11091 3722 11100 3756
rect 11288 3730 11338 3763
rect 11288 3729 11298 3730
rect 9454 3668 9575 3702
rect 9454 3657 9541 3668
rect 11254 3696 11298 3729
rect 11332 3696 11338 3730
rect 11254 3695 11338 3696
rect 11288 3661 11338 3695
rect 8476 3596 8522 3620
rect 9454 3623 9465 3657
rect 9499 3623 9537 3657
rect 9571 3623 9575 3634
rect 9454 3618 9575 3623
rect 10555 3643 10824 3659
rect 8476 3546 8482 3596
rect 8516 3546 8522 3596
rect 8476 3526 8522 3546
rect 8476 3472 8482 3526
rect 8516 3472 8522 3526
rect 10555 3609 10636 3643
rect 10674 3609 10774 3643
rect 10812 3609 10824 3643
rect 11254 3656 11338 3661
rect 11254 3627 11298 3656
rect 10555 3523 10621 3609
rect 11288 3622 11298 3627
rect 11332 3622 11338 3656
rect 19967 3818 20013 3824
rect 19967 3784 19973 3818
rect 20007 3790 20013 3818
rect 19967 3756 19975 3784
rect 20009 3756 20013 3790
rect 19967 3745 20013 3756
rect 19967 3711 19973 3745
rect 20007 3722 20013 3745
rect 19967 3688 19975 3711
rect 20009 3688 20013 3722
rect 19967 3672 20013 3688
rect 19967 3638 19973 3672
rect 20007 3654 20013 3672
rect 11288 3593 11338 3622
rect 11552 3598 11576 3632
rect 11610 3598 11645 3632
rect 11679 3598 11714 3632
rect 11748 3598 11783 3632
rect 11817 3598 11852 3632
rect 11886 3598 11921 3632
rect 11955 3598 11990 3632
rect 12024 3598 12059 3632
rect 12093 3598 12128 3632
rect 12162 3598 12197 3632
rect 12231 3598 12266 3632
rect 12300 3598 12335 3632
rect 12369 3598 12404 3632
rect 12438 3598 12473 3632
rect 12507 3598 12542 3632
rect 12576 3598 12611 3632
rect 12645 3598 12680 3632
rect 12714 3598 12749 3632
rect 12783 3598 12818 3632
rect 12852 3598 12887 3632
rect 12921 3598 12956 3632
rect 12990 3598 13025 3632
rect 13059 3598 13094 3632
rect 13128 3598 13163 3632
rect 13197 3598 13232 3632
rect 13266 3598 13301 3632
rect 13335 3598 13370 3632
rect 13404 3598 13439 3632
rect 13473 3598 13508 3632
rect 13542 3598 13577 3632
rect 13611 3598 13646 3632
rect 13680 3598 13715 3632
rect 13749 3598 13784 3632
rect 13818 3598 13853 3632
rect 13887 3598 13922 3632
rect 13956 3598 13991 3632
rect 14025 3598 14059 3632
rect 14093 3598 14127 3632
rect 14161 3598 14195 3632
rect 14229 3598 14263 3632
rect 14297 3598 14331 3632
rect 14365 3598 14399 3632
rect 14433 3598 14467 3632
rect 14501 3598 14535 3632
rect 14569 3598 14603 3632
rect 14637 3598 14671 3632
rect 14705 3598 14739 3632
rect 14773 3598 14807 3632
rect 14841 3598 14875 3632
rect 14909 3598 14943 3632
rect 14977 3598 15011 3632
rect 15045 3598 15079 3632
rect 15113 3598 15147 3632
rect 15181 3598 15215 3632
rect 15249 3598 15283 3632
rect 15317 3598 15351 3632
rect 15385 3598 15419 3632
rect 15453 3598 15487 3632
rect 15521 3598 15555 3632
rect 15589 3598 15623 3632
rect 15657 3598 15691 3632
rect 15725 3598 15759 3632
rect 15793 3598 15827 3632
rect 15861 3598 15895 3632
rect 15929 3598 15963 3632
rect 15997 3598 16031 3632
rect 16065 3598 16099 3632
rect 16133 3598 16167 3632
rect 16201 3598 16235 3632
rect 16269 3598 16303 3632
rect 16337 3598 16371 3632
rect 16405 3598 16439 3632
rect 16473 3598 16507 3632
rect 16541 3598 16575 3632
rect 16609 3598 16643 3632
rect 16677 3598 16711 3632
rect 16745 3598 16779 3632
rect 16813 3598 16847 3632
rect 16881 3598 16915 3632
rect 16949 3598 16983 3632
rect 17017 3598 17051 3632
rect 17085 3598 17119 3632
rect 17153 3598 17187 3632
rect 17221 3598 17255 3632
rect 17289 3598 17323 3632
rect 17357 3598 17391 3632
rect 17425 3598 17459 3632
rect 17493 3598 17527 3632
rect 17561 3598 17595 3632
rect 17629 3598 17663 3632
rect 17697 3598 17731 3632
rect 17765 3598 17799 3632
rect 17833 3598 17867 3632
rect 17901 3598 17935 3632
rect 17969 3598 18003 3632
rect 18037 3598 18071 3632
rect 18105 3598 18139 3632
rect 18173 3598 18207 3632
rect 18241 3598 18275 3632
rect 18309 3598 18343 3632
rect 18377 3598 18411 3632
rect 18445 3598 18479 3632
rect 18513 3598 18547 3632
rect 18581 3598 18615 3632
rect 18649 3598 18683 3632
rect 18717 3598 18751 3632
rect 18785 3598 18819 3632
rect 18853 3598 18887 3632
rect 18921 3598 18955 3632
rect 18989 3598 19023 3632
rect 19057 3598 19091 3632
rect 19125 3598 19159 3632
rect 19193 3598 19227 3632
rect 19261 3598 19295 3632
rect 19329 3598 19363 3632
rect 19397 3598 19431 3632
rect 19465 3598 19499 3632
rect 19533 3598 19567 3632
rect 19601 3598 19635 3632
rect 19669 3598 19703 3632
rect 19737 3598 19761 3632
rect 19967 3620 19975 3638
rect 20009 3620 20013 3654
rect 19967 3599 20013 3620
rect 11254 3582 11338 3593
rect 8939 3475 8961 3509
rect 9007 3475 9033 3509
rect 9075 3475 9105 3509
rect 9143 3475 9177 3509
rect 9211 3475 9245 3509
rect 9283 3475 9313 3509
rect 9355 3475 9381 3509
rect 9427 3475 9449 3509
rect 9499 3475 9517 3509
rect 9571 3475 9585 3509
rect 9643 3475 9653 3509
rect 9715 3475 9721 3509
rect 9787 3475 9789 3509
rect 9823 3475 9825 3509
rect 10555 3489 10579 3523
rect 10613 3489 10621 3523
rect 10555 3473 10621 3489
rect 10835 3532 10891 3566
rect 10925 3532 10963 3566
rect 11254 3559 11298 3582
rect 10835 3523 10937 3532
rect 10869 3489 10937 3523
rect 10835 3473 10937 3489
rect 11288 3548 11298 3559
rect 11332 3548 11338 3582
rect 11288 3525 11338 3548
rect 11254 3504 11338 3525
rect 11254 3491 11298 3504
rect 8476 3456 8522 3472
rect 8476 3398 8482 3456
rect 8516 3398 8522 3456
rect 8476 3386 8522 3398
rect 8476 3324 8482 3386
rect 8516 3324 8522 3386
rect 9941 3455 9975 3464
rect 9941 3355 9975 3414
rect 11288 3470 11298 3491
rect 11332 3470 11338 3504
rect 11288 3457 11338 3470
rect 11254 3393 11338 3457
rect 8476 3316 8522 3324
rect 8939 3319 8961 3353
rect 9007 3319 9033 3353
rect 9075 3319 9105 3353
rect 9143 3319 9177 3353
rect 9211 3319 9245 3353
rect 9283 3319 9313 3353
rect 9355 3319 9381 3353
rect 9427 3319 9449 3353
rect 9499 3319 9517 3353
rect 9571 3319 9585 3353
rect 9643 3319 9653 3353
rect 9715 3319 9721 3353
rect 9787 3319 9789 3353
rect 9823 3319 9825 3353
rect 8476 3250 8482 3316
rect 8516 3250 8522 3316
rect 8476 3246 8522 3250
rect 8476 3212 8482 3246
rect 8516 3212 8522 3246
rect 8476 3210 8522 3212
rect 8476 3142 8482 3210
rect 8516 3142 8522 3210
rect 9941 3258 9975 3319
rect 9941 3208 9975 3220
rect 10070 3337 10104 3351
rect 10220 3336 10222 3370
rect 10256 3336 10258 3370
rect 10324 3336 10330 3370
rect 10392 3336 10402 3370
rect 10460 3336 10474 3370
rect 10528 3336 10546 3370
rect 10596 3336 10618 3370
rect 10664 3336 10690 3370
rect 10732 3336 10762 3370
rect 10800 3336 10834 3370
rect 10868 3336 10902 3370
rect 10940 3336 10970 3370
rect 11012 3336 11038 3370
rect 11084 3336 11106 3370
rect 11254 3359 11298 3393
rect 11332 3382 11338 3393
rect 19967 3565 19973 3599
rect 20007 3586 20013 3599
rect 19967 3552 19975 3565
rect 20009 3552 20013 3586
rect 19967 3526 20013 3552
rect 19967 3492 19973 3526
rect 20007 3518 20013 3526
rect 19967 3484 19975 3492
rect 20009 3484 20013 3518
rect 19967 3454 20013 3484
rect 19967 3420 19973 3454
rect 20007 3450 20013 3454
rect 19967 3416 19975 3420
rect 20009 3416 20013 3450
rect 19967 3382 20013 3416
rect 11254 3348 11322 3359
rect 11356 3348 11390 3382
rect 11424 3348 11458 3382
rect 11492 3348 11526 3382
rect 11560 3377 11594 3382
rect 11628 3377 11662 3382
rect 11696 3377 11730 3382
rect 11764 3377 11798 3382
rect 11832 3377 11866 3382
rect 11900 3377 11934 3382
rect 11560 3348 11565 3377
rect 11628 3348 11638 3377
rect 11696 3348 11711 3377
rect 11764 3348 11784 3377
rect 11832 3348 11857 3377
rect 11900 3348 11930 3377
rect 11968 3348 12002 3382
rect 12036 3377 12070 3382
rect 12104 3377 12138 3382
rect 12172 3377 12206 3382
rect 12240 3377 12274 3382
rect 12308 3377 12342 3382
rect 12376 3377 12410 3382
rect 12444 3377 12478 3382
rect 12037 3348 12070 3377
rect 12110 3348 12138 3377
rect 12183 3348 12206 3377
rect 12256 3348 12274 3377
rect 12329 3348 12342 3377
rect 12402 3348 12410 3377
rect 12475 3348 12478 3377
rect 12512 3377 12546 3382
rect 12580 3377 12614 3382
rect 12648 3377 12682 3382
rect 12716 3377 12750 3382
rect 12784 3377 12818 3382
rect 12852 3377 12886 3382
rect 12920 3377 12954 3382
rect 12512 3348 12514 3377
rect 12580 3348 12587 3377
rect 12648 3348 12660 3377
rect 12716 3348 12733 3377
rect 12784 3348 12806 3377
rect 12852 3348 12879 3377
rect 12920 3348 12952 3377
rect 12988 3348 13022 3382
rect 13056 3377 13090 3382
rect 13124 3377 13158 3382
rect 13192 3377 13226 3382
rect 13260 3377 13294 3382
rect 13328 3377 13362 3382
rect 13396 3377 13430 3382
rect 13464 3377 13498 3382
rect 13059 3348 13090 3377
rect 13132 3348 13158 3377
rect 13205 3348 13226 3377
rect 13278 3348 13294 3377
rect 13351 3348 13362 3377
rect 13424 3348 13430 3377
rect 13497 3348 13498 3377
rect 13532 3377 13566 3382
rect 13600 3377 13634 3382
rect 13668 3377 13702 3382
rect 13736 3377 13770 3382
rect 13804 3377 13838 3382
rect 13872 3377 13906 3382
rect 13532 3348 13536 3377
rect 13600 3348 13609 3377
rect 13668 3348 13682 3377
rect 13736 3348 13755 3377
rect 13804 3348 13828 3377
rect 13872 3348 13901 3377
rect 13940 3348 13974 3382
rect 14008 3348 14042 3382
rect 14076 3377 14110 3382
rect 14144 3377 14178 3382
rect 14212 3377 14246 3382
rect 14280 3377 14314 3382
rect 14348 3377 14382 3382
rect 14416 3377 14450 3382
rect 14081 3348 14110 3377
rect 14154 3348 14178 3377
rect 14227 3348 14246 3377
rect 14300 3348 14314 3377
rect 14373 3348 14382 3377
rect 14446 3348 14450 3377
rect 14484 3377 14518 3382
rect 14552 3377 14586 3382
rect 14620 3377 14654 3382
rect 14688 3377 14722 3382
rect 14756 3377 14790 3382
rect 14824 3377 14858 3382
rect 14892 3377 14926 3382
rect 14960 3377 14994 3382
rect 14484 3348 14485 3377
rect 14552 3348 14558 3377
rect 14620 3348 14631 3377
rect 14688 3348 14704 3377
rect 14756 3348 14777 3377
rect 14824 3348 14849 3377
rect 14892 3348 14921 3377
rect 14960 3348 14993 3377
rect 15028 3348 15062 3382
rect 15096 3377 15130 3382
rect 15164 3377 15198 3382
rect 15232 3377 15266 3382
rect 15300 3377 15334 3382
rect 15368 3377 15402 3382
rect 15436 3377 15470 3382
rect 15504 3377 15538 3382
rect 15572 3377 15606 3382
rect 15099 3348 15130 3377
rect 15171 3348 15198 3377
rect 15243 3348 15266 3377
rect 15315 3348 15334 3377
rect 15387 3348 15402 3377
rect 15459 3348 15470 3377
rect 15531 3348 15538 3377
rect 15603 3348 15606 3377
rect 15640 3377 15674 3382
rect 15708 3377 15742 3382
rect 15776 3377 15810 3382
rect 15844 3377 15878 3382
rect 15912 3377 15946 3382
rect 15980 3377 16014 3382
rect 16048 3377 16082 3382
rect 16116 3377 16150 3382
rect 16184 3377 16218 3382
rect 15640 3348 15641 3377
rect 15708 3348 15713 3377
rect 15776 3348 15785 3377
rect 15844 3348 15857 3377
rect 15912 3348 15929 3377
rect 15980 3348 16001 3377
rect 16048 3348 16073 3377
rect 16116 3348 16145 3377
rect 16184 3348 16217 3377
rect 16252 3348 16286 3382
rect 16320 3377 16354 3382
rect 16388 3377 16422 3382
rect 16456 3377 16490 3382
rect 16524 3377 16558 3382
rect 16592 3377 16626 3382
rect 16660 3377 16694 3382
rect 16728 3377 16762 3382
rect 16796 3377 16830 3382
rect 16323 3348 16354 3377
rect 16395 3348 16422 3377
rect 16467 3348 16490 3377
rect 16539 3348 16558 3377
rect 16611 3348 16626 3377
rect 16683 3348 16694 3377
rect 16755 3348 16762 3377
rect 16827 3348 16830 3377
rect 16864 3377 16898 3382
rect 16932 3377 16966 3382
rect 17000 3377 17034 3382
rect 17068 3377 17102 3382
rect 17136 3377 17170 3382
rect 17204 3377 17238 3382
rect 17272 3377 17306 3382
rect 17340 3377 17374 3382
rect 17408 3377 17442 3382
rect 16864 3348 16865 3377
rect 16932 3348 16937 3377
rect 17000 3348 17009 3377
rect 17068 3348 17081 3377
rect 17136 3348 17153 3377
rect 17204 3348 17225 3377
rect 17272 3348 17297 3377
rect 17340 3348 17369 3377
rect 17408 3348 17441 3377
rect 17476 3348 17510 3382
rect 17544 3377 17578 3382
rect 17612 3377 17646 3382
rect 17680 3377 17714 3382
rect 17748 3377 17782 3382
rect 17816 3377 17850 3382
rect 17884 3377 17918 3382
rect 17952 3377 17986 3382
rect 18020 3377 18054 3382
rect 17547 3348 17578 3377
rect 17619 3348 17646 3377
rect 17691 3348 17714 3377
rect 17763 3348 17782 3377
rect 17835 3348 17850 3377
rect 17907 3348 17918 3377
rect 17979 3348 17986 3377
rect 18051 3348 18054 3377
rect 18088 3377 18122 3382
rect 18156 3377 18190 3382
rect 18224 3377 18258 3382
rect 18292 3377 18326 3382
rect 18360 3377 18394 3382
rect 18428 3377 18462 3382
rect 18496 3377 18530 3382
rect 18564 3377 18598 3382
rect 18632 3377 18666 3382
rect 18088 3348 18089 3377
rect 18156 3348 18161 3377
rect 18224 3348 18233 3377
rect 18292 3348 18305 3377
rect 18360 3348 18377 3377
rect 18428 3348 18449 3377
rect 18496 3348 18521 3377
rect 18564 3348 18593 3377
rect 18632 3348 18665 3377
rect 18700 3348 18734 3382
rect 18768 3377 18802 3382
rect 18836 3377 18870 3382
rect 18904 3377 18938 3382
rect 18972 3377 19006 3382
rect 19040 3377 19074 3382
rect 19108 3377 19142 3382
rect 19176 3377 19210 3382
rect 19244 3377 19278 3382
rect 18771 3348 18802 3377
rect 18843 3348 18870 3377
rect 18915 3348 18938 3377
rect 18987 3348 19006 3377
rect 19059 3348 19074 3377
rect 19131 3348 19142 3377
rect 19203 3348 19210 3377
rect 19275 3348 19278 3377
rect 19312 3377 19346 3382
rect 19380 3377 19414 3382
rect 19448 3377 19482 3382
rect 19516 3377 19550 3382
rect 19584 3377 19618 3382
rect 19652 3377 19686 3382
rect 19720 3377 19754 3382
rect 19788 3377 19822 3382
rect 19856 3377 19890 3382
rect 19312 3348 19313 3377
rect 19380 3348 19385 3377
rect 19448 3348 19457 3377
rect 19516 3348 19529 3377
rect 19584 3348 19601 3377
rect 19652 3348 19673 3377
rect 19720 3348 19745 3377
rect 19788 3348 19817 3377
rect 19856 3348 19889 3377
rect 19924 3348 20013 3382
rect 10070 3267 10104 3301
rect 10070 3217 10104 3231
rect 11254 3315 11338 3348
rect 11599 3343 11638 3348
rect 11672 3343 11711 3348
rect 11745 3343 11784 3348
rect 11818 3343 11857 3348
rect 11891 3343 11930 3348
rect 11964 3343 12003 3348
rect 12037 3343 12076 3348
rect 12110 3343 12149 3348
rect 12183 3343 12222 3348
rect 12256 3343 12295 3348
rect 12329 3343 12368 3348
rect 12402 3343 12441 3348
rect 12475 3343 12514 3348
rect 12548 3343 12587 3348
rect 12621 3343 12660 3348
rect 12694 3343 12733 3348
rect 12767 3343 12806 3348
rect 12840 3343 12879 3348
rect 12913 3343 12952 3348
rect 12986 3343 13025 3348
rect 13059 3343 13098 3348
rect 13132 3343 13171 3348
rect 13205 3343 13244 3348
rect 13278 3343 13317 3348
rect 13351 3343 13390 3348
rect 13424 3343 13463 3348
rect 13497 3343 13536 3348
rect 13570 3343 13609 3348
rect 13643 3343 13682 3348
rect 13716 3343 13755 3348
rect 13789 3343 13828 3348
rect 13862 3343 13901 3348
rect 13935 3343 13974 3348
rect 14008 3343 14047 3348
rect 14081 3343 14120 3348
rect 14154 3343 14193 3348
rect 14227 3343 14266 3348
rect 14300 3343 14339 3348
rect 14373 3343 14412 3348
rect 14446 3343 14485 3348
rect 14519 3343 14558 3348
rect 14592 3343 14631 3348
rect 14665 3343 14704 3348
rect 14738 3343 14777 3348
rect 14811 3343 14849 3348
rect 14883 3343 14921 3348
rect 14955 3343 14993 3348
rect 15027 3343 15065 3348
rect 15099 3343 15137 3348
rect 15171 3343 15209 3348
rect 15243 3343 15281 3348
rect 15315 3343 15353 3348
rect 15387 3343 15425 3348
rect 15459 3343 15497 3348
rect 15531 3343 15569 3348
rect 15603 3343 15641 3348
rect 15675 3343 15713 3348
rect 15747 3343 15785 3348
rect 15819 3343 15857 3348
rect 15891 3343 15929 3348
rect 15963 3343 16001 3348
rect 16035 3343 16073 3348
rect 16107 3343 16145 3348
rect 16179 3343 16217 3348
rect 16251 3343 16289 3348
rect 16323 3343 16361 3348
rect 16395 3343 16433 3348
rect 16467 3343 16505 3348
rect 16539 3343 16577 3348
rect 16611 3343 16649 3348
rect 16683 3343 16721 3348
rect 16755 3343 16793 3348
rect 16827 3343 16865 3348
rect 16899 3343 16937 3348
rect 16971 3343 17009 3348
rect 17043 3343 17081 3348
rect 17115 3343 17153 3348
rect 17187 3343 17225 3348
rect 17259 3343 17297 3348
rect 17331 3343 17369 3348
rect 17403 3343 17441 3348
rect 17475 3343 17513 3348
rect 17547 3343 17585 3348
rect 17619 3343 17657 3348
rect 17691 3343 17729 3348
rect 17763 3343 17801 3348
rect 17835 3343 17873 3348
rect 17907 3343 17945 3348
rect 17979 3343 18017 3348
rect 18051 3343 18089 3348
rect 18123 3343 18161 3348
rect 18195 3343 18233 3348
rect 18267 3343 18305 3348
rect 18339 3343 18377 3348
rect 18411 3343 18449 3348
rect 18483 3343 18521 3348
rect 18555 3343 18593 3348
rect 18627 3343 18665 3348
rect 18699 3343 18737 3348
rect 18771 3343 18809 3348
rect 18843 3343 18881 3348
rect 18915 3343 18953 3348
rect 18987 3343 19025 3348
rect 19059 3343 19097 3348
rect 19131 3343 19169 3348
rect 19203 3343 19241 3348
rect 19275 3343 19313 3348
rect 19347 3343 19385 3348
rect 19419 3343 19457 3348
rect 19491 3343 19529 3348
rect 19563 3343 19601 3348
rect 19635 3343 19673 3348
rect 19707 3343 19745 3348
rect 19779 3343 19817 3348
rect 19851 3343 19889 3348
rect 11254 3314 11298 3315
rect 11254 3280 11261 3314
rect 11295 3281 11298 3314
rect 11332 3281 11338 3315
rect 11295 3280 11338 3281
rect 11254 3237 11338 3280
rect 18900 3305 18934 3343
rect 19923 3342 20013 3348
rect 11254 3231 11298 3237
rect 8939 3163 8961 3197
rect 9007 3163 9033 3197
rect 9075 3163 9105 3197
rect 9143 3163 9177 3197
rect 9211 3163 9245 3197
rect 9283 3163 9313 3197
rect 9355 3163 9381 3197
rect 9427 3163 9449 3197
rect 9499 3163 9517 3197
rect 9571 3163 9585 3197
rect 9643 3163 9653 3197
rect 9715 3163 9721 3197
rect 9787 3163 9789 3197
rect 9823 3163 9825 3197
rect 10220 3180 10222 3214
rect 10256 3180 10258 3214
rect 10324 3180 10330 3214
rect 10392 3180 10402 3214
rect 10460 3180 10474 3214
rect 10528 3180 10546 3214
rect 10596 3180 10618 3214
rect 10664 3180 10690 3214
rect 10732 3180 10762 3214
rect 10800 3180 10834 3214
rect 10868 3180 10902 3214
rect 10940 3180 10970 3214
rect 11012 3180 11038 3214
rect 11084 3180 11106 3214
rect 11254 3197 11261 3231
rect 11295 3203 11298 3231
rect 11332 3203 11338 3237
rect 11295 3197 11338 3203
rect 8476 3136 8522 3142
rect 3418 3077 3456 3094
rect 3490 3077 3528 3094
rect 3562 3077 3600 3094
rect 3634 3077 3672 3094
rect 3706 3077 3744 3094
rect 3778 3077 3850 3094
rect 8476 3072 8482 3136
rect 8516 3072 8522 3136
rect 11254 3159 11338 3197
rect 17033 3195 17049 3229
rect 17083 3216 17117 3229
rect 17083 3195 17104 3216
rect 17151 3195 17185 3229
rect 17219 3216 17253 3229
rect 17287 3216 17321 3229
rect 17223 3195 17253 3216
rect 17307 3195 17321 3216
rect 17355 3216 17389 3229
rect 17423 3216 17457 3229
rect 17355 3195 17357 3216
rect 17423 3195 17441 3216
rect 17491 3195 17525 3229
rect 17559 3195 17575 3229
rect 17798 3216 17832 3232
rect 17138 3182 17189 3195
rect 17223 3182 17273 3195
rect 17307 3182 17357 3195
rect 17391 3182 17441 3195
rect 17475 3182 17525 3195
rect 11254 3148 11298 3159
rect 11254 3114 11261 3148
rect 11295 3125 11298 3148
rect 11332 3125 11338 3159
rect 11295 3114 11338 3125
rect 11254 3094 11338 3114
rect 10295 3093 11338 3094
rect 8476 3062 8522 3072
rect 8476 3002 8482 3062
rect 8516 3002 8522 3062
rect 10284 3087 11338 3093
rect 10284 3053 10362 3087
rect 10396 3053 10401 3087
rect 10468 3053 10474 3087
rect 10540 3053 10547 3087
rect 10612 3053 10620 3087
rect 10684 3053 10692 3087
rect 10756 3053 10764 3087
rect 10828 3053 10836 3087
rect 10900 3053 10908 3087
rect 10972 3053 10980 3087
rect 11044 3053 11052 3087
rect 11116 3053 11124 3087
rect 11188 3053 11196 3087
rect 11260 3053 11338 3087
rect 17619 3130 17653 3134
rect 10284 3046 11338 3053
rect 10284 3002 10337 3046
rect 17033 3019 17049 3053
rect 17083 3019 17117 3053
rect 17151 3019 17185 3053
rect 17219 3047 17253 3053
rect 17241 3019 17253 3047
rect 17287 3047 17321 3053
rect 17355 3047 17389 3053
rect 17287 3019 17291 3047
rect 17355 3019 17374 3047
rect 17423 3019 17457 3053
rect 17491 3019 17525 3053
rect 17559 3019 17575 3053
rect 17619 3050 17653 3066
rect 17798 3178 17832 3182
rect 17798 3106 17832 3114
rect 17798 3030 17832 3046
rect 17954 3216 17988 3241
rect 18900 3233 18934 3271
rect 19967 3294 20013 3342
rect 19967 3248 20042 3294
rect 17954 3148 17988 3169
rect 17954 3080 17988 3114
rect 17954 3030 17988 3046
rect 18110 3216 18144 3232
rect 18110 3148 18144 3182
rect 18110 3080 18144 3114
rect 18110 3030 18144 3042
rect 18282 3216 18316 3232
rect 18282 3148 18316 3182
rect 18282 3080 18316 3114
rect 18282 3030 18316 3042
rect 18438 3216 18472 3232
rect 18438 3148 18472 3174
rect 18438 3080 18472 3102
rect 18594 3216 18628 3232
rect 18594 3148 18628 3182
rect 18594 3080 18628 3114
rect 18594 3030 18628 3042
rect 18744 3216 18778 3232
rect 18744 3148 18778 3182
rect 18744 3080 18778 3114
rect 18744 3030 18778 3042
rect 18900 3148 18934 3182
rect 18900 3080 18934 3114
rect 18900 3030 18934 3046
rect 19056 3216 19090 3232
rect 19056 3148 19090 3182
rect 19056 3080 19090 3114
rect 19056 3030 19090 3042
rect 19996 3216 20042 3248
rect 19996 3182 20002 3216
rect 20036 3182 20042 3216
rect 19996 3143 20042 3182
rect 19996 3109 20002 3143
rect 20036 3109 20042 3143
rect 19996 3070 20042 3109
rect 19996 3036 20002 3070
rect 20036 3036 20042 3070
rect 17241 3013 17291 3019
rect 17325 3013 17374 3019
rect 17408 3013 17457 3019
rect 8476 2988 8550 3002
rect 8476 2954 8482 2988
rect 8516 2968 8550 2988
rect 8584 2968 8619 3002
rect 8653 2968 8688 3002
rect 8722 2968 8757 3002
rect 8791 2968 8826 3002
rect 8860 2968 8867 3002
rect 8929 2968 8942 3002
rect 8998 2968 9017 3002
rect 9067 2968 9092 3002
rect 9136 2968 9167 3002
rect 9205 2968 9240 3002
rect 9276 2968 9309 3002
rect 9351 2968 9378 3002
rect 9426 2968 9447 3002
rect 9501 2968 9516 3002
rect 9576 2968 9585 3002
rect 9651 2968 9654 3002
rect 9688 2968 9692 3002
rect 9757 2968 9767 3002
rect 9826 2968 9842 3002
rect 9895 2968 9917 3002
rect 9963 2968 9992 3002
rect 10031 2968 10065 3002
rect 10101 2968 10133 3002
rect 10176 2968 10201 3002
rect 10251 2968 10269 3002
rect 10325 2968 10337 3002
rect 19996 2998 20042 3036
rect 8516 2954 8522 2968
rect 8476 2914 8522 2954
rect 17889 2942 17954 2976
rect 17988 2942 18053 2976
rect 18373 2942 18438 2976
rect 18472 2942 18537 2976
rect 18835 2942 18900 2976
rect 18934 2942 18999 2976
rect 19996 2964 20002 2998
rect 20036 2964 20042 2998
rect 8476 2880 8482 2914
rect 8516 2880 8522 2914
rect 19996 2926 20042 2964
rect 19996 2892 20002 2926
rect 20036 2892 20042 2926
rect 8476 2840 8522 2880
rect 8476 2806 8482 2840
rect 8516 2806 8522 2840
rect 10522 2855 10568 2856
rect 10602 2855 10647 2856
rect 10681 2855 10726 2856
rect 10760 2855 10805 2856
rect 10839 2855 10884 2856
rect 10918 2855 10963 2856
rect 10997 2855 11042 2856
rect 11076 2855 11121 2856
rect 11155 2855 11200 2856
rect 11234 2855 11279 2856
rect 10522 2822 10562 2855
rect 10602 2822 10630 2855
rect 10681 2822 10698 2855
rect 10760 2822 10766 2855
rect 10488 2821 10562 2822
rect 10596 2821 10630 2822
rect 10664 2821 10698 2822
rect 10732 2821 10766 2822
rect 10800 2822 10805 2855
rect 10868 2822 10884 2855
rect 10936 2822 10963 2855
rect 10800 2821 10834 2822
rect 10868 2821 10902 2822
rect 10936 2821 10970 2822
rect 11004 2821 11038 2855
rect 11076 2822 11106 2855
rect 11155 2822 11174 2855
rect 11234 2822 11242 2855
rect 11072 2821 11106 2822
rect 11140 2821 11174 2822
rect 11208 2821 11242 2822
rect 11276 2822 11279 2855
rect 11276 2821 11310 2822
rect 11344 2821 11378 2855
rect 11412 2821 11446 2855
rect 11480 2821 11514 2855
rect 11548 2821 11582 2855
rect 11616 2821 11650 2855
rect 11684 2821 11718 2855
rect 11752 2821 11786 2855
rect 11820 2821 11854 2855
rect 11888 2821 11922 2855
rect 11956 2821 11990 2855
rect 12024 2821 12058 2855
rect 12092 2821 12126 2855
rect 12160 2821 12194 2855
rect 12228 2849 12262 2855
rect 12296 2849 12330 2855
rect 12364 2849 12398 2855
rect 12228 2821 12253 2849
rect 12296 2821 12325 2849
rect 12364 2821 12397 2849
rect 12432 2821 12466 2855
rect 12500 2849 12534 2855
rect 12568 2849 12602 2855
rect 12636 2849 12670 2855
rect 12704 2849 12738 2855
rect 12772 2849 12806 2855
rect 12840 2849 12874 2855
rect 12908 2849 12942 2855
rect 12503 2821 12534 2849
rect 12576 2821 12602 2849
rect 12649 2821 12670 2849
rect 12722 2821 12738 2849
rect 12795 2821 12806 2849
rect 12868 2821 12874 2849
rect 12941 2821 12942 2849
rect 12976 2849 13010 2855
rect 13044 2849 13078 2855
rect 13112 2849 13146 2855
rect 13180 2849 13214 2855
rect 13248 2849 13282 2855
rect 13316 2849 13350 2855
rect 12976 2821 12980 2849
rect 13044 2821 13053 2849
rect 13112 2821 13126 2849
rect 13180 2821 13199 2849
rect 13248 2821 13272 2849
rect 13316 2821 13345 2849
rect 13384 2821 13418 2855
rect 13452 2821 13486 2855
rect 13520 2849 13554 2855
rect 13588 2849 13622 2855
rect 13656 2849 13690 2855
rect 13724 2849 13758 2855
rect 13792 2849 13826 2855
rect 13860 2849 13894 2855
rect 13525 2821 13554 2849
rect 13598 2821 13622 2849
rect 13671 2821 13690 2849
rect 13744 2821 13758 2849
rect 13817 2821 13826 2849
rect 13890 2821 13894 2849
rect 13928 2849 13962 2855
rect 13996 2849 14030 2855
rect 14064 2849 14098 2855
rect 14132 2849 14166 2855
rect 14200 2849 14234 2855
rect 14268 2849 14302 2855
rect 14336 2849 14370 2855
rect 13928 2821 13929 2849
rect 13996 2821 14002 2849
rect 14064 2821 14075 2849
rect 14132 2821 14148 2849
rect 14200 2821 14221 2849
rect 14268 2821 14294 2849
rect 14336 2821 14367 2849
rect 14404 2821 14438 2855
rect 14472 2849 14506 2855
rect 14540 2849 14574 2855
rect 14608 2849 14642 2855
rect 14676 2849 14710 2855
rect 14744 2849 14778 2855
rect 14812 2849 14846 2855
rect 14880 2849 14914 2855
rect 14474 2821 14506 2849
rect 14547 2821 14574 2849
rect 14620 2821 14642 2849
rect 14693 2821 14710 2849
rect 14766 2821 14778 2849
rect 14839 2821 14846 2849
rect 14912 2821 14914 2849
rect 14948 2849 14982 2855
rect 15016 2849 15050 2855
rect 15084 2849 15118 2855
rect 15152 2849 15186 2855
rect 15220 2849 15254 2855
rect 15288 2849 15322 2855
rect 15356 2849 15390 2855
rect 14948 2821 14951 2849
rect 15016 2821 15024 2849
rect 15084 2821 15097 2849
rect 15152 2821 15170 2849
rect 15220 2821 15243 2849
rect 15288 2821 15316 2849
rect 15356 2821 15389 2849
rect 15424 2821 15458 2855
rect 15492 2849 15526 2855
rect 15560 2849 15594 2855
rect 15628 2849 15662 2855
rect 15696 2849 15730 2855
rect 15764 2849 15798 2855
rect 15832 2849 15866 2855
rect 15496 2821 15526 2849
rect 15569 2821 15594 2849
rect 15642 2821 15662 2849
rect 15715 2821 15730 2849
rect 15788 2821 15798 2849
rect 15861 2821 15866 2849
rect 15900 2849 15934 2855
rect 8476 2766 8522 2806
rect 8476 2732 8482 2766
rect 8516 2732 8522 2766
rect 8476 2691 8522 2732
rect 8476 2657 8482 2691
rect 8516 2657 8522 2691
rect 8476 2616 8522 2657
rect 8476 2582 8482 2616
rect 8516 2582 8522 2616
rect 574 2518 582 2552
rect 632 2518 660 2552
rect 702 2518 738 2552
rect 772 2518 808 2552
rect 849 2518 878 2552
rect 926 2518 948 2552
rect 1003 2518 1019 2552
rect 1080 2518 1090 2552
rect 1157 2518 1161 2552
rect 1195 2518 1200 2552
rect 1266 2518 1277 2552
rect 1337 2518 1354 2552
rect 1408 2518 1431 2552
rect 1479 2518 1508 2552
rect 1550 2518 1574 2552
rect 8476 2544 8522 2582
rect 9716 2778 10412 2812
rect 9716 2744 9723 2778
rect 9757 2744 9795 2778
rect 9829 2744 9867 2778
rect 9901 2744 9939 2778
rect 9973 2744 10011 2778
rect 10045 2744 10083 2778
rect 10117 2744 10155 2778
rect 10189 2744 10227 2778
rect 10261 2744 10299 2778
rect 10333 2744 10371 2778
rect 10405 2744 10412 2778
rect 9716 2705 10412 2744
rect 9716 2671 9723 2705
rect 9757 2671 9795 2705
rect 9829 2671 9867 2705
rect 9901 2671 9939 2705
rect 9973 2671 10011 2705
rect 10045 2671 10083 2705
rect 10117 2671 10155 2705
rect 10189 2671 10227 2705
rect 10261 2671 10299 2705
rect 10333 2671 10371 2705
rect 10405 2671 10412 2705
rect 9716 2632 10412 2671
rect 9716 2598 9723 2632
rect 9757 2598 9795 2632
rect 9829 2598 9867 2632
rect 9901 2598 9939 2632
rect 9973 2598 10011 2632
rect 10045 2598 10083 2632
rect 10117 2598 10155 2632
rect 10189 2598 10227 2632
rect 10261 2598 10299 2632
rect 10333 2598 10371 2632
rect 10405 2598 10412 2632
rect 9716 2558 10412 2598
rect 9716 2524 9723 2558
rect 9757 2524 9795 2558
rect 9829 2524 9867 2558
rect 9901 2524 9939 2558
rect 9973 2524 10011 2558
rect 10045 2524 10083 2558
rect 10117 2524 10155 2558
rect 10189 2524 10227 2558
rect 10261 2524 10299 2558
rect 10333 2524 10371 2558
rect 10405 2524 10412 2558
rect 2207 2499 8472 2505
rect 2151 2465 2245 2499
rect 2305 2465 2323 2499
rect 2373 2465 2400 2499
rect 2441 2465 2475 2499
rect 2509 2465 2510 2499
rect 2577 2465 2583 2499
rect 2645 2465 2656 2499
rect 2713 2465 2729 2499
rect 2781 2465 2802 2499
rect 2849 2465 2875 2499
rect 2917 2465 2948 2499
rect 2985 2465 3019 2499
rect 3055 2465 3087 2499
rect 3128 2465 3155 2499
rect 3201 2465 3223 2499
rect 3274 2465 3291 2499
rect 3347 2465 3359 2499
rect 3420 2465 3427 2499
rect 3493 2465 3495 2499
rect 3529 2465 3532 2499
rect 3597 2465 3605 2499
rect 3665 2465 3678 2499
rect 3733 2465 3751 2499
rect 3801 2465 3824 2499
rect 3869 2465 3897 2499
rect 3937 2465 3970 2499
rect 4005 2465 4039 2499
rect 4077 2465 4107 2499
rect 4150 2465 4175 2499
rect 4223 2465 4243 2499
rect 4296 2465 4311 2499
rect 4369 2465 4379 2499
rect 4442 2465 4447 2499
rect 4549 2465 4554 2499
rect 4617 2465 4627 2499
rect 4685 2465 4700 2499
rect 4753 2465 4773 2499
rect 4821 2465 4846 2499
rect 4889 2465 4919 2499
rect 4957 2465 4991 2499
rect 5026 2465 5059 2499
rect 5099 2465 5127 2499
rect 5172 2465 5195 2499
rect 5245 2465 5263 2499
rect 5318 2465 5331 2499
rect 5391 2465 5399 2499
rect 5464 2465 5467 2499
rect 5501 2465 5503 2499
rect 5569 2465 5576 2499
rect 5637 2465 5649 2499
rect 5705 2465 5722 2499
rect 5773 2465 5795 2499
rect 5841 2465 5868 2499
rect 5909 2465 5941 2499
rect 5977 2465 6011 2499
rect 6048 2465 6079 2499
rect 6121 2465 6147 2499
rect 6194 2465 6215 2499
rect 6267 2465 6283 2499
rect 6340 2465 6351 2499
rect 6413 2465 6419 2499
rect 6486 2465 6487 2499
rect 6521 2465 6525 2499
rect 6589 2465 6598 2499
rect 6657 2465 6671 2499
rect 6725 2465 6744 2499
rect 6793 2465 6816 2499
rect 6861 2465 6888 2499
rect 6929 2465 6960 2499
rect 6997 2465 7031 2499
rect 7066 2465 7099 2499
rect 7138 2465 7167 2499
rect 7210 2465 7235 2499
rect 7282 2465 7303 2499
rect 7354 2465 7371 2499
rect 7426 2465 7439 2499
rect 7498 2465 7507 2499
rect 7570 2465 7575 2499
rect 7642 2465 7643 2499
rect 7677 2465 7680 2499
rect 7745 2465 7752 2499
rect 7813 2465 7824 2499
rect 7881 2465 7896 2499
rect 7949 2465 7968 2499
rect 8017 2465 8040 2499
rect 8085 2465 8112 2499
rect 8153 2465 8184 2499
rect 8221 2465 8255 2499
rect 8290 2465 8323 2499
rect 8362 2465 8391 2499
rect 8434 2465 8459 2499
rect 8493 2465 8527 2499
rect 8561 2465 8595 2499
rect 8629 2465 8663 2499
rect 8697 2465 8731 2499
rect 8765 2465 8799 2499
rect 8833 2465 8867 2499
rect 8901 2465 8935 2499
rect 8969 2465 9003 2499
rect 9037 2465 9071 2499
rect 9105 2465 9139 2499
rect 9173 2465 9207 2499
rect 9241 2465 9275 2499
rect 9309 2465 9343 2499
rect 9377 2465 9445 2499
rect 2151 2440 2185 2465
rect 2207 2459 8472 2465
rect 466 2369 500 2407
rect 620 2399 642 2433
rect 688 2399 714 2433
rect 756 2399 786 2433
rect 824 2399 858 2433
rect 892 2399 926 2433
rect 964 2399 994 2433
rect 1036 2399 1062 2433
rect 1108 2399 1130 2433
rect 1180 2399 1198 2433
rect 1252 2399 1266 2433
rect 1324 2399 1334 2433
rect 1396 2399 1402 2433
rect 1468 2399 1470 2433
rect 1504 2399 1506 2433
rect 2145 2431 2191 2440
rect 466 2297 500 2335
rect 1622 2381 1656 2397
rect 1622 2313 1656 2346
rect 466 2225 500 2263
rect 620 2243 642 2277
rect 688 2243 714 2277
rect 756 2243 786 2277
rect 824 2243 858 2277
rect 892 2243 926 2277
rect 964 2243 994 2277
rect 1036 2243 1062 2277
rect 1108 2243 1130 2277
rect 1180 2243 1198 2277
rect 1252 2243 1266 2277
rect 1324 2243 1334 2277
rect 1396 2243 1402 2277
rect 1468 2243 1470 2277
rect 1504 2243 1506 2277
rect 1622 2263 1656 2274
rect 2145 2368 2151 2431
rect 2185 2368 2191 2431
rect 2145 2363 2191 2368
rect 2145 2261 2151 2363
rect 2185 2261 2191 2363
rect 2145 2256 2191 2261
rect 466 2153 500 2191
rect 2145 2193 2151 2256
rect 2185 2193 2191 2256
rect 9411 2375 9445 2465
rect 9411 2307 9445 2341
rect 2428 2231 2452 2253
rect 2428 2197 2443 2231
rect 2486 2219 2521 2253
rect 2555 2231 2590 2253
rect 2569 2219 2590 2231
rect 2624 2231 2659 2253
rect 2624 2219 2627 2231
rect 2693 2219 2728 2253
rect 2762 2219 2797 2253
rect 2831 2219 2866 2253
rect 2900 2219 2935 2253
rect 2969 2219 3004 2253
rect 3038 2219 3073 2253
rect 3107 2231 3142 2253
rect 3107 2219 3138 2231
rect 3176 2219 3211 2253
rect 3245 2219 3280 2253
rect 3314 2231 3349 2253
rect 3383 2231 3418 2253
rect 3452 2231 3487 2253
rect 3521 2231 3556 2253
rect 3590 2231 3625 2253
rect 3659 2231 3694 2253
rect 3728 2231 3762 2253
rect 3796 2231 3830 2253
rect 3318 2219 3349 2231
rect 3391 2219 3418 2231
rect 3464 2219 3487 2231
rect 3537 2219 3556 2231
rect 3610 2219 3625 2231
rect 3683 2219 3694 2231
rect 3756 2219 3762 2231
rect 3829 2219 3830 2231
rect 3864 2231 3898 2253
rect 3932 2231 3966 2253
rect 4000 2231 4034 2253
rect 4068 2231 4102 2253
rect 4136 2231 4170 2253
rect 4204 2231 4238 2253
rect 3864 2219 3868 2231
rect 3932 2219 3941 2231
rect 4000 2219 4014 2231
rect 4068 2219 4087 2231
rect 4136 2219 4160 2231
rect 4204 2219 4233 2231
rect 4272 2219 4306 2253
rect 4340 2219 4374 2253
rect 4408 2231 4442 2253
rect 4476 2231 4510 2253
rect 4544 2231 4578 2253
rect 4612 2231 4646 2253
rect 4680 2231 4714 2253
rect 4748 2231 4782 2253
rect 4413 2219 4442 2231
rect 4486 2219 4510 2231
rect 4559 2219 4578 2231
rect 4632 2219 4646 2231
rect 4705 2219 4714 2231
rect 4778 2219 4782 2231
rect 4816 2231 4850 2253
rect 4884 2231 4918 2253
rect 4952 2231 4986 2253
rect 5020 2231 5054 2253
rect 5088 2231 5122 2253
rect 5156 2231 5190 2253
rect 5224 2231 5258 2253
rect 4816 2219 4817 2231
rect 4884 2219 4890 2231
rect 4952 2219 4963 2231
rect 5020 2219 5036 2231
rect 5088 2219 5109 2231
rect 5156 2219 5182 2231
rect 5224 2219 5255 2231
rect 5292 2219 5326 2253
rect 5360 2231 5394 2253
rect 5428 2231 5462 2253
rect 5496 2231 5530 2253
rect 5564 2231 5598 2253
rect 5632 2231 5666 2253
rect 5700 2231 5734 2253
rect 5768 2231 5802 2253
rect 5362 2219 5394 2231
rect 5435 2219 5462 2231
rect 5508 2219 5530 2231
rect 5581 2219 5598 2231
rect 5654 2219 5666 2231
rect 5727 2219 5734 2231
rect 5800 2219 5802 2231
rect 5836 2231 5870 2253
rect 5904 2231 5938 2253
rect 5972 2231 6006 2253
rect 6040 2231 6074 2253
rect 6108 2231 6142 2253
rect 6176 2231 6210 2253
rect 6244 2231 6278 2253
rect 5836 2219 5839 2231
rect 5904 2219 5912 2231
rect 5972 2219 5985 2231
rect 6040 2219 6058 2231
rect 6108 2219 6131 2231
rect 6176 2219 6204 2231
rect 6244 2219 6277 2231
rect 6312 2219 6346 2253
rect 6380 2231 6414 2253
rect 6448 2231 6482 2253
rect 6516 2231 6550 2253
rect 6584 2231 6618 2253
rect 6652 2231 6686 2253
rect 6720 2231 6754 2253
rect 6788 2231 6822 2253
rect 6384 2219 6414 2231
rect 6457 2219 6482 2231
rect 6530 2219 6550 2231
rect 6603 2219 6618 2231
rect 6675 2219 6686 2231
rect 6747 2219 6754 2231
rect 6819 2219 6822 2231
rect 6856 2231 6890 2253
rect 6924 2231 6958 2253
rect 6856 2219 6857 2231
rect 6924 2219 6929 2231
rect 6992 2219 7016 2253
rect 2477 2197 2535 2219
rect 2569 2197 2627 2219
rect 2661 2197 2790 2219
rect 2145 2182 2191 2193
rect 2718 2185 2790 2197
rect 2824 2185 2882 2219
rect 2916 2185 2974 2219
rect 3008 2197 3138 2219
rect 3172 2197 3211 2219
rect 3245 2197 3284 2219
rect 3318 2197 3357 2219
rect 3391 2197 3430 2219
rect 3464 2197 3503 2219
rect 3537 2197 3576 2219
rect 3610 2197 3649 2219
rect 3683 2197 3722 2219
rect 3756 2197 3795 2219
rect 3829 2197 3868 2219
rect 3902 2197 3941 2219
rect 3975 2197 4014 2219
rect 4048 2197 4087 2219
rect 4121 2197 4160 2219
rect 4194 2197 4233 2219
rect 4267 2197 4306 2219
rect 4340 2197 4379 2219
rect 4413 2197 4452 2219
rect 4486 2197 4525 2219
rect 4559 2197 4598 2219
rect 4632 2197 4671 2219
rect 4705 2197 4744 2219
rect 4778 2197 4817 2219
rect 4851 2197 4890 2219
rect 4924 2197 4963 2219
rect 4997 2197 5036 2219
rect 5070 2197 5109 2219
rect 5143 2197 5182 2219
rect 5216 2197 5255 2219
rect 5289 2197 5328 2219
rect 5362 2197 5401 2219
rect 5435 2197 5474 2219
rect 5508 2197 5547 2219
rect 5581 2197 5620 2219
rect 5654 2197 5693 2219
rect 5727 2197 5766 2219
rect 5800 2197 5839 2219
rect 5873 2197 5912 2219
rect 5946 2197 5985 2219
rect 6019 2197 6058 2219
rect 6092 2197 6131 2219
rect 6165 2197 6204 2219
rect 6238 2197 6277 2219
rect 6311 2197 6350 2219
rect 6384 2197 6423 2219
rect 6457 2197 6496 2219
rect 6530 2197 6569 2219
rect 6603 2197 6641 2219
rect 6675 2197 6713 2219
rect 6747 2197 6785 2219
rect 6819 2197 6857 2219
rect 6891 2197 6929 2219
rect 6963 2197 7016 2219
rect 7499 2203 7515 2237
rect 7549 2203 7583 2237
rect 7617 2203 7651 2237
rect 7701 2203 7719 2237
rect 7778 2203 7787 2237
rect 7889 2203 7898 2237
rect 7957 2203 7975 2237
rect 8025 2203 8052 2237
rect 8093 2203 8127 2237
rect 8163 2203 8195 2237
rect 8240 2203 8263 2237
rect 8317 2203 8331 2237
rect 8393 2203 8399 2237
rect 8433 2203 8435 2237
rect 8555 2211 8613 2245
rect 8647 2211 8689 2245
rect 3008 2185 3100 2197
rect 466 2081 500 2119
rect 466 2009 500 2047
rect 466 1937 500 1975
rect 574 2162 598 2164
rect 632 2162 669 2164
rect 703 2162 740 2164
rect 774 2162 811 2164
rect 845 2162 882 2164
rect 916 2162 953 2164
rect 987 2162 1024 2164
rect 1058 2162 1095 2164
rect 1129 2162 1166 2164
rect 632 2130 648 2162
rect 703 2130 722 2162
rect 774 2130 796 2162
rect 845 2130 870 2162
rect 916 2130 944 2162
rect 987 2130 1017 2162
rect 1058 2130 1090 2162
rect 1129 2130 1163 2162
rect 1200 2130 1236 2164
rect 1270 2130 1306 2164
rect 1340 2162 1376 2164
rect 1410 2162 1446 2164
rect 1480 2162 1516 2164
rect 1550 2162 1574 2164
rect 1343 2130 1376 2162
rect 1416 2130 1446 2162
rect 1489 2130 1516 2162
rect 608 2128 648 2130
rect 682 2128 722 2130
rect 756 2128 796 2130
rect 830 2128 870 2130
rect 904 2128 944 2130
rect 978 2128 1017 2130
rect 1051 2128 1090 2130
rect 1124 2128 1163 2130
rect 1197 2128 1236 2130
rect 1270 2128 1309 2130
rect 1343 2128 1382 2130
rect 1416 2128 1455 2130
rect 1489 2128 1528 2130
rect 1562 2128 1574 2162
rect 574 2096 1574 2128
rect 574 2062 598 2096
rect 632 2062 669 2096
rect 703 2062 740 2096
rect 774 2062 811 2096
rect 845 2062 882 2096
rect 916 2062 953 2096
rect 987 2062 1024 2096
rect 1058 2062 1095 2096
rect 1129 2062 1166 2096
rect 1200 2062 1236 2096
rect 1270 2062 1306 2096
rect 1340 2062 1376 2096
rect 1410 2062 1446 2096
rect 1480 2062 1516 2096
rect 1550 2062 1574 2096
rect 608 2028 648 2062
rect 682 2028 722 2062
rect 756 2028 796 2062
rect 830 2028 870 2062
rect 904 2028 944 2062
rect 978 2028 1017 2062
rect 1051 2028 1090 2062
rect 1124 2028 1163 2062
rect 1197 2028 1236 2062
rect 1270 2028 1309 2062
rect 1343 2028 1382 2062
rect 1416 2028 1455 2062
rect 1489 2028 1528 2062
rect 1562 2028 1574 2062
rect 574 1994 598 2028
rect 632 1994 669 2028
rect 703 1994 740 2028
rect 774 1994 811 2028
rect 845 1994 882 2028
rect 916 1994 953 2028
rect 987 1994 1024 2028
rect 1058 1994 1095 2028
rect 1129 1994 1166 2028
rect 1200 1994 1236 2028
rect 1270 1994 1306 2028
rect 1340 1994 1376 2028
rect 1410 1994 1446 2028
rect 1480 1994 1516 2028
rect 1550 1994 1574 2028
rect 574 1962 1574 1994
rect 608 1960 648 1962
rect 682 1960 722 1962
rect 756 1960 796 1962
rect 830 1960 870 1962
rect 904 1960 944 1962
rect 978 1960 1017 1962
rect 1051 1960 1090 1962
rect 1124 1960 1163 1962
rect 1197 1960 1236 1962
rect 1270 1960 1309 1962
rect 1343 1960 1382 1962
rect 1416 1960 1455 1962
rect 1489 1960 1528 1962
rect 632 1928 648 1960
rect 703 1928 722 1960
rect 774 1928 796 1960
rect 845 1928 870 1960
rect 916 1928 944 1960
rect 987 1928 1017 1960
rect 1058 1928 1090 1960
rect 1129 1928 1163 1960
rect 574 1926 598 1928
rect 632 1926 669 1928
rect 703 1926 740 1928
rect 774 1926 811 1928
rect 845 1926 882 1928
rect 916 1926 953 1928
rect 987 1926 1024 1928
rect 1058 1926 1095 1928
rect 1129 1926 1166 1928
rect 1200 1926 1236 1960
rect 1270 1926 1306 1960
rect 1343 1928 1376 1960
rect 1416 1928 1446 1960
rect 1489 1928 1516 1960
rect 1562 1928 1574 1962
rect 1340 1926 1376 1928
rect 1410 1926 1446 1928
rect 1480 1926 1516 1928
rect 1550 1926 1574 1928
rect 2145 2125 2151 2182
rect 2185 2125 2191 2182
rect 8555 2173 8689 2211
rect 8555 2158 8613 2173
rect 8647 2158 8689 2173
rect 2145 2108 2191 2125
rect 2145 2057 2151 2108
rect 2185 2057 2191 2108
rect 2470 2103 2492 2137
rect 2538 2103 2564 2137
rect 2606 2103 2636 2137
rect 2674 2103 2708 2137
rect 2742 2103 2776 2137
rect 2814 2103 2844 2137
rect 2886 2103 2912 2137
rect 2958 2103 2980 2137
rect 3030 2103 3048 2137
rect 3102 2103 3116 2137
rect 3174 2103 3184 2137
rect 3246 2103 3252 2137
rect 3318 2103 3320 2137
rect 3354 2103 3356 2137
rect 3422 2103 3428 2137
rect 3490 2103 3500 2137
rect 3558 2103 3572 2137
rect 3626 2103 3644 2137
rect 3694 2103 3716 2137
rect 3762 2103 3788 2137
rect 3830 2103 3860 2137
rect 3898 2103 3932 2137
rect 3966 2103 4000 2137
rect 4038 2103 4068 2137
rect 4110 2103 4136 2137
rect 4182 2103 4204 2137
rect 4254 2103 4272 2137
rect 4326 2103 4340 2137
rect 4746 2103 4760 2137
rect 4814 2103 4832 2137
rect 4882 2103 4904 2137
rect 4950 2103 4976 2137
rect 5018 2103 5048 2137
rect 5086 2103 5120 2137
rect 5154 2103 5188 2137
rect 5226 2103 5256 2137
rect 5298 2103 5324 2137
rect 5370 2103 5392 2137
rect 5442 2103 5460 2137
rect 5514 2103 5528 2137
rect 5586 2103 5596 2137
rect 5658 2103 5664 2137
rect 5730 2103 5732 2137
rect 5766 2103 5768 2137
rect 5834 2103 5840 2137
rect 5902 2103 5912 2137
rect 5970 2103 5984 2137
rect 6038 2103 6056 2137
rect 6106 2103 6128 2137
rect 6174 2103 6200 2137
rect 6242 2103 6272 2137
rect 6310 2103 6344 2137
rect 6378 2103 6412 2137
rect 6450 2103 6480 2137
rect 6522 2103 6548 2137
rect 6594 2103 6616 2137
rect 8555 2124 8571 2158
rect 8605 2139 8613 2158
rect 8605 2124 8639 2139
rect 8673 2124 8689 2158
rect 9411 2239 9445 2273
rect 9411 2171 9445 2205
rect 9411 2103 9445 2137
rect 2145 2034 2191 2057
rect 2145 1989 2151 2034
rect 2185 1989 2191 2034
rect 2145 1960 2191 1989
rect 466 1865 500 1903
rect 2145 1921 2151 1960
rect 2185 1921 2191 1960
rect 2145 1887 2191 1921
rect 4472 2082 4506 2092
rect 4472 2008 4506 2042
rect 4472 1940 4506 1971
rect 2145 1852 2151 1887
rect 2185 1852 2191 1887
rect 2470 1867 2492 1901
rect 2538 1867 2564 1901
rect 2606 1867 2636 1901
rect 2674 1867 2708 1901
rect 2742 1867 2776 1901
rect 2814 1867 2844 1901
rect 2886 1867 2912 1901
rect 2958 1867 2980 1901
rect 3030 1867 3048 1901
rect 3102 1867 3116 1901
rect 3174 1867 3184 1901
rect 3246 1867 3252 1901
rect 3318 1867 3320 1901
rect 3354 1867 3356 1901
rect 3422 1867 3428 1901
rect 3490 1867 3500 1901
rect 3558 1867 3572 1901
rect 3626 1867 3644 1901
rect 3694 1867 3716 1901
rect 3762 1867 3788 1901
rect 3830 1867 3860 1901
rect 3898 1867 3932 1901
rect 3966 1867 4000 1901
rect 4038 1867 4068 1901
rect 4110 1867 4136 1901
rect 4182 1867 4204 1901
rect 4254 1867 4272 1901
rect 4326 1867 4340 1901
rect 4472 1872 4506 1894
rect 466 1793 500 1831
rect 620 1807 642 1841
rect 688 1807 714 1841
rect 756 1807 786 1841
rect 824 1807 858 1841
rect 892 1807 926 1841
rect 964 1807 994 1841
rect 1036 1807 1062 1841
rect 1108 1807 1130 1841
rect 1180 1807 1198 1841
rect 1252 1807 1266 1841
rect 1324 1807 1334 1841
rect 1396 1807 1402 1841
rect 1468 1807 1470 1841
rect 1504 1807 1506 1841
rect 2145 1819 2191 1852
rect 1622 1780 1656 1796
rect 466 1721 500 1759
rect 1100 1764 1622 1773
rect 1100 1730 1114 1764
rect 1148 1730 1186 1764
rect 1220 1746 1622 1764
rect 1220 1730 1656 1746
rect 1100 1719 1656 1730
rect 466 1649 500 1687
rect 1622 1685 1656 1719
rect 620 1651 642 1685
rect 688 1651 714 1685
rect 756 1651 786 1685
rect 824 1651 858 1685
rect 892 1651 926 1685
rect 964 1651 994 1685
rect 1036 1651 1062 1685
rect 1108 1651 1130 1685
rect 1180 1651 1198 1685
rect 1252 1651 1266 1685
rect 1324 1651 1334 1685
rect 1396 1651 1402 1685
rect 1468 1651 1470 1685
rect 1504 1651 1506 1685
rect 1622 1617 1656 1651
rect 466 1577 500 1615
rect 1100 1607 1656 1617
rect 1100 1573 1114 1607
rect 1148 1573 1186 1607
rect 1220 1590 1656 1607
rect 1220 1573 1622 1590
rect 1100 1563 1622 1573
rect 466 1505 500 1543
rect 1622 1540 1656 1556
rect 2145 1778 2151 1819
rect 2185 1778 2191 1819
rect 2145 1751 2191 1778
rect 2145 1704 2151 1751
rect 2185 1704 2191 1751
rect 2145 1683 2191 1704
rect 2145 1630 2151 1683
rect 2185 1630 2191 1683
rect 4472 1804 4506 1817
rect 4472 1736 4506 1740
rect 4472 1697 4506 1702
rect 4580 2077 4614 2092
rect 7549 2047 7571 2081
rect 7617 2047 7643 2081
rect 7685 2047 7715 2081
rect 7753 2047 7787 2081
rect 7821 2047 7855 2081
rect 7893 2047 7923 2081
rect 7965 2047 7991 2081
rect 8037 2047 8059 2081
rect 8109 2047 8127 2081
rect 8181 2047 8195 2081
rect 8253 2047 8263 2081
rect 8325 2047 8331 2081
rect 8397 2047 8399 2081
rect 8433 2047 8435 2081
rect 4580 2006 4614 2042
rect 9411 2035 9445 2069
rect 9405 2001 9411 2019
rect 9716 2484 10412 2524
rect 9716 2450 9723 2484
rect 9757 2450 9795 2484
rect 9829 2450 9867 2484
rect 9901 2450 9939 2484
rect 9973 2450 10011 2484
rect 10045 2450 10083 2484
rect 10117 2450 10155 2484
rect 10189 2450 10227 2484
rect 10261 2450 10299 2484
rect 10333 2450 10371 2484
rect 10405 2450 10412 2484
rect 9716 2410 10412 2450
rect 9716 2376 9723 2410
rect 9757 2376 9795 2410
rect 9829 2376 9867 2410
rect 9901 2376 9939 2410
rect 9973 2376 10011 2410
rect 10045 2376 10083 2410
rect 10117 2376 10155 2410
rect 10189 2376 10227 2410
rect 10261 2376 10299 2410
rect 10333 2376 10371 2410
rect 10405 2376 10412 2410
rect 9716 2336 10412 2376
rect 9716 2302 9723 2336
rect 9757 2302 9795 2336
rect 9829 2302 9867 2336
rect 9901 2302 9939 2336
rect 9973 2302 10011 2336
rect 10045 2302 10083 2336
rect 10117 2302 10155 2336
rect 10189 2302 10227 2336
rect 10261 2302 10299 2336
rect 10333 2302 10371 2336
rect 10405 2302 10412 2336
rect 9716 2262 10412 2302
rect 9716 2228 9723 2262
rect 9757 2228 9795 2262
rect 9829 2228 9867 2262
rect 9901 2228 9939 2262
rect 9973 2228 10011 2262
rect 10045 2228 10083 2262
rect 10117 2228 10155 2262
rect 10189 2228 10227 2262
rect 10261 2228 10299 2262
rect 10333 2228 10371 2262
rect 10405 2228 10412 2262
rect 9716 2188 10412 2228
rect 9716 2154 9723 2188
rect 9757 2154 9795 2188
rect 9829 2154 9867 2188
rect 9901 2154 9939 2188
rect 9973 2154 10011 2188
rect 10045 2154 10083 2188
rect 10117 2154 10155 2188
rect 10189 2154 10227 2188
rect 10261 2154 10299 2188
rect 10333 2154 10371 2188
rect 10405 2154 10412 2188
rect 9716 2114 10412 2154
rect 9716 2080 9723 2114
rect 9757 2080 9795 2114
rect 9829 2080 9867 2114
rect 9901 2080 9939 2114
rect 9973 2080 10011 2114
rect 10045 2080 10083 2114
rect 10117 2080 10155 2114
rect 10189 2080 10227 2114
rect 10261 2080 10299 2114
rect 10333 2080 10371 2114
rect 10405 2080 10412 2114
rect 9716 2040 10412 2080
rect 9445 2001 9451 2019
rect 9405 1987 9451 2001
rect 4580 1936 4614 1955
rect 4580 1900 4614 1902
rect 4746 1867 4760 1901
rect 4814 1867 4832 1901
rect 4882 1867 4904 1901
rect 4950 1867 4976 1901
rect 5018 1867 5048 1901
rect 5086 1867 5120 1901
rect 5154 1867 5188 1901
rect 5226 1867 5256 1901
rect 5298 1867 5324 1901
rect 5370 1867 5392 1901
rect 5442 1867 5460 1901
rect 5514 1867 5528 1901
rect 5586 1867 5596 1901
rect 5658 1867 5664 1901
rect 5730 1867 5732 1901
rect 5766 1867 5768 1901
rect 5834 1867 5840 1901
rect 5902 1867 5912 1901
rect 5970 1867 5984 1901
rect 6038 1867 6056 1901
rect 6106 1867 6128 1901
rect 6174 1867 6200 1901
rect 6242 1867 6272 1901
rect 6310 1867 6344 1901
rect 6378 1867 6412 1901
rect 6450 1867 6480 1901
rect 6522 1867 6548 1901
rect 6594 1867 6616 1901
rect 6829 1886 6863 1908
rect 8485 1886 8519 1908
rect 9405 1933 9411 1987
rect 9445 1933 9451 1987
rect 9405 1908 9451 1933
rect 9405 1865 9411 1908
rect 9445 1865 9451 1908
rect 4580 1811 4614 1832
rect 9405 1831 9451 1865
rect 7001 1822 7043 1823
rect 7077 1822 7119 1823
rect 7153 1822 7195 1823
rect 7229 1822 7271 1823
rect 7305 1822 7347 1823
rect 7381 1822 7423 1823
rect 7457 1822 7499 1823
rect 7533 1822 7575 1823
rect 7609 1822 7651 1823
rect 7685 1822 7726 1823
rect 7760 1822 7801 1823
rect 7835 1822 7876 1823
rect 7910 1822 7951 1823
rect 7985 1822 8026 1823
rect 8060 1822 8101 1823
rect 8135 1822 8176 1823
rect 8210 1822 8251 1823
rect 8285 1822 8326 1823
rect 8360 1822 8401 1823
rect 6893 1788 6909 1822
rect 6943 1789 6967 1822
rect 7011 1789 7043 1822
rect 6943 1788 6977 1789
rect 7011 1788 7045 1789
rect 7079 1788 7113 1822
rect 7153 1789 7181 1822
rect 7229 1789 7249 1822
rect 7305 1789 7317 1822
rect 7381 1789 7385 1822
rect 7147 1788 7181 1789
rect 7215 1788 7249 1789
rect 7283 1788 7317 1789
rect 7351 1788 7385 1789
rect 7419 1789 7423 1822
rect 7487 1789 7499 1822
rect 7555 1789 7575 1822
rect 7623 1789 7651 1822
rect 7419 1788 7453 1789
rect 7487 1788 7521 1789
rect 7555 1788 7589 1789
rect 7623 1788 7657 1789
rect 7691 1788 7725 1822
rect 7760 1789 7793 1822
rect 7835 1789 7862 1822
rect 7910 1789 7931 1822
rect 7985 1789 8000 1822
rect 8060 1789 8069 1822
rect 8135 1789 8138 1822
rect 7759 1788 7793 1789
rect 7827 1788 7862 1789
rect 7896 1788 7931 1789
rect 7965 1788 8000 1789
rect 8034 1788 8069 1789
rect 8103 1788 8138 1789
rect 8172 1789 8176 1822
rect 8241 1789 8251 1822
rect 8310 1789 8326 1822
rect 8379 1789 8401 1822
rect 8172 1788 8207 1789
rect 8241 1788 8276 1789
rect 8310 1788 8345 1789
rect 8379 1788 8414 1789
rect 8448 1788 8464 1822
rect 9405 1795 9411 1831
rect 9445 1795 9451 1831
rect 4580 1726 4614 1762
rect 9405 1763 9451 1795
rect 4580 1676 4614 1688
rect 6829 1702 6863 1724
rect 2470 1631 2492 1665
rect 2538 1631 2564 1665
rect 2606 1631 2636 1665
rect 2674 1631 2708 1665
rect 2742 1631 2776 1665
rect 2814 1631 2844 1665
rect 2886 1631 2912 1665
rect 2958 1631 2980 1665
rect 3030 1631 3048 1665
rect 3102 1631 3116 1665
rect 3174 1631 3184 1665
rect 3246 1631 3252 1665
rect 3318 1631 3320 1665
rect 3354 1631 3356 1665
rect 3422 1631 3428 1665
rect 3490 1631 3500 1665
rect 3558 1631 3572 1665
rect 3626 1631 3644 1665
rect 3694 1631 3716 1665
rect 3762 1631 3788 1665
rect 3830 1631 3860 1665
rect 3898 1631 3932 1665
rect 3966 1631 4000 1665
rect 4038 1631 4068 1665
rect 4110 1631 4136 1665
rect 4182 1631 4204 1665
rect 4254 1631 4272 1665
rect 4326 1631 4340 1665
rect 2145 1615 2191 1630
rect 2145 1556 2151 1615
rect 2185 1556 2191 1615
rect 2145 1547 2191 1556
rect 620 1495 642 1529
rect 688 1495 714 1529
rect 756 1495 786 1529
rect 824 1495 858 1529
rect 892 1495 926 1529
rect 964 1495 994 1529
rect 1036 1495 1062 1529
rect 1108 1495 1130 1529
rect 1180 1495 1198 1529
rect 1252 1495 1266 1529
rect 1324 1495 1334 1529
rect 1396 1495 1402 1529
rect 1468 1495 1470 1529
rect 1504 1495 1506 1529
rect 466 1433 500 1471
rect 2145 1482 2151 1547
rect 2185 1482 2191 1547
rect 2145 1479 2191 1482
rect 2145 1445 2151 1479
rect 2185 1445 2191 1479
rect 2145 1442 2191 1445
rect 466 1361 500 1399
rect 574 1367 597 1401
rect 632 1367 668 1401
rect 709 1367 738 1401
rect 787 1367 808 1401
rect 865 1367 878 1401
rect 943 1367 948 1401
rect 982 1367 987 1401
rect 1053 1367 1065 1401
rect 1124 1367 1143 1401
rect 1195 1367 1220 1401
rect 1266 1367 1297 1401
rect 1337 1367 1374 1401
rect 1408 1367 1445 1401
rect 1485 1367 1516 1401
rect 1562 1367 1574 1401
rect 2145 1377 2151 1442
rect 2185 1377 2191 1442
rect 4472 1619 4506 1634
rect 4746 1631 4760 1665
rect 4814 1631 4832 1665
rect 4882 1631 4904 1665
rect 4950 1631 4976 1665
rect 5018 1631 5048 1665
rect 5086 1631 5120 1665
rect 5154 1631 5188 1665
rect 5226 1631 5256 1665
rect 5298 1631 5324 1665
rect 5370 1631 5392 1665
rect 5442 1631 5460 1665
rect 5514 1631 5528 1665
rect 5586 1631 5596 1665
rect 5658 1631 5664 1665
rect 5730 1631 5732 1665
rect 5766 1631 5768 1665
rect 5834 1631 5840 1665
rect 5902 1631 5912 1665
rect 5970 1631 5984 1665
rect 6038 1631 6056 1665
rect 6106 1631 6128 1665
rect 6174 1631 6200 1665
rect 6242 1631 6272 1665
rect 6310 1631 6344 1665
rect 6378 1631 6412 1665
rect 6450 1631 6480 1665
rect 6522 1631 6548 1665
rect 6594 1631 6616 1665
rect 8485 1702 8519 1724
rect 9405 1716 9411 1763
rect 9445 1716 9451 1763
rect 9405 1695 9451 1716
rect 9405 1637 9411 1695
rect 9445 1637 9451 1695
rect 4472 1541 4506 1565
rect 4472 1461 4506 1496
rect 9405 1627 9451 1637
rect 9405 1593 9411 1627
rect 9445 1593 9451 1627
rect 9405 1592 9451 1593
rect 9716 2006 9723 2040
rect 9757 2006 9795 2040
rect 9829 2006 9867 2040
rect 9901 2006 9939 2040
rect 9973 2006 10011 2040
rect 10045 2006 10083 2040
rect 10117 2006 10155 2040
rect 10189 2006 10227 2040
rect 10261 2006 10299 2040
rect 10333 2006 10371 2040
rect 10405 2006 10412 2040
rect 10488 2787 10522 2821
rect 12287 2815 12325 2821
rect 12359 2815 12397 2821
rect 12431 2815 12469 2821
rect 12503 2815 12542 2821
rect 12576 2815 12615 2821
rect 12649 2815 12688 2821
rect 12722 2815 12761 2821
rect 12795 2815 12834 2821
rect 12868 2815 12907 2821
rect 12941 2815 12980 2821
rect 13014 2815 13053 2821
rect 13087 2815 13126 2821
rect 13160 2815 13199 2821
rect 13233 2815 13272 2821
rect 13306 2815 13345 2821
rect 13379 2815 13418 2821
rect 13452 2815 13491 2821
rect 13525 2815 13564 2821
rect 13598 2815 13637 2821
rect 13671 2815 13710 2821
rect 13744 2815 13783 2821
rect 13817 2815 13856 2821
rect 13890 2815 13929 2821
rect 13963 2815 14002 2821
rect 14036 2815 14075 2821
rect 14109 2815 14148 2821
rect 14182 2815 14221 2821
rect 14255 2815 14294 2821
rect 14328 2815 14367 2821
rect 14401 2815 14440 2821
rect 14474 2815 14513 2821
rect 14547 2815 14586 2821
rect 14620 2815 14659 2821
rect 14693 2815 14732 2821
rect 14766 2815 14805 2821
rect 14839 2815 14878 2821
rect 14912 2815 14951 2821
rect 14985 2815 15024 2821
rect 15058 2815 15097 2821
rect 15131 2815 15170 2821
rect 15204 2815 15243 2821
rect 15277 2815 15316 2821
rect 15350 2815 15389 2821
rect 15423 2815 15462 2821
rect 15496 2815 15535 2821
rect 15569 2815 15608 2821
rect 15642 2815 15681 2821
rect 15715 2815 15754 2821
rect 15788 2815 15827 2821
rect 15861 2815 15900 2821
rect 15968 2849 16002 2855
rect 16036 2849 16070 2855
rect 16104 2849 16138 2855
rect 16172 2849 16206 2855
rect 16240 2849 16274 2855
rect 16308 2849 16342 2855
rect 15968 2821 15973 2849
rect 16036 2821 16046 2849
rect 16104 2821 16119 2849
rect 16172 2821 16192 2849
rect 16240 2821 16265 2849
rect 16308 2821 16338 2849
rect 16376 2821 16444 2855
rect 18140 2849 18156 2883
rect 18190 2849 18224 2883
rect 18258 2849 18292 2883
rect 18326 2849 18360 2883
rect 18394 2849 18417 2883
rect 18462 2849 18496 2883
rect 18531 2849 18564 2883
rect 18611 2849 18632 2883
rect 18691 2849 18700 2883
rect 18734 2849 18737 2883
rect 18802 2849 18817 2883
rect 18870 2849 18897 2883
rect 18938 2849 18972 2883
rect 19011 2849 19040 2883
rect 19996 2854 20042 2892
rect 15934 2815 15973 2821
rect 16007 2815 16046 2821
rect 16080 2815 16119 2821
rect 16153 2815 16192 2821
rect 16226 2815 16265 2821
rect 16299 2815 16338 2821
rect 16372 2815 16444 2821
rect 10488 2719 10522 2753
rect 16410 2776 16444 2815
rect 19996 2820 20002 2854
rect 20036 2820 20042 2854
rect 17916 2768 17932 2802
rect 17966 2778 18000 2802
rect 18034 2778 18050 2802
rect 17969 2768 18000 2778
rect 18041 2768 18050 2778
rect 19996 2782 20042 2820
rect 17969 2744 18007 2768
rect 19996 2748 20002 2782
rect 20036 2748 20042 2782
rect 10488 2651 10522 2685
rect 10488 2583 10522 2617
rect 10612 2710 10719 2728
rect 10612 2676 10637 2710
rect 10671 2676 10719 2710
rect 10612 2618 10719 2676
rect 10612 2584 10613 2618
rect 10647 2584 10685 2618
rect 10612 2572 10719 2584
rect 16410 2727 16444 2742
rect 16410 2659 16444 2669
rect 16410 2591 16444 2596
rect 10488 2515 10522 2549
rect 10488 2357 10522 2481
rect 10488 2289 10522 2323
rect 10488 2221 10522 2255
rect 16410 2484 16444 2489
rect 16410 2411 16444 2421
rect 16410 2338 16444 2353
rect 16410 2265 16444 2285
rect 10488 2153 10522 2187
rect 10647 2188 10685 2213
rect 10668 2179 10685 2188
rect 10613 2154 10634 2179
rect 10668 2154 10719 2179
rect 10613 2138 10719 2154
rect 16410 2192 16444 2217
rect 10488 2047 10522 2119
rect 16410 2119 16444 2149
rect 16410 2047 16444 2081
rect 10488 2013 10500 2047
rect 10534 2013 10556 2047
rect 10607 2013 10624 2047
rect 10680 2013 10692 2047
rect 10753 2013 10760 2047
rect 10826 2013 10828 2047
rect 10862 2013 10865 2047
rect 10930 2013 10938 2047
rect 10998 2013 11010 2047
rect 11066 2013 11082 2047
rect 11134 2013 11154 2047
rect 11202 2013 11226 2047
rect 11270 2013 11298 2047
rect 11338 2013 11370 2047
rect 11406 2013 11440 2047
rect 11476 2013 11508 2047
rect 11548 2013 11576 2047
rect 11620 2013 11644 2047
rect 11692 2013 11712 2047
rect 11764 2013 11780 2047
rect 11836 2013 11848 2047
rect 11908 2013 11916 2047
rect 11980 2013 11984 2047
rect 12086 2013 12090 2047
rect 12154 2013 12162 2047
rect 12222 2013 12234 2047
rect 12290 2013 12306 2047
rect 12358 2013 12378 2047
rect 12426 2013 12450 2047
rect 12494 2013 12522 2047
rect 12562 2013 12594 2047
rect 12630 2013 12664 2047
rect 12700 2013 12732 2047
rect 12772 2013 12800 2047
rect 12844 2013 12868 2047
rect 12916 2013 12936 2047
rect 12988 2013 13004 2047
rect 13060 2013 13072 2047
rect 13132 2013 13140 2047
rect 13204 2013 13208 2047
rect 13310 2013 13314 2047
rect 13378 2013 13386 2047
rect 13446 2013 13458 2047
rect 13514 2013 13530 2047
rect 13582 2013 13602 2047
rect 13650 2013 13674 2047
rect 13718 2013 13746 2047
rect 13786 2013 13818 2047
rect 13854 2013 13888 2047
rect 13924 2013 13956 2047
rect 13996 2013 14024 2047
rect 14068 2013 14092 2047
rect 14140 2013 14160 2047
rect 14212 2013 14228 2047
rect 14284 2013 14296 2047
rect 14356 2013 14364 2047
rect 14428 2013 14432 2047
rect 14534 2013 14538 2047
rect 14602 2013 14610 2047
rect 14670 2013 14682 2047
rect 14738 2013 14754 2047
rect 14806 2013 14826 2047
rect 14874 2013 14898 2047
rect 14942 2013 14970 2047
rect 15010 2013 15042 2047
rect 15078 2013 15112 2047
rect 15148 2013 15180 2047
rect 15220 2013 15248 2047
rect 15292 2013 15316 2047
rect 15364 2013 15384 2047
rect 15436 2013 15452 2047
rect 15508 2013 15520 2047
rect 15580 2013 15588 2047
rect 15652 2013 15656 2047
rect 15758 2013 15762 2047
rect 15826 2013 15834 2047
rect 15894 2013 15906 2047
rect 15962 2013 15978 2047
rect 16030 2013 16050 2047
rect 16098 2013 16122 2047
rect 16166 2013 16194 2047
rect 16234 2013 16266 2047
rect 16302 2013 16336 2047
rect 16372 2013 16444 2047
rect 16563 2579 17258 2694
rect 18140 2693 18156 2727
rect 18190 2693 18224 2727
rect 18258 2693 18292 2727
rect 18326 2693 18360 2727
rect 18394 2693 18428 2727
rect 18464 2693 18496 2727
rect 18543 2693 18564 2727
rect 18622 2693 18632 2727
rect 18734 2693 18744 2727
rect 18802 2693 18822 2727
rect 18870 2693 18900 2727
rect 18938 2693 18972 2727
rect 19012 2693 19040 2727
rect 19996 2710 20042 2748
rect 19996 2676 20002 2710
rect 20036 2676 20042 2710
rect 19996 2638 20042 2676
rect 16563 2545 16601 2579
rect 16635 2545 16675 2579
rect 16709 2545 16749 2579
rect 16783 2545 16823 2579
rect 16857 2545 16897 2579
rect 16931 2545 16971 2579
rect 17005 2545 17045 2579
rect 17079 2545 17119 2579
rect 17153 2545 17192 2579
rect 17226 2545 17258 2579
rect 17793 2572 17805 2606
rect 17851 2572 17878 2606
rect 17923 2572 17951 2606
rect 17995 2572 18024 2606
rect 18067 2572 18097 2606
rect 18139 2572 18170 2606
rect 18210 2572 18243 2606
rect 18281 2572 18316 2606
rect 18352 2572 18389 2606
rect 18423 2572 18460 2606
rect 18496 2572 18531 2606
rect 18569 2572 18602 2606
rect 18642 2572 18673 2606
rect 18714 2572 18744 2606
rect 18786 2572 18815 2606
rect 18858 2572 18886 2606
rect 18930 2572 18957 2606
rect 19002 2572 19028 2606
rect 19074 2572 19086 2606
rect 19996 2604 20002 2638
rect 20036 2604 20042 2638
rect 16563 2507 17258 2545
rect 16563 2473 16601 2507
rect 16635 2473 16675 2507
rect 16709 2473 16749 2507
rect 16783 2473 16823 2507
rect 16857 2473 16897 2507
rect 16931 2473 16971 2507
rect 17005 2473 17045 2507
rect 17079 2473 17119 2507
rect 17153 2473 17192 2507
rect 17226 2473 17258 2507
rect 16563 2435 17258 2473
rect 16563 2401 16601 2435
rect 16635 2401 16675 2435
rect 16709 2401 16749 2435
rect 16783 2401 16823 2435
rect 16857 2401 16897 2435
rect 16931 2401 16971 2435
rect 17005 2401 17045 2435
rect 17079 2401 17119 2435
rect 17153 2401 17192 2435
rect 17226 2410 17258 2435
rect 19996 2566 20042 2604
rect 19996 2532 20002 2566
rect 20036 2532 20042 2566
rect 19996 2494 20042 2532
rect 19996 2460 20002 2494
rect 20036 2460 20042 2494
rect 19996 2422 20042 2460
rect 17226 2401 19045 2410
rect 16563 2376 19045 2401
rect 19996 2388 20002 2422
rect 20036 2388 20042 2422
rect 19996 2350 20042 2388
rect 19996 2316 20002 2350
rect 20036 2316 20042 2350
rect 19045 2293 19585 2294
rect 19045 2259 19079 2293
rect 19113 2259 19152 2293
rect 19186 2259 19225 2293
rect 19259 2259 19298 2293
rect 19332 2259 19371 2293
rect 19405 2259 19444 2293
rect 19478 2259 19517 2293
rect 19551 2259 19585 2293
rect 19045 2219 19585 2259
rect 19045 2185 19079 2219
rect 19113 2185 19152 2219
rect 19186 2185 19225 2219
rect 19259 2185 19298 2219
rect 19332 2185 19371 2219
rect 19405 2185 19444 2219
rect 19478 2185 19517 2219
rect 19551 2185 19585 2219
rect 19045 2145 19585 2185
rect 19045 2111 19079 2145
rect 19113 2111 19152 2145
rect 19186 2111 19225 2145
rect 19259 2111 19298 2145
rect 19332 2111 19371 2145
rect 19405 2111 19444 2145
rect 19478 2111 19517 2145
rect 19551 2111 19585 2145
rect 19045 2071 19585 2111
rect 19045 2070 19079 2071
rect 16563 2066 16590 2070
rect 16624 2066 16662 2070
rect 16696 2066 16734 2070
rect 16768 2066 16806 2070
rect 16840 2066 19079 2070
rect 16563 2037 19079 2066
rect 19113 2037 19152 2071
rect 19186 2037 19225 2071
rect 19259 2037 19298 2071
rect 19332 2037 19371 2071
rect 19405 2037 19444 2071
rect 19478 2037 19517 2071
rect 19551 2037 19585 2071
rect 16563 2035 19585 2037
rect 9716 1966 10412 2006
rect 9716 1932 9723 1966
rect 9757 1932 9795 1966
rect 9829 1932 9867 1966
rect 9901 1932 9939 1966
rect 9973 1932 10011 1966
rect 10045 1932 10083 1966
rect 10117 1932 10155 1966
rect 10189 1932 10227 1966
rect 10261 1932 10299 1966
rect 10333 1932 10371 1966
rect 10405 1932 10412 1966
rect 16597 2012 16631 2035
rect 16665 2012 16699 2035
rect 16624 2001 16631 2012
rect 16696 2001 16699 2012
rect 16733 2012 16767 2035
rect 16801 2012 16835 2035
rect 16733 2001 16734 2012
rect 16801 2001 16806 2012
rect 16869 2001 16903 2035
rect 16937 2001 16971 2035
rect 17005 2001 17039 2035
rect 17073 2001 17107 2035
rect 17141 2001 17175 2035
rect 17209 2001 17243 2035
rect 17277 2001 17311 2035
rect 17345 2001 17379 2035
rect 17413 2001 17447 2035
rect 17481 2001 17515 2035
rect 17549 2001 17583 2035
rect 17617 2001 17651 2035
rect 17685 2001 17719 2035
rect 17753 2001 17787 2035
rect 17821 2001 17855 2035
rect 17889 2001 17923 2035
rect 17957 2001 17991 2035
rect 18025 2001 18059 2035
rect 18093 2001 18127 2035
rect 18161 2001 18195 2035
rect 18229 2001 18263 2035
rect 18297 2001 18331 2035
rect 18365 2001 18399 2035
rect 18433 2001 18467 2035
rect 18501 2001 18535 2035
rect 18569 2001 18603 2035
rect 18637 2001 18671 2035
rect 18705 2001 18739 2035
rect 18773 2001 18807 2035
rect 18841 2001 18875 2035
rect 18909 2001 18943 2035
rect 18977 2001 19011 2035
rect 19045 2001 19585 2035
rect 16563 1978 16590 2001
rect 16624 1978 16662 2001
rect 16696 1978 16734 2001
rect 16768 1978 16806 2001
rect 16840 1997 19585 2001
rect 16840 1978 19079 1997
rect 16563 1966 19079 1978
rect 9716 1921 10412 1932
rect 9716 1918 12405 1921
rect 9716 1884 9734 1918
rect 9768 1898 9808 1918
rect 9842 1898 9882 1918
rect 9916 1898 9956 1918
rect 9990 1898 10030 1918
rect 10064 1898 10104 1918
rect 10138 1898 10178 1918
rect 10212 1898 10252 1918
rect 10286 1898 10326 1918
rect 10360 1898 10400 1918
rect 10434 1898 10473 1918
rect 10507 1898 10546 1918
rect 10580 1898 10619 1918
rect 10653 1898 10692 1918
rect 10726 1898 10765 1918
rect 10799 1898 10838 1918
rect 10872 1898 10911 1918
rect 10945 1898 10984 1918
rect 11018 1898 11057 1918
rect 11091 1898 11130 1918
rect 11164 1898 11203 1918
rect 11237 1898 11276 1918
rect 11310 1898 11349 1918
rect 11383 1898 11422 1918
rect 11456 1898 11495 1918
rect 11529 1898 11568 1918
rect 11602 1898 11641 1918
rect 11675 1898 11714 1918
rect 11748 1898 11787 1918
rect 11821 1898 11860 1918
rect 11894 1898 11933 1918
rect 11967 1898 12006 1918
rect 12040 1898 12079 1918
rect 12113 1898 12152 1918
rect 12186 1898 12225 1918
rect 12259 1898 12298 1918
rect 12332 1898 12371 1918
rect 12756 1911 16563 1938
rect 19045 1963 19079 1966
rect 19113 1963 19152 1997
rect 19186 1963 19225 1997
rect 19259 1963 19298 1997
rect 19332 1963 19371 1997
rect 19405 1963 19444 1997
rect 19478 1963 19517 1997
rect 19551 1963 19585 1997
rect 19045 1932 19585 1963
rect 19011 1923 19585 1932
rect 19996 2278 20042 2316
rect 19996 2244 20002 2278
rect 20036 2244 20042 2278
rect 19996 2206 20042 2244
rect 19996 2172 20002 2206
rect 20036 2172 20042 2206
rect 19996 2134 20042 2172
rect 19996 2100 20002 2134
rect 20036 2100 20042 2134
rect 19996 2062 20042 2100
rect 19996 2028 20002 2062
rect 20036 2028 20042 2062
rect 19996 1990 20042 2028
rect 24079 1991 24121 2025
rect 24155 1991 24197 2025
rect 24231 1991 24273 2025
rect 24307 1991 24349 2025
rect 24383 1991 24424 2025
rect 24458 1991 24499 2025
rect 24533 1991 24574 2025
rect 24608 1991 24649 2025
rect 19996 1956 20002 1990
rect 20036 1956 20042 1990
rect 19996 1924 20042 1956
rect 12790 1898 12830 1911
rect 12864 1898 12904 1911
rect 12938 1898 12978 1911
rect 13012 1898 13052 1911
rect 13086 1898 13126 1911
rect 13160 1898 13200 1911
rect 13234 1898 13274 1911
rect 13308 1898 13348 1911
rect 13382 1898 13422 1911
rect 13456 1898 13496 1911
rect 13530 1898 13569 1911
rect 13603 1898 13642 1911
rect 13676 1898 13715 1911
rect 13749 1898 13788 1911
rect 13822 1898 13861 1911
rect 13895 1898 13934 1911
rect 13968 1898 14007 1911
rect 14041 1898 14080 1911
rect 14114 1898 14153 1911
rect 14187 1898 14226 1911
rect 14260 1898 14299 1911
rect 14333 1898 14372 1911
rect 14406 1898 14445 1911
rect 14479 1898 14518 1911
rect 14552 1898 14591 1911
rect 14625 1898 14664 1911
rect 14698 1898 14737 1911
rect 14771 1898 14810 1911
rect 14844 1898 14883 1911
rect 14917 1898 14956 1911
rect 14990 1898 15029 1911
rect 15063 1898 15102 1911
rect 15136 1898 15175 1911
rect 15209 1898 15248 1911
rect 15282 1898 15321 1911
rect 15355 1898 15394 1911
rect 15428 1898 15467 1911
rect 15501 1898 15540 1911
rect 15574 1898 15613 1911
rect 15647 1898 15686 1911
rect 15720 1898 15759 1911
rect 15793 1898 15832 1911
rect 15866 1898 15905 1911
rect 15939 1898 15978 1911
rect 16012 1898 16051 1911
rect 16085 1898 16124 1911
rect 16158 1898 16197 1911
rect 16231 1898 16270 1911
rect 16304 1898 16343 1911
rect 16377 1898 16416 1911
rect 16450 1898 16489 1911
rect 16523 1898 16562 1911
rect 9784 1884 9808 1898
rect 9853 1884 9882 1898
rect 9922 1884 9956 1898
rect 9716 1864 9750 1884
rect 9784 1864 9819 1884
rect 9853 1864 9888 1884
rect 9922 1864 9957 1884
rect 9991 1864 10026 1898
rect 10064 1884 10095 1898
rect 10138 1884 10164 1898
rect 10212 1884 10233 1898
rect 10286 1884 10302 1898
rect 10360 1884 10371 1898
rect 10434 1884 10440 1898
rect 10507 1884 10509 1898
rect 10060 1864 10095 1884
rect 10129 1864 10164 1884
rect 10198 1864 10233 1884
rect 10267 1864 10302 1884
rect 10336 1864 10371 1884
rect 10405 1864 10440 1884
rect 10474 1864 10509 1884
rect 10543 1884 10546 1898
rect 10612 1884 10619 1898
rect 10681 1884 10692 1898
rect 10750 1884 10765 1898
rect 10819 1884 10838 1898
rect 10888 1884 10911 1898
rect 10957 1884 10984 1898
rect 11026 1884 11057 1898
rect 10543 1864 10578 1884
rect 10612 1864 10647 1884
rect 10681 1864 10716 1884
rect 10750 1864 10785 1884
rect 10819 1864 10854 1884
rect 10888 1864 10923 1884
rect 10957 1864 10992 1884
rect 11026 1864 11061 1884
rect 11095 1864 11130 1898
rect 11164 1864 11199 1898
rect 11237 1884 11268 1898
rect 11310 1884 11337 1898
rect 11383 1884 11406 1898
rect 11456 1884 11475 1898
rect 11529 1884 11544 1898
rect 11602 1884 11613 1898
rect 11675 1884 11682 1898
rect 11748 1884 11751 1898
rect 11233 1864 11268 1884
rect 11302 1864 11337 1884
rect 11371 1864 11406 1884
rect 11440 1864 11475 1884
rect 11509 1864 11544 1884
rect 11578 1864 11613 1884
rect 11647 1864 11682 1884
rect 11716 1864 11751 1884
rect 11785 1884 11787 1898
rect 11854 1884 11860 1898
rect 11923 1884 11933 1898
rect 11992 1884 12006 1898
rect 12061 1884 12079 1898
rect 12130 1884 12152 1898
rect 12199 1884 12225 1898
rect 12268 1884 12298 1898
rect 12337 1884 12371 1898
rect 11785 1864 11820 1884
rect 11854 1864 11889 1884
rect 11923 1864 11958 1884
rect 11992 1864 12027 1884
rect 12061 1864 12096 1884
rect 12130 1864 12165 1884
rect 12199 1864 12234 1884
rect 12268 1864 12303 1884
rect 12337 1864 12372 1884
rect 12406 1864 12441 1898
rect 12475 1864 12510 1898
rect 12544 1864 12579 1898
rect 12613 1864 12648 1898
rect 12682 1864 12717 1898
rect 12751 1877 12756 1898
rect 12820 1877 12830 1898
rect 12889 1877 12904 1898
rect 12958 1877 12978 1898
rect 19011 1902 19079 1923
rect 19113 1902 19152 1923
rect 12751 1864 12786 1877
rect 12820 1864 12855 1877
rect 12889 1864 12924 1877
rect 12958 1864 12993 1877
rect 19041 1868 19079 1902
rect 19113 1868 19151 1902
rect 19186 1889 19225 1923
rect 19259 1889 19298 1923
rect 19332 1889 19371 1923
rect 19405 1889 19444 1923
rect 19478 1889 19517 1923
rect 19551 1889 19585 1923
rect 19185 1868 19585 1889
rect 9716 1836 12993 1864
rect 9716 1802 9734 1836
rect 9768 1830 9808 1836
rect 9842 1830 9882 1836
rect 9916 1830 9956 1836
rect 9990 1830 10030 1836
rect 10064 1830 10104 1836
rect 10138 1830 10178 1836
rect 10212 1830 10252 1836
rect 10286 1830 10326 1836
rect 10360 1830 10400 1836
rect 10434 1830 10473 1836
rect 10507 1830 10546 1836
rect 10580 1830 10619 1836
rect 10653 1830 10692 1836
rect 10726 1830 10765 1836
rect 10799 1830 10838 1836
rect 10872 1830 10911 1836
rect 10945 1830 10984 1836
rect 11018 1830 11057 1836
rect 11091 1830 11130 1836
rect 11164 1830 11203 1836
rect 11237 1830 11276 1836
rect 11310 1830 11349 1836
rect 11383 1830 11422 1836
rect 11456 1830 11495 1836
rect 11529 1830 11568 1836
rect 11602 1830 11641 1836
rect 11675 1830 11714 1836
rect 11748 1830 11787 1836
rect 11821 1830 11860 1836
rect 11894 1830 11933 1836
rect 11967 1830 12006 1836
rect 12040 1830 12079 1836
rect 12113 1830 12152 1836
rect 12186 1830 12225 1836
rect 12259 1830 12298 1836
rect 12332 1830 12371 1836
rect 12405 1830 12993 1836
rect 9784 1802 9808 1830
rect 9853 1802 9882 1830
rect 9922 1802 9956 1830
rect 9716 1796 9750 1802
rect 9784 1796 9819 1802
rect 9853 1796 9888 1802
rect 9922 1796 9957 1802
rect 9991 1796 10026 1830
rect 10064 1802 10095 1830
rect 10138 1802 10164 1830
rect 10212 1802 10233 1830
rect 10286 1802 10302 1830
rect 10360 1802 10371 1830
rect 10434 1802 10440 1830
rect 10507 1802 10509 1830
rect 10060 1796 10095 1802
rect 10129 1796 10164 1802
rect 10198 1796 10233 1802
rect 10267 1796 10302 1802
rect 10336 1796 10371 1802
rect 10405 1796 10440 1802
rect 10474 1796 10509 1802
rect 10543 1802 10546 1830
rect 10612 1802 10619 1830
rect 10681 1802 10692 1830
rect 10750 1802 10765 1830
rect 10819 1802 10838 1830
rect 10888 1802 10911 1830
rect 10957 1802 10984 1830
rect 11026 1802 11057 1830
rect 10543 1796 10578 1802
rect 10612 1796 10647 1802
rect 10681 1796 10716 1802
rect 10750 1796 10785 1802
rect 10819 1796 10854 1802
rect 10888 1796 10923 1802
rect 10957 1796 10992 1802
rect 11026 1796 11061 1802
rect 11095 1796 11130 1830
rect 11164 1796 11199 1830
rect 11237 1802 11268 1830
rect 11310 1802 11337 1830
rect 11383 1802 11406 1830
rect 11456 1802 11475 1830
rect 11529 1802 11544 1830
rect 11602 1802 11613 1830
rect 11675 1802 11682 1830
rect 11748 1802 11751 1830
rect 11233 1796 11268 1802
rect 11302 1796 11337 1802
rect 11371 1796 11406 1802
rect 11440 1796 11475 1802
rect 11509 1796 11544 1802
rect 11578 1796 11613 1802
rect 11647 1796 11682 1802
rect 11716 1796 11751 1802
rect 11785 1802 11787 1830
rect 11854 1802 11860 1830
rect 11923 1802 11933 1830
rect 11992 1802 12006 1830
rect 12061 1802 12079 1830
rect 12130 1802 12152 1830
rect 12199 1802 12225 1830
rect 12268 1802 12298 1830
rect 12337 1802 12371 1830
rect 11785 1796 11820 1802
rect 11854 1796 11889 1802
rect 11923 1796 11958 1802
rect 11992 1796 12027 1802
rect 12061 1796 12096 1802
rect 12130 1796 12165 1802
rect 12199 1796 12234 1802
rect 12268 1796 12303 1802
rect 12337 1796 12372 1802
rect 12406 1796 12441 1830
rect 12475 1796 12510 1830
rect 12544 1796 12579 1830
rect 12613 1796 12648 1830
rect 12682 1796 12717 1830
rect 12751 1796 12786 1830
rect 12820 1796 12855 1830
rect 12889 1796 12924 1830
rect 12958 1796 12993 1830
rect 19011 1849 19585 1868
rect 19011 1816 19079 1849
rect 19113 1816 19152 1849
rect 9716 1762 12993 1796
rect 19041 1782 19079 1816
rect 19113 1782 19151 1816
rect 19186 1815 19225 1849
rect 19259 1815 19298 1849
rect 19332 1815 19371 1849
rect 19405 1815 19444 1849
rect 19478 1815 19517 1849
rect 19551 1815 19585 1849
rect 19185 1782 19585 1815
rect 9716 1754 9750 1762
rect 9784 1754 9819 1762
rect 9853 1754 9888 1762
rect 9922 1754 9957 1762
rect 9716 1720 9734 1754
rect 9784 1728 9808 1754
rect 9853 1728 9882 1754
rect 9922 1728 9956 1754
rect 9991 1728 10026 1762
rect 10060 1754 10095 1762
rect 10129 1754 10164 1762
rect 10198 1754 10233 1762
rect 10267 1754 10302 1762
rect 10336 1754 10371 1762
rect 10405 1754 10440 1762
rect 10474 1754 10509 1762
rect 10064 1728 10095 1754
rect 10138 1728 10164 1754
rect 10212 1728 10233 1754
rect 10286 1728 10302 1754
rect 10360 1728 10371 1754
rect 10434 1728 10440 1754
rect 10507 1728 10509 1754
rect 10543 1754 10578 1762
rect 10612 1754 10647 1762
rect 10681 1754 10716 1762
rect 10750 1754 10785 1762
rect 10819 1754 10854 1762
rect 10888 1754 10923 1762
rect 10957 1754 10992 1762
rect 11026 1754 11061 1762
rect 10543 1728 10546 1754
rect 10612 1728 10619 1754
rect 10681 1728 10692 1754
rect 10750 1728 10765 1754
rect 10819 1728 10838 1754
rect 10888 1728 10911 1754
rect 10957 1728 10984 1754
rect 11026 1728 11057 1754
rect 11095 1728 11130 1762
rect 11164 1728 11199 1762
rect 11233 1754 11268 1762
rect 11302 1754 11337 1762
rect 11371 1754 11406 1762
rect 11440 1754 11475 1762
rect 11509 1754 11544 1762
rect 11578 1754 11613 1762
rect 11647 1754 11682 1762
rect 11716 1754 11751 1762
rect 11237 1728 11268 1754
rect 11310 1728 11337 1754
rect 11383 1728 11406 1754
rect 11456 1728 11475 1754
rect 11529 1728 11544 1754
rect 11602 1728 11613 1754
rect 11675 1728 11682 1754
rect 11748 1728 11751 1754
rect 11785 1754 11820 1762
rect 11854 1754 11889 1762
rect 11923 1754 11958 1762
rect 11992 1754 12027 1762
rect 12061 1754 12096 1762
rect 12130 1754 12165 1762
rect 12199 1754 12234 1762
rect 12268 1754 12303 1762
rect 12337 1754 12372 1762
rect 11785 1728 11787 1754
rect 11854 1728 11860 1754
rect 11923 1728 11933 1754
rect 11992 1728 12006 1754
rect 12061 1728 12079 1754
rect 12130 1728 12152 1754
rect 12199 1728 12225 1754
rect 12268 1728 12298 1754
rect 12337 1728 12371 1754
rect 12406 1728 12441 1762
rect 12475 1728 12510 1762
rect 12544 1728 12579 1762
rect 12613 1728 12648 1762
rect 12682 1728 12717 1762
rect 12751 1728 12786 1762
rect 12820 1728 12855 1762
rect 12889 1728 12924 1762
rect 12958 1728 12993 1762
rect 19011 1775 19585 1782
rect 19011 1741 19079 1775
rect 19113 1741 19152 1775
rect 19186 1741 19225 1775
rect 19259 1741 19298 1775
rect 19332 1741 19371 1775
rect 19405 1741 19444 1775
rect 19478 1741 19517 1775
rect 19551 1741 19585 1775
rect 19011 1730 19585 1741
rect 9768 1720 9808 1728
rect 9842 1720 9882 1728
rect 9916 1720 9956 1728
rect 9990 1720 10030 1728
rect 10064 1720 10104 1728
rect 10138 1720 10178 1728
rect 10212 1720 10252 1728
rect 10286 1720 10326 1728
rect 10360 1720 10400 1728
rect 10434 1720 10473 1728
rect 10507 1720 10546 1728
rect 10580 1720 10619 1728
rect 10653 1720 10692 1728
rect 10726 1720 10765 1728
rect 10799 1720 10838 1728
rect 10872 1720 10911 1728
rect 10945 1720 10984 1728
rect 11018 1720 11057 1728
rect 11091 1720 11130 1728
rect 11164 1720 11203 1728
rect 11237 1720 11276 1728
rect 11310 1720 11349 1728
rect 11383 1720 11422 1728
rect 11456 1720 11495 1728
rect 11529 1720 11568 1728
rect 11602 1720 11641 1728
rect 11675 1720 11714 1728
rect 11748 1720 11787 1728
rect 11821 1720 11860 1728
rect 11894 1720 11933 1728
rect 11967 1720 12006 1728
rect 12040 1720 12079 1728
rect 12113 1720 12152 1728
rect 12186 1720 12225 1728
rect 12259 1720 12298 1728
rect 12332 1720 12371 1728
rect 12405 1720 12993 1728
rect 9716 1694 12993 1720
rect 19041 1696 19079 1730
rect 19113 1696 19151 1730
rect 19185 1701 19585 1730
rect 9716 1672 9750 1694
rect 9784 1672 9819 1694
rect 9853 1672 9888 1694
rect 9922 1672 9957 1694
rect 9716 1638 9734 1672
rect 9784 1660 9808 1672
rect 9853 1660 9882 1672
rect 9922 1660 9956 1672
rect 9991 1660 10026 1694
rect 10060 1672 10095 1694
rect 10129 1672 10164 1694
rect 10198 1672 10233 1694
rect 10267 1672 10302 1694
rect 10336 1672 10371 1694
rect 10405 1672 10440 1694
rect 10474 1672 10509 1694
rect 10064 1660 10095 1672
rect 10138 1660 10164 1672
rect 10212 1660 10233 1672
rect 10286 1660 10302 1672
rect 10360 1660 10371 1672
rect 10434 1660 10440 1672
rect 10507 1660 10509 1672
rect 10543 1672 10578 1694
rect 10612 1672 10647 1694
rect 10681 1672 10716 1694
rect 10750 1672 10785 1694
rect 10819 1672 10854 1694
rect 10888 1672 10923 1694
rect 10957 1672 10992 1694
rect 11026 1672 11061 1694
rect 10543 1660 10546 1672
rect 10612 1660 10619 1672
rect 10681 1660 10692 1672
rect 10750 1660 10765 1672
rect 10819 1660 10838 1672
rect 10888 1660 10911 1672
rect 10957 1660 10984 1672
rect 11026 1660 11057 1672
rect 11095 1660 11130 1694
rect 11164 1660 11199 1694
rect 11233 1672 11268 1694
rect 11302 1672 11337 1694
rect 11371 1672 11406 1694
rect 11440 1672 11475 1694
rect 11509 1672 11544 1694
rect 11578 1672 11613 1694
rect 11647 1672 11682 1694
rect 11716 1672 11751 1694
rect 11237 1660 11268 1672
rect 11310 1660 11337 1672
rect 11383 1660 11406 1672
rect 11456 1660 11475 1672
rect 11529 1660 11544 1672
rect 11602 1660 11613 1672
rect 11675 1660 11682 1672
rect 11748 1660 11751 1672
rect 11785 1672 11820 1694
rect 11854 1672 11889 1694
rect 11923 1672 11958 1694
rect 11992 1672 12027 1694
rect 12061 1672 12096 1694
rect 12130 1672 12165 1694
rect 12199 1672 12234 1694
rect 12268 1672 12303 1694
rect 12337 1672 12372 1694
rect 11785 1660 11787 1672
rect 11854 1660 11860 1672
rect 11923 1660 11933 1672
rect 11992 1660 12006 1672
rect 12061 1660 12079 1672
rect 12130 1660 12152 1672
rect 12199 1660 12225 1672
rect 12268 1660 12298 1672
rect 12337 1660 12371 1672
rect 12406 1660 12441 1694
rect 12475 1660 12510 1694
rect 12544 1660 12579 1694
rect 12613 1660 12648 1694
rect 12682 1660 12717 1694
rect 12751 1660 12786 1694
rect 12820 1660 12855 1694
rect 12889 1660 12924 1694
rect 12958 1660 12993 1694
rect 9768 1638 9808 1660
rect 9842 1638 9882 1660
rect 9916 1638 9956 1660
rect 9990 1638 10030 1660
rect 10064 1638 10104 1660
rect 10138 1638 10178 1660
rect 10212 1638 10252 1660
rect 10286 1638 10326 1660
rect 10360 1638 10400 1660
rect 10434 1638 10473 1660
rect 10507 1638 10546 1660
rect 10580 1638 10619 1660
rect 10653 1638 10692 1660
rect 10726 1638 10765 1660
rect 10799 1638 10838 1660
rect 10872 1638 10911 1660
rect 10945 1638 10984 1660
rect 11018 1638 11057 1660
rect 11091 1638 11130 1660
rect 11164 1638 11203 1660
rect 11237 1638 11276 1660
rect 11310 1638 11349 1660
rect 11383 1638 11422 1660
rect 11456 1638 11495 1660
rect 11529 1638 11568 1660
rect 11602 1638 11641 1660
rect 11675 1638 11714 1660
rect 11748 1638 11787 1660
rect 11821 1638 11860 1660
rect 11894 1638 11933 1660
rect 11967 1638 12006 1660
rect 12040 1638 12079 1660
rect 12113 1638 12152 1660
rect 12186 1638 12225 1660
rect 12259 1638 12298 1660
rect 12332 1638 12371 1660
rect 12405 1638 12993 1660
rect 19011 1667 19079 1696
rect 19113 1667 19152 1696
rect 19186 1667 19225 1701
rect 19259 1667 19298 1701
rect 19332 1667 19371 1701
rect 19405 1667 19444 1701
rect 19478 1667 19517 1701
rect 19551 1667 19585 1701
rect 19011 1644 19585 1667
rect 9716 1626 12993 1638
rect 9716 1592 9750 1626
rect 9784 1592 9819 1626
rect 9853 1592 9888 1626
rect 9922 1592 9957 1626
rect 9991 1592 10026 1626
rect 10060 1592 10095 1626
rect 10129 1592 10164 1626
rect 10198 1592 10233 1626
rect 10267 1592 10302 1626
rect 10336 1592 10371 1626
rect 10405 1592 10440 1626
rect 10474 1592 10509 1626
rect 10543 1592 10578 1626
rect 10612 1592 10647 1626
rect 10681 1592 10716 1626
rect 10750 1592 10785 1626
rect 10819 1592 10854 1626
rect 10888 1592 10923 1626
rect 10957 1592 10992 1626
rect 11026 1592 11061 1626
rect 11095 1592 11130 1626
rect 11164 1592 11199 1626
rect 11233 1592 11268 1626
rect 11302 1592 11337 1626
rect 11371 1592 11406 1626
rect 11440 1592 11475 1626
rect 11509 1592 11544 1626
rect 11578 1592 11613 1626
rect 11647 1592 11682 1626
rect 11716 1592 11751 1626
rect 11785 1592 11820 1626
rect 11854 1592 11889 1626
rect 11923 1592 11958 1626
rect 11992 1592 12027 1626
rect 12061 1592 12096 1626
rect 12130 1592 12165 1626
rect 12199 1592 12234 1626
rect 12268 1592 12303 1626
rect 12337 1592 12372 1626
rect 12406 1592 12441 1626
rect 12475 1592 12510 1626
rect 12544 1592 12579 1626
rect 12613 1592 12648 1626
rect 12682 1592 12717 1626
rect 12751 1592 12786 1626
rect 12820 1592 12855 1626
rect 12889 1592 12924 1626
rect 12958 1592 12993 1626
rect 19041 1610 19079 1644
rect 19113 1610 19151 1644
rect 19185 1627 19585 1644
rect 19011 1593 19079 1610
rect 19113 1593 19152 1610
rect 19186 1593 19225 1627
rect 19259 1593 19298 1627
rect 19332 1593 19371 1627
rect 19405 1593 19444 1627
rect 19478 1593 19517 1627
rect 19551 1593 19585 1627
rect 19011 1592 19585 1593
rect 19967 1878 20042 1924
rect 19967 1846 20013 1878
rect 19967 1812 19973 1846
rect 20007 1812 20013 1846
rect 19967 1768 20013 1812
rect 25343 1794 25381 1828
rect 28031 1795 28065 1829
rect 19967 1734 19973 1768
rect 20007 1734 20013 1768
rect 25787 1761 25821 1785
rect 19967 1690 20013 1734
rect 19967 1656 19973 1690
rect 20007 1656 20013 1690
rect 25413 1674 25471 1740
rect 19967 1612 20013 1656
rect 9405 1525 9411 1592
rect 9445 1525 9451 1592
rect 9734 1590 12405 1592
rect 9768 1556 9808 1590
rect 9842 1556 9882 1590
rect 9916 1556 9956 1590
rect 9990 1556 10030 1590
rect 10064 1556 10104 1590
rect 10138 1556 10178 1590
rect 10212 1556 10252 1590
rect 10286 1556 10326 1590
rect 10360 1556 10400 1590
rect 10434 1556 10473 1590
rect 10507 1556 10546 1590
rect 10580 1556 10619 1590
rect 10653 1556 10692 1590
rect 10726 1556 10765 1590
rect 10799 1556 10838 1590
rect 10872 1556 10911 1590
rect 10945 1556 10984 1590
rect 11018 1556 11057 1590
rect 11091 1556 11130 1590
rect 11164 1556 11203 1590
rect 11237 1556 11276 1590
rect 11310 1556 11349 1590
rect 11383 1556 11422 1590
rect 11456 1556 11495 1590
rect 11529 1556 11568 1590
rect 11602 1556 11641 1590
rect 11675 1556 11714 1590
rect 11748 1556 11787 1590
rect 11821 1556 11860 1590
rect 11894 1556 11933 1590
rect 11967 1556 12006 1590
rect 12040 1556 12079 1590
rect 12113 1556 12152 1590
rect 12186 1556 12225 1590
rect 12259 1556 12298 1590
rect 12332 1556 12371 1590
rect 9734 1553 12405 1556
rect 19967 1578 19973 1612
rect 20007 1578 20013 1612
rect 9405 1513 9451 1525
rect 2470 1395 2492 1429
rect 2538 1395 2564 1429
rect 2606 1395 2636 1429
rect 2674 1395 2708 1429
rect 2742 1395 2776 1429
rect 2814 1395 2844 1429
rect 2886 1395 2912 1429
rect 2958 1395 2980 1429
rect 3030 1395 3048 1429
rect 3102 1395 3116 1429
rect 3174 1395 3184 1429
rect 3246 1395 3252 1429
rect 3318 1395 3320 1429
rect 3354 1395 3356 1429
rect 3422 1395 3428 1429
rect 3490 1395 3500 1429
rect 3558 1395 3572 1429
rect 3626 1395 3644 1429
rect 3694 1395 3716 1429
rect 3762 1395 3788 1429
rect 3830 1395 3860 1429
rect 3898 1395 3932 1429
rect 3966 1395 4000 1429
rect 4038 1395 4068 1429
rect 4110 1395 4136 1429
rect 4182 1395 4204 1429
rect 4254 1395 4272 1429
rect 4326 1395 4340 1429
rect 7469 1439 7485 1473
rect 7545 1439 7562 1473
rect 7596 1439 7601 1473
rect 7635 1439 7639 1473
rect 7673 1439 7691 1473
rect 7750 1439 7781 1473
rect 7827 1439 7843 1473
rect 9405 1457 9411 1513
rect 9445 1457 9451 1513
rect 9405 1434 9451 1457
rect 2145 1368 2191 1377
rect 466 1289 500 1327
rect 2145 1309 2151 1368
rect 2185 1309 2191 1368
rect 2145 1294 2191 1309
rect 466 1217 500 1255
rect 620 1245 642 1279
rect 688 1245 714 1279
rect 756 1245 786 1279
rect 824 1245 858 1279
rect 892 1245 926 1279
rect 964 1245 994 1279
rect 1036 1245 1062 1279
rect 1108 1245 1130 1279
rect 1180 1245 1198 1279
rect 1252 1245 1266 1279
rect 1324 1245 1334 1279
rect 1396 1245 1402 1279
rect 1468 1245 1470 1279
rect 1504 1245 1506 1279
rect 2145 1241 2151 1294
rect 2185 1241 2191 1294
rect 466 1145 500 1183
rect 1622 1218 1656 1234
rect 1622 1123 1656 1170
rect 466 1073 500 1111
rect 620 1089 642 1123
rect 688 1089 714 1123
rect 756 1089 786 1123
rect 824 1089 858 1123
rect 892 1089 926 1123
rect 964 1089 994 1123
rect 1036 1089 1062 1123
rect 1108 1089 1130 1123
rect 1180 1089 1198 1123
rect 1252 1089 1266 1123
rect 1324 1089 1334 1123
rect 1396 1089 1402 1123
rect 1468 1089 1470 1123
rect 1504 1089 1506 1123
rect 466 1001 500 1039
rect 1622 1033 1656 1085
rect 1622 978 1656 994
rect 2145 1220 2191 1241
rect 2145 1173 2151 1220
rect 2185 1173 2191 1220
rect 4472 1392 4506 1427
rect 4746 1395 4760 1429
rect 4814 1395 4832 1429
rect 4882 1395 4904 1429
rect 4950 1395 4976 1429
rect 5018 1395 5048 1429
rect 5086 1395 5120 1429
rect 5154 1395 5188 1429
rect 5226 1395 5256 1429
rect 5298 1395 5324 1429
rect 5370 1395 5392 1429
rect 5442 1395 5460 1429
rect 5514 1395 5528 1429
rect 5586 1395 5596 1429
rect 5658 1395 5664 1429
rect 5730 1395 5732 1429
rect 5766 1395 5768 1429
rect 5834 1395 5840 1429
rect 5902 1395 5912 1429
rect 5970 1395 5984 1429
rect 6038 1395 6056 1429
rect 6106 1395 6128 1429
rect 6174 1395 6200 1429
rect 6242 1395 6272 1429
rect 6310 1395 6344 1429
rect 6378 1395 6412 1429
rect 6450 1395 6480 1429
rect 6522 1395 6548 1429
rect 6594 1395 6616 1429
rect 9405 1389 9411 1434
rect 9445 1389 9451 1434
rect 4506 1368 4614 1384
rect 4506 1358 4580 1368
rect 4472 1355 4580 1358
rect 4472 1323 4486 1355
rect 4520 1321 4558 1355
rect 4592 1321 4614 1334
rect 4506 1289 4614 1321
rect 4472 1273 4614 1289
rect 4472 1254 4486 1273
rect 4520 1239 4558 1273
rect 4592 1254 4614 1273
rect 4506 1220 4580 1239
rect 4472 1204 4614 1220
rect 7424 1329 7458 1355
rect 7424 1261 7458 1283
rect 7424 1193 7458 1211
rect 2145 1146 2191 1173
rect 2470 1159 2492 1193
rect 2538 1159 2564 1193
rect 2606 1159 2636 1193
rect 2674 1159 2708 1193
rect 2742 1159 2776 1193
rect 2814 1159 2844 1193
rect 2886 1159 2912 1193
rect 2958 1159 2980 1193
rect 3030 1159 3048 1193
rect 3102 1159 3116 1193
rect 3174 1159 3184 1193
rect 3246 1159 3252 1193
rect 3318 1159 3320 1193
rect 3354 1159 3356 1193
rect 3422 1159 3428 1193
rect 3490 1159 3500 1193
rect 3558 1159 3572 1193
rect 3626 1159 3644 1193
rect 3694 1159 3716 1193
rect 3762 1159 3788 1193
rect 3830 1159 3860 1193
rect 3898 1159 3932 1193
rect 3966 1159 4000 1193
rect 4038 1159 4068 1193
rect 4110 1159 4136 1193
rect 4182 1159 4204 1193
rect 4254 1159 4272 1193
rect 4326 1159 4340 1193
rect 4746 1159 4760 1193
rect 4814 1159 4832 1193
rect 4882 1159 4904 1193
rect 4950 1159 4976 1193
rect 5018 1159 5048 1193
rect 5086 1159 5120 1193
rect 5154 1159 5188 1193
rect 5226 1159 5256 1193
rect 5298 1159 5324 1193
rect 5370 1159 5392 1193
rect 5442 1159 5460 1193
rect 5514 1159 5528 1193
rect 5586 1159 5596 1193
rect 5658 1159 5664 1193
rect 5730 1159 5732 1193
rect 5766 1159 5768 1193
rect 5834 1159 5840 1193
rect 5902 1159 5912 1193
rect 5970 1159 5984 1193
rect 6038 1159 6056 1193
rect 6106 1159 6128 1193
rect 6174 1159 6200 1193
rect 6242 1159 6272 1193
rect 6310 1159 6344 1193
rect 6378 1159 6412 1193
rect 6450 1159 6480 1193
rect 6522 1159 6548 1193
rect 6594 1159 6616 1193
rect 2145 1105 2151 1146
rect 2185 1105 2191 1146
rect 2145 1072 2191 1105
rect 7424 1125 7458 1139
rect 2145 1037 2151 1072
rect 2185 1037 2191 1072
rect 2451 1064 2466 1098
rect 2501 1064 2539 1098
rect 2583 1064 2611 1098
rect 2666 1064 2683 1098
rect 2749 1064 2755 1098
rect 2789 1064 2797 1098
rect 2861 1064 2879 1098
rect 2932 1064 2961 1098
rect 3003 1064 3019 1098
rect 3075 1064 3091 1098
rect 3128 1064 3162 1098
rect 3211 1064 3233 1098
rect 3293 1064 3305 1098
rect 3339 1064 3341 1098
rect 3375 1064 3377 1098
rect 3411 1064 3423 1098
rect 3483 1064 3505 1098
rect 3555 1064 3587 1098
rect 3627 1064 3643 1098
rect 3823 1064 3839 1098
rect 3876 1064 3933 1098
rect 3968 1064 4023 1098
rect 4063 1064 4079 1098
rect 4135 1097 4151 1098
rect 4135 1064 4147 1097
rect 4185 1064 4246 1098
rect 4280 1097 4341 1098
rect 4375 1097 4391 1098
rect 4286 1064 4341 1097
rect 4181 1063 4252 1064
rect 4286 1063 4357 1064
rect 4447 1064 4463 1098
rect 4497 1064 4547 1098
rect 2145 1003 2191 1037
rect 466 929 500 967
rect 620 933 642 967
rect 688 933 714 967
rect 756 933 786 967
rect 824 933 858 967
rect 892 933 926 967
rect 964 933 994 967
rect 1036 933 1062 967
rect 1108 933 1130 967
rect 1180 933 1198 967
rect 1252 933 1266 967
rect 1324 933 1334 967
rect 1396 933 1402 967
rect 1468 933 1470 967
rect 1504 933 1506 967
rect 2145 964 2151 1003
rect 2185 964 2191 1003
rect 4447 982 4547 1064
rect 4603 1097 4619 1098
rect 4653 1097 4714 1098
rect 4653 1064 4677 1097
rect 4637 1063 4677 1064
rect 4711 1064 4714 1097
rect 4748 1097 4809 1098
rect 4843 1097 4859 1098
rect 4748 1064 4751 1097
rect 4711 1063 4751 1064
rect 4785 1064 4809 1097
rect 4785 1063 4825 1064
rect 4915 1064 4931 1098
rect 4965 1064 5015 1098
rect 4915 982 5015 1064
rect 5071 1097 5087 1098
rect 5121 1097 5157 1098
rect 5191 1097 5226 1098
rect 5260 1097 5295 1098
rect 5329 1097 5364 1098
rect 5121 1064 5144 1097
rect 5191 1064 5217 1097
rect 5260 1064 5289 1097
rect 5329 1064 5361 1097
rect 5398 1064 5433 1098
rect 5467 1064 5483 1098
rect 5713 1064 5729 1098
rect 5764 1064 5807 1098
rect 5858 1064 5884 1098
rect 5918 1064 5919 1098
rect 5953 1064 5969 1098
rect 6025 1064 6041 1098
rect 6075 1064 6136 1098
rect 6170 1064 6226 1098
rect 6265 1064 6298 1098
rect 6445 1096 6461 1098
rect 6495 1096 6544 1098
rect 6578 1096 6627 1098
rect 6495 1064 6516 1096
rect 6578 1064 6590 1096
rect 5105 1063 5144 1064
rect 5178 1063 5217 1064
rect 5251 1063 5289 1064
rect 5323 1063 5361 1064
rect 5395 1063 5433 1064
rect 6476 1062 6516 1064
rect 6550 1062 6590 1064
rect 6624 1064 6627 1096
rect 6661 1096 6709 1098
rect 6743 1096 6791 1098
rect 6661 1064 6663 1096
rect 6624 1062 6663 1064
rect 6697 1064 6709 1096
rect 6770 1064 6791 1096
rect 6825 1064 6841 1098
rect 6897 1064 6913 1098
rect 6947 1090 6983 1098
rect 6959 1064 6983 1090
rect 7017 1064 7033 1098
rect 6697 1062 6736 1064
rect 6925 1014 6959 1056
rect 2145 935 2191 964
rect 1622 895 1724 922
rect 466 857 500 895
rect 1427 889 1724 895
rect 1461 855 1499 889
rect 1533 872 1724 889
rect 1533 855 1622 872
rect 1427 849 1622 855
rect 466 785 500 823
rect 1656 838 1690 872
rect 1622 822 1724 838
rect 2145 890 2151 935
rect 2185 890 2191 935
rect 2145 867 2191 890
rect 2145 816 2151 867
rect 2185 816 2191 867
rect 620 777 642 811
rect 688 777 714 811
rect 756 777 786 811
rect 824 777 858 811
rect 892 777 926 811
rect 964 777 994 811
rect 1036 777 1062 811
rect 1108 777 1130 811
rect 1180 777 1198 811
rect 1252 777 1266 811
rect 1324 777 1334 811
rect 1396 777 1402 811
rect 1468 777 1470 811
rect 1504 777 1506 811
rect 2145 799 2191 816
rect 466 713 500 751
rect 466 641 500 679
rect 1622 750 1656 766
rect 1622 655 1656 702
rect 620 621 642 655
rect 688 621 714 655
rect 756 621 786 655
rect 824 621 858 655
rect 892 621 926 655
rect 964 621 994 655
rect 1036 621 1062 655
rect 1108 621 1130 655
rect 1180 621 1198 655
rect 1252 621 1266 655
rect 1324 621 1334 655
rect 1396 621 1402 655
rect 1468 621 1470 655
rect 1504 621 1506 655
rect 466 569 500 607
rect 466 497 500 535
rect 1622 560 1656 606
rect 2145 742 2151 799
rect 2185 742 2191 799
rect 2145 731 2191 742
rect 2145 668 2151 731
rect 2185 668 2191 731
rect 2145 663 2191 668
rect 2145 629 2151 663
rect 2185 629 2191 663
rect 2145 628 2191 629
rect 2145 561 2151 628
rect 2185 561 2191 628
rect 2145 554 2191 561
rect 620 465 642 499
rect 688 465 714 499
rect 756 465 786 499
rect 824 465 858 499
rect 892 465 926 499
rect 964 465 994 499
rect 1036 465 1062 499
rect 1108 465 1130 499
rect 1180 465 1198 499
rect 1252 465 1266 499
rect 1324 465 1334 499
rect 1396 465 1402 499
rect 1468 465 1470 499
rect 1504 465 1506 499
rect 2145 493 2151 554
rect 2185 493 2191 554
rect 2145 480 2191 493
rect 466 425 500 463
rect 1622 427 1724 454
rect 466 353 500 391
rect 1427 421 1724 427
rect 1461 387 1499 421
rect 1533 404 1724 421
rect 1533 387 1622 404
rect 1427 381 1622 387
rect 1656 370 1690 404
rect 1622 354 1724 370
rect 2145 425 2151 480
rect 2185 425 2191 480
rect 2145 406 2191 425
rect 2145 357 2151 406
rect 2185 357 2191 406
rect 466 281 500 319
rect 620 309 642 343
rect 688 309 714 343
rect 756 309 786 343
rect 824 309 858 343
rect 892 309 926 343
rect 964 309 994 343
rect 1036 309 1062 343
rect 1108 309 1130 343
rect 1180 309 1198 343
rect 1252 309 1266 343
rect 1324 309 1334 343
rect 1396 309 1402 343
rect 1468 309 1470 343
rect 1504 309 1506 343
rect 2145 332 2191 357
rect 466 209 500 247
rect 1622 282 1656 298
rect 1622 187 1656 234
rect 466 137 500 175
rect 620 153 642 187
rect 688 153 714 187
rect 756 153 786 187
rect 824 153 858 187
rect 892 153 926 187
rect 964 153 994 187
rect 1036 153 1062 187
rect 1108 153 1130 187
rect 1180 153 1198 187
rect 1252 153 1266 187
rect 1324 153 1334 187
rect 1396 153 1402 187
rect 1468 153 1470 187
rect 1504 153 1506 187
rect 466 65 500 103
rect 1622 92 1656 138
rect 2145 289 2151 332
rect 2185 289 2191 332
rect 2145 258 2191 289
rect 2145 221 2151 258
rect 2185 221 2191 258
rect 2145 187 2191 221
rect 2145 150 2151 187
rect 2185 150 2191 187
rect 2145 119 2191 150
rect 2145 76 2151 119
rect 2185 76 2191 119
rect 2145 51 2191 76
rect 466 -7 500 31
rect 620 -3 642 31
rect 688 -3 714 31
rect 756 -3 786 31
rect 824 -3 858 31
rect 892 -3 926 31
rect 964 -3 994 31
rect 1036 -3 1062 31
rect 1108 -3 1130 31
rect 1180 -3 1198 31
rect 1252 -3 1266 31
rect 1324 -3 1334 31
rect 1396 -3 1402 31
rect 1468 -3 1470 31
rect 1504 -3 1506 31
rect 2145 2 2151 51
rect 2185 2 2191 51
rect 2406 946 2440 948
rect 2406 910 2440 912
rect 2406 838 2440 844
rect 2406 766 2440 776
rect 2406 694 2440 708
rect 2406 622 2440 640
rect 2406 550 2440 572
rect 2406 478 2440 504
rect 2406 406 2440 436
rect 2406 334 2440 368
rect 2406 266 2440 300
rect 2406 198 2440 228
rect 2406 130 2440 156
rect 2406 62 2440 84
rect 2562 946 2596 948
rect 2562 910 2596 912
rect 2562 838 2596 844
rect 2562 766 2596 776
rect 2562 694 2596 708
rect 2562 622 2596 640
rect 2562 550 2596 572
rect 2562 478 2596 504
rect 2562 406 2596 436
rect 2562 334 2596 368
rect 2562 266 2596 300
rect 2562 198 2596 228
rect 2562 130 2596 156
rect 2562 62 2596 84
rect 2718 946 2752 948
rect 2718 910 2752 912
rect 2718 838 2752 844
rect 2718 766 2752 776
rect 2718 694 2752 708
rect 2718 622 2752 640
rect 2718 550 2752 572
rect 2718 478 2752 504
rect 2718 406 2752 436
rect 2718 334 2752 368
rect 2718 266 2752 300
rect 2718 198 2752 228
rect 2718 130 2752 156
rect 2718 62 2752 84
rect 2874 946 2908 948
rect 2874 910 2908 912
rect 2874 838 2908 844
rect 2874 766 2908 776
rect 2874 694 2908 708
rect 2874 622 2908 640
rect 2874 550 2908 572
rect 2874 478 2908 504
rect 2874 406 2908 436
rect 2874 334 2908 368
rect 2874 266 2908 300
rect 2874 198 2908 228
rect 2874 130 2908 156
rect 2874 62 2908 84
rect 3030 946 3064 948
rect 3030 910 3064 912
rect 3030 838 3064 844
rect 3030 766 3064 776
rect 3030 694 3064 708
rect 3030 622 3064 640
rect 3030 550 3064 572
rect 3030 478 3064 504
rect 3030 406 3064 436
rect 3030 334 3064 368
rect 3030 266 3064 300
rect 3030 198 3064 228
rect 3030 130 3064 156
rect 3030 62 3064 84
rect 3186 946 3220 948
rect 3186 910 3220 912
rect 3186 838 3220 844
rect 3186 766 3220 776
rect 3186 694 3220 708
rect 3186 622 3220 640
rect 3186 550 3220 572
rect 3186 478 3220 504
rect 3186 406 3220 436
rect 3186 334 3220 368
rect 3186 266 3220 300
rect 3186 198 3220 228
rect 3186 130 3220 156
rect 3186 62 3220 84
rect 3342 946 3376 948
rect 3342 910 3376 912
rect 3342 838 3376 844
rect 3342 766 3376 776
rect 3342 694 3376 708
rect 3342 622 3376 640
rect 3342 550 3376 572
rect 3342 478 3376 504
rect 3342 406 3376 436
rect 3342 334 3376 368
rect 3342 266 3376 300
rect 3342 198 3376 228
rect 3342 130 3376 156
rect 3342 62 3376 84
rect 3498 946 3532 948
rect 3498 910 3532 912
rect 3498 838 3532 844
rect 3498 766 3532 776
rect 3498 694 3532 708
rect 3498 622 3532 640
rect 3498 550 3532 572
rect 3498 478 3532 504
rect 3498 406 3532 436
rect 3498 334 3532 368
rect 3498 266 3532 300
rect 3498 198 3532 228
rect 3498 130 3532 156
rect 3498 62 3532 84
rect 3654 946 3688 948
rect 3654 910 3688 912
rect 3654 838 3688 844
rect 3654 766 3688 776
rect 3654 694 3688 708
rect 3654 622 3688 640
rect 3654 550 3688 572
rect 3654 478 3688 504
rect 3654 406 3688 436
rect 3654 334 3688 368
rect 3654 266 3688 300
rect 3654 198 3688 228
rect 3654 130 3688 156
rect 3654 62 3688 84
rect 3778 946 3812 948
rect 3778 910 3812 912
rect 3778 838 3812 844
rect 3778 766 3812 776
rect 3778 694 3812 708
rect 3778 622 3812 640
rect 3778 550 3812 572
rect 3778 478 3812 504
rect 3778 406 3812 436
rect 3778 334 3812 368
rect 3778 266 3812 300
rect 3778 198 3812 228
rect 3778 130 3812 156
rect 3778 62 3812 84
rect 3934 946 3968 948
rect 3934 910 3968 912
rect 3934 838 3968 844
rect 3934 766 3968 776
rect 3934 694 3968 708
rect 3934 622 3968 640
rect 3934 550 3968 572
rect 3934 478 3968 504
rect 3934 406 3968 436
rect 3934 334 3968 368
rect 3934 266 3968 300
rect 3934 198 3968 228
rect 3934 130 3968 156
rect 3934 62 3968 84
rect 4090 946 4124 948
rect 4090 910 4124 912
rect 4090 838 4124 844
rect 4090 766 4124 776
rect 4090 694 4124 708
rect 4090 622 4124 640
rect 4090 550 4124 572
rect 4090 478 4124 504
rect 4090 406 4124 436
rect 4090 334 4124 368
rect 4090 266 4124 300
rect 4090 198 4124 228
rect 4090 130 4124 156
rect 4090 62 4124 84
rect 4246 946 4280 948
rect 4246 910 4280 912
rect 4246 838 4280 844
rect 4246 766 4280 776
rect 4246 694 4280 708
rect 4246 622 4280 640
rect 4246 550 4280 572
rect 4246 478 4280 504
rect 4246 406 4280 436
rect 4246 334 4280 368
rect 4246 266 4280 300
rect 4246 198 4280 228
rect 4246 130 4280 156
rect 4246 62 4280 84
rect 4436 948 4558 982
rect 4402 946 4592 948
rect 4436 912 4558 946
rect 4402 910 4592 912
rect 4436 844 4558 910
rect 4402 838 4592 844
rect 4436 776 4558 838
rect 4402 766 4592 776
rect 4436 708 4558 766
rect 4402 694 4592 708
rect 4436 640 4558 694
rect 4402 622 4592 640
rect 4436 572 4558 622
rect 4402 550 4592 572
rect 4436 504 4558 550
rect 4402 478 4592 504
rect 4436 436 4558 478
rect 4402 406 4592 436
rect 4436 368 4558 406
rect 4402 334 4592 368
rect 4436 300 4558 334
rect 4402 266 4592 300
rect 4436 228 4558 266
rect 4402 198 4592 228
rect 4436 156 4558 198
rect 4402 130 4592 156
rect 4436 84 4558 130
rect 4402 62 4592 84
rect 4436 12 4558 62
rect 4714 946 4748 948
rect 4714 910 4748 912
rect 4714 838 4748 844
rect 4714 766 4748 776
rect 4714 694 4748 708
rect 4714 622 4748 640
rect 4714 550 4748 572
rect 4714 478 4748 504
rect 4714 406 4748 436
rect 4714 334 4748 368
rect 4714 266 4748 300
rect 4714 198 4748 228
rect 4714 130 4748 156
rect 4714 62 4748 84
rect 4904 948 5026 982
rect 4870 946 5060 948
rect 4904 912 5026 946
rect 4870 910 5060 912
rect 4904 844 5026 910
rect 4870 838 5060 844
rect 4904 776 5026 838
rect 4870 766 5060 776
rect 4904 708 5026 766
rect 4870 694 5060 708
rect 4904 640 5026 694
rect 4870 622 5060 640
rect 4904 572 5026 622
rect 4870 550 5060 572
rect 4904 504 5026 550
rect 4870 478 5060 504
rect 4904 436 5026 478
rect 4870 406 5060 436
rect 4904 368 5026 406
rect 4870 334 5060 368
rect 4904 300 5026 334
rect 4870 266 5060 300
rect 4904 228 5026 266
rect 4870 198 5060 228
rect 4904 156 5026 198
rect 4870 130 5060 156
rect 4904 84 5026 130
rect 4870 62 5060 84
rect 4904 12 5026 62
rect 5182 946 5216 948
rect 5182 910 5216 912
rect 5182 838 5216 844
rect 5182 766 5216 776
rect 5182 694 5216 708
rect 5182 622 5216 640
rect 5182 550 5216 572
rect 5182 478 5216 504
rect 5182 406 5216 436
rect 5182 334 5216 368
rect 5182 266 5216 300
rect 5182 198 5216 228
rect 5182 130 5216 156
rect 5182 62 5216 84
rect 5338 946 5372 948
rect 5338 910 5372 912
rect 5338 838 5372 844
rect 5338 766 5372 776
rect 5338 694 5372 708
rect 5338 622 5372 640
rect 5338 550 5372 572
rect 5338 478 5372 504
rect 5338 406 5372 436
rect 5338 334 5372 368
rect 5338 266 5372 300
rect 5338 198 5372 228
rect 5338 130 5372 156
rect 5338 62 5372 84
rect 5494 946 5528 948
rect 5494 910 5528 912
rect 5494 838 5528 844
rect 5494 766 5528 776
rect 5494 694 5528 708
rect 5494 622 5528 640
rect 5494 550 5528 572
rect 5494 478 5528 504
rect 5494 406 5528 436
rect 5494 334 5528 368
rect 5494 266 5528 300
rect 5494 198 5528 228
rect 5494 130 5528 156
rect 5494 62 5528 84
rect 5668 946 5702 948
rect 5668 910 5702 912
rect 5668 838 5702 844
rect 5668 766 5702 776
rect 5668 694 5702 708
rect 5668 622 5702 640
rect 5668 550 5702 572
rect 5668 478 5702 504
rect 5668 406 5702 436
rect 5668 334 5702 368
rect 5668 266 5702 300
rect 5668 198 5702 228
rect 5668 130 5702 156
rect 5668 62 5702 84
rect 5824 946 5858 948
rect 5824 910 5858 912
rect 5824 838 5858 844
rect 5824 766 5858 776
rect 5824 694 5858 708
rect 5824 622 5858 640
rect 5824 550 5858 572
rect 5824 478 5858 504
rect 5824 406 5858 436
rect 5824 334 5858 368
rect 5824 266 5858 300
rect 5824 198 5858 228
rect 5824 130 5858 156
rect 5824 62 5858 84
rect 5980 946 6014 948
rect 5980 910 6014 912
rect 5980 838 6014 844
rect 5980 766 6014 776
rect 5980 694 6014 708
rect 5980 622 6014 640
rect 5980 550 6014 572
rect 5980 478 6014 504
rect 5980 406 6014 436
rect 5980 334 6014 368
rect 5980 266 6014 300
rect 5980 198 6014 228
rect 5980 130 6014 156
rect 5980 62 6014 84
rect 6136 946 6170 948
rect 6136 910 6170 912
rect 6136 838 6170 844
rect 6136 766 6170 776
rect 6136 694 6170 708
rect 6136 622 6170 640
rect 6136 550 6170 572
rect 6136 478 6170 504
rect 6136 406 6170 436
rect 6136 334 6170 368
rect 6136 266 6170 300
rect 6136 198 6170 228
rect 6136 130 6170 156
rect 6136 62 6170 84
rect 6292 946 6326 948
rect 6292 910 6326 912
rect 6292 838 6326 844
rect 6292 766 6326 776
rect 6292 694 6326 708
rect 6292 622 6326 640
rect 6292 550 6326 572
rect 6292 478 6326 504
rect 6292 406 6326 436
rect 6292 334 6326 368
rect 6292 266 6326 300
rect 6292 198 6326 228
rect 6292 130 6326 156
rect 6292 62 6326 84
rect 6416 946 6450 948
rect 6416 910 6450 912
rect 6416 838 6450 844
rect 6416 766 6450 776
rect 6416 694 6450 708
rect 6416 622 6450 640
rect 6416 550 6450 572
rect 6416 478 6450 504
rect 6416 406 6450 436
rect 6416 334 6450 368
rect 6416 266 6450 300
rect 6416 198 6450 228
rect 6416 130 6450 156
rect 6416 62 6450 84
rect 6572 946 6606 948
rect 6572 910 6606 912
rect 6572 838 6606 844
rect 6572 766 6606 776
rect 6572 694 6606 708
rect 6572 622 6606 640
rect 6572 550 6606 572
rect 6572 478 6606 504
rect 6572 406 6606 436
rect 6572 334 6606 368
rect 6572 266 6606 300
rect 6572 198 6606 228
rect 6572 130 6606 156
rect 6572 62 6606 84
rect 6696 946 6730 948
rect 6696 910 6730 912
rect 6696 838 6730 844
rect 6696 766 6730 776
rect 6696 694 6730 708
rect 6696 622 6730 640
rect 6696 550 6730 572
rect 6696 478 6730 504
rect 6696 406 6730 436
rect 6696 334 6730 368
rect 6696 266 6730 300
rect 6696 198 6730 228
rect 6696 130 6730 156
rect 6696 62 6730 84
rect 7424 1057 7458 1067
rect 7424 989 7458 995
rect 6852 946 6886 948
rect 6852 910 6886 912
rect 6852 838 6886 844
rect 6852 766 6886 776
rect 6852 694 6886 708
rect 6852 622 6886 640
rect 6852 550 6886 572
rect 6852 478 6886 504
rect 6852 406 6886 436
rect 6852 334 6886 368
rect 6852 266 6886 300
rect 6852 198 6886 228
rect 6852 130 6886 156
rect 6852 62 6886 84
rect 7008 946 7042 948
rect 7008 910 7042 912
rect 7008 838 7042 844
rect 7008 766 7042 776
rect 7008 694 7042 708
rect 7008 622 7042 640
rect 7008 550 7042 572
rect 7008 478 7042 504
rect 7008 406 7042 436
rect 7008 334 7042 368
rect 7008 266 7042 300
rect 7008 198 7042 228
rect 7008 130 7042 156
rect 7008 62 7042 84
rect 7424 921 7458 923
rect 7424 885 7458 887
rect 7424 813 7458 819
rect 7424 741 7458 751
rect 7424 669 7458 683
rect 7424 597 7458 615
rect 7424 525 7458 547
rect 7424 453 7458 479
rect 7424 381 7458 411
rect 7424 309 7458 343
rect 7424 241 7458 275
rect 7424 173 7458 203
rect 7424 105 7458 131
rect 7424 37 7458 59
rect 1622 -41 1724 -14
rect 466 -79 500 -41
rect 1427 -47 1724 -41
rect 1461 -81 1499 -47
rect 1533 -64 1724 -47
rect 1533 -81 1622 -64
rect 1427 -87 1622 -81
rect 466 -151 500 -113
rect 1656 -98 1690 -64
rect 1622 -114 1724 -98
rect 2145 -17 2191 2
rect 7510 1329 7544 1355
rect 7510 1261 7544 1283
rect 7510 1193 7544 1211
rect 7510 1125 7544 1139
rect 7510 1057 7544 1067
rect 7510 989 7544 995
rect 7510 921 7544 923
rect 7510 885 7544 887
rect 7510 813 7544 819
rect 7510 741 7544 751
rect 7510 669 7544 683
rect 7510 597 7544 615
rect 7510 525 7544 547
rect 7510 453 7544 479
rect 7510 381 7544 411
rect 7510 309 7544 343
rect 7510 241 7544 275
rect 7510 173 7544 203
rect 7510 105 7544 131
rect 7510 37 7544 59
rect 7596 1329 7630 1355
rect 7596 1261 7630 1283
rect 7596 1193 7630 1211
rect 7596 1125 7630 1139
rect 7596 1057 7630 1067
rect 7596 989 7630 995
rect 7596 921 7630 923
rect 7596 885 7630 887
rect 7596 813 7630 819
rect 7596 741 7630 751
rect 7596 669 7630 683
rect 7596 597 7630 615
rect 7596 525 7630 547
rect 7596 453 7630 479
rect 7596 381 7630 411
rect 7596 309 7630 343
rect 7596 241 7630 275
rect 7596 173 7630 203
rect 7596 105 7630 131
rect 7596 37 7630 59
rect 7682 1329 7716 1355
rect 7682 1261 7716 1283
rect 7682 1193 7716 1211
rect 7682 1125 7716 1139
rect 7682 1057 7716 1067
rect 7682 989 7716 995
rect 7682 921 7716 923
rect 7682 885 7716 887
rect 7682 813 7716 819
rect 7682 741 7716 751
rect 7682 669 7716 683
rect 7682 597 7716 615
rect 7682 525 7716 547
rect 7682 453 7716 479
rect 7682 381 7716 411
rect 7682 309 7716 343
rect 7682 241 7716 275
rect 7682 173 7716 203
rect 7682 105 7716 131
rect 7682 37 7716 59
rect 7768 1329 7802 1355
rect 7768 1261 7802 1283
rect 7768 1193 7802 1211
rect 7768 1125 7802 1139
rect 7768 1057 7802 1067
rect 7768 989 7802 995
rect 7768 921 7802 923
rect 7768 885 7802 887
rect 7768 813 7802 819
rect 7768 741 7802 751
rect 7768 669 7802 683
rect 7768 597 7802 615
rect 7768 525 7802 547
rect 7768 453 7802 479
rect 7768 381 7802 411
rect 7768 309 7802 343
rect 7768 241 7802 275
rect 7768 173 7802 203
rect 7768 105 7802 131
rect 7768 37 7802 59
rect 7854 1329 7888 1355
rect 9405 1361 9451 1389
rect 19967 1534 20013 1578
rect 19967 1500 19973 1534
rect 20007 1500 20013 1534
rect 19967 1456 20013 1500
rect 25277 1496 25315 1530
rect 19967 1422 19973 1456
rect 20007 1422 20013 1456
rect 19967 1378 20013 1422
rect 9405 1355 12386 1361
rect 13494 1360 18903 1361
rect 13494 1355 19023 1360
rect 9405 1321 9479 1355
rect 9517 1321 9547 1355
rect 9590 1321 9615 1355
rect 9663 1321 9683 1355
rect 9736 1321 9751 1355
rect 9809 1321 9819 1355
rect 9882 1321 9887 1355
rect 9989 1321 9994 1355
rect 10057 1321 10067 1355
rect 10125 1321 10140 1355
rect 10193 1321 10213 1355
rect 10261 1321 10286 1355
rect 10329 1321 10359 1355
rect 10397 1321 10431 1355
rect 10466 1321 10499 1355
rect 10539 1321 10567 1355
rect 10612 1321 10635 1355
rect 10685 1321 10703 1355
rect 10758 1321 10771 1355
rect 10831 1321 10839 1355
rect 10904 1321 10907 1355
rect 10941 1321 10943 1355
rect 11009 1321 11016 1355
rect 11077 1321 11089 1355
rect 11145 1321 11162 1355
rect 11213 1321 11235 1355
rect 11281 1321 11308 1355
rect 11349 1321 11381 1355
rect 11417 1321 11451 1355
rect 11488 1321 11519 1355
rect 11561 1321 11587 1355
rect 11634 1321 11655 1355
rect 11706 1321 11723 1355
rect 11778 1321 11791 1355
rect 11850 1321 11859 1355
rect 11922 1321 11927 1355
rect 11994 1321 11995 1355
rect 12029 1321 12032 1355
rect 12097 1321 12104 1355
rect 12165 1321 12176 1355
rect 12233 1321 12248 1355
rect 12301 1321 12320 1355
rect 12369 1321 12403 1355
rect 12437 1321 12471 1355
rect 12505 1321 12539 1355
rect 12573 1321 12607 1355
rect 12641 1321 12675 1355
rect 12709 1321 12743 1355
rect 12777 1321 12811 1355
rect 12845 1321 12879 1355
rect 12913 1321 12947 1355
rect 12981 1321 13015 1355
rect 13049 1321 13083 1355
rect 13117 1321 13151 1355
rect 13185 1321 13219 1355
rect 13253 1321 13287 1355
rect 13321 1321 13355 1355
rect 13389 1321 13423 1355
rect 13457 1321 13491 1355
rect 13525 1321 13526 1355
rect 13593 1321 13599 1355
rect 13661 1321 13672 1355
rect 13729 1321 13745 1355
rect 13797 1321 13818 1355
rect 13865 1321 13891 1355
rect 13933 1321 13964 1355
rect 14001 1321 14035 1355
rect 14071 1321 14103 1355
rect 14144 1321 14171 1355
rect 14217 1321 14239 1355
rect 14289 1321 14307 1355
rect 14361 1321 14375 1355
rect 14433 1321 14443 1355
rect 14505 1321 14511 1355
rect 14577 1321 14579 1355
rect 14613 1321 14615 1355
rect 14681 1321 14687 1355
rect 14749 1321 14759 1355
rect 14817 1321 14831 1355
rect 14885 1321 14903 1355
rect 14953 1321 14975 1355
rect 15021 1321 15047 1355
rect 15089 1321 15119 1355
rect 15157 1321 15191 1355
rect 15225 1321 15259 1355
rect 15297 1321 15327 1355
rect 15369 1321 15395 1355
rect 15441 1321 15463 1355
rect 15513 1321 15531 1355
rect 15585 1321 15599 1355
rect 15657 1321 15667 1355
rect 15729 1321 15735 1355
rect 15801 1321 15803 1355
rect 15837 1321 15839 1355
rect 15905 1321 15911 1355
rect 15973 1321 15983 1355
rect 16041 1321 16055 1355
rect 16109 1321 16127 1355
rect 16177 1321 16199 1355
rect 16245 1321 16271 1355
rect 16313 1321 16343 1355
rect 16381 1321 16415 1355
rect 16449 1321 16483 1355
rect 16521 1321 16551 1355
rect 16593 1321 16619 1355
rect 16665 1321 16687 1355
rect 16737 1321 16755 1355
rect 16809 1321 16823 1355
rect 16881 1321 16891 1355
rect 16953 1321 16959 1355
rect 17025 1321 17027 1355
rect 17061 1321 17063 1355
rect 17129 1321 17135 1355
rect 17197 1321 17207 1355
rect 17265 1321 17279 1355
rect 17333 1321 17351 1355
rect 17401 1321 17423 1355
rect 17469 1321 17495 1355
rect 17537 1321 17567 1355
rect 17605 1321 17639 1355
rect 17673 1321 17707 1355
rect 17745 1321 17775 1355
rect 17817 1321 17843 1355
rect 17889 1321 17911 1355
rect 17961 1321 17979 1355
rect 18033 1321 18047 1355
rect 18105 1321 18115 1355
rect 18177 1321 18183 1355
rect 18249 1321 18251 1355
rect 18285 1321 18287 1355
rect 18353 1321 18359 1355
rect 18421 1321 18431 1355
rect 18489 1321 18503 1355
rect 18557 1321 18575 1355
rect 18625 1321 18647 1355
rect 18693 1321 18719 1355
rect 18761 1321 18791 1355
rect 18829 1321 19023 1355
rect 9405 1315 12386 1321
rect 13494 1315 19023 1321
rect 7854 1261 7888 1283
rect 7854 1193 7888 1211
rect 18850 1250 19023 1315
rect 18850 1214 18863 1250
rect 18897 1214 19023 1250
rect 18850 1180 19023 1214
rect 18850 1146 18863 1180
rect 18897 1150 19023 1180
rect 19967 1344 19973 1378
rect 20007 1344 20013 1378
rect 19967 1300 20013 1344
rect 19967 1266 19973 1300
rect 20007 1266 20013 1300
rect 19967 1222 20013 1266
rect 20252 1433 20286 1452
rect 25415 1410 25471 1674
rect 25787 1690 25821 1727
rect 25787 1619 25821 1656
rect 25787 1548 25821 1585
rect 25787 1476 25821 1514
rect 20252 1325 20286 1394
rect 25787 1404 25821 1442
rect 25277 1320 25315 1354
rect 25787 1332 25821 1370
rect 20252 1252 20286 1276
rect 25787 1260 25821 1298
rect 19967 1188 19973 1222
rect 20007 1188 20013 1222
rect 25787 1202 25821 1226
rect 28031 1727 28065 1761
rect 28031 1659 28065 1693
rect 28031 1591 28065 1625
rect 28031 1523 28065 1557
rect 28031 1455 28065 1489
rect 28031 1387 28065 1421
rect 28031 1319 28065 1353
rect 28031 1251 28065 1285
rect 19967 1150 20013 1188
rect 18897 1146 20013 1150
rect 18850 1144 20013 1146
rect 7854 1125 7888 1139
rect 15116 1135 15572 1141
rect 7854 1057 7888 1067
rect 12868 1042 12902 1080
rect 15116 1101 15219 1135
rect 15253 1101 15411 1135
rect 15445 1101 15506 1135
rect 15540 1101 15644 1135
rect 15678 1101 15736 1135
rect 15770 1101 15861 1135
rect 15116 1095 15606 1101
rect 8386 1030 8431 1033
rect 8465 1030 8510 1033
rect 8544 1030 8589 1033
rect 8623 1030 8668 1033
rect 8329 996 8345 1030
rect 8386 999 8416 1030
rect 8465 999 8487 1030
rect 8544 999 8559 1030
rect 8623 999 8631 1030
rect 8379 996 8416 999
rect 8450 996 8487 999
rect 8521 996 8559 999
rect 8593 996 8631 999
rect 8665 999 8668 1030
rect 8702 1030 8747 1033
rect 8781 1030 8825 1033
rect 13122 1035 13144 1069
rect 13190 1035 13216 1069
rect 13258 1035 13288 1069
rect 13326 1035 13360 1069
rect 13394 1035 13428 1069
rect 13466 1035 13496 1069
rect 13538 1035 13564 1069
rect 13610 1035 13632 1069
rect 13682 1035 13700 1069
rect 13754 1035 13768 1069
rect 13826 1035 13836 1069
rect 13898 1035 13904 1069
rect 13970 1035 13972 1069
rect 14006 1035 14008 1069
rect 14074 1035 14080 1069
rect 14142 1035 14152 1069
rect 14210 1035 14224 1069
rect 14278 1035 14296 1069
rect 14346 1035 14368 1069
rect 14414 1035 14440 1069
rect 14482 1035 14512 1069
rect 14550 1035 14584 1069
rect 14618 1035 14652 1069
rect 14690 1035 14720 1069
rect 14762 1035 14788 1069
rect 14834 1035 14856 1069
rect 14906 1035 14924 1069
rect 14978 1035 14992 1069
rect 15116 1057 15162 1095
rect 8702 999 8703 1030
rect 8665 996 8703 999
rect 8737 999 8747 1030
rect 8809 999 8825 1030
rect 8737 996 8775 999
rect 8809 996 8847 999
rect 8881 996 8897 1030
rect 8953 996 8967 1030
rect 9003 996 9041 1030
rect 9077 996 9115 1030
rect 9150 996 9189 1030
rect 9223 996 9262 1030
rect 9297 996 9335 1030
rect 9371 996 9408 1030
rect 9445 996 9481 1030
rect 9519 996 9554 1030
rect 9592 996 9627 1030
rect 9665 996 9677 1030
rect 9733 996 9745 1030
rect 9783 996 9819 1030
rect 9856 996 9893 1030
rect 9929 996 9967 1030
rect 10002 996 10041 1030
rect 10075 996 10114 1030
rect 10150 996 10187 1030
rect 10225 996 10260 1030
rect 10300 996 10333 1030
rect 10375 996 10407 1030
rect 10450 996 10457 1030
rect 7854 989 7888 995
rect 10788 996 10804 1030
rect 10839 996 10875 1030
rect 10911 996 10946 1030
rect 10983 996 11017 1030
rect 11055 996 11088 1030
rect 11127 996 11159 1030
rect 11199 996 11230 1030
rect 11271 996 11301 1030
rect 11343 996 11372 1030
rect 11415 996 11443 1030
rect 11487 996 11514 1030
rect 11559 996 11585 1030
rect 11631 996 11656 1030
rect 11703 996 11727 1030
rect 11775 996 11798 1030
rect 11847 996 11869 1030
rect 11919 996 11940 1030
rect 11991 996 12010 1030
rect 12063 996 12080 1030
rect 12135 996 12150 1030
rect 12207 996 12220 1030
rect 12279 996 12290 1030
rect 12324 996 12360 1030
rect 12394 996 12430 1030
rect 12464 996 12500 1030
rect 12534 996 12550 1030
rect 12828 996 12844 1030
rect 12902 1008 12912 1030
rect 12878 996 12912 1008
rect 12946 996 12962 1030
rect 15116 1023 15122 1057
rect 15156 1023 15162 1057
rect 15311 1063 15357 1095
rect 15116 1008 15162 1023
rect 7854 921 7888 923
rect 7854 885 7888 887
rect 7854 813 7888 819
rect 7854 741 7888 751
rect 7854 669 7888 683
rect 7854 597 7888 615
rect 7854 525 7888 547
rect 7854 453 7888 479
rect 7854 381 7888 411
rect 7854 309 7888 343
rect 7854 241 7888 275
rect 7854 173 7888 203
rect 7854 105 7888 131
rect 7854 37 7888 59
rect 8168 942 8202 966
rect 10604 936 10638 977
rect 15116 979 15124 1008
rect 8168 880 8177 908
rect 8168 870 8211 880
rect 8202 838 8211 870
rect 8168 804 8177 836
rect 8168 798 8211 804
rect 8202 764 8211 798
rect 8168 762 8211 764
rect 8168 728 8177 762
rect 8168 726 8211 728
rect 8202 692 8211 726
rect 8168 686 8211 692
rect 8168 654 8177 686
rect 8202 620 8211 652
rect 8168 610 8211 620
rect 8168 582 8177 610
rect 8202 548 8211 576
rect 8168 533 8211 548
rect 8168 510 8177 533
rect 8202 476 8211 499
rect 8168 456 8211 476
rect 8168 438 8177 456
rect 8202 404 8211 422
rect 8168 379 8211 404
rect 8168 366 8177 379
rect 8202 332 8211 345
rect 8168 302 8211 332
rect 8168 294 8177 302
rect 8202 260 8211 268
rect 8168 225 8211 260
rect 8168 222 8177 225
rect 8202 188 8211 191
rect 8168 150 8211 188
rect 8202 148 8211 150
rect 8168 114 8177 116
rect 8168 78 8211 114
rect 8202 71 8211 78
rect 8168 37 8177 44
rect 8168 6 8211 37
rect 8202 -6 8211 6
rect 2145 -72 2151 -17
rect 2185 -72 2191 -17
rect 8168 -40 8177 -28
rect 8284 878 8318 880
rect 8284 842 8318 844
rect 8284 770 8318 776
rect 8284 698 8318 708
rect 8284 626 8318 640
rect 8284 554 8318 572
rect 8284 482 8318 504
rect 8284 410 8318 436
rect 8284 338 8318 368
rect 8284 266 8318 300
rect 8284 198 8318 232
rect 8284 130 8318 160
rect 8284 62 8318 88
rect 8284 -6 8318 16
rect 8168 -52 8202 -40
rect 8440 878 8474 880
rect 8440 842 8474 844
rect 8440 770 8474 776
rect 8440 698 8474 708
rect 8440 626 8474 640
rect 8440 554 8474 572
rect 8440 482 8474 504
rect 8440 410 8474 436
rect 8440 338 8474 368
rect 8440 266 8474 300
rect 8440 198 8474 232
rect 8440 130 8474 160
rect 8440 62 8474 88
rect 8440 -6 8474 16
rect 8596 878 8630 880
rect 8596 842 8630 844
rect 8596 770 8630 776
rect 8596 698 8630 708
rect 8596 626 8630 640
rect 8596 554 8630 572
rect 8596 482 8630 504
rect 8596 410 8630 436
rect 8596 338 8630 368
rect 8596 266 8630 300
rect 8596 198 8630 232
rect 8596 130 8630 160
rect 8596 62 8630 88
rect 8596 -6 8630 16
rect 8752 878 8786 880
rect 8752 842 8786 844
rect 8752 770 8786 776
rect 8752 698 8786 708
rect 8752 626 8786 640
rect 8752 554 8786 572
rect 8752 482 8786 504
rect 8752 410 8786 436
rect 8752 338 8786 368
rect 8752 266 8786 300
rect 8752 198 8786 232
rect 8752 130 8786 160
rect 8752 62 8786 88
rect 8752 -6 8786 16
rect 8908 878 8942 880
rect 8908 842 8942 844
rect 8908 770 8942 776
rect 8908 698 8942 708
rect 8908 626 8942 640
rect 8908 554 8942 572
rect 8908 482 8942 504
rect 8908 410 8942 436
rect 8908 338 8942 368
rect 8908 266 8942 300
rect 8908 198 8942 232
rect 8908 130 8942 160
rect 8908 62 8942 88
rect 8908 -6 8942 16
rect 9064 878 9098 880
rect 9064 842 9098 844
rect 9064 770 9098 776
rect 9064 698 9098 708
rect 9064 626 9098 640
rect 9064 554 9098 572
rect 9064 482 9098 504
rect 9064 410 9098 436
rect 9064 338 9098 368
rect 9064 266 9098 300
rect 9064 198 9098 232
rect 9064 130 9098 160
rect 9064 62 9098 88
rect 9064 -6 9098 16
rect 9220 878 9254 880
rect 9220 842 9254 844
rect 9220 770 9254 776
rect 9220 698 9254 708
rect 9220 626 9254 640
rect 9220 554 9254 572
rect 9220 482 9254 504
rect 9220 410 9254 436
rect 9220 338 9254 368
rect 9220 266 9254 300
rect 9220 198 9254 232
rect 9220 130 9254 160
rect 9220 62 9254 88
rect 9220 -6 9254 16
rect 9376 878 9410 880
rect 9376 842 9410 844
rect 9376 770 9410 776
rect 9376 698 9410 708
rect 9376 626 9410 640
rect 9376 554 9410 572
rect 9376 482 9410 504
rect 9376 410 9410 436
rect 9376 338 9410 368
rect 9376 266 9410 300
rect 9376 198 9410 232
rect 9376 130 9410 160
rect 9376 62 9410 88
rect 9376 -6 9410 16
rect 9532 878 9566 880
rect 9532 842 9566 844
rect 9532 770 9566 776
rect 9532 698 9566 708
rect 9532 626 9566 640
rect 9532 554 9566 572
rect 9532 482 9566 504
rect 9532 410 9566 436
rect 9532 338 9566 368
rect 9532 266 9566 300
rect 9532 198 9566 232
rect 9532 130 9566 160
rect 9532 62 9566 88
rect 9532 -6 9566 16
rect 9688 878 9722 880
rect 9688 842 9722 844
rect 9688 770 9722 776
rect 9688 698 9722 708
rect 9688 626 9722 640
rect 9688 554 9722 572
rect 9688 482 9722 504
rect 9688 410 9722 436
rect 9688 338 9722 368
rect 9688 266 9722 300
rect 9688 198 9722 232
rect 9688 130 9722 160
rect 9688 62 9722 88
rect 9688 -6 9722 16
rect 9844 878 9878 880
rect 9844 842 9878 844
rect 9844 770 9878 776
rect 9844 698 9878 708
rect 9844 626 9878 640
rect 9844 554 9878 572
rect 9844 482 9878 504
rect 9844 410 9878 436
rect 9844 338 9878 368
rect 9844 266 9878 300
rect 9844 198 9878 232
rect 9844 130 9878 160
rect 9844 62 9878 88
rect 9844 -6 9878 16
rect 10000 878 10034 880
rect 10000 842 10034 844
rect 10000 770 10034 776
rect 10000 698 10034 708
rect 10000 626 10034 640
rect 10000 554 10034 572
rect 10000 482 10034 504
rect 10000 410 10034 436
rect 10000 338 10034 368
rect 10000 266 10034 300
rect 10000 198 10034 232
rect 10000 130 10034 160
rect 10000 62 10034 88
rect 10000 -6 10034 16
rect 10156 878 10190 880
rect 10156 842 10190 844
rect 10156 770 10190 776
rect 10156 698 10190 708
rect 10156 626 10190 640
rect 10156 554 10190 572
rect 10156 482 10190 504
rect 10156 410 10190 436
rect 10156 338 10190 368
rect 10156 266 10190 300
rect 10156 198 10190 232
rect 10156 130 10190 160
rect 10156 62 10190 88
rect 10156 -6 10190 16
rect 10312 878 10346 880
rect 10312 842 10346 844
rect 10312 770 10346 776
rect 10312 698 10346 708
rect 10312 626 10346 640
rect 10312 554 10346 572
rect 10312 482 10346 504
rect 10312 410 10346 436
rect 10312 338 10346 368
rect 10312 266 10346 300
rect 10312 198 10346 232
rect 10312 130 10346 160
rect 10312 62 10346 88
rect 10312 -6 10346 16
rect 10468 878 10502 880
rect 10468 842 10502 844
rect 10468 770 10502 776
rect 10468 698 10502 708
rect 10468 626 10502 640
rect 10468 554 10502 572
rect 10468 482 10502 504
rect 10468 410 10502 436
rect 10468 338 10502 368
rect 10468 266 10502 300
rect 10468 198 10502 232
rect 10468 130 10502 160
rect 10468 62 10502 88
rect 10468 -6 10502 16
rect 12783 930 12817 946
rect 10604 861 10638 890
rect 10604 786 10638 820
rect 10604 714 10638 750
rect 10604 644 10638 676
rect 10604 574 10638 600
rect 10604 503 10638 524
rect 10604 432 10638 448
rect 10604 361 10638 372
rect 10604 290 10638 296
rect 10604 254 10638 256
rect 10604 219 10638 220
rect 10604 178 10638 185
rect 10604 102 10638 114
rect 10604 26 10638 43
rect 10604 -50 10638 -28
rect 2145 -85 2191 -72
rect 620 -159 642 -125
rect 688 -159 714 -125
rect 756 -159 786 -125
rect 824 -159 858 -125
rect 892 -159 926 -125
rect 964 -159 994 -125
rect 1036 -159 1062 -125
rect 1108 -159 1130 -125
rect 1180 -159 1198 -125
rect 1252 -159 1266 -125
rect 1324 -159 1334 -125
rect 1396 -159 1402 -125
rect 1468 -159 1470 -125
rect 1504 -159 1506 -125
rect 2145 -146 2151 -85
rect 2185 -146 2191 -85
rect 2398 -92 2410 -58
rect 2456 -92 2483 -58
rect 2525 -92 2556 -58
rect 2594 -92 2629 -58
rect 2663 -92 2698 -58
rect 2736 -92 2767 -58
rect 2809 -92 2836 -58
rect 2882 -92 2905 -58
rect 2955 -92 2974 -58
rect 3028 -92 3043 -58
rect 3101 -92 3112 -58
rect 3174 -92 3181 -58
rect 3247 -92 3250 -58
rect 3284 -92 3286 -58
rect 3353 -92 3359 -58
rect 3422 -92 3432 -58
rect 3491 -92 3505 -58
rect 3560 -92 3578 -58
rect 3629 -92 3651 -58
rect 3698 -92 3724 -58
rect 3767 -92 3797 -58
rect 3836 -92 3870 -58
rect 3905 -92 3940 -58
rect 3977 -92 4008 -58
rect 4050 -92 4076 -58
rect 4123 -92 4144 -58
rect 4195 -92 4212 -58
rect 4267 -92 4280 -58
rect 4339 -92 4348 -58
rect 4411 -92 4416 -58
rect 4483 -92 4484 -58
rect 4518 -92 4521 -58
rect 4586 -92 4593 -58
rect 4654 -92 4665 -58
rect 4722 -92 4737 -58
rect 4790 -92 4809 -58
rect 4858 -92 4881 -58
rect 4926 -92 4953 -58
rect 4994 -92 5025 -58
rect 5062 -92 5096 -58
rect 5131 -92 5164 -58
rect 5203 -92 5232 -58
rect 5275 -92 5300 -58
rect 5347 -92 5368 -58
rect 5419 -92 5436 -58
rect 5491 -92 5504 -58
rect 5563 -92 5572 -58
rect 5635 -92 5640 -58
rect 5674 -92 5686 -58
rect 5742 -92 5760 -58
rect 5810 -92 5834 -58
rect 5878 -92 5908 -58
rect 5946 -92 5980 -58
rect 6016 -92 6048 -58
rect 6090 -92 6116 -58
rect 6163 -92 6184 -58
rect 6236 -92 6252 -58
rect 6309 -92 6320 -58
rect 6382 -92 6388 -58
rect 6455 -92 6456 -58
rect 6490 -92 6494 -58
rect 6558 -92 6567 -58
rect 6626 -92 6640 -58
rect 6694 -92 6713 -58
rect 6762 -92 6786 -58
rect 6830 -92 6859 -58
rect 6898 -92 6922 -58
rect 10737 878 10771 880
rect 10737 842 10771 844
rect 10737 770 10771 776
rect 10737 698 10771 708
rect 10737 626 10771 640
rect 10737 554 10771 572
rect 10737 482 10771 504
rect 10737 410 10771 436
rect 10737 338 10771 368
rect 10737 266 10771 300
rect 10737 198 10771 232
rect 10737 130 10771 160
rect 10737 62 10771 88
rect 10737 -6 10771 16
rect 11193 878 11227 880
rect 11193 842 11227 844
rect 11193 770 11227 776
rect 11193 698 11227 708
rect 11193 626 11227 640
rect 11193 554 11227 572
rect 11193 482 11227 504
rect 11193 410 11227 436
rect 11193 338 11227 368
rect 11193 266 11227 300
rect 11193 198 11227 232
rect 11193 130 11227 160
rect 11193 62 11227 88
rect 11193 -6 11227 16
rect 11649 878 11683 880
rect 11649 842 11683 844
rect 11649 770 11683 776
rect 11649 698 11683 708
rect 11649 626 11683 640
rect 11649 554 11683 572
rect 11649 482 11683 504
rect 11649 410 11683 436
rect 11649 338 11683 368
rect 11649 266 11683 300
rect 11649 198 11683 232
rect 11649 130 11683 160
rect 11649 62 11683 88
rect 11649 -6 11683 16
rect 12105 878 12139 880
rect 12105 842 12139 844
rect 12105 770 12139 776
rect 12105 698 12139 708
rect 12105 626 12139 640
rect 12105 554 12139 572
rect 12105 482 12139 504
rect 12105 410 12139 436
rect 12105 338 12139 368
rect 12105 266 12139 300
rect 12105 198 12139 232
rect 12105 130 12139 160
rect 12105 62 12139 88
rect 12105 -6 12139 16
rect 12561 878 12595 880
rect 12561 842 12595 844
rect 12561 770 12595 776
rect 12783 862 12817 893
rect 12783 805 12817 828
rect 12783 744 12817 760
rect 12959 930 12993 946
rect 12959 862 12993 893
rect 15116 945 15122 979
rect 15158 974 15162 1008
rect 15156 945 15162 974
rect 15116 940 15162 945
rect 15116 906 15124 940
rect 15158 906 15162 940
rect 15116 901 15162 906
rect 15116 867 15122 901
rect 15156 872 15162 901
rect 15116 838 15124 867
rect 15158 838 15162 872
rect 12959 805 12993 828
rect 13122 799 13144 833
rect 13190 799 13216 833
rect 13258 799 13288 833
rect 13326 799 13360 833
rect 13394 799 13428 833
rect 13466 799 13496 833
rect 13538 799 13564 833
rect 13610 799 13632 833
rect 13682 799 13700 833
rect 13754 799 13768 833
rect 13826 799 13836 833
rect 13898 799 13904 833
rect 13970 799 13972 833
rect 14006 799 14008 833
rect 14074 799 14080 833
rect 14142 799 14152 833
rect 14210 799 14224 833
rect 14278 799 14296 833
rect 14346 799 14368 833
rect 14414 799 14440 833
rect 14482 799 14512 833
rect 14550 799 14584 833
rect 14618 799 14652 833
rect 14690 799 14720 833
rect 14762 799 14788 833
rect 14834 799 14856 833
rect 14906 799 14924 833
rect 14978 799 14992 833
rect 15116 823 15162 838
rect 15223 966 15257 988
rect 15223 894 15257 920
rect 15223 836 15257 852
rect 15311 1029 15317 1063
rect 15351 1029 15357 1063
rect 15572 1058 15606 1095
rect 15311 983 15357 1029
rect 15311 949 15317 983
rect 15351 949 15357 983
rect 15311 903 15357 949
rect 15311 869 15317 903
rect 15351 869 15357 903
rect 12959 744 12993 760
rect 15116 789 15122 823
rect 15156 804 15162 823
rect 15116 770 15124 789
rect 15158 778 15162 804
rect 15311 823 15357 869
rect 15459 966 15493 988
rect 15459 894 15493 920
rect 15459 836 15493 852
rect 15827 1063 15861 1101
rect 18850 1112 18937 1144
rect 15572 981 15606 1024
rect 15572 904 15606 947
rect 15311 789 15317 823
rect 15351 789 15357 823
rect 15311 778 15357 789
rect 15572 826 15606 870
rect 15695 966 15729 988
rect 15695 894 15729 920
rect 15695 836 15729 852
rect 16344 1073 16394 1085
rect 15827 988 15861 1029
rect 15827 913 15861 954
rect 15827 839 15861 879
rect 15572 778 15606 792
rect 15931 966 15965 988
rect 15931 894 15965 920
rect 15931 836 15965 852
rect 16049 978 16083 1017
rect 16049 905 16083 944
rect 15827 778 15861 805
rect 16049 832 16083 871
rect 16167 966 16201 988
rect 16167 894 16201 920
rect 16167 836 16201 852
rect 16344 1027 16352 1073
rect 16386 1027 16394 1073
rect 16344 999 16394 1027
rect 16344 940 16352 999
rect 16386 940 16394 999
rect 16344 925 16394 940
rect 16344 891 16352 925
rect 16386 891 16394 925
rect 16344 887 16394 891
rect 16344 853 16352 887
rect 16386 853 16394 887
rect 16344 851 16394 853
rect 16049 778 16083 798
rect 16344 817 16352 851
rect 16386 817 16394 851
rect 16344 800 16394 817
rect 15158 770 15284 778
rect 15116 745 15284 770
rect 12561 698 12595 708
rect 15116 711 15122 745
rect 15156 744 15284 745
rect 15318 744 15353 778
rect 15387 744 15422 778
rect 15456 744 15491 778
rect 15525 744 15560 778
rect 15594 748 15629 778
rect 15606 744 15629 748
rect 15663 744 15698 778
rect 15732 744 15766 778
rect 15800 765 15834 778
rect 15800 744 15827 765
rect 15868 744 15902 778
rect 15936 744 15970 778
rect 16004 744 16038 778
rect 16072 759 16106 778
rect 16083 744 16106 759
rect 16140 744 16156 778
rect 15156 736 15162 744
rect 15116 702 15124 711
rect 15158 702 15162 736
rect 15116 668 15162 702
rect 15311 743 15357 744
rect 15311 709 15317 743
rect 15351 709 15357 743
rect 15116 667 15124 668
rect 12561 626 12595 640
rect 12561 554 12595 572
rect 12561 482 12595 504
rect 12561 410 12595 436
rect 12561 338 12595 368
rect 12561 266 12595 300
rect 12561 198 12595 232
rect 12561 130 12595 160
rect 12561 62 12595 88
rect 12561 -6 12595 16
rect 12678 636 12712 644
rect 15116 633 15122 667
rect 15158 634 15162 668
rect 15156 633 15162 634
rect 15116 599 15162 633
rect 12678 560 12712 586
rect 13122 563 13144 597
rect 13190 563 13216 597
rect 13258 563 13288 597
rect 13326 563 13360 597
rect 13394 563 13428 597
rect 13466 563 13496 597
rect 13538 563 13564 597
rect 13610 563 13632 597
rect 13682 563 13700 597
rect 13754 563 13768 597
rect 13826 563 13836 597
rect 13898 563 13904 597
rect 13970 563 13972 597
rect 14006 563 14008 597
rect 14074 563 14080 597
rect 14142 563 14152 597
rect 14210 563 14224 597
rect 14278 563 14296 597
rect 14346 563 14368 597
rect 14414 563 14440 597
rect 14482 563 14512 597
rect 14550 563 14584 597
rect 14618 563 14652 597
rect 14690 563 14720 597
rect 14762 563 14788 597
rect 14834 563 14856 597
rect 14906 563 14924 597
rect 14978 563 14992 597
rect 15116 589 15124 599
rect 15116 555 15122 589
rect 15158 565 15162 599
rect 15156 555 15162 565
rect 15116 530 15162 555
rect 15116 522 15124 530
rect 12678 484 12712 513
rect 12678 408 12712 440
rect 12784 516 15124 522
rect 12784 482 12816 516
rect 12850 482 12889 516
rect 12923 482 12962 516
rect 12784 444 12962 482
rect 12784 410 12816 444
rect 12850 410 12889 444
rect 12923 410 12962 444
rect 15084 511 15124 516
rect 15084 477 15122 511
rect 15158 496 15162 530
rect 15156 477 15162 496
rect 15084 461 15162 477
rect 15223 661 15257 677
rect 15223 593 15257 619
rect 15223 525 15257 547
rect 15311 663 15357 709
rect 15311 629 15317 663
rect 15351 629 15357 663
rect 15311 584 15357 629
rect 15311 550 15317 584
rect 15351 550 15357 584
rect 15311 505 15357 550
rect 15084 433 15124 461
rect 15084 410 15122 433
rect 15158 427 15162 461
rect 12784 404 15122 410
rect 12678 332 12712 367
rect 15116 399 15122 404
rect 15156 399 15162 427
rect 15116 398 15162 399
rect 15311 471 15317 505
rect 15351 471 15357 505
rect 15459 661 15493 677
rect 15459 593 15493 619
rect 15459 525 15493 547
rect 15572 670 15606 714
rect 15827 691 15861 731
rect 15572 592 15606 636
rect 15572 514 15606 558
rect 15311 426 15357 471
rect 15311 398 15317 426
rect 15351 398 15357 426
rect 15572 436 15606 480
rect 15695 661 15729 677
rect 15695 593 15729 619
rect 15695 525 15729 547
rect 16049 686 16083 725
rect 15827 617 15861 657
rect 15827 543 15861 583
rect 15572 398 15606 402
rect 15827 469 15861 509
rect 15931 661 15965 677
rect 15931 593 15965 619
rect 15931 525 15965 547
rect 16344 743 16352 800
rect 16386 743 16394 800
rect 16344 713 16394 743
rect 16049 613 16083 652
rect 16049 540 16083 579
rect 15827 398 15861 435
rect 16049 467 16083 506
rect 16167 661 16201 677
rect 16167 593 16201 619
rect 16167 525 16201 547
rect 16344 669 16352 713
rect 16386 669 16394 713
rect 16344 629 16394 669
rect 16344 592 16352 629
rect 16386 592 16394 629
rect 16344 555 16394 592
rect 16344 505 16352 555
rect 16386 505 16394 555
rect 16344 481 16394 505
rect 16049 398 16083 433
rect 16344 418 16352 481
rect 16386 418 16394 481
rect 16344 407 16394 418
rect 15116 392 15284 398
rect 15351 392 15353 398
rect 13122 327 13144 361
rect 13190 327 13216 361
rect 13258 327 13288 361
rect 13326 327 13360 361
rect 13394 327 13428 361
rect 13466 327 13496 361
rect 13538 327 13564 361
rect 13610 327 13632 361
rect 13682 327 13700 361
rect 13754 327 13768 361
rect 13826 327 13836 361
rect 13898 327 13904 361
rect 13970 327 13972 361
rect 14006 327 14008 361
rect 14074 327 14080 361
rect 14142 327 14152 361
rect 14210 327 14224 361
rect 14278 327 14296 361
rect 14346 327 14368 361
rect 14414 327 14440 361
rect 14482 327 14512 361
rect 14550 327 14584 361
rect 14618 327 14652 361
rect 14690 327 14720 361
rect 14762 327 14788 361
rect 14834 327 14856 361
rect 14906 327 14924 361
rect 14978 327 14992 361
rect 15116 358 15124 392
rect 15158 364 15284 392
rect 15318 364 15353 392
rect 15387 364 15422 398
rect 15456 364 15491 398
rect 15525 364 15560 398
rect 15594 364 15629 398
rect 15663 364 15698 398
rect 15732 364 15766 398
rect 15800 364 15834 398
rect 15868 395 15902 398
rect 15868 364 15899 395
rect 15936 364 15970 398
rect 16004 395 16038 398
rect 16008 364 16038 395
rect 16072 364 16106 398
rect 16140 364 16156 398
rect 16344 373 16352 407
rect 16386 373 16394 407
rect 16344 365 16394 373
rect 15158 358 15162 364
rect 15311 360 15357 364
rect 15116 354 15162 358
rect 12678 256 12712 294
rect 12678 182 12712 221
rect 15116 320 15122 354
rect 15156 323 15162 354
rect 15116 289 15124 320
rect 15158 289 15162 323
rect 15572 358 15606 364
rect 15827 361 15899 364
rect 15933 361 15974 364
rect 16008 361 16083 364
rect 15116 275 15162 289
rect 15116 241 15122 275
rect 15156 254 15162 275
rect 15116 220 15124 241
rect 15158 220 15162 254
rect 15116 209 15162 220
rect 15223 226 15257 248
rect 12678 109 12712 146
rect 15124 185 15158 209
rect 15124 135 15158 151
rect 15223 154 15257 180
rect 13122 91 13144 125
rect 13190 91 13216 125
rect 13258 91 13288 125
rect 13326 91 13360 125
rect 13394 91 13428 125
rect 13466 91 13496 125
rect 13538 91 13564 125
rect 13610 91 13632 125
rect 13682 91 13700 125
rect 13754 91 13768 125
rect 13826 91 13836 125
rect 13898 91 13904 125
rect 13970 91 13972 125
rect 14006 91 14008 125
rect 14074 91 14080 125
rect 14142 91 14152 125
rect 14210 91 14224 125
rect 14278 91 14296 125
rect 14346 91 14368 125
rect 14414 91 14440 125
rect 14482 91 14512 125
rect 14550 91 14584 125
rect 14618 91 14652 125
rect 14690 91 14720 125
rect 14762 91 14788 125
rect 14834 91 14856 125
rect 14906 91 14924 125
rect 14978 91 14992 125
rect 15223 96 15257 112
rect 15459 226 15493 248
rect 15459 154 15493 180
rect 15572 280 15606 324
rect 16344 299 16352 365
rect 16386 299 16394 365
rect 18850 1078 18863 1112
rect 18897 1110 18937 1112
rect 18971 1110 19011 1144
rect 19045 1110 19085 1144
rect 19119 1110 19159 1144
rect 19193 1110 19233 1144
rect 19267 1110 19307 1144
rect 19341 1110 19381 1144
rect 19415 1110 19455 1144
rect 19489 1110 19529 1144
rect 19563 1110 19603 1144
rect 19637 1110 19677 1144
rect 19711 1110 19751 1144
rect 19785 1110 19826 1144
rect 19860 1110 19901 1144
rect 19935 1110 20013 1144
rect 18897 1104 20013 1110
rect 28031 1183 28065 1217
rect 28031 1115 28065 1149
rect 18897 1078 19023 1104
rect 18850 1072 19023 1078
rect 18850 1010 18863 1072
rect 18897 1010 19023 1072
rect 18850 995 19023 1010
rect 18850 942 18863 995
rect 18897 942 19023 995
rect 18850 918 19023 942
rect 18850 874 18863 918
rect 18897 874 19023 918
rect 18850 842 19023 874
rect 18850 806 18863 842
rect 18897 806 19023 842
rect 18850 772 19023 806
rect 18850 732 18863 772
rect 18897 732 19023 772
rect 18850 704 19023 732
rect 18850 656 18863 704
rect 18897 656 19023 704
rect 18850 636 19023 656
rect 18850 580 18863 636
rect 18897 580 19023 636
rect 18850 568 19023 580
rect 18850 504 18863 568
rect 18897 504 19023 568
rect 18850 500 19023 504
rect 18850 466 18863 500
rect 18897 466 19023 500
rect 18850 462 19023 466
rect 18850 398 18863 462
rect 18897 398 19023 462
rect 18850 386 19023 398
rect 18416 338 18454 341
rect 18448 307 18454 338
rect 18398 304 18414 307
rect 18448 304 18482 307
rect 18516 304 18550 338
rect 18584 304 18600 338
rect 18850 330 18863 386
rect 18897 330 19023 386
rect 18850 310 19023 330
rect 15572 202 15606 246
rect 16344 278 16394 299
rect 15695 226 15729 248
rect 15895 225 15911 259
rect 15945 225 15979 259
rect 16017 225 16029 259
rect 16085 225 16097 259
rect 16135 225 16169 259
rect 16207 225 16219 259
rect 16344 225 16352 278
rect 16386 225 16394 278
rect 18850 262 18863 310
rect 18897 262 19023 310
rect 15459 96 15493 112
rect 15695 154 15729 180
rect 16344 191 16394 225
rect 18628 223 18644 257
rect 18681 223 18712 257
rect 18753 223 18762 257
rect 18850 234 19023 262
rect 16344 151 16352 191
rect 16386 151 16394 191
rect 18850 194 18863 234
rect 18897 194 19023 234
rect 15695 96 15729 112
rect 15884 107 15918 109
rect 12678 36 12712 70
rect 12678 -37 12712 -7
rect 15884 71 15918 73
rect 15884 -1 15918 5
rect 13180 -37 13219 -36
rect 13253 -37 13292 -36
rect 13326 -37 13365 -36
rect 13399 -37 13438 -36
rect 13472 -37 13511 -36
rect 13545 -37 13584 -36
rect 13618 -37 13657 -36
rect 13691 -37 13730 -36
rect 13764 -37 13803 -36
rect 13837 -37 13876 -36
rect 13910 -37 13949 -36
rect 13983 -37 14022 -36
rect 14056 -37 14095 -36
rect 14129 -37 14168 -36
rect 14202 -37 14241 -36
rect 14275 -37 14314 -36
rect 14348 -37 14387 -36
rect 14421 -37 14460 -36
rect 14494 -37 14533 -36
rect 14567 -37 14606 -36
rect 14640 -37 14679 -36
rect 14713 -37 14752 -36
rect 14786 -37 14825 -36
rect 14859 -37 14898 -36
rect 14932 -37 14971 -36
rect 15005 -37 15043 -36
rect 15077 -37 15115 -36
rect 15149 -37 15187 -36
rect 15221 -37 15259 -36
rect 15293 -37 15331 -36
rect 15365 -37 15403 -36
rect 15437 -37 15475 -36
rect 15509 -37 15547 -36
rect 15581 -37 15619 -36
rect 13118 -71 13142 -37
rect 13180 -70 13211 -37
rect 13253 -70 13280 -37
rect 13326 -70 13349 -37
rect 13399 -70 13418 -37
rect 13472 -70 13486 -37
rect 13545 -70 13554 -37
rect 13618 -70 13622 -37
rect 13176 -71 13211 -70
rect 13245 -71 13280 -70
rect 13314 -71 13349 -70
rect 13383 -71 13418 -70
rect 13452 -71 13486 -70
rect 13520 -71 13554 -70
rect 13588 -71 13622 -70
rect 13656 -70 13657 -37
rect 13724 -70 13730 -37
rect 13792 -70 13803 -37
rect 13860 -70 13876 -37
rect 13928 -70 13949 -37
rect 13996 -70 14022 -37
rect 14064 -70 14095 -37
rect 13656 -71 13690 -70
rect 13724 -71 13758 -70
rect 13792 -71 13826 -70
rect 13860 -71 13894 -70
rect 13928 -71 13962 -70
rect 13996 -71 14030 -70
rect 14064 -71 14098 -70
rect 14132 -71 14166 -37
rect 14202 -70 14234 -37
rect 14275 -70 14302 -37
rect 14348 -70 14370 -37
rect 14421 -70 14438 -37
rect 14494 -70 14506 -37
rect 14567 -70 14574 -37
rect 14640 -70 14642 -37
rect 14200 -71 14234 -70
rect 14268 -71 14302 -70
rect 14336 -71 14370 -70
rect 14404 -71 14438 -70
rect 14472 -71 14506 -70
rect 14540 -71 14574 -70
rect 14608 -71 14642 -70
rect 14676 -70 14679 -37
rect 14744 -70 14752 -37
rect 14812 -70 14825 -37
rect 14880 -70 14898 -37
rect 14948 -70 14971 -37
rect 15016 -70 15043 -37
rect 15084 -70 15115 -37
rect 14676 -71 14710 -70
rect 14744 -71 14778 -70
rect 14812 -71 14846 -70
rect 14880 -71 14914 -70
rect 14948 -71 14982 -70
rect 15016 -71 15050 -70
rect 15084 -71 15118 -70
rect 15152 -71 15186 -37
rect 15221 -70 15254 -37
rect 15293 -70 15322 -37
rect 15365 -70 15390 -37
rect 15437 -70 15458 -37
rect 15509 -70 15526 -37
rect 15581 -70 15594 -37
rect 15653 -70 15662 -37
rect 15220 -71 15254 -70
rect 15288 -71 15322 -70
rect 15356 -71 15390 -70
rect 15424 -71 15458 -70
rect 15492 -71 15526 -70
rect 15560 -71 15594 -70
rect 15628 -71 15662 -70
rect 15696 -69 15730 -37
rect 15764 -69 15821 -37
rect 15696 -71 15709 -69
rect 15764 -71 15781 -69
rect 12678 -95 12712 -84
rect 466 -223 500 -185
rect 466 -295 500 -257
rect 1622 -186 1656 -170
rect 1622 -281 1656 -234
rect 620 -315 642 -281
rect 688 -315 714 -281
rect 756 -315 786 -281
rect 824 -315 858 -281
rect 892 -315 926 -281
rect 964 -315 994 -281
rect 1036 -315 1062 -281
rect 1108 -315 1130 -281
rect 1180 -315 1198 -281
rect 1252 -315 1266 -281
rect 1324 -315 1334 -281
rect 1396 -315 1402 -281
rect 1468 -315 1470 -281
rect 1504 -315 1506 -281
rect 466 -368 500 -329
rect 466 -441 500 -402
rect 1622 -371 1656 -319
rect 2145 -186 2191 -146
rect 2145 -220 2151 -186
rect 2185 -220 2191 -186
rect 2145 -234 2191 -220
rect 2145 -294 2151 -234
rect 2185 -294 2191 -234
rect 2145 -326 2191 -294
rect 15703 -103 15709 -71
rect 15743 -103 15781 -71
rect 15815 -103 15821 -69
rect 15703 -142 15821 -103
rect 15703 -176 15709 -142
rect 15743 -176 15781 -142
rect 15815 -176 15821 -142
rect 15703 -215 15821 -176
rect 15703 -249 15709 -215
rect 15743 -249 15781 -215
rect 15815 -249 15821 -215
rect 15703 -288 15821 -249
rect 15703 -322 15709 -288
rect 15743 -322 15781 -288
rect 15815 -322 15821 -288
rect 2145 -360 2219 -326
rect 2253 -332 2287 -326
rect 2321 -332 2355 -326
rect 2389 -332 2423 -326
rect 2457 -332 2491 -326
rect 2261 -360 2287 -332
rect 2337 -360 2355 -332
rect 2413 -360 2423 -332
rect 2489 -360 2491 -332
rect 2525 -332 2559 -326
rect 2593 -332 2627 -326
rect 2661 -332 2695 -326
rect 2729 -332 2763 -326
rect 2525 -360 2531 -332
rect 2593 -360 2607 -332
rect 2661 -360 2683 -332
rect 2729 -360 2759 -332
rect 2797 -360 2831 -326
rect 2865 -332 2899 -326
rect 2933 -332 2967 -326
rect 3001 -332 3035 -326
rect 3069 -332 3103 -326
rect 2869 -360 2899 -332
rect 2945 -360 2967 -332
rect 3021 -360 3035 -332
rect 3097 -360 3103 -332
rect 3137 -332 3171 -326
rect 3205 -332 3239 -326
rect 3273 -332 3307 -326
rect 3137 -360 3140 -332
rect 3205 -360 3217 -332
rect 3273 -360 3294 -332
rect 3341 -360 15632 -326
rect 2145 -366 2227 -360
rect 2261 -366 2303 -360
rect 2337 -366 2379 -360
rect 2413 -366 2455 -360
rect 2489 -366 2531 -360
rect 2565 -366 2607 -360
rect 2641 -366 2683 -360
rect 2717 -366 2759 -360
rect 2793 -366 2835 -360
rect 2869 -366 2911 -360
rect 2945 -366 2987 -360
rect 3021 -366 3063 -360
rect 3097 -366 3140 -360
rect 3174 -366 3217 -360
rect 3251 -366 3294 -360
rect 3328 -366 3386 -360
rect 2145 -372 3386 -366
rect 1622 -426 1656 -410
rect 620 -471 642 -437
rect 688 -471 714 -437
rect 756 -471 786 -437
rect 824 -471 858 -437
rect 892 -471 926 -437
rect 964 -471 994 -437
rect 1036 -471 1062 -437
rect 1108 -471 1130 -437
rect 1180 -471 1198 -437
rect 1252 -471 1266 -437
rect 1324 -471 1334 -437
rect 1396 -471 1402 -437
rect 1468 -471 1470 -437
rect 1504 -471 1506 -437
rect 466 -514 500 -475
rect 1622 -509 1724 -482
rect 466 -587 500 -548
rect 1427 -515 1724 -509
rect 1461 -549 1499 -515
rect 1533 -532 1724 -515
rect 1533 -549 1622 -532
rect 1427 -555 1622 -549
rect 1656 -566 1690 -532
rect 1622 -582 1724 -566
rect 1782 -531 1882 -519
rect 1782 -565 1802 -531
rect 1836 -565 1882 -531
rect 466 -660 500 -621
rect 620 -627 642 -593
rect 688 -627 714 -593
rect 756 -627 786 -593
rect 824 -627 858 -593
rect 892 -627 926 -593
rect 964 -627 994 -593
rect 1036 -627 1062 -593
rect 1108 -627 1130 -593
rect 1180 -627 1198 -593
rect 1252 -627 1266 -593
rect 1324 -627 1334 -593
rect 1396 -627 1402 -593
rect 1468 -627 1470 -593
rect 1504 -627 1506 -593
rect 1782 -603 1882 -565
rect 1782 -637 1802 -603
rect 1836 -637 1882 -603
rect 1782 -638 1882 -637
rect 466 -733 500 -694
rect 1622 -688 1882 -638
rect 1656 -722 1690 -688
rect 1724 -722 1882 -688
rect 1622 -738 1882 -722
rect 466 -806 500 -767
rect 570 -783 586 -749
rect 620 -783 654 -749
rect 688 -783 722 -749
rect 756 -783 790 -749
rect 824 -783 836 -749
rect 892 -783 911 -749
rect 960 -783 986 -749
rect 1028 -783 1061 -749
rect 1096 -783 1130 -749
rect 1170 -783 1198 -749
rect 1244 -783 1266 -749
rect 1318 -783 1334 -749
rect 1392 -783 1402 -749
rect 1466 -783 1470 -749
rect 1504 -783 1506 -749
rect 466 -879 500 -840
rect 466 -952 500 -913
rect 574 -917 598 -883
rect 632 -886 668 -883
rect 632 -917 666 -886
rect 702 -917 738 -883
rect 772 -886 808 -883
rect 842 -886 878 -883
rect 912 -886 948 -883
rect 982 -886 1019 -883
rect 1053 -886 1090 -883
rect 1124 -886 1161 -883
rect 776 -917 808 -886
rect 852 -917 878 -886
rect 928 -917 948 -886
rect 1004 -917 1019 -886
rect 1080 -917 1090 -886
rect 1156 -917 1161 -886
rect 1195 -886 1232 -883
rect 1195 -917 1198 -886
rect 700 -920 742 -917
rect 776 -920 818 -917
rect 852 -920 894 -917
rect 928 -920 970 -917
rect 1004 -920 1046 -917
rect 1080 -920 1122 -917
rect 1156 -920 1198 -917
rect 1266 -886 1303 -883
rect 1337 -886 1374 -883
rect 1408 -886 1445 -883
rect 1479 -886 1516 -883
rect 1266 -917 1274 -886
rect 1337 -917 1350 -886
rect 1408 -917 1426 -886
rect 1479 -917 1502 -886
rect 1550 -917 1574 -883
rect 1232 -920 1274 -917
rect 1308 -920 1350 -917
rect 1384 -920 1426 -917
rect 1460 -920 1502 -917
rect 466 -1025 500 -986
rect 466 -1098 500 -1059
rect 570 -1068 586 -1034
rect 620 -1068 654 -1034
rect 688 -1068 722 -1034
rect 756 -1068 790 -1034
rect 824 -1068 858 -1034
rect 892 -1068 926 -1034
rect 960 -1068 994 -1034
rect 1028 -1068 1062 -1034
rect 1096 -1068 1103 -1034
rect 1164 -1068 1183 -1034
rect 1232 -1068 1263 -1034
rect 1300 -1068 1334 -1034
rect 1377 -1068 1402 -1034
rect 1457 -1068 1470 -1034
rect 466 -1171 500 -1132
rect 1622 -1095 1656 -1079
rect 1622 -1190 1656 -1143
rect 466 -1244 500 -1205
rect 620 -1224 642 -1190
rect 688 -1224 714 -1190
rect 756 -1224 786 -1190
rect 824 -1224 858 -1190
rect 892 -1224 926 -1190
rect 964 -1224 994 -1190
rect 1036 -1224 1062 -1190
rect 1108 -1224 1130 -1190
rect 1180 -1224 1198 -1190
rect 1252 -1224 1266 -1190
rect 1324 -1224 1334 -1190
rect 1396 -1224 1402 -1190
rect 1468 -1224 1470 -1190
rect 1504 -1224 1506 -1190
rect 466 -1317 500 -1278
rect 1622 -1231 1656 -1224
rect 15598 -1200 15632 -360
rect 15703 -361 15821 -322
rect 15703 -395 15709 -361
rect 15743 -395 15781 -361
rect 15815 -395 15821 -361
rect 15703 -434 15821 -395
rect 15703 -468 15709 -434
rect 15743 -468 15781 -434
rect 15815 -468 15821 -434
rect 15703 -507 15821 -468
rect 15703 -541 15709 -507
rect 15743 -541 15781 -507
rect 15815 -541 15821 -507
rect 15703 -580 15821 -541
rect 15703 -614 15709 -580
rect 15743 -614 15781 -580
rect 15815 -614 15821 -580
rect 15703 -653 15821 -614
rect 15703 -687 15709 -653
rect 15743 -687 15781 -653
rect 15815 -687 15821 -653
rect 15703 -727 15821 -687
rect 15703 -761 15709 -727
rect 15743 -761 15781 -727
rect 15815 -761 15821 -727
rect 15703 -801 15821 -761
rect 15703 -835 15709 -801
rect 15743 -835 15781 -801
rect 15815 -835 15821 -801
rect 15884 -73 15918 -63
rect 15884 -145 15918 -131
rect 15884 -217 15918 -199
rect 15884 -289 15918 -267
rect 15884 -361 15918 -335
rect 15884 -433 15918 -403
rect 15884 -505 15918 -471
rect 15884 -573 15918 -539
rect 15884 -641 15918 -611
rect 15884 -709 15918 -683
rect 15884 -777 15918 -755
rect 16040 107 16074 109
rect 16040 71 16074 73
rect 16040 -1 16074 5
rect 16040 -73 16074 -63
rect 16040 -145 16074 -131
rect 16040 -217 16074 -199
rect 16040 -289 16074 -267
rect 16040 -361 16074 -335
rect 16040 -433 16074 -403
rect 16040 -505 16074 -471
rect 16040 -573 16074 -539
rect 16040 -641 16074 -611
rect 16040 -709 16074 -683
rect 16040 -777 16074 -755
rect 16196 107 16230 109
rect 16196 71 16230 73
rect 16196 -1 16230 5
rect 16196 -73 16230 -63
rect 16196 -145 16230 -131
rect 16196 -217 16230 -199
rect 16196 -289 16230 -267
rect 16196 -361 16230 -335
rect 16196 -433 16230 -403
rect 16196 -505 16230 -471
rect 16196 -573 16230 -539
rect 16196 -641 16230 -611
rect 16196 -709 16230 -683
rect 16196 -777 16230 -755
rect 16344 111 16394 151
rect 18398 148 18414 182
rect 18448 148 18482 182
rect 18516 148 18550 182
rect 18588 148 18600 182
rect 18850 160 19023 194
rect 16344 70 16352 111
rect 16386 70 16394 111
rect 18850 126 18863 160
rect 18897 126 19023 160
rect 18628 71 18644 105
rect 18681 71 18712 105
rect 18753 71 18762 105
rect 18850 92 19023 126
rect 16344 37 16394 70
rect 16344 -17 16352 37
rect 16386 -17 16394 37
rect 18850 58 18863 92
rect 18897 86 19023 92
rect 18897 58 18953 86
rect 18850 52 18953 58
rect 18987 52 19023 86
rect 18398 -8 18414 26
rect 18448 -8 18482 26
rect 18516 -8 18550 26
rect 18588 -8 18600 26
rect 18850 24 19023 52
rect 16344 -38 16394 -17
rect 16344 -104 16352 -38
rect 16386 -104 16394 -38
rect 16344 -113 16394 -104
rect 16344 -147 16352 -113
rect 16386 -147 16394 -113
rect 16344 -157 16394 -147
rect 16344 -222 16352 -157
rect 16386 -222 16394 -157
rect 16344 -245 16394 -222
rect 16344 -297 16352 -245
rect 16386 -297 16394 -245
rect 16344 -333 16394 -297
rect 16344 -372 16352 -333
rect 16386 -372 16394 -333
rect 16344 -413 16394 -372
rect 16344 -455 16352 -413
rect 16386 -455 16394 -413
rect 16344 -488 16394 -455
rect 16344 -543 16352 -488
rect 16386 -543 16394 -488
rect 16344 -563 16394 -543
rect 16344 -631 16352 -563
rect 16386 -631 16394 -563
rect 16344 -638 16394 -631
rect 16344 -672 16352 -638
rect 16386 -672 16394 -638
rect 16344 -685 16394 -672
rect 16344 -747 16352 -685
rect 16386 -747 16394 -685
rect 16344 -773 16394 -747
rect 16344 -822 16352 -773
rect 16386 -822 16394 -773
rect 15703 -867 15821 -835
rect 16344 -861 16394 -822
rect 16344 -897 16352 -861
rect 16386 -897 16394 -861
rect 16344 -929 16394 -897
rect 15874 -935 16394 -929
rect 15874 -937 15917 -935
rect 15874 -971 15898 -937
rect 15951 -969 15990 -935
rect 16024 -937 16063 -935
rect 16097 -937 16136 -935
rect 16025 -969 16063 -937
rect 16118 -969 16136 -937
rect 16170 -937 16208 -935
rect 16242 -937 16280 -935
rect 16170 -969 16176 -937
rect 16242 -969 16268 -937
rect 16314 -969 16394 -935
rect 15932 -971 15991 -969
rect 16025 -971 16084 -969
rect 16118 -971 16176 -969
rect 16210 -971 16268 -969
rect 16302 -971 16394 -969
rect 15874 -979 16394 -971
rect 18850 -10 18863 24
rect 18897 12 19023 24
rect 18897 -10 18953 12
rect 18850 -22 18953 -10
rect 18987 -22 19023 12
rect 18850 -44 19023 -22
rect 18850 -78 18863 -44
rect 18897 -62 19023 -44
rect 18897 -78 18953 -62
rect 18850 -96 18953 -78
rect 18987 -96 19023 -62
rect 18850 -112 19023 -96
rect 18850 -146 18863 -112
rect 18897 -136 19023 -112
rect 18897 -146 18953 -136
rect 18850 -170 18953 -146
rect 18987 -170 19023 -136
rect 18850 -180 19023 -170
rect 18850 -214 18863 -180
rect 18897 -210 19023 -180
rect 18897 -214 18953 -210
rect 18850 -244 18953 -214
rect 18987 -244 19023 -210
rect 18850 -248 19023 -244
rect 18850 -282 18863 -248
rect 18897 -282 19023 -248
rect 18850 -284 19023 -282
rect 18850 -316 18953 -284
rect 18850 -350 18863 -316
rect 18897 -318 18953 -316
rect 18987 -318 19023 -284
rect 18897 -350 19023 -318
rect 18850 -358 19023 -350
rect 18850 -384 18953 -358
rect 18850 -418 18863 -384
rect 18897 -392 18953 -384
rect 18987 -392 19023 -358
rect 18897 -418 19023 -392
rect 18850 -432 19023 -418
rect 18850 -452 18953 -432
rect 18850 -486 18863 -452
rect 18897 -466 18953 -452
rect 18987 -466 19023 -432
rect 18897 -486 19023 -466
rect 18850 -506 19023 -486
rect 18850 -520 18953 -506
rect 18850 -554 18863 -520
rect 18897 -540 18953 -520
rect 18987 -540 19023 -506
rect 18897 -554 19023 -540
rect 18850 -580 19023 -554
rect 18850 -588 18953 -580
rect 18850 -622 18863 -588
rect 18897 -614 18953 -588
rect 18987 -614 19023 -580
rect 18897 -622 19023 -614
rect 18850 -653 19023 -622
rect 18850 -656 18953 -653
rect 18850 -690 18863 -656
rect 18897 -687 18953 -656
rect 18987 -687 19023 -653
rect 18897 -690 19023 -687
rect 18850 -724 19023 -690
rect 18850 -758 18863 -724
rect 18897 -726 19023 -724
rect 18897 -758 18953 -726
rect 18850 -760 18953 -758
rect 18987 -760 19023 -726
rect 18850 -792 19023 -760
rect 18850 -826 18863 -792
rect 18897 -799 19023 -792
rect 18897 -826 18953 -799
rect 18850 -833 18953 -826
rect 18987 -833 19023 -799
rect 18850 -860 19023 -833
rect 18850 -894 18863 -860
rect 18897 -872 19023 -860
rect 18897 -894 18953 -872
rect 18850 -906 18953 -894
rect 18987 -906 19023 -872
rect 18850 -928 19023 -906
rect 18850 -962 18863 -928
rect 18897 -945 19023 -928
rect 18897 -962 18953 -945
rect 18850 -979 18953 -962
rect 18987 -979 19023 -945
rect 18850 -996 19023 -979
rect 18850 -1030 18863 -996
rect 18897 -1018 19023 -996
rect 18897 -1030 18953 -1018
rect 18850 -1052 18953 -1030
rect 18987 -1052 19023 -1018
rect 18850 -1064 19023 -1052
rect 18850 -1098 18863 -1064
rect 18897 -1091 19023 -1064
rect 18897 -1098 18953 -1091
rect 18850 -1125 18953 -1098
rect 18987 -1125 19023 -1091
rect 18850 -1132 19023 -1125
rect 18850 -1166 18863 -1132
rect 18897 -1164 19023 -1132
rect 18897 -1166 18953 -1164
rect 18850 -1198 18953 -1166
rect 18987 -1198 19023 -1164
rect 18850 -1200 19023 -1198
rect 15598 -1234 18016 -1200
rect 18050 -1234 18096 -1200
rect 18130 -1234 18176 -1200
rect 18210 -1234 18255 -1200
rect 18289 -1234 18334 -1200
rect 18368 -1234 18413 -1200
rect 18447 -1234 18530 -1200
rect 18564 -1234 18598 -1200
rect 18632 -1234 18666 -1200
rect 18700 -1234 18734 -1200
rect 18768 -1234 19023 -1200
rect 1622 -1285 1656 -1265
rect 1622 -1335 1656 -1319
rect 17913 -1237 19023 -1234
rect 17913 -1252 18953 -1237
rect 17913 -1286 17961 -1252
rect 17995 -1286 18037 -1252
rect 18071 -1286 18113 -1252
rect 18147 -1286 18189 -1252
rect 18223 -1286 18265 -1252
rect 18299 -1286 18341 -1252
rect 18375 -1286 18417 -1252
rect 18451 -1271 18953 -1252
rect 18987 -1271 19023 -1237
rect 18451 -1286 19023 -1271
rect 17913 -1310 19023 -1286
rect 17913 -1332 18953 -1310
rect 466 -1390 500 -1351
rect 620 -1380 642 -1346
rect 688 -1380 714 -1346
rect 756 -1380 786 -1346
rect 824 -1380 858 -1346
rect 892 -1380 926 -1346
rect 964 -1380 994 -1346
rect 1036 -1380 1062 -1346
rect 1108 -1380 1130 -1346
rect 1180 -1380 1198 -1346
rect 1252 -1380 1266 -1346
rect 1324 -1380 1334 -1346
rect 1396 -1380 1402 -1346
rect 1468 -1380 1470 -1346
rect 1504 -1380 1506 -1346
rect 17913 -1366 17961 -1332
rect 17995 -1366 18037 -1332
rect 18071 -1366 18113 -1332
rect 18147 -1366 18189 -1332
rect 18223 -1366 18265 -1332
rect 18299 -1366 18341 -1332
rect 18375 -1366 18417 -1332
rect 18451 -1344 18953 -1332
rect 18987 -1344 19023 -1310
rect 18451 -1366 19023 -1344
rect 17913 -1383 19023 -1366
rect 466 -1463 500 -1424
rect 466 -1536 500 -1497
rect 1622 -1407 1656 -1391
rect 1622 -1502 1656 -1441
rect 17913 -1412 18953 -1383
rect 17913 -1446 17961 -1412
rect 17995 -1446 18037 -1412
rect 18071 -1446 18113 -1412
rect 18147 -1446 18189 -1412
rect 18223 -1446 18265 -1412
rect 18299 -1446 18341 -1412
rect 18375 -1446 18417 -1412
rect 18451 -1417 18953 -1412
rect 18987 -1417 19023 -1383
rect 18451 -1446 19023 -1417
rect 17913 -1456 19023 -1446
rect 28031 1047 28065 1081
rect 28031 979 28065 1013
rect 28031 911 28065 945
rect 28031 843 28065 877
rect 28031 775 28065 809
rect 28031 707 28065 741
rect 28031 639 28065 673
rect 28031 571 28065 605
rect 28031 503 28065 537
rect 28031 435 28065 469
rect 28031 367 28065 401
rect 28031 299 28065 333
rect 28031 231 28065 265
rect 28031 163 28065 197
rect 28031 95 28065 129
rect 28031 27 28065 61
rect 28031 -41 28065 -7
rect 28031 -109 28065 -75
rect 28031 -177 28065 -143
rect 28031 -245 28065 -211
rect 28031 -313 28065 -279
rect 28031 -381 28065 -347
rect 28031 -449 28065 -415
rect 28031 -517 28065 -483
rect 28031 -585 28065 -551
rect 28031 -653 28065 -619
rect 28031 -721 28065 -687
rect 28031 -789 28065 -755
rect 28031 -857 28065 -823
rect 28031 -925 28065 -891
rect 28031 -993 28065 -959
rect 28031 -1061 28065 -1027
rect 28031 -1129 28065 -1095
rect 28031 -1197 28065 -1163
rect 28031 -1265 28065 -1231
rect 28031 -1333 28065 -1299
rect 28031 -1401 28065 -1367
rect 620 -1536 642 -1502
rect 688 -1536 714 -1502
rect 756 -1536 786 -1502
rect 824 -1536 858 -1502
rect 892 -1536 926 -1502
rect 964 -1536 994 -1502
rect 1036 -1536 1062 -1502
rect 1108 -1536 1130 -1502
rect 1180 -1536 1198 -1502
rect 1252 -1536 1266 -1502
rect 1324 -1536 1334 -1502
rect 1396 -1536 1402 -1502
rect 1468 -1536 1470 -1502
rect 1504 -1536 1506 -1502
rect 466 -1609 500 -1570
rect 466 -1682 500 -1643
rect 1622 -1592 1656 -1541
rect 1622 -1647 1656 -1631
rect 28031 -1469 28065 -1435
rect 28031 -1537 28065 -1503
rect 28031 -1605 28065 -1571
rect 620 -1692 642 -1658
rect 688 -1692 714 -1658
rect 756 -1692 786 -1658
rect 824 -1692 858 -1658
rect 892 -1692 926 -1658
rect 964 -1692 994 -1658
rect 1036 -1692 1062 -1658
rect 1108 -1692 1130 -1658
rect 1180 -1692 1198 -1658
rect 1252 -1692 1266 -1658
rect 1324 -1692 1334 -1658
rect 1396 -1692 1402 -1658
rect 1468 -1692 1470 -1658
rect 1504 -1692 1506 -1658
rect 28031 -1673 28065 -1639
rect 466 -1755 500 -1716
rect 466 -1828 500 -1789
rect 1622 -1719 1656 -1703
rect 1622 -1814 1656 -1767
rect 620 -1848 642 -1814
rect 688 -1848 714 -1814
rect 756 -1848 786 -1814
rect 824 -1848 858 -1814
rect 892 -1848 926 -1814
rect 964 -1848 994 -1814
rect 1036 -1848 1062 -1814
rect 1108 -1848 1130 -1814
rect 1180 -1848 1198 -1814
rect 1252 -1848 1266 -1814
rect 1324 -1848 1334 -1814
rect 1396 -1848 1402 -1814
rect 1468 -1848 1470 -1814
rect 1504 -1848 1506 -1814
rect 466 -1901 500 -1862
rect 466 -1974 500 -1935
rect 1622 -1904 1656 -1852
rect 1622 -1959 1656 -1943
rect 28031 -1741 28065 -1707
rect 28031 -1809 28065 -1775
rect 28031 -1877 28065 -1843
rect 28031 -1945 28065 -1911
rect 620 -2004 642 -1970
rect 688 -2004 714 -1970
rect 756 -2004 786 -1970
rect 824 -2004 858 -1970
rect 892 -2004 926 -1970
rect 964 -2004 994 -1970
rect 1036 -2004 1062 -1970
rect 1108 -2004 1130 -1970
rect 1180 -2004 1198 -1970
rect 1252 -2004 1266 -1970
rect 1324 -2004 1334 -1970
rect 1396 -2004 1402 -1970
rect 1468 -2004 1470 -1970
rect 1504 -2004 1506 -1970
rect 466 -2047 500 -2008
rect 28031 -2013 28065 -1979
rect 466 -2120 500 -2081
rect 1622 -2031 1656 -2015
rect 1622 -2126 1656 -2079
rect 620 -2160 644 -2126
rect 688 -2160 718 -2126
rect 756 -2160 790 -2126
rect 826 -2160 858 -2126
rect 899 -2160 926 -2126
rect 972 -2160 994 -2126
rect 1045 -2160 1062 -2126
rect 1096 -2160 1130 -2126
rect 1164 -2160 1198 -2126
rect 1232 -2160 1266 -2126
rect 1300 -2160 1334 -2126
rect 1368 -2160 1402 -2126
rect 1436 -2160 1470 -2126
rect 1504 -2160 1520 -2126
rect 1622 -2216 1656 -2164
rect 1622 -2271 1656 -2255
rect 28031 -2081 28065 -2047
rect 28031 -2149 28065 -2115
rect 28031 -2217 28065 -2183
rect 620 -2316 642 -2282
rect 688 -2316 714 -2282
rect 756 -2316 786 -2282
rect 824 -2316 858 -2282
rect 892 -2316 926 -2282
rect 964 -2316 994 -2282
rect 1036 -2316 1062 -2282
rect 1108 -2316 1130 -2282
rect 1180 -2316 1198 -2282
rect 1252 -2316 1266 -2282
rect 1324 -2316 1334 -2282
rect 1396 -2316 1402 -2282
rect 1468 -2316 1470 -2282
rect 1504 -2316 1506 -2282
rect 28031 -2285 28065 -2251
rect 28031 -2353 28065 -2319
rect 631 -2398 675 -2397
rect 709 -2398 753 -2397
rect 787 -2398 831 -2397
rect 865 -2398 909 -2397
rect 943 -2398 987 -2397
rect 1021 -2398 1065 -2397
rect 1099 -2398 1143 -2397
rect 1177 -2398 1220 -2397
rect 1254 -2398 1297 -2397
rect 1331 -2398 1374 -2397
rect 1408 -2398 1451 -2397
rect 1485 -2398 1528 -2397
rect 574 -2431 597 -2398
rect 574 -2432 598 -2431
rect 632 -2432 668 -2398
rect 709 -2431 738 -2398
rect 787 -2431 808 -2398
rect 865 -2431 878 -2398
rect 943 -2431 948 -2398
rect 702 -2432 738 -2431
rect 772 -2432 808 -2431
rect 842 -2432 878 -2431
rect 912 -2432 948 -2431
rect 982 -2431 987 -2398
rect 1053 -2431 1065 -2398
rect 1124 -2431 1143 -2398
rect 1195 -2431 1220 -2398
rect 1266 -2431 1297 -2398
rect 982 -2432 1019 -2431
rect 1053 -2432 1090 -2431
rect 1124 -2432 1161 -2431
rect 1195 -2432 1232 -2431
rect 1266 -2432 1303 -2431
rect 1337 -2432 1374 -2398
rect 1408 -2432 1445 -2398
rect 1485 -2431 1516 -2398
rect 1562 -2431 1574 -2398
rect 1479 -2432 1516 -2431
rect 1550 -2432 1574 -2431
rect 28031 -2421 28065 -2387
rect 28031 -2489 28065 -2455
rect 28031 -2557 28065 -2523
rect 28031 -2625 28065 -2591
rect 28031 -2693 28065 -2659
rect 28031 -2761 28065 -2727
rect 28031 -2829 28065 -2795
rect 28031 -2897 28065 -2863
rect 28031 -2965 28065 -2931
rect 28031 -3033 28065 -2999
rect 28031 -3101 28065 -3067
rect 28031 -3169 28065 -3135
rect 406 -3243 495 -3231
rect 406 -3277 407 -3243
rect 441 -3265 495 -3243
rect 529 -3265 563 -3231
rect 597 -3265 631 -3231
rect 665 -3265 699 -3231
rect 734 -3265 767 -3231
rect 811 -3265 835 -3231
rect 869 -3265 903 -3231
rect 937 -3265 971 -3231
rect 1005 -3241 1073 -3231
rect 1005 -3265 1039 -3241
rect 406 -3299 441 -3277
rect 440 -3316 441 -3299
rect 406 -3350 407 -3333
rect 406 -3367 441 -3350
rect 440 -3389 441 -3367
rect 1039 -3313 1073 -3275
rect 406 -3423 407 -3401
rect 880 -3369 946 -3368
rect 880 -3403 890 -3369
rect 930 -3403 946 -3369
rect 1039 -3385 1073 -3355
rect 406 -3435 441 -3423
rect 440 -3462 441 -3435
rect 406 -3496 407 -3469
rect 890 -3441 924 -3403
rect 1039 -3457 1073 -3423
rect 406 -3503 441 -3496
rect 440 -3535 441 -3503
rect 406 -3569 407 -3537
rect 406 -3571 441 -3569
rect 440 -3605 441 -3571
rect 406 -3608 441 -3605
rect 406 -3639 407 -3608
rect 440 -3673 441 -3642
rect 406 -3681 441 -3673
rect 406 -3715 407 -3681
rect 406 -3746 441 -3715
rect 440 -3754 441 -3746
rect 406 -3788 407 -3780
rect 406 -3814 441 -3788
rect 440 -3827 441 -3814
rect 406 -3861 407 -3848
rect 406 -3882 441 -3861
rect 440 -3900 441 -3882
rect 406 -3934 407 -3916
rect 406 -3950 441 -3934
rect 440 -3973 441 -3950
rect 406 -4007 407 -3984
rect 406 -4018 441 -4007
rect 440 -4046 441 -4018
rect 406 -4080 407 -4052
rect 406 -4086 441 -4080
rect 440 -4119 441 -4086
rect 406 -4153 407 -4120
rect 406 -4154 441 -4153
rect 440 -4188 441 -4154
rect 406 -4192 441 -4188
rect 406 -4222 407 -4192
rect 440 -4256 441 -4226
rect 406 -4265 441 -4256
rect 406 -4290 407 -4265
rect 440 -4324 441 -4299
rect 406 -4338 441 -4324
rect 406 -4358 407 -4338
rect 440 -4392 441 -4372
rect 406 -4411 441 -4392
rect 406 -4426 407 -4411
rect 440 -4460 441 -4445
rect 406 -4484 441 -4460
rect 406 -4494 407 -4484
rect 440 -4528 441 -4518
rect 406 -4557 441 -4528
rect 406 -4562 407 -4557
rect 440 -4596 441 -4591
rect 406 -4630 441 -4596
rect 406 -4698 441 -4664
rect 440 -4703 441 -4698
rect 406 -4737 407 -4732
rect 406 -4766 441 -4737
rect 440 -4775 441 -4766
rect 406 -4809 407 -4800
rect 406 -4834 441 -4809
rect 440 -4847 441 -4834
rect 406 -4881 407 -4868
rect 406 -4902 441 -4881
rect 440 -4919 441 -4902
rect 406 -4953 407 -4936
rect 406 -4970 441 -4953
rect 440 -4991 441 -4970
rect 406 -5025 407 -5004
rect 406 -5038 441 -5025
rect 440 -5063 441 -5038
rect 406 -5097 407 -5072
rect 406 -5106 441 -5097
rect 440 -5135 441 -5106
rect 406 -5169 407 -5140
rect 406 -5174 441 -5169
rect 440 -5207 441 -5174
rect 406 -5241 407 -5208
rect 406 -5242 441 -5241
rect 440 -5276 441 -5242
rect 406 -5279 441 -5276
rect 406 -5310 407 -5279
rect 440 -5344 441 -5313
rect 406 -5351 441 -5344
rect 406 -5378 407 -5351
rect 440 -5412 441 -5385
rect 406 -5423 441 -5412
rect 406 -5446 407 -5423
rect 440 -5480 441 -5457
rect 406 -5495 441 -5480
rect 406 -5514 407 -5495
rect 440 -5548 441 -5529
rect 406 -5567 441 -5548
rect 406 -5582 407 -5567
rect 440 -5616 441 -5601
rect 406 -5639 441 -5616
rect 406 -5650 407 -5639
rect 440 -5684 441 -5673
rect 406 -5711 441 -5684
rect 406 -5718 407 -5711
rect 440 -5752 441 -5745
rect 406 -5783 441 -5752
rect 406 -5786 407 -5783
rect 440 -5820 441 -5817
rect 406 -5854 441 -5820
rect 440 -5855 441 -5854
rect 406 -5889 407 -5888
rect 406 -5922 441 -5889
rect 440 -5927 441 -5922
rect 406 -5961 407 -5956
rect 406 -5990 441 -5961
rect 440 -5999 441 -5990
rect 406 -6033 407 -6024
rect 406 -6058 441 -6033
rect 440 -6071 441 -6058
rect 406 -6105 407 -6092
rect 406 -6126 441 -6105
rect 440 -6143 441 -6126
rect 406 -6177 407 -6160
rect 406 -6194 441 -6177
rect 440 -6215 441 -6194
rect 406 -6249 407 -6228
rect 406 -6262 441 -6249
rect 440 -6287 441 -6262
rect 406 -6321 407 -6296
rect 406 -6330 441 -6321
rect 440 -6359 441 -6330
rect 406 -6393 407 -6364
rect 406 -6398 441 -6393
rect 440 -6431 441 -6398
rect 406 -6465 407 -6432
rect 406 -6466 441 -6465
rect 440 -6500 441 -6466
rect 406 -6503 441 -6500
rect 406 -6534 407 -6503
rect 440 -6568 441 -6537
rect 406 -6575 441 -6568
rect 406 -6602 407 -6575
rect 440 -6636 441 -6609
rect 406 -6647 441 -6636
rect 406 -6670 407 -6647
rect 440 -6704 441 -6681
rect 406 -6719 441 -6704
rect 406 -6738 407 -6719
rect 440 -6772 441 -6753
rect 406 -6791 441 -6772
rect 406 -6806 407 -6791
rect 440 -6840 441 -6825
rect 406 -6863 441 -6840
rect 406 -6874 407 -6863
rect 440 -6908 441 -6897
rect 406 -6935 441 -6908
rect 406 -6942 407 -6935
rect 440 -6976 441 -6969
rect 406 -7007 441 -6976
rect 406 -7010 407 -7007
rect 440 -7044 441 -7041
rect 406 -7078 441 -7044
rect 440 -7079 441 -7078
rect 406 -7113 407 -7112
rect 406 -7146 441 -7113
rect 440 -7151 441 -7146
rect 406 -7185 407 -7180
rect 406 -7214 441 -7185
rect 440 -7223 441 -7214
rect 406 -7257 407 -7248
rect 406 -7282 441 -7257
rect 440 -7295 441 -7282
rect 406 -7329 407 -7316
rect 406 -7350 441 -7329
rect 440 -7367 441 -7350
rect 406 -7401 407 -7384
rect 406 -7418 441 -7401
rect 440 -7439 441 -7418
rect 406 -7473 407 -7452
rect 406 -7486 441 -7473
rect 440 -7511 441 -7486
rect 406 -7545 407 -7520
rect 406 -7554 441 -7545
rect 440 -7583 441 -7554
rect 406 -7617 407 -7588
rect 406 -7622 441 -7617
rect 440 -7655 441 -7622
rect 406 -7689 407 -7656
rect 406 -7690 441 -7689
rect 440 -7724 441 -7690
rect 406 -7727 441 -7724
rect 406 -7758 407 -7727
rect 440 -7792 441 -7761
rect 406 -7799 441 -7792
rect 406 -7826 407 -7799
rect 440 -7860 441 -7833
rect 406 -7871 441 -7860
rect 406 -7894 407 -7871
rect 440 -7928 441 -7905
rect 406 -7943 441 -7928
rect 406 -7962 407 -7943
rect 440 -7996 441 -7977
rect 406 -8015 441 -7996
rect 406 -8030 407 -8015
rect 440 -8064 441 -8049
rect 406 -8087 441 -8064
rect 406 -8098 407 -8087
rect 440 -8132 441 -8121
rect 406 -8159 441 -8132
rect 406 -8166 407 -8159
rect 440 -8200 441 -8193
rect 406 -8231 441 -8200
rect 406 -8234 407 -8231
rect 440 -8268 441 -8265
rect 406 -8302 441 -8268
rect 440 -8303 441 -8302
rect 406 -8337 407 -8336
rect 406 -8370 441 -8337
rect 440 -8375 441 -8370
rect 406 -8409 407 -8404
rect 406 -8438 441 -8409
rect 440 -8447 441 -8438
rect 406 -8481 407 -8472
rect 406 -8506 441 -8481
rect 440 -8519 441 -8506
rect 406 -8553 407 -8540
rect 406 -8574 441 -8553
rect 440 -8591 441 -8574
rect 406 -8625 407 -8608
rect 406 -8642 441 -8625
rect 440 -8663 441 -8642
rect 406 -8697 407 -8676
rect 406 -8710 441 -8697
rect 440 -8735 441 -8710
rect 406 -8769 407 -8744
rect 406 -8778 441 -8769
rect 440 -8807 441 -8778
rect 406 -8841 407 -8812
rect 406 -8846 441 -8841
rect 440 -8879 441 -8846
rect 406 -8913 407 -8880
rect 406 -8914 441 -8913
rect 440 -8948 441 -8914
rect 406 -8951 441 -8948
rect 406 -8982 407 -8951
rect 440 -9016 441 -8985
rect 406 -9023 441 -9016
rect 406 -9050 407 -9023
rect 440 -9084 441 -9057
rect 406 -9095 441 -9084
rect 406 -9118 407 -9095
rect 440 -9152 441 -9129
rect 406 -9167 441 -9152
rect 406 -9186 407 -9167
rect 440 -9220 441 -9201
rect 406 -9239 441 -9220
rect 406 -9254 407 -9239
rect 440 -9288 441 -9273
rect 406 -9311 441 -9288
rect 406 -9322 407 -9311
rect 440 -9356 441 -9345
rect 406 -9383 441 -9356
rect 406 -9390 407 -9383
rect 440 -9424 441 -9417
rect 406 -9455 441 -9424
rect 406 -9458 407 -9455
rect 440 -9492 441 -9489
rect 406 -9526 441 -9492
rect 440 -9527 441 -9526
rect 406 -9561 407 -9560
rect 406 -9594 441 -9561
rect 440 -9599 441 -9594
rect 406 -9633 407 -9628
rect 406 -9662 441 -9633
rect 440 -9671 441 -9662
rect 406 -9705 407 -9696
rect 406 -9730 441 -9705
rect 440 -9743 441 -9730
rect 406 -9777 407 -9764
rect 406 -9798 441 -9777
rect 440 -9815 441 -9798
rect 406 -9849 407 -9832
rect 406 -9866 441 -9849
rect 440 -9887 441 -9866
rect 406 -9921 407 -9900
rect 406 -9934 441 -9921
rect 440 -9959 441 -9934
rect 406 -9993 407 -9968
rect 406 -10002 441 -9993
rect 440 -10031 441 -10002
rect 406 -10065 407 -10036
rect 406 -10070 441 -10065
rect 440 -10103 441 -10070
rect 406 -10137 407 -10104
rect 406 -10138 441 -10137
rect 440 -10172 441 -10138
rect 406 -10175 441 -10172
rect 406 -10206 407 -10175
rect 440 -10240 441 -10209
rect 406 -10247 441 -10240
rect 406 -10274 407 -10247
rect 440 -10308 441 -10281
rect 406 -10319 441 -10308
rect 406 -10342 407 -10319
rect 440 -10376 441 -10353
rect 406 -10391 441 -10376
rect 406 -10410 407 -10391
rect 440 -10444 441 -10425
rect 406 -10463 441 -10444
rect 406 -10478 407 -10463
rect 440 -10512 441 -10497
rect 406 -10535 441 -10512
rect 406 -10546 407 -10535
rect 440 -10580 441 -10569
rect 406 -10607 441 -10580
rect 406 -10614 407 -10607
rect 440 -10648 441 -10641
rect 406 -10679 441 -10648
rect 406 -10682 407 -10679
rect 440 -10716 441 -10713
rect 406 -10750 441 -10716
rect 440 -10751 441 -10750
rect 406 -10785 407 -10784
rect 406 -10818 441 -10785
rect 440 -10823 441 -10818
rect 1039 -3525 1073 -3491
rect 1039 -3593 1073 -3563
rect 1039 -3661 1073 -3635
rect 1039 -3729 1073 -3707
rect 1039 -3797 1073 -3779
rect 1039 -3865 1073 -3851
rect 1039 -3933 1073 -3923
rect 1039 -4001 1073 -3995
rect 1039 -4069 1073 -4067
rect 1039 -4105 1073 -4103
rect 1039 -4177 1073 -4171
rect 1039 -4249 1073 -4239
rect 1039 -4321 1073 -4307
rect 1039 -4393 1073 -4375
rect 1039 -4465 1073 -4443
rect 1039 -4537 1073 -4511
rect 1039 -4609 1073 -4579
rect 1039 -4681 1073 -4647
rect 1039 -4749 1073 -4715
rect 1039 -4817 1073 -4787
rect 1039 -4885 1073 -4859
rect 1039 -4953 1073 -4931
rect 1039 -5021 1073 -5003
rect 1039 -5089 1073 -5075
rect 1039 -5157 1073 -5147
rect 1039 -5225 1073 -5219
rect 1039 -5293 1073 -5291
rect 1039 -5329 1073 -5327
rect 1039 -5401 1073 -5395
rect 1039 -5473 1073 -5463
rect 1039 -5545 1073 -5531
rect 1039 -5617 1073 -5599
rect 1039 -5689 1073 -5667
rect 1039 -5761 1073 -5735
rect 1039 -5833 1073 -5803
rect 1039 -5905 1073 -5871
rect 1039 -5973 1073 -5939
rect 1039 -6041 1073 -6011
rect 1039 -6109 1073 -6083
rect 1039 -6177 1073 -6155
rect 1039 -6245 1073 -6227
rect 1039 -6313 1073 -6299
rect 1039 -6381 1073 -6371
rect 1039 -6449 1073 -6443
rect 1039 -6517 1073 -6515
rect 1039 -6553 1073 -6551
rect 1039 -6625 1073 -6619
rect 1039 -6697 1073 -6687
rect 1039 -6769 1073 -6755
rect 1039 -6841 1073 -6823
rect 1039 -6913 1073 -6891
rect 1039 -6985 1073 -6959
rect 1039 -7057 1073 -7027
rect 1039 -7129 1073 -7095
rect 1039 -7197 1073 -7163
rect 1039 -7265 1073 -7235
rect 1039 -7333 1073 -7307
rect 1039 -7401 1073 -7379
rect 1039 -7469 1073 -7451
rect 1039 -7537 1073 -7523
rect 1039 -7605 1073 -7595
rect 1039 -7673 1073 -7667
rect 1039 -7741 1073 -7739
rect 1039 -7777 1073 -7775
rect 1039 -7849 1073 -7843
rect 1039 -7921 1073 -7911
rect 1039 -7993 1073 -7979
rect 1039 -8065 1073 -8047
rect 1039 -8137 1073 -8115
rect 1039 -8209 1073 -8183
rect 1039 -8281 1073 -8251
rect 1039 -8353 1073 -8319
rect 1039 -8421 1073 -8387
rect 1039 -8489 1073 -8459
rect 1039 -8557 1073 -8531
rect 1039 -8625 1073 -8603
rect 1039 -8693 1073 -8675
rect 1039 -8761 1073 -8747
rect 1039 -8829 1073 -8819
rect 1039 -8897 1073 -8891
rect 1039 -8965 1073 -8963
rect 1039 -9001 1073 -8999
rect 1039 -9073 1073 -9067
rect 1039 -9145 1073 -9135
rect 1039 -9217 1073 -9203
rect 1039 -9289 1073 -9271
rect 1039 -9361 1073 -9339
rect 1039 -9433 1073 -9407
rect 1039 -9506 1073 -9475
rect 1039 -9577 1073 -9543
rect 1039 -9645 1073 -9613
rect 28031 -3237 28065 -3203
rect 28031 -3305 28065 -3271
rect 28031 -3373 28065 -3339
rect 28031 -3441 28065 -3407
rect 28031 -3509 28065 -3475
rect 28031 -3577 28065 -3543
rect 28031 -3645 28065 -3611
rect 28031 -3713 28065 -3679
rect 28031 -3781 28065 -3747
rect 28031 -3849 28065 -3815
rect 28031 -3917 28065 -3883
rect 28031 -3985 28065 -3951
rect 28031 -4053 28065 -4019
rect 28031 -4121 28065 -4087
rect 28031 -4189 28065 -4155
rect 28031 -4257 28065 -4223
rect 28031 -4325 28065 -4291
rect 28031 -4393 28065 -4359
rect 28031 -4461 28065 -4427
rect 28031 -4529 28065 -4495
rect 28031 -4597 28065 -4563
rect 28031 -4665 28065 -4631
rect 28031 -4733 28065 -4699
rect 28031 -4801 28065 -4767
rect 28031 -4869 28065 -4835
rect 28031 -4937 28065 -4903
rect 28031 -5005 28065 -4971
rect 28031 -5073 28065 -5039
rect 28031 -5141 28065 -5107
rect 28031 -5209 28065 -5175
rect 28031 -5277 28065 -5243
rect 28031 -5345 28065 -5311
rect 28031 -5413 28065 -5379
rect 28031 -5481 28065 -5447
rect 28031 -5549 28065 -5515
rect 28031 -5617 28065 -5583
rect 28031 -5685 28065 -5651
rect 28031 -5753 28065 -5719
rect 28031 -5821 28065 -5787
rect 28031 -5889 28065 -5855
rect 28031 -5957 28065 -5923
rect 28031 -6025 28065 -5991
rect 28031 -6093 28065 -6059
rect 28031 -6161 28065 -6127
rect 28031 -6229 28065 -6195
rect 28031 -6297 28065 -6263
rect 28031 -6365 28065 -6331
rect 28031 -6433 28065 -6399
rect 28031 -6501 28065 -6467
rect 28031 -6569 28065 -6535
rect 28031 -6637 28065 -6603
rect 28031 -6705 28065 -6671
rect 28031 -6773 28065 -6739
rect 28031 -6841 28065 -6807
rect 28031 -6909 28065 -6875
rect 28031 -6977 28065 -6943
rect 28031 -7045 28065 -7011
rect 28031 -7113 28065 -7079
rect 28031 -7181 28065 -7147
rect 28031 -7249 28065 -7215
rect 28031 -7317 28065 -7283
rect 28031 -7385 28065 -7351
rect 28031 -7453 28065 -7419
rect 28031 -7521 28065 -7487
rect 28031 -7589 28065 -7555
rect 28031 -7657 28065 -7623
rect 28031 -7725 28065 -7691
rect 28031 -7793 28065 -7759
rect 28031 -7861 28065 -7827
rect 28031 -7929 28065 -7895
rect 28031 -7997 28065 -7963
rect 28031 -8065 28065 -8031
rect 28031 -8133 28065 -8099
rect 28031 -8201 28065 -8167
rect 28031 -8269 28065 -8235
rect 28031 -8337 28065 -8303
rect 28031 -8405 28065 -8371
rect 28031 -8473 28065 -8439
rect 28031 -8541 28065 -8507
rect 28031 -8609 28065 -8575
rect 28031 -8677 28065 -8643
rect 28031 -8745 28065 -8711
rect 28031 -8813 28065 -8779
rect 28031 -8881 28065 -8847
rect 28031 -8949 28065 -8915
rect 28031 -9017 28065 -8983
rect 28031 -9085 28065 -9051
rect 28031 -9153 28065 -9119
rect 28031 -9221 28065 -9187
rect 28031 -9289 28065 -9255
rect 28031 -9357 28065 -9323
rect 28031 -9425 28065 -9391
rect 28031 -9493 28065 -9459
rect 28031 -9561 28065 -9527
rect 1039 -9713 1073 -9686
rect 1039 -9781 1073 -9759
rect 1039 -9849 1073 -9832
rect 1039 -9917 1073 -9905
rect 1039 -9985 1073 -9978
rect 1039 -10053 1073 -10051
rect 1039 -10090 1073 -10087
rect 1039 -10163 1073 -10155
rect 2624 -9662 2658 -9658
rect 2624 -9698 2658 -9696
rect 2624 -9772 2658 -9764
rect 2624 -9846 2658 -9832
rect 2624 -9920 2658 -9900
rect 2624 -9994 2658 -9968
rect 2624 -10068 2658 -10036
rect 2624 -10138 2658 -10104
rect 2624 -10188 2658 -10176
rect 2780 -9662 2814 -9658
rect 2780 -9698 2814 -9696
rect 2780 -9772 2814 -9764
rect 2780 -9846 2814 -9832
rect 2780 -9920 2814 -9900
rect 2780 -9994 2814 -9968
rect 2780 -10068 2814 -10036
rect 2780 -10138 2814 -10104
rect 2780 -10188 2814 -10176
rect 2936 -9662 2970 -9658
rect 2936 -9698 2970 -9696
rect 2936 -9772 2970 -9764
rect 2936 -9846 2970 -9832
rect 2936 -9920 2970 -9900
rect 2936 -9994 2970 -9968
rect 2936 -10068 2970 -10036
rect 2936 -10138 2970 -10104
rect 2936 -10188 2970 -10176
rect 28031 -9629 28065 -9595
rect 28031 -9697 28065 -9663
rect 28031 -9765 28065 -9731
rect 28031 -9833 28065 -9799
rect 28031 -9901 28065 -9867
rect 28031 -9969 28065 -9935
rect 28031 -10037 28065 -10003
rect 28031 -10105 28065 -10071
rect 28031 -10173 28065 -10139
rect 1039 -10236 1073 -10223
rect 2669 -10266 2681 -10232
rect 2719 -10266 2780 -10232
rect 2814 -10266 2875 -10232
rect 2913 -10266 2925 -10232
rect 28031 -10241 28065 -10207
rect 1039 -10309 1073 -10291
rect 1039 -10382 1073 -10359
rect 1039 -10455 1073 -10427
rect 1039 -10528 1073 -10495
rect 1039 -10597 1073 -10563
rect 28031 -10309 28065 -10275
rect 28031 -10377 28065 -10343
rect 28031 -10445 28065 -10411
rect 28031 -10608 28065 -10479
rect 1039 -10665 1073 -10635
rect 23953 -10642 23987 -10608
rect 24021 -10642 24055 -10608
rect 24089 -10642 24123 -10608
rect 24157 -10642 24191 -10608
rect 24225 -10642 24259 -10608
rect 24293 -10642 24327 -10608
rect 24361 -10642 24395 -10608
rect 24429 -10642 24463 -10608
rect 24497 -10642 24531 -10608
rect 24565 -10642 24599 -10608
rect 24633 -10642 24667 -10608
rect 24701 -10642 24735 -10608
rect 24769 -10642 24803 -10608
rect 24837 -10642 24871 -10608
rect 24905 -10642 24939 -10608
rect 24973 -10642 25007 -10608
rect 25041 -10642 25075 -10608
rect 25109 -10642 25143 -10608
rect 25177 -10642 25211 -10608
rect 25245 -10642 25279 -10608
rect 25313 -10642 25347 -10608
rect 25381 -10642 25415 -10608
rect 25449 -10642 25483 -10608
rect 25517 -10642 25551 -10608
rect 25585 -10642 25619 -10608
rect 25653 -10642 25687 -10608
rect 25721 -10642 25755 -10608
rect 25789 -10642 25823 -10608
rect 25857 -10642 25891 -10608
rect 25925 -10642 25959 -10608
rect 25993 -10642 26027 -10608
rect 26061 -10642 26095 -10608
rect 26129 -10642 26163 -10608
rect 26197 -10642 26231 -10608
rect 26265 -10642 26299 -10608
rect 26333 -10642 26367 -10608
rect 26401 -10642 26435 -10608
rect 26469 -10642 26503 -10608
rect 26537 -10642 26571 -10608
rect 26605 -10642 26639 -10608
rect 26673 -10642 26707 -10608
rect 26741 -10642 26775 -10608
rect 26809 -10642 26843 -10608
rect 26877 -10642 26911 -10608
rect 26945 -10642 26979 -10608
rect 27013 -10642 27047 -10608
rect 27081 -10642 27115 -10608
rect 27149 -10642 27183 -10608
rect 27217 -10642 27251 -10608
rect 27285 -10642 27319 -10608
rect 27353 -10642 27387 -10608
rect 27421 -10642 27455 -10608
rect 27489 -10642 27523 -10608
rect 27557 -10642 27591 -10608
rect 27625 -10642 27659 -10608
rect 27693 -10642 27727 -10608
rect 27761 -10642 27795 -10608
rect 27829 -10642 27863 -10608
rect 27897 -10642 27931 -10608
rect 27965 -10642 28065 -10608
rect 1039 -10733 1073 -10708
rect 1039 -10801 1073 -10781
rect 406 -10857 407 -10852
rect 406 -10886 441 -10857
rect 440 -10895 441 -10886
rect 406 -10929 407 -10920
rect 548 -10918 582 -10880
rect 1039 -10869 1073 -10854
rect 406 -10954 441 -10929
rect 440 -10967 441 -10954
rect 532 -10956 548 -10922
rect 582 -10956 598 -10922
rect 1039 -10937 1073 -10927
rect 406 -11001 407 -10988
rect 406 -11039 441 -11001
rect 406 -11073 407 -11039
rect 1039 -11005 1073 -11000
rect 406 -11107 474 -11073
rect 508 -11107 542 -11073
rect 576 -11107 610 -11073
rect 644 -11107 678 -11073
rect 712 -11107 746 -11073
rect 780 -11107 814 -11073
rect 848 -11107 882 -11073
rect 916 -11107 950 -11073
rect 984 -11107 1073 -11073
rect 407 -11111 441 -11107
rect 1039 -11111 1073 -11107
rect 407 -11145 479 -11111
rect 513 -11145 559 -11111
rect 593 -11145 639 -11111
rect 673 -11145 719 -11111
rect 753 -11145 799 -11111
rect 833 -11145 879 -11111
rect 913 -11145 959 -11111
rect 993 -11145 1073 -11111
rect 18751 -11604 18923 -11593
rect 18751 -11638 18762 -11604
rect 18796 -11617 18923 -11604
rect 18796 -11638 18870 -11617
rect 18751 -11651 18870 -11638
rect 18904 -11651 18923 -11617
rect 18751 -11685 18923 -11651
rect 18751 -11692 18870 -11685
rect 18751 -11726 18762 -11692
rect 18796 -11719 18870 -11692
rect 18904 -11719 18923 -11685
rect 18796 -11726 18923 -11719
rect 18751 -11743 18923 -11726
rect 18874 -12867 18908 -12831
rect 18874 -12935 18908 -12901
rect 18874 -12985 18908 -12974
rect 3114 -17018 3179 -17011
rect 3213 -17018 3278 -17011
rect 3068 -17045 3080 -17018
rect 3068 -17052 3084 -17045
rect 3118 -17052 3179 -17018
rect 3213 -17052 3274 -17018
rect 3312 -17045 3324 -17018
rect 3308 -17052 3324 -17045
rect 3023 -17112 3057 -17096
rect 3023 -17180 3057 -17146
rect 3023 -17248 3057 -17214
rect 3023 -17316 3057 -17282
rect 3023 -17384 3057 -17350
rect 3023 -17428 3057 -17418
rect 3023 -17501 3057 -17486
rect 3023 -17575 3057 -17554
rect 3023 -17649 3057 -17622
rect 3179 -17112 3213 -17096
rect 3179 -17180 3213 -17146
rect 3179 -17248 3213 -17214
rect 3179 -17316 3213 -17282
rect 3179 -17384 3213 -17350
rect 3179 -17431 3213 -17418
rect 3179 -17503 3213 -17486
rect 3179 -17576 3213 -17554
rect 3179 -17649 3213 -17622
rect 3335 -17112 3369 -17096
rect 3335 -17180 3369 -17146
rect 3335 -17248 3369 -17214
rect 3335 -17316 3369 -17282
rect 3335 -17384 3369 -17350
rect 3335 -17428 3369 -17418
rect 3335 -17501 3369 -17486
rect 3335 -17575 3369 -17554
rect 3335 -17649 3369 -17622
rect 2625 -17867 2637 -17833
rect 2675 -17867 2736 -17833
rect 2771 -17867 2831 -17833
rect 2870 -17867 2881 -17833
rect 2580 -17985 2614 -17969
rect 2580 -18053 2614 -18019
rect 2580 -18114 2614 -18087
rect 2580 -18189 2614 -18155
rect 2580 -18257 2614 -18228
rect 2580 -18325 2614 -18308
rect 2580 -18393 2614 -18388
rect 2580 -18435 2614 -18427
rect 2580 -18516 2614 -18495
rect 2580 -18597 2614 -18563
rect 2580 -18665 2614 -18631
rect 2580 -18733 2614 -18712
rect 2580 -18801 2614 -18767
rect 2580 -18869 2614 -18835
rect 2580 -18919 2614 -18903
rect 2736 -17985 2770 -17969
rect 2736 -18053 2770 -18019
rect 2736 -18121 2770 -18087
rect 2736 -18189 2770 -18155
rect 2736 -18257 2770 -18248
rect 2736 -18325 2770 -18321
rect 2736 -18360 2770 -18359
rect 2736 -18433 2770 -18427
rect 2736 -18506 2770 -18495
rect 2736 -18579 2770 -18563
rect 2736 -18652 2770 -18631
rect 2736 -18725 2770 -18699
rect 2736 -18799 2770 -18767
rect 2736 -18869 2770 -18835
rect 2736 -18919 2770 -18907
rect 2892 -17985 2926 -17969
rect 2892 -18053 2926 -18019
rect 2892 -18114 2926 -18087
rect 2892 -18187 2926 -18155
rect 2892 -18257 2926 -18223
rect 2892 -18325 2926 -18294
rect 2892 -18393 2926 -18367
rect 2892 -18461 2926 -18440
rect 2892 -18529 2926 -18513
rect 2892 -18597 2926 -18586
rect 2892 -18665 2926 -18659
rect 2892 -18773 2926 -18767
rect 2892 -18869 2926 -18835
rect 2892 -18919 2926 -18903
<< viali >>
rect 539 4960 573 4994
rect 611 4971 645 4994
rect 683 4971 717 4994
rect 755 4971 789 4994
rect 827 4971 861 4994
rect 899 4971 933 4994
rect 971 4971 1005 4994
rect 1043 4971 1077 4994
rect 1115 4971 1149 4994
rect 1187 4971 1221 4994
rect 1259 4971 1293 4994
rect 1331 4971 1365 4994
rect 1403 4971 1437 4994
rect 1475 4971 1509 4994
rect 1547 4971 1581 4994
rect 1619 4971 1653 4994
rect 1691 4971 1725 4994
rect 1763 4971 1797 4994
rect 1835 4971 1869 4994
rect 1907 4971 1941 4994
rect 1979 4971 2013 4994
rect 2051 4971 2085 4994
rect 2123 4971 2157 4994
rect 2195 4971 2229 4994
rect 2267 4971 2301 4994
rect 2339 4971 2373 4994
rect 2411 4971 2445 4994
rect 2483 4971 2517 4994
rect 2555 4971 2589 4994
rect 2627 4971 2661 4994
rect 2699 4971 2733 4994
rect 2771 4971 2805 4994
rect 2843 4971 2877 4994
rect 2915 4971 2949 4994
rect 2987 4971 3021 4994
rect 3059 4971 3093 4994
rect 3131 4971 3165 4994
rect 3203 4971 3237 4994
rect 3275 4971 3309 4994
rect 3347 4971 3381 4994
rect 3419 4971 3453 4994
rect 3491 4971 3525 4994
rect 3563 4971 3597 4994
rect 3635 4971 3669 4994
rect 3707 4971 3741 4994
rect 3779 4971 3813 4994
rect 3851 4971 3885 4994
rect 3923 4971 3957 4994
rect 3995 4971 4029 4994
rect 4067 4971 4101 4994
rect 4139 4971 4173 4994
rect 4211 4971 4245 4994
rect 4283 4971 4317 4994
rect 4355 4971 4389 4994
rect 4427 4971 4461 4994
rect 4499 4971 4533 4994
rect 4571 4971 4605 4994
rect 4643 4971 4677 4994
rect 4715 4971 4749 4994
rect 4787 4971 4821 4994
rect 4859 4971 4893 4994
rect 4931 4971 4965 4994
rect 5003 4971 5037 4994
rect 5075 4971 5109 4994
rect 5147 4971 5181 4994
rect 5219 4971 5253 4994
rect 5291 4971 5325 4994
rect 5363 4971 5397 4994
rect 5435 4971 5469 4994
rect 5507 4971 5541 4994
rect 5579 4971 5613 4994
rect 5651 4971 5685 4994
rect 5723 4971 5757 4994
rect 5795 4971 5829 4994
rect 5868 4971 5902 4994
rect 5941 4971 5975 4994
rect 6014 4971 6048 4994
rect 6087 4971 6121 4994
rect 6160 4971 6194 4994
rect 6233 4971 6267 4994
rect 6306 4971 6340 4994
rect 6379 4971 6413 4994
rect 6452 4971 6486 4994
rect 6525 4971 6559 4994
rect 6598 4971 6632 4994
rect 6671 4971 6705 4994
rect 611 4960 624 4971
rect 624 4960 645 4971
rect 683 4960 692 4971
rect 692 4960 717 4971
rect 755 4960 760 4971
rect 760 4960 789 4971
rect 827 4960 828 4971
rect 828 4960 861 4971
rect 899 4960 930 4971
rect 930 4960 933 4971
rect 971 4960 998 4971
rect 998 4960 1005 4971
rect 1043 4960 1066 4971
rect 1066 4960 1077 4971
rect 1115 4960 1134 4971
rect 1134 4960 1149 4971
rect 1187 4960 1202 4971
rect 1202 4960 1221 4971
rect 1259 4960 1270 4971
rect 1270 4960 1293 4971
rect 1331 4960 1338 4971
rect 1338 4960 1365 4971
rect 1403 4960 1406 4971
rect 1406 4960 1437 4971
rect 1475 4960 1508 4971
rect 1508 4960 1509 4971
rect 1547 4960 1576 4971
rect 1576 4960 1581 4971
rect 1619 4960 1644 4971
rect 1644 4960 1653 4971
rect 1691 4960 1712 4971
rect 1712 4960 1725 4971
rect 1763 4960 1780 4971
rect 1780 4960 1797 4971
rect 1835 4960 1848 4971
rect 1848 4960 1869 4971
rect 1907 4960 1916 4971
rect 1916 4960 1941 4971
rect 1979 4960 1984 4971
rect 1984 4960 2013 4971
rect 2051 4960 2052 4971
rect 2052 4960 2085 4971
rect 2123 4960 2154 4971
rect 2154 4960 2157 4971
rect 2195 4960 2222 4971
rect 2222 4960 2229 4971
rect 2267 4960 2290 4971
rect 2290 4960 2301 4971
rect 2339 4960 2358 4971
rect 2358 4960 2373 4971
rect 2411 4960 2426 4971
rect 2426 4960 2445 4971
rect 2483 4960 2494 4971
rect 2494 4960 2517 4971
rect 2555 4960 2562 4971
rect 2562 4960 2589 4971
rect 2627 4960 2630 4971
rect 2630 4960 2661 4971
rect 2699 4960 2732 4971
rect 2732 4960 2733 4971
rect 2771 4960 2800 4971
rect 2800 4960 2805 4971
rect 2843 4960 2868 4971
rect 2868 4960 2877 4971
rect 2915 4960 2936 4971
rect 2936 4960 2949 4971
rect 2987 4960 3004 4971
rect 3004 4960 3021 4971
rect 3059 4960 3072 4971
rect 3072 4960 3093 4971
rect 3131 4960 3140 4971
rect 3140 4960 3165 4971
rect 3203 4960 3208 4971
rect 3208 4960 3237 4971
rect 3275 4960 3276 4971
rect 3276 4960 3309 4971
rect 3347 4960 3378 4971
rect 3378 4960 3381 4971
rect 3419 4960 3446 4971
rect 3446 4960 3453 4971
rect 3491 4960 3514 4971
rect 3514 4960 3525 4971
rect 3563 4960 3582 4971
rect 3582 4960 3597 4971
rect 3635 4960 3650 4971
rect 3650 4960 3669 4971
rect 3707 4960 3718 4971
rect 3718 4960 3741 4971
rect 3779 4960 3786 4971
rect 3786 4960 3813 4971
rect 3851 4960 3854 4971
rect 3854 4960 3885 4971
rect 3923 4960 3956 4971
rect 3956 4960 3957 4971
rect 3995 4960 4024 4971
rect 4024 4960 4029 4971
rect 4067 4960 4092 4971
rect 4092 4960 4101 4971
rect 4139 4960 4160 4971
rect 4160 4960 4173 4971
rect 4211 4960 4228 4971
rect 4228 4960 4245 4971
rect 4283 4960 4296 4971
rect 4296 4960 4317 4971
rect 4355 4960 4364 4971
rect 4364 4960 4389 4971
rect 4427 4960 4432 4971
rect 4432 4960 4461 4971
rect 4499 4960 4500 4971
rect 4500 4960 4533 4971
rect 4571 4960 4602 4971
rect 4602 4960 4605 4971
rect 4643 4960 4670 4971
rect 4670 4960 4677 4971
rect 4715 4960 4738 4971
rect 4738 4960 4749 4971
rect 4787 4960 4806 4971
rect 4806 4960 4821 4971
rect 4859 4960 4874 4971
rect 4874 4960 4893 4971
rect 4931 4960 4942 4971
rect 4942 4960 4965 4971
rect 5003 4960 5010 4971
rect 5010 4960 5037 4971
rect 5075 4960 5078 4971
rect 5078 4960 5109 4971
rect 5147 4960 5180 4971
rect 5180 4960 5181 4971
rect 5219 4960 5248 4971
rect 5248 4960 5253 4971
rect 5291 4960 5316 4971
rect 5316 4960 5325 4971
rect 5363 4960 5384 4971
rect 5384 4960 5397 4971
rect 5435 4960 5452 4971
rect 5452 4960 5469 4971
rect 5507 4960 5520 4971
rect 5520 4960 5541 4971
rect 5579 4960 5588 4971
rect 5588 4960 5613 4971
rect 5651 4960 5656 4971
rect 5656 4960 5685 4971
rect 5723 4960 5724 4971
rect 5724 4960 5757 4971
rect 5795 4960 5826 4971
rect 5826 4960 5829 4971
rect 5868 4960 5894 4971
rect 5894 4960 5902 4971
rect 5941 4960 5962 4971
rect 5962 4960 5975 4971
rect 6014 4960 6030 4971
rect 6030 4960 6048 4971
rect 6087 4960 6098 4971
rect 6098 4960 6121 4971
rect 6160 4960 6166 4971
rect 6166 4960 6194 4971
rect 6233 4960 6234 4971
rect 6234 4960 6267 4971
rect 6306 4960 6336 4971
rect 6336 4960 6340 4971
rect 6379 4960 6404 4971
rect 6404 4960 6413 4971
rect 6452 4960 6472 4971
rect 6472 4960 6486 4971
rect 6525 4960 6540 4971
rect 6540 4960 6559 4971
rect 6598 4960 6608 4971
rect 6608 4960 6632 4971
rect 6671 4960 6676 4971
rect 6676 4960 6705 4971
rect 6744 4960 6778 4994
rect 6817 4971 6851 4994
rect 6890 4971 6924 4994
rect 6963 4971 6997 4994
rect 7036 4971 7070 4994
rect 7109 4971 7143 4994
rect 7182 4971 7216 4994
rect 7255 4971 7289 4994
rect 7328 4971 7362 4994
rect 7401 4971 7435 4994
rect 7474 4971 7508 4994
rect 7547 4971 7581 4994
rect 7620 4971 7654 4994
rect 7693 4971 7727 4994
rect 6817 4960 6846 4971
rect 6846 4960 6851 4971
rect 6890 4960 6914 4971
rect 6914 4960 6924 4971
rect 6963 4960 6982 4971
rect 6982 4960 6997 4971
rect 7036 4960 7050 4971
rect 7050 4960 7070 4971
rect 7109 4960 7118 4971
rect 7118 4960 7143 4971
rect 7182 4960 7186 4971
rect 7186 4960 7216 4971
rect 7255 4960 7288 4971
rect 7288 4960 7289 4971
rect 7328 4960 7356 4971
rect 7356 4960 7362 4971
rect 7401 4960 7424 4971
rect 7424 4960 7435 4971
rect 7474 4960 7492 4971
rect 7492 4960 7508 4971
rect 7547 4960 7560 4971
rect 7560 4960 7581 4971
rect 7620 4960 7628 4971
rect 7628 4960 7654 4971
rect 7693 4960 7696 4971
rect 7696 4960 7727 4971
rect 7766 4960 7800 4994
rect 467 4888 501 4922
rect 467 4813 501 4847
rect 7838 4903 7872 4920
rect 7838 4886 7872 4903
rect 7838 4835 7872 4846
rect 663 4791 697 4823
rect 467 4738 501 4772
rect 663 4789 679 4791
rect 679 4789 697 4791
rect 663 4721 697 4740
rect 467 4663 501 4697
rect 663 4706 679 4721
rect 679 4706 697 4721
rect 871 4807 905 4823
rect 871 4789 905 4807
rect 871 4717 905 4751
rect 1727 4807 1761 4823
rect 1727 4789 1761 4807
rect 1727 4717 1761 4751
rect 1983 4807 2017 4823
rect 1983 4789 2017 4807
rect 1983 4717 2017 4751
rect 2239 4807 2273 4823
rect 2239 4789 2273 4807
rect 2239 4717 2273 4751
rect 2495 4807 2529 4823
rect 2495 4789 2529 4807
rect 2495 4717 2529 4751
rect 2751 4807 2785 4823
rect 2751 4789 2785 4807
rect 2751 4717 2785 4751
rect 3007 4807 3041 4823
rect 3007 4789 3041 4807
rect 3007 4717 3041 4751
rect 3263 4807 3297 4823
rect 3263 4789 3297 4807
rect 3263 4717 3297 4751
rect 3519 4807 3553 4823
rect 3519 4789 3553 4807
rect 3519 4717 3553 4751
rect 3775 4807 3809 4823
rect 3775 4789 3809 4807
rect 3775 4717 3809 4751
rect 4031 4807 4065 4823
rect 4031 4789 4065 4807
rect 4031 4717 4065 4751
rect 4287 4807 4321 4823
rect 4287 4789 4321 4807
rect 4287 4717 4321 4751
rect 4543 4807 4577 4823
rect 4543 4789 4577 4807
rect 4543 4717 4577 4751
rect 4799 4807 4833 4823
rect 4799 4789 4833 4807
rect 4799 4717 4833 4751
rect 5055 4807 5089 4823
rect 5055 4789 5089 4807
rect 5055 4717 5089 4751
rect 5311 4807 5345 4823
rect 5311 4789 5345 4807
rect 5311 4717 5345 4751
rect 5567 4807 5601 4823
rect 5567 4789 5601 4807
rect 5567 4717 5601 4751
rect 5823 4807 5857 4823
rect 5823 4789 5857 4807
rect 5823 4717 5857 4751
rect 6079 4807 6113 4823
rect 6079 4789 6113 4807
rect 6079 4717 6113 4751
rect 6335 4807 6369 4823
rect 6335 4789 6369 4807
rect 6335 4717 6369 4751
rect 6591 4807 6625 4823
rect 6591 4789 6625 4807
rect 6591 4717 6625 4751
rect 6847 4807 6881 4823
rect 6847 4789 6881 4807
rect 6847 4717 6881 4751
rect 7703 4807 7737 4823
rect 7703 4789 7737 4807
rect 7703 4717 7737 4751
rect 7838 4812 7872 4835
rect 7838 4767 7872 4772
rect 7838 4738 7872 4767
rect 7838 4665 7872 4698
rect 7838 4664 7872 4665
rect 663 4651 697 4657
rect 467 4588 501 4622
rect 663 4623 679 4651
rect 679 4623 697 4651
rect 928 4627 932 4652
rect 932 4627 962 4652
rect 1006 4627 1037 4652
rect 1037 4627 1040 4652
rect 1084 4627 1108 4652
rect 1108 4627 1118 4652
rect 1162 4627 1179 4652
rect 1179 4627 1196 4652
rect 1239 4627 1250 4652
rect 1250 4627 1273 4652
rect 1316 4627 1321 4652
rect 1321 4627 1350 4652
rect 928 4618 962 4627
rect 1006 4618 1040 4627
rect 1084 4618 1118 4627
rect 1162 4618 1196 4627
rect 1239 4618 1273 4627
rect 1316 4618 1350 4627
rect 1393 4618 1427 4652
rect 1470 4627 1500 4652
rect 1500 4627 1504 4652
rect 1547 4627 1571 4652
rect 1571 4627 1581 4652
rect 1624 4627 1642 4652
rect 1642 4627 1658 4652
rect 2051 4627 2078 4661
rect 2078 4627 2085 4661
rect 2130 4627 2146 4661
rect 2146 4627 2164 4661
rect 2342 4627 2350 4661
rect 2350 4627 2376 4661
rect 2421 4627 2452 4661
rect 2452 4627 2455 4661
rect 2500 4627 2520 4661
rect 2520 4627 2534 4661
rect 2578 4627 2588 4661
rect 2588 4627 2612 4661
rect 2656 4627 2690 4661
rect 2837 4627 2860 4661
rect 2860 4627 2871 4661
rect 2922 4627 2928 4661
rect 2928 4627 2956 4661
rect 3007 4627 3030 4661
rect 3030 4627 3041 4661
rect 3091 4627 3098 4661
rect 3098 4627 3125 4661
rect 3175 4627 3202 4661
rect 3202 4627 3209 4661
rect 3385 4627 3419 4661
rect 3462 4627 3492 4661
rect 3492 4627 3496 4661
rect 3576 4627 3580 4661
rect 3580 4627 3610 4661
rect 3691 4627 3716 4661
rect 3716 4627 3725 4661
rect 3858 4627 3886 4661
rect 3886 4627 3892 4661
rect 3945 4627 3954 4661
rect 3954 4627 3979 4661
rect 4032 4627 4056 4661
rect 4056 4627 4066 4661
rect 4119 4627 4124 4661
rect 4124 4627 4153 4661
rect 4206 4627 4226 4661
rect 4226 4627 4240 4661
rect 4371 4627 4396 4661
rect 4396 4627 4405 4661
rect 4457 4627 4464 4661
rect 4464 4627 4491 4661
rect 4543 4627 4566 4661
rect 4566 4627 4577 4661
rect 4629 4627 4634 4661
rect 4634 4627 4663 4661
rect 4715 4627 4736 4661
rect 4736 4627 4749 4661
rect 4881 4627 4906 4661
rect 4906 4627 4915 4661
rect 4955 4627 4974 4661
rect 4974 4627 4989 4661
rect 5029 4627 5042 4661
rect 5042 4627 5063 4661
rect 5102 4627 5110 4661
rect 5110 4627 5136 4661
rect 5175 4627 5178 4661
rect 5178 4627 5209 4661
rect 5248 4627 5280 4661
rect 5280 4627 5282 4661
rect 5321 4627 5348 4661
rect 5348 4627 5355 4661
rect 5394 4627 5416 4661
rect 5416 4627 5428 4661
rect 5467 4627 5484 4661
rect 5484 4627 5501 4661
rect 5540 4627 5552 4661
rect 5552 4627 5574 4661
rect 5613 4627 5620 4661
rect 5620 4627 5647 4661
rect 5686 4627 5688 4661
rect 5688 4627 5720 4661
rect 5759 4627 5790 4661
rect 5790 4627 5793 4661
rect 5832 4627 5858 4661
rect 5858 4627 5866 4661
rect 5905 4627 5926 4661
rect 5926 4627 5939 4661
rect 5978 4627 5994 4661
rect 5994 4627 6012 4661
rect 6051 4627 6062 4661
rect 6062 4627 6085 4661
rect 6124 4627 6130 4661
rect 6130 4627 6158 4661
rect 6197 4627 6199 4661
rect 6199 4627 6231 4661
rect 6270 4627 6303 4661
rect 6303 4627 6304 4661
rect 6343 4627 6372 4661
rect 6372 4627 6377 4661
rect 6416 4627 6441 4661
rect 6441 4627 6450 4661
rect 6489 4627 6510 4661
rect 6510 4627 6523 4661
rect 7066 4627 7080 4652
rect 7080 4627 7100 4652
rect 7150 4627 7184 4652
rect 7235 4627 7254 4652
rect 7254 4627 7269 4652
rect 7320 4627 7324 4652
rect 7324 4627 7354 4652
rect 7405 4627 7430 4652
rect 7430 4627 7439 4652
rect 7490 4627 7500 4652
rect 7500 4627 7524 4652
rect 1470 4618 1504 4627
rect 1547 4618 1581 4627
rect 1624 4618 1658 4627
rect 7066 4618 7100 4627
rect 7150 4618 7184 4627
rect 7235 4618 7269 4627
rect 7320 4618 7354 4627
rect 7405 4618 7439 4627
rect 7490 4618 7524 4627
rect 467 4513 501 4547
rect 467 4438 501 4472
rect 7838 4597 7872 4624
rect 7838 4590 7872 4597
rect 7838 4529 7872 4550
rect 7838 4516 7872 4529
rect 660 4477 679 4486
rect 679 4477 694 4486
rect 928 4483 962 4492
rect 1006 4483 1040 4492
rect 1084 4483 1118 4492
rect 1162 4483 1196 4492
rect 1239 4483 1273 4492
rect 1316 4483 1350 4492
rect 1393 4483 1427 4492
rect 1470 4483 1504 4492
rect 1547 4483 1581 4492
rect 1624 4483 1658 4492
rect 1789 4483 1823 4486
rect 1865 4483 1899 4486
rect 1941 4483 1975 4486
rect 2017 4483 2051 4486
rect 2093 4483 2127 4486
rect 2169 4483 2203 4486
rect 2244 4483 2278 4486
rect 2319 4483 2353 4486
rect 2394 4483 2428 4486
rect 2469 4483 2503 4486
rect 2544 4483 2578 4486
rect 2619 4483 2653 4486
rect 2694 4483 2728 4486
rect 2769 4483 2803 4486
rect 2844 4483 2878 4486
rect 2919 4483 2953 4486
rect 3095 4483 3129 4486
rect 3173 4483 3207 4486
rect 3251 4483 3285 4486
rect 3329 4483 3363 4486
rect 3407 4483 3441 4486
rect 3485 4483 3519 4486
rect 3563 4483 3597 4486
rect 3641 4483 3675 4486
rect 3718 4483 3752 4486
rect 3832 4483 3866 4486
rect 660 4452 694 4477
rect 928 4458 932 4483
rect 932 4458 962 4483
rect 1006 4458 1040 4483
rect 1084 4458 1114 4483
rect 1114 4458 1118 4483
rect 1162 4458 1188 4483
rect 1188 4458 1196 4483
rect 1239 4458 1262 4483
rect 1262 4458 1273 4483
rect 1316 4458 1335 4483
rect 1335 4458 1350 4483
rect 1393 4458 1408 4483
rect 1408 4458 1427 4483
rect 1470 4458 1481 4483
rect 1481 4458 1504 4483
rect 1547 4458 1554 4483
rect 1554 4458 1581 4483
rect 1624 4458 1627 4483
rect 1627 4458 1658 4483
rect 1789 4452 1822 4483
rect 1822 4452 1823 4483
rect 1865 4452 1890 4483
rect 1890 4452 1899 4483
rect 1941 4452 1958 4483
rect 1958 4452 1975 4483
rect 2017 4452 2026 4483
rect 2026 4452 2051 4483
rect 2093 4452 2094 4483
rect 2094 4452 2127 4483
rect 2169 4452 2196 4483
rect 2196 4452 2203 4483
rect 2244 4452 2265 4483
rect 2265 4452 2278 4483
rect 2319 4452 2334 4483
rect 2334 4452 2353 4483
rect 2394 4452 2403 4483
rect 2403 4452 2428 4483
rect 2469 4452 2472 4483
rect 2472 4452 2503 4483
rect 2544 4452 2575 4483
rect 2575 4452 2578 4483
rect 2619 4452 2644 4483
rect 2644 4452 2653 4483
rect 2694 4452 2713 4483
rect 2713 4452 2728 4483
rect 2769 4452 2782 4483
rect 2782 4452 2803 4483
rect 2844 4452 2851 4483
rect 2851 4452 2878 4483
rect 2919 4452 2920 4483
rect 2920 4452 2953 4483
rect 3095 4452 3127 4483
rect 3127 4452 3129 4483
rect 3173 4452 3196 4483
rect 3196 4452 3207 4483
rect 3251 4452 3265 4483
rect 3265 4452 3285 4483
rect 3329 4452 3334 4483
rect 3334 4452 3363 4483
rect 3407 4452 3438 4483
rect 3438 4452 3441 4483
rect 3485 4452 3507 4483
rect 3507 4452 3519 4483
rect 3563 4452 3576 4483
rect 3576 4452 3597 4483
rect 3641 4452 3645 4483
rect 3645 4452 3675 4483
rect 3718 4452 3748 4483
rect 3748 4452 3752 4483
rect 3832 4452 3836 4483
rect 3836 4452 3866 4483
rect 3929 4452 3963 4486
rect 4133 4452 4167 4486
rect 4230 4483 4264 4486
rect 4344 4483 4378 4486
rect 4451 4483 4485 4486
rect 4600 4483 4634 4486
rect 4675 4483 4709 4486
rect 4750 4483 4784 4486
rect 4825 4483 4859 4486
rect 4900 4483 4934 4486
rect 4975 4483 5009 4486
rect 5050 4483 5084 4486
rect 5125 4483 5159 4486
rect 5199 4483 5233 4486
rect 5273 4483 5307 4486
rect 5347 4483 5381 4486
rect 5421 4483 5455 4486
rect 5495 4483 5529 4486
rect 5569 4483 5603 4486
rect 5643 4483 5677 4486
rect 5717 4483 5751 4486
rect 5791 4483 5825 4486
rect 5865 4483 5899 4486
rect 5939 4483 5973 4486
rect 4230 4452 4260 4483
rect 4260 4452 4264 4483
rect 4344 4452 4348 4483
rect 4348 4452 4378 4483
rect 4451 4452 4482 4483
rect 4482 4452 4485 4483
rect 4600 4452 4604 4483
rect 4604 4452 4634 4483
rect 4675 4452 4706 4483
rect 4706 4452 4709 4483
rect 4750 4452 4774 4483
rect 4774 4452 4784 4483
rect 4825 4452 4842 4483
rect 4842 4452 4859 4483
rect 4900 4452 4910 4483
rect 4910 4452 4934 4483
rect 4975 4452 4978 4483
rect 4978 4452 5009 4483
rect 5050 4452 5082 4483
rect 5082 4452 5084 4483
rect 5125 4452 5151 4483
rect 5151 4452 5159 4483
rect 5199 4452 5220 4483
rect 5220 4452 5233 4483
rect 5273 4452 5289 4483
rect 5289 4452 5307 4483
rect 5347 4452 5358 4483
rect 5358 4452 5381 4483
rect 5421 4452 5427 4483
rect 5427 4452 5455 4483
rect 5495 4452 5496 4483
rect 5496 4452 5529 4483
rect 5569 4452 5599 4483
rect 5599 4452 5603 4483
rect 5643 4452 5668 4483
rect 5668 4452 5677 4483
rect 5717 4452 5737 4483
rect 5737 4452 5751 4483
rect 5791 4452 5806 4483
rect 5806 4452 5825 4483
rect 5865 4452 5875 4483
rect 5875 4452 5899 4483
rect 5939 4452 5944 4483
rect 5944 4452 5973 4483
rect 6013 4452 6047 4486
rect 6087 4483 6121 4486
rect 6161 4483 6195 4486
rect 6235 4483 6269 4486
rect 6309 4483 6343 4486
rect 6383 4483 6417 4486
rect 6457 4483 6491 4486
rect 6531 4483 6565 4486
rect 7066 4483 7100 4492
rect 7138 4483 7172 4492
rect 7210 4483 7244 4492
rect 7282 4483 7316 4492
rect 7355 4483 7389 4492
rect 7428 4483 7462 4492
rect 7501 4483 7535 4492
rect 7574 4483 7608 4492
rect 7647 4483 7681 4492
rect 6087 4452 6117 4483
rect 6117 4452 6121 4483
rect 6161 4452 6186 4483
rect 6186 4452 6195 4483
rect 6235 4452 6255 4483
rect 6255 4452 6269 4483
rect 6309 4452 6324 4483
rect 6324 4452 6343 4483
rect 6383 4452 6393 4483
rect 6393 4452 6417 4483
rect 6457 4452 6462 4483
rect 6462 4452 6491 4483
rect 6531 4452 6565 4483
rect 7066 4458 7074 4483
rect 7074 4458 7100 4483
rect 7138 4458 7145 4483
rect 7145 4458 7172 4483
rect 7210 4458 7216 4483
rect 7216 4458 7244 4483
rect 7282 4458 7287 4483
rect 7287 4458 7316 4483
rect 7355 4458 7358 4483
rect 7358 4458 7389 4483
rect 7428 4458 7429 4483
rect 7429 4458 7462 4483
rect 7501 4458 7534 4483
rect 7534 4458 7535 4483
rect 7574 4458 7605 4483
rect 7605 4458 7608 4483
rect 7647 4458 7676 4483
rect 7676 4458 7681 4483
rect 7838 4461 7872 4475
rect 467 4363 501 4397
rect 660 4371 694 4404
rect 7838 4441 7872 4461
rect 7838 4393 7872 4400
rect 467 4288 501 4322
rect 660 4370 679 4371
rect 679 4370 694 4371
rect 660 4301 694 4321
rect 660 4287 679 4301
rect 679 4287 694 4301
rect 871 4359 905 4393
rect 871 4303 905 4321
rect 871 4287 905 4303
rect 1727 4359 1761 4393
rect 1727 4303 1761 4321
rect 1727 4287 1761 4303
rect 1983 4359 2017 4393
rect 1983 4303 2017 4321
rect 1983 4287 2017 4303
rect 2239 4359 2273 4393
rect 2239 4303 2273 4321
rect 2239 4287 2273 4303
rect 2495 4359 2529 4393
rect 2495 4303 2529 4321
rect 2495 4287 2529 4303
rect 2751 4359 2785 4393
rect 2751 4303 2785 4321
rect 2751 4287 2785 4303
rect 3007 4359 3041 4393
rect 3007 4303 3041 4321
rect 3007 4287 3041 4303
rect 3263 4359 3297 4393
rect 3263 4303 3297 4321
rect 3263 4287 3297 4303
rect 3519 4359 3553 4393
rect 3519 4303 3553 4321
rect 3519 4287 3553 4303
rect 3775 4359 3809 4393
rect 3775 4303 3809 4321
rect 3775 4287 3809 4303
rect 4031 4359 4065 4393
rect 4031 4303 4065 4321
rect 4031 4287 4065 4303
rect 4287 4359 4321 4393
rect 4287 4303 4321 4321
rect 4287 4287 4321 4303
rect 4543 4359 4577 4393
rect 4543 4303 4577 4321
rect 4543 4287 4577 4303
rect 4799 4359 4833 4393
rect 4799 4303 4833 4321
rect 4799 4287 4833 4303
rect 5055 4359 5089 4393
rect 5055 4303 5089 4321
rect 5055 4287 5089 4303
rect 5311 4359 5345 4393
rect 5311 4303 5345 4321
rect 5311 4287 5345 4303
rect 5567 4359 5601 4393
rect 5567 4303 5601 4321
rect 5567 4287 5601 4303
rect 5823 4359 5857 4393
rect 5823 4303 5857 4321
rect 5823 4287 5857 4303
rect 6079 4359 6113 4393
rect 6079 4303 6113 4321
rect 6079 4287 6113 4303
rect 6335 4359 6369 4393
rect 6335 4303 6369 4321
rect 6335 4287 6369 4303
rect 6591 4359 6625 4393
rect 6591 4303 6625 4321
rect 6591 4287 6625 4303
rect 6847 4359 6881 4393
rect 6847 4303 6881 4321
rect 6847 4287 6881 4303
rect 7703 4359 7737 4393
rect 7703 4303 7737 4321
rect 7703 4287 7737 4303
rect 7838 4366 7872 4393
rect 7838 4291 7872 4325
rect 467 4213 501 4247
rect 467 4138 501 4172
rect 467 4063 501 4097
rect 467 3988 501 4022
rect 467 3913 501 3947
rect 467 3838 501 3872
rect 7838 4223 7872 4250
rect 7838 4216 7872 4223
rect 7838 4155 7872 4175
rect 7838 4141 7872 4155
rect 7838 4087 7872 4100
rect 7838 4066 7872 4087
rect 7838 4019 7872 4025
rect 7838 3991 7872 4019
rect 7838 3917 7872 3950
rect 7838 3916 7872 3917
rect 7838 3849 7872 3875
rect 7838 3841 7872 3849
rect 467 3763 501 3797
rect 660 3806 694 3813
rect 660 3779 679 3806
rect 679 3779 694 3806
rect 467 3688 501 3722
rect 660 3701 679 3731
rect 679 3701 694 3731
rect 871 3797 905 3813
rect 871 3779 905 3797
rect 871 3707 905 3741
rect 1727 3797 1761 3813
rect 1727 3779 1761 3797
rect 1727 3707 1761 3741
rect 1983 3797 2017 3813
rect 1983 3779 2017 3797
rect 1983 3707 2017 3741
rect 2239 3797 2273 3813
rect 2239 3779 2273 3797
rect 2239 3707 2273 3741
rect 2495 3797 2529 3813
rect 2495 3779 2529 3797
rect 2495 3707 2529 3741
rect 2751 3797 2785 3813
rect 2751 3779 2785 3797
rect 2751 3707 2785 3741
rect 3007 3797 3041 3813
rect 3007 3779 3041 3797
rect 3007 3707 3041 3741
rect 3263 3797 3297 3813
rect 3263 3779 3297 3797
rect 3263 3707 3297 3741
rect 3519 3797 3553 3813
rect 3519 3779 3553 3797
rect 3519 3707 3553 3741
rect 3775 3797 3809 3813
rect 3775 3779 3809 3797
rect 3775 3707 3809 3741
rect 4031 3797 4065 3813
rect 4031 3779 4065 3797
rect 4031 3707 4065 3741
rect 4287 3797 4321 3813
rect 4287 3779 4321 3797
rect 4287 3707 4321 3741
rect 4543 3797 4577 3813
rect 4543 3779 4577 3797
rect 4543 3707 4577 3741
rect 4799 3797 4833 3813
rect 4799 3779 4833 3797
rect 4799 3707 4833 3741
rect 5055 3797 5089 3813
rect 5055 3779 5089 3797
rect 5055 3707 5089 3741
rect 5311 3797 5345 3813
rect 5311 3779 5345 3797
rect 5311 3707 5345 3741
rect 5567 3797 5601 3813
rect 5567 3779 5601 3797
rect 5567 3707 5601 3741
rect 5823 3797 5857 3813
rect 5823 3779 5857 3797
rect 5823 3707 5857 3741
rect 6079 3797 6113 3813
rect 6079 3779 6113 3797
rect 6079 3707 6113 3741
rect 6335 3797 6369 3813
rect 6335 3779 6369 3797
rect 6335 3707 6369 3741
rect 6591 3797 6625 3813
rect 6591 3779 6625 3797
rect 6591 3707 6625 3741
rect 6847 3797 6881 3813
rect 6847 3779 6881 3797
rect 6847 3707 6881 3741
rect 7703 3797 7737 3813
rect 7703 3779 7737 3797
rect 7703 3707 7737 3741
rect 7838 3781 7872 3800
rect 7838 3766 7872 3781
rect 660 3697 694 3701
rect 467 3613 501 3647
rect 7838 3691 7872 3725
rect 660 3630 679 3648
rect 679 3630 694 3648
rect 660 3614 694 3630
rect 928 3617 932 3642
rect 932 3617 962 3642
rect 1006 3617 1037 3642
rect 1037 3617 1040 3642
rect 1084 3617 1108 3642
rect 1108 3617 1118 3642
rect 1162 3617 1179 3642
rect 1179 3617 1196 3642
rect 1239 3617 1250 3642
rect 1250 3617 1273 3642
rect 1316 3617 1321 3642
rect 1321 3617 1350 3642
rect 928 3608 962 3617
rect 1006 3608 1040 3617
rect 1084 3608 1118 3617
rect 1162 3608 1196 3617
rect 1239 3608 1273 3617
rect 1316 3608 1350 3617
rect 1393 3608 1427 3642
rect 1470 3617 1500 3642
rect 1500 3617 1504 3642
rect 1547 3617 1571 3642
rect 1571 3617 1581 3642
rect 1624 3617 1642 3642
rect 1642 3617 1658 3642
rect 2557 3617 2590 3645
rect 2590 3617 2591 3645
rect 2633 3617 2659 3645
rect 2659 3617 2667 3645
rect 2709 3617 2728 3645
rect 2728 3617 2743 3645
rect 2785 3617 2797 3645
rect 2797 3617 2819 3645
rect 2861 3617 2866 3645
rect 2866 3617 2895 3645
rect 2936 3617 2969 3645
rect 2969 3617 2970 3645
rect 3011 3617 3038 3645
rect 3038 3617 3045 3645
rect 3086 3617 3107 3645
rect 3107 3617 3120 3645
rect 3161 3617 3176 3645
rect 3176 3617 3195 3645
rect 3236 3617 3245 3645
rect 3245 3617 3270 3645
rect 3311 3617 3314 3645
rect 3314 3617 3345 3645
rect 3386 3617 3418 3645
rect 3418 3617 3420 3645
rect 3461 3617 3487 3645
rect 3487 3617 3495 3645
rect 3536 3617 3556 3645
rect 3556 3617 3570 3645
rect 3611 3617 3625 3645
rect 3625 3617 3645 3645
rect 3686 3617 3694 3645
rect 3694 3617 3720 3645
rect 3761 3617 3763 3645
rect 3763 3617 3795 3645
rect 3836 3617 3866 3645
rect 3866 3617 3870 3645
rect 3911 3617 3935 3645
rect 3935 3617 3945 3645
rect 3986 3617 4004 3645
rect 4004 3617 4020 3645
rect 4088 3617 4092 3648
rect 4092 3617 4122 3648
rect 4195 3617 4226 3648
rect 4226 3617 4229 3648
rect 4332 3617 4348 3645
rect 4348 3617 4366 3645
rect 1470 3608 1504 3617
rect 1547 3608 1581 3617
rect 1624 3608 1658 3617
rect 2557 3611 2591 3617
rect 2633 3611 2667 3617
rect 2709 3611 2743 3617
rect 2785 3611 2819 3617
rect 2861 3611 2895 3617
rect 2936 3611 2970 3617
rect 3011 3611 3045 3617
rect 3086 3611 3120 3617
rect 3161 3611 3195 3617
rect 3236 3611 3270 3617
rect 3311 3611 3345 3617
rect 3386 3611 3420 3617
rect 3461 3611 3495 3617
rect 3536 3611 3570 3617
rect 3611 3611 3645 3617
rect 3686 3611 3720 3617
rect 3761 3611 3795 3617
rect 3836 3611 3870 3617
rect 3911 3611 3945 3617
rect 3986 3611 4020 3617
rect 4088 3614 4122 3617
rect 4195 3614 4229 3617
rect 4332 3611 4366 3617
rect 4445 3611 4479 3645
rect 4641 3614 4675 3648
rect 4742 3617 4772 3648
rect 4772 3617 4776 3648
rect 4844 3617 4860 3645
rect 4860 3617 4878 3645
rect 4916 3617 4929 3645
rect 4929 3617 4950 3645
rect 4988 3617 4998 3645
rect 4998 3617 5022 3645
rect 5060 3617 5067 3645
rect 5067 3617 5094 3645
rect 5132 3617 5136 3645
rect 5136 3617 5166 3645
rect 5204 3617 5205 3645
rect 5205 3617 5238 3645
rect 5276 3617 5308 3645
rect 5308 3617 5310 3645
rect 5348 3617 5377 3645
rect 5377 3617 5382 3645
rect 5420 3617 5446 3645
rect 5446 3617 5454 3645
rect 5492 3617 5515 3645
rect 5515 3617 5526 3645
rect 5564 3617 5584 3645
rect 5584 3617 5598 3645
rect 4742 3614 4776 3617
rect 4844 3611 4878 3617
rect 4916 3611 4950 3617
rect 4988 3611 5022 3617
rect 5060 3611 5094 3617
rect 5132 3611 5166 3617
rect 5204 3611 5238 3617
rect 5276 3611 5310 3617
rect 5348 3611 5382 3617
rect 5420 3611 5454 3617
rect 5492 3611 5526 3617
rect 5564 3611 5598 3617
rect 5655 3611 5689 3645
rect 5729 3617 5760 3645
rect 5760 3617 5763 3645
rect 5803 3617 5830 3645
rect 5830 3617 5837 3645
rect 5877 3617 5900 3645
rect 5900 3617 5911 3645
rect 5951 3617 5970 3645
rect 5970 3617 5985 3645
rect 6025 3617 6040 3645
rect 6040 3617 6059 3645
rect 6099 3617 6110 3645
rect 6110 3617 6133 3645
rect 6173 3617 6180 3645
rect 6180 3617 6207 3645
rect 6247 3617 6250 3645
rect 6250 3617 6281 3645
rect 6416 3617 6424 3645
rect 6424 3617 6450 3645
rect 6535 3617 6564 3645
rect 6564 3617 6569 3645
rect 6992 3617 7003 3642
rect 7003 3617 7026 3642
rect 7064 3617 7074 3642
rect 7074 3617 7098 3642
rect 7136 3617 7145 3642
rect 7145 3617 7170 3642
rect 7208 3617 7216 3642
rect 7216 3617 7242 3642
rect 7280 3617 7287 3642
rect 7287 3617 7314 3642
rect 7353 3617 7358 3642
rect 7358 3617 7387 3642
rect 7426 3617 7429 3642
rect 7429 3617 7460 3642
rect 7499 3617 7500 3642
rect 7500 3617 7533 3642
rect 7838 3640 7872 3650
rect 5729 3611 5763 3617
rect 5803 3611 5837 3617
rect 5877 3611 5911 3617
rect 5951 3611 5985 3617
rect 6025 3611 6059 3617
rect 6099 3611 6133 3617
rect 6173 3611 6207 3617
rect 6247 3611 6281 3617
rect 6416 3611 6450 3617
rect 6535 3611 6569 3617
rect 6992 3608 7026 3617
rect 7064 3608 7098 3617
rect 7136 3608 7170 3617
rect 7208 3608 7242 3617
rect 7280 3608 7314 3617
rect 7353 3608 7387 3617
rect 7426 3608 7460 3617
rect 7499 3608 7533 3617
rect 7838 3616 7872 3640
rect 467 3538 501 3572
rect 467 3464 501 3498
rect 7838 3572 7872 3575
rect 7838 3541 7872 3572
rect 660 3451 694 3476
rect 928 3473 962 3482
rect 1006 3473 1040 3482
rect 1084 3473 1118 3482
rect 1162 3473 1196 3482
rect 1239 3473 1273 3482
rect 1316 3473 1350 3482
rect 1393 3473 1427 3482
rect 1470 3473 1504 3482
rect 1547 3473 1581 3482
rect 1624 3473 1658 3482
rect 1785 3473 1819 3476
rect 1859 3473 1893 3476
rect 1932 3473 1966 3476
rect 2005 3473 2039 3476
rect 2078 3473 2112 3476
rect 2151 3473 2185 3476
rect 2224 3473 2258 3476
rect 2297 3473 2331 3476
rect 2370 3473 2404 3476
rect 2443 3473 2477 3476
rect 2516 3473 2550 3476
rect 2589 3473 2623 3476
rect 2662 3473 2696 3476
rect 2735 3473 2769 3476
rect 2808 3473 2842 3476
rect 2881 3473 2915 3476
rect 2954 3473 2988 3476
rect 3027 3473 3061 3476
rect 3100 3473 3134 3476
rect 3173 3473 3207 3476
rect 3246 3473 3280 3476
rect 3319 3473 3353 3476
rect 3392 3473 3426 3476
rect 3465 3473 3499 3476
rect 3538 3473 3572 3476
rect 3611 3473 3645 3476
rect 3684 3473 3718 3476
rect 3861 3473 3895 3476
rect 3946 3473 3980 3476
rect 4031 3473 4065 3476
rect 4116 3473 4150 3476
rect 4201 3473 4235 3476
rect 4373 3473 4407 3476
rect 4458 3473 4492 3476
rect 4543 3473 4577 3476
rect 4628 3473 4662 3476
rect 4713 3473 4747 3476
rect 4885 3473 4919 3476
rect 4998 3473 5032 3476
rect 5112 3473 5146 3476
rect 5192 3473 5226 3476
rect 5272 3473 5306 3476
rect 5352 3473 5386 3476
rect 5431 3473 5465 3476
rect 5510 3473 5544 3476
rect 5624 3473 5658 3476
rect 5700 3473 5734 3476
rect 5776 3473 5810 3476
rect 5852 3473 5886 3476
rect 5928 3473 5962 3476
rect 6004 3473 6038 3476
rect 6080 3473 6114 3476
rect 6156 3473 6190 3476
rect 6232 3473 6266 3476
rect 6308 3473 6342 3476
rect 6384 3473 6418 3476
rect 6459 3473 6493 3476
rect 6534 3473 6568 3476
rect 6992 3473 7026 3482
rect 7064 3473 7098 3482
rect 7136 3473 7170 3482
rect 7208 3473 7242 3482
rect 7280 3473 7314 3482
rect 7353 3473 7387 3482
rect 7426 3473 7460 3482
rect 7499 3473 7533 3482
rect 467 3390 501 3424
rect 660 3442 679 3451
rect 679 3442 694 3451
rect 928 3448 932 3473
rect 932 3448 962 3473
rect 1006 3448 1040 3473
rect 1084 3448 1114 3473
rect 1114 3448 1118 3473
rect 1162 3448 1188 3473
rect 1188 3448 1196 3473
rect 1239 3448 1262 3473
rect 1262 3448 1273 3473
rect 1316 3448 1335 3473
rect 1335 3448 1350 3473
rect 1393 3448 1408 3473
rect 1408 3448 1427 3473
rect 1470 3448 1481 3473
rect 1481 3448 1504 3473
rect 1547 3448 1554 3473
rect 1554 3448 1581 3473
rect 1624 3448 1627 3473
rect 1627 3448 1658 3473
rect 1785 3442 1788 3473
rect 1788 3442 1819 3473
rect 1859 3442 1890 3473
rect 1890 3442 1893 3473
rect 1932 3442 1958 3473
rect 1958 3442 1966 3473
rect 2005 3442 2026 3473
rect 2026 3442 2039 3473
rect 2078 3442 2094 3473
rect 2094 3442 2112 3473
rect 2151 3442 2162 3473
rect 2162 3442 2185 3473
rect 2224 3442 2230 3473
rect 2230 3442 2258 3473
rect 2297 3442 2298 3473
rect 2298 3442 2331 3473
rect 2370 3442 2400 3473
rect 2400 3442 2404 3473
rect 2443 3442 2468 3473
rect 2468 3442 2477 3473
rect 2516 3442 2536 3473
rect 2536 3442 2550 3473
rect 2589 3442 2604 3473
rect 2604 3442 2623 3473
rect 2662 3442 2672 3473
rect 2672 3442 2696 3473
rect 2735 3442 2740 3473
rect 2740 3442 2769 3473
rect 2808 3442 2842 3473
rect 2881 3442 2910 3473
rect 2910 3442 2915 3473
rect 2954 3442 2978 3473
rect 2978 3442 2988 3473
rect 3027 3442 3046 3473
rect 3046 3442 3061 3473
rect 3100 3442 3114 3473
rect 3114 3442 3134 3473
rect 3173 3442 3182 3473
rect 3182 3442 3207 3473
rect 3246 3442 3250 3473
rect 3250 3442 3280 3473
rect 3319 3442 3352 3473
rect 3352 3442 3353 3473
rect 3392 3442 3420 3473
rect 3420 3442 3426 3473
rect 3465 3442 3488 3473
rect 3488 3442 3499 3473
rect 3538 3442 3556 3473
rect 3556 3442 3572 3473
rect 3611 3442 3624 3473
rect 3624 3442 3645 3473
rect 3684 3442 3692 3473
rect 3692 3442 3718 3473
rect 3861 3442 3862 3473
rect 3862 3442 3895 3473
rect 3946 3442 3964 3473
rect 3964 3442 3980 3473
rect 4031 3442 4032 3473
rect 4032 3442 4065 3473
rect 4116 3442 4134 3473
rect 4134 3442 4150 3473
rect 4201 3442 4202 3473
rect 4202 3442 4235 3473
rect 4373 3442 4407 3473
rect 4458 3442 4476 3473
rect 4476 3442 4492 3473
rect 4543 3442 4545 3473
rect 4545 3442 4577 3473
rect 4628 3442 4649 3473
rect 4649 3442 4662 3473
rect 4713 3442 4718 3473
rect 4718 3442 4747 3473
rect 4885 3442 4890 3473
rect 4890 3442 4919 3473
rect 4998 3442 5028 3473
rect 5028 3442 5032 3473
rect 5112 3442 5116 3473
rect 5116 3442 5146 3473
rect 5192 3442 5194 3473
rect 5194 3442 5226 3473
rect 5272 3442 5306 3473
rect 5352 3442 5384 3473
rect 5384 3442 5386 3473
rect 5431 3442 5462 3473
rect 5462 3442 5465 3473
rect 5510 3442 5540 3473
rect 5540 3442 5544 3473
rect 5624 3442 5628 3473
rect 5628 3442 5658 3473
rect 5700 3442 5731 3473
rect 5731 3442 5734 3473
rect 5776 3442 5800 3473
rect 5800 3442 5810 3473
rect 5852 3442 5869 3473
rect 5869 3442 5886 3473
rect 5928 3442 5938 3473
rect 5938 3442 5962 3473
rect 6004 3442 6007 3473
rect 6007 3442 6038 3473
rect 6080 3442 6111 3473
rect 6111 3442 6114 3473
rect 6156 3442 6180 3473
rect 6180 3442 6190 3473
rect 6232 3442 6250 3473
rect 6250 3442 6266 3473
rect 6308 3442 6320 3473
rect 6320 3442 6342 3473
rect 6384 3442 6390 3473
rect 6390 3442 6418 3473
rect 6459 3442 6460 3473
rect 6460 3442 6493 3473
rect 6534 3442 6564 3473
rect 6564 3442 6568 3473
rect 6992 3448 7003 3473
rect 7003 3448 7026 3473
rect 7064 3448 7074 3473
rect 7074 3448 7098 3473
rect 7136 3448 7145 3473
rect 7145 3448 7170 3473
rect 7208 3448 7216 3473
rect 7216 3448 7242 3473
rect 7280 3448 7287 3473
rect 7287 3448 7314 3473
rect 7353 3448 7358 3473
rect 7358 3448 7387 3473
rect 7426 3448 7429 3473
rect 7429 3448 7460 3473
rect 7499 3448 7500 3473
rect 7500 3448 7533 3473
rect 7838 3470 7872 3500
rect 7838 3466 7872 3470
rect 660 3380 694 3394
rect 7838 3402 7872 3425
rect 7838 3391 7872 3402
rect 467 3316 501 3350
rect 660 3360 679 3380
rect 679 3360 694 3380
rect 660 3309 694 3311
rect 467 3242 501 3276
rect 660 3277 679 3309
rect 679 3277 694 3309
rect 871 3349 905 3383
rect 871 3293 905 3311
rect 871 3277 905 3293
rect 1727 3349 1761 3383
rect 1727 3293 1761 3311
rect 1727 3277 1761 3293
rect 1983 3349 2017 3383
rect 1983 3293 2017 3311
rect 1983 3277 2017 3293
rect 2239 3349 2273 3383
rect 2239 3293 2273 3311
rect 2239 3277 2273 3293
rect 2495 3349 2529 3383
rect 2495 3293 2529 3311
rect 2495 3277 2529 3293
rect 2751 3349 2785 3383
rect 2751 3293 2785 3311
rect 2751 3277 2785 3293
rect 3007 3349 3041 3383
rect 3007 3293 3041 3311
rect 3007 3277 3041 3293
rect 3263 3349 3297 3383
rect 3263 3293 3297 3311
rect 3263 3277 3297 3293
rect 3519 3349 3553 3383
rect 3519 3293 3553 3311
rect 3519 3277 3553 3293
rect 3775 3349 3809 3383
rect 3775 3293 3809 3311
rect 3775 3277 3809 3293
rect 4031 3349 4065 3383
rect 4031 3293 4065 3311
rect 4031 3277 4065 3293
rect 4287 3349 4321 3383
rect 4287 3293 4321 3311
rect 4287 3277 4321 3293
rect 4543 3349 4577 3383
rect 4543 3293 4577 3311
rect 4543 3277 4577 3293
rect 4799 3349 4833 3383
rect 4799 3293 4833 3311
rect 4799 3277 4833 3293
rect 5055 3349 5089 3383
rect 5055 3293 5089 3311
rect 5055 3277 5089 3293
rect 5311 3349 5345 3383
rect 5311 3293 5345 3311
rect 5311 3277 5345 3293
rect 5567 3349 5601 3383
rect 5567 3293 5601 3311
rect 5567 3277 5601 3293
rect 5823 3349 5857 3383
rect 5823 3293 5857 3311
rect 5823 3277 5857 3293
rect 6079 3349 6113 3383
rect 6079 3293 6113 3311
rect 6079 3277 6113 3293
rect 6335 3349 6369 3383
rect 6335 3293 6369 3311
rect 6335 3277 6369 3293
rect 6591 3349 6625 3383
rect 6591 3293 6625 3311
rect 6591 3277 6625 3293
rect 6847 3349 6881 3383
rect 6847 3293 6881 3311
rect 6847 3277 6881 3293
rect 7703 3349 7737 3383
rect 7703 3293 7737 3311
rect 7703 3277 7737 3293
rect 7838 3334 7872 3350
rect 7838 3316 7872 3334
rect 467 3168 501 3202
rect 7838 3266 7872 3275
rect 7838 3241 7872 3266
rect 7838 3198 7872 3200
rect 7838 3166 7872 3198
rect 482 3094 516 3128
rect 1077 3094 1106 3111
rect 1106 3094 1111 3111
rect 1150 3094 1174 3111
rect 1174 3094 1184 3111
rect 1223 3094 1242 3111
rect 1242 3094 1257 3111
rect 1296 3094 1310 3111
rect 1310 3094 1330 3111
rect 1368 3094 1378 3111
rect 1378 3094 1402 3111
rect 1440 3094 1446 3111
rect 1446 3094 1474 3111
rect 1512 3094 1514 3111
rect 1514 3094 1546 3111
rect 1584 3094 1616 3111
rect 1616 3094 1618 3111
rect 1656 3094 1684 3111
rect 1684 3094 1690 3111
rect 1728 3094 1752 3111
rect 1752 3094 1762 3111
rect 1800 3094 1820 3111
rect 1820 3094 1834 3111
rect 1872 3094 1888 3111
rect 1888 3094 1906 3111
rect 1944 3094 1956 3111
rect 1956 3094 1978 3111
rect 2016 3094 2024 3111
rect 2024 3094 2050 3111
rect 2088 3094 2092 3111
rect 2092 3094 2122 3111
rect 1077 3077 1111 3094
rect 1150 3077 1184 3094
rect 1223 3077 1257 3094
rect 1296 3077 1330 3094
rect 1368 3077 1402 3094
rect 1440 3077 1474 3094
rect 1512 3077 1546 3094
rect 1584 3077 1618 3094
rect 1656 3077 1690 3094
rect 1728 3077 1762 3094
rect 1800 3077 1834 3094
rect 1872 3077 1906 3094
rect 1944 3077 1978 3094
rect 2016 3077 2050 3094
rect 2088 3077 2122 3094
rect 2160 3077 2194 3111
rect 2232 3094 2262 3111
rect 2262 3094 2266 3111
rect 2304 3094 2330 3111
rect 2330 3094 2338 3111
rect 2376 3094 2398 3111
rect 2398 3094 2410 3111
rect 2448 3094 2466 3111
rect 2466 3094 2482 3111
rect 2520 3094 2534 3111
rect 2534 3094 2554 3111
rect 2592 3094 2602 3111
rect 2602 3094 2626 3111
rect 2664 3094 2670 3111
rect 2670 3094 2698 3111
rect 2736 3094 2738 3111
rect 2738 3094 2770 3111
rect 2808 3094 2840 3111
rect 2840 3094 2842 3111
rect 2880 3094 2908 3111
rect 2908 3094 2914 3111
rect 2952 3094 2976 3111
rect 2976 3094 2986 3111
rect 3024 3094 3044 3111
rect 3044 3094 3058 3111
rect 3096 3094 3112 3111
rect 3112 3094 3130 3111
rect 3168 3094 3180 3111
rect 3180 3094 3202 3111
rect 3240 3094 3248 3111
rect 3248 3094 3274 3111
rect 3312 3094 3316 3111
rect 3316 3094 3346 3111
rect 2232 3077 2266 3094
rect 2304 3077 2338 3094
rect 2376 3077 2410 3094
rect 2448 3077 2482 3094
rect 2520 3077 2554 3094
rect 2592 3077 2626 3094
rect 2664 3077 2698 3094
rect 2736 3077 2770 3094
rect 2808 3077 2842 3094
rect 2880 3077 2914 3094
rect 2952 3077 2986 3094
rect 3024 3077 3058 3094
rect 3096 3077 3130 3094
rect 3168 3077 3202 3094
rect 3240 3077 3274 3094
rect 3312 3077 3346 3094
rect 3384 3077 3418 3111
rect 3456 3094 3486 3111
rect 3486 3094 3490 3111
rect 3528 3094 3554 3111
rect 3554 3094 3562 3111
rect 3600 3094 3622 3111
rect 3622 3094 3634 3111
rect 3672 3094 3690 3111
rect 3690 3094 3706 3111
rect 3744 3094 3758 3111
rect 3758 3094 3778 3111
rect 3888 3094 3894 3128
rect 3894 3094 3922 3128
rect 3962 3094 3996 3128
rect 4036 3094 4064 3128
rect 4064 3094 4070 3128
rect 4110 3094 4132 3128
rect 4132 3094 4144 3128
rect 4184 3094 4200 3128
rect 4200 3094 4218 3128
rect 4258 3094 4268 3128
rect 4268 3094 4292 3128
rect 4332 3094 4336 3128
rect 4336 3094 4366 3128
rect 4406 3094 4438 3128
rect 4438 3094 4440 3128
rect 4480 3094 4506 3128
rect 4506 3094 4514 3128
rect 4553 3094 4574 3128
rect 4574 3094 4587 3128
rect 4626 3094 4642 3128
rect 4642 3094 4660 3128
rect 4699 3094 4710 3128
rect 4710 3094 4733 3128
rect 4772 3094 4778 3128
rect 4778 3094 4806 3128
rect 4845 3094 4846 3128
rect 4846 3094 4879 3128
rect 4918 3094 4948 3128
rect 4948 3094 4952 3128
rect 4991 3094 5016 3128
rect 5016 3094 5025 3128
rect 5064 3094 5084 3128
rect 5084 3094 5098 3128
rect 5137 3094 5152 3128
rect 5152 3094 5171 3128
rect 5210 3094 5220 3128
rect 5220 3094 5244 3128
rect 5283 3094 5288 3128
rect 5288 3094 5317 3128
rect 5356 3094 5390 3128
rect 5429 3094 5458 3128
rect 5458 3094 5463 3128
rect 5502 3094 5526 3128
rect 5526 3094 5536 3128
rect 5575 3094 5594 3128
rect 5594 3094 5609 3128
rect 5648 3094 5662 3128
rect 5662 3094 5682 3128
rect 5721 3094 5730 3128
rect 5730 3094 5755 3128
rect 5794 3094 5798 3128
rect 5798 3094 5828 3128
rect 5867 3094 5900 3128
rect 5900 3094 5901 3128
rect 5940 3094 5968 3128
rect 5968 3094 5974 3128
rect 6013 3094 6036 3128
rect 6036 3094 6047 3128
rect 6086 3094 6104 3128
rect 6104 3094 6120 3128
rect 6159 3094 6172 3128
rect 6172 3094 6193 3128
rect 6232 3094 6240 3128
rect 6240 3094 6266 3128
rect 6305 3094 6308 3128
rect 6308 3094 6339 3128
rect 6378 3094 6410 3128
rect 6410 3094 6412 3128
rect 6451 3094 6478 3128
rect 6478 3094 6485 3128
rect 6524 3094 6546 3128
rect 6546 3094 6558 3128
rect 6597 3094 6614 3128
rect 6614 3094 6631 3128
rect 6670 3094 6682 3128
rect 6682 3094 6704 3128
rect 6743 3094 6750 3128
rect 6750 3094 6777 3128
rect 6816 3094 6818 3128
rect 6818 3094 6850 3128
rect 6889 3094 6920 3128
rect 6920 3094 6923 3128
rect 6962 3094 6988 3128
rect 6988 3094 6996 3128
rect 7035 3094 7056 3128
rect 7056 3094 7069 3128
rect 7108 3094 7124 3128
rect 7124 3094 7142 3128
rect 7181 3094 7192 3128
rect 7192 3094 7215 3128
rect 7254 3094 7260 3128
rect 7260 3094 7288 3128
rect 7327 3094 7328 3128
rect 7328 3094 7361 3128
rect 7400 3094 7430 3128
rect 7430 3094 7434 3128
rect 7473 3094 7498 3128
rect 7498 3094 7507 3128
rect 7546 3094 7566 3128
rect 7566 3094 7580 3128
rect 7619 3094 7634 3128
rect 7634 3094 7653 3128
rect 7692 3094 7702 3128
rect 7702 3094 7726 3128
rect 7765 3094 7770 3128
rect 7770 3094 7799 3128
rect 8554 4883 8584 4912
rect 8584 4883 8588 4912
rect 8627 4883 8654 4912
rect 8654 4883 8661 4912
rect 8700 4883 8724 4912
rect 8724 4883 8734 4912
rect 8773 4883 8794 4912
rect 8794 4883 8807 4912
rect 8846 4883 8864 4912
rect 8864 4883 8880 4912
rect 8919 4883 8934 4912
rect 8934 4883 8953 4912
rect 8992 4883 9004 4912
rect 9004 4883 9026 4912
rect 9065 4883 9074 4912
rect 9074 4883 9099 4912
rect 9138 4883 9144 4912
rect 9144 4883 9172 4912
rect 9211 4883 9214 4912
rect 9214 4883 9245 4912
rect 8554 4878 8588 4883
rect 8627 4878 8661 4883
rect 8700 4878 8734 4883
rect 8773 4878 8807 4883
rect 8846 4878 8880 4883
rect 8919 4878 8953 4883
rect 8992 4878 9026 4883
rect 9065 4878 9099 4883
rect 9138 4878 9172 4883
rect 9211 4878 9245 4883
rect 9284 4878 9318 4912
rect 9357 4883 9390 4912
rect 9390 4883 9391 4912
rect 9430 4883 9460 4912
rect 9460 4883 9464 4912
rect 9503 4883 9530 4912
rect 9530 4883 9537 4912
rect 9576 4883 9599 4912
rect 9599 4883 9610 4912
rect 9649 4883 9668 4912
rect 9668 4883 9683 4912
rect 9722 4883 9737 4912
rect 9737 4883 9756 4912
rect 9795 4883 9806 4912
rect 9806 4883 9829 4912
rect 9868 4883 9875 4912
rect 9875 4883 9902 4912
rect 9941 4883 9944 4912
rect 9944 4883 9975 4912
rect 10014 4883 10047 4912
rect 10047 4883 10048 4912
rect 10087 4883 10116 4912
rect 10116 4883 10121 4912
rect 10160 4883 10185 4912
rect 10185 4883 10194 4912
rect 10233 4883 10254 4912
rect 10254 4883 10267 4912
rect 10306 4883 10323 4912
rect 10323 4883 10340 4912
rect 10379 4883 10392 4912
rect 10392 4883 10413 4912
rect 10452 4883 10461 4912
rect 10461 4883 10486 4912
rect 10525 4883 10530 4912
rect 10530 4883 10559 4912
rect 10598 4883 10599 4912
rect 10599 4883 10632 4912
rect 10671 4883 10703 4912
rect 10703 4883 10705 4912
rect 10744 4883 10772 4912
rect 10772 4883 10778 4912
rect 10817 4883 10841 4912
rect 10841 4883 10851 4912
rect 10890 4883 10910 4912
rect 10910 4883 10924 4912
rect 10963 4883 10979 4912
rect 10979 4883 10997 4912
rect 11036 4883 11048 4912
rect 11048 4883 11070 4912
rect 11109 4883 11117 4912
rect 11117 4883 11143 4912
rect 11182 4883 11186 4912
rect 11186 4883 11216 4912
rect 9357 4878 9391 4883
rect 9430 4878 9464 4883
rect 9503 4878 9537 4883
rect 9576 4878 9610 4883
rect 9649 4878 9683 4883
rect 9722 4878 9756 4883
rect 9795 4878 9829 4883
rect 9868 4878 9902 4883
rect 9941 4878 9975 4883
rect 10014 4878 10048 4883
rect 10087 4878 10121 4883
rect 10160 4878 10194 4883
rect 10233 4878 10267 4883
rect 10306 4878 10340 4883
rect 10379 4878 10413 4883
rect 10452 4878 10486 4883
rect 10525 4878 10559 4883
rect 10598 4878 10632 4883
rect 10671 4878 10705 4883
rect 10744 4878 10778 4883
rect 10817 4878 10851 4883
rect 10890 4878 10924 4883
rect 10963 4878 10997 4883
rect 11036 4878 11070 4883
rect 11109 4878 11143 4883
rect 11182 4878 11216 4883
rect 11255 4878 11289 4912
rect 11328 4883 11356 4912
rect 11356 4883 11362 4912
rect 11401 4883 11425 4912
rect 11425 4883 11435 4912
rect 11474 4883 11494 4912
rect 11494 4883 11508 4912
rect 11547 4883 11563 4912
rect 11563 4883 11581 4912
rect 11620 4883 11632 4912
rect 11632 4883 11654 4912
rect 11693 4883 11701 4912
rect 11701 4883 11727 4912
rect 11765 4883 11770 4912
rect 11770 4883 11799 4912
rect 11837 4883 11839 4912
rect 11839 4883 11871 4912
rect 11328 4878 11362 4883
rect 11401 4878 11435 4883
rect 11474 4878 11508 4883
rect 11547 4878 11581 4883
rect 11620 4878 11654 4883
rect 11693 4878 11727 4883
rect 11765 4878 11799 4883
rect 11837 4878 11871 4883
rect 11909 4878 11943 4912
rect 11981 4883 12012 4912
rect 12012 4883 12015 4912
rect 12053 4883 12081 4912
rect 12081 4883 12087 4912
rect 12125 4883 12150 4912
rect 12150 4883 12159 4912
rect 12197 4883 12219 4912
rect 12219 4883 12231 4912
rect 12269 4883 12288 4912
rect 12288 4883 12303 4912
rect 12341 4883 12357 4912
rect 12357 4883 12375 4912
rect 12413 4883 12426 4912
rect 12426 4883 12447 4912
rect 12485 4883 12495 4912
rect 12495 4883 12519 4912
rect 12557 4883 12563 4912
rect 12563 4883 12591 4912
rect 12629 4883 12631 4912
rect 12631 4883 12663 4912
rect 12701 4883 12733 4912
rect 12733 4883 12735 4912
rect 12773 4883 12801 4912
rect 12801 4883 12807 4912
rect 12845 4883 12869 4912
rect 12869 4883 12879 4912
rect 12917 4883 12937 4912
rect 12937 4883 12951 4912
rect 12989 4883 13005 4912
rect 13005 4883 13023 4912
rect 13061 4883 13073 4912
rect 13073 4883 13095 4912
rect 13133 4883 13141 4912
rect 13141 4883 13167 4912
rect 13205 4883 13209 4912
rect 13209 4883 13239 4912
rect 11981 4878 12015 4883
rect 12053 4878 12087 4883
rect 12125 4878 12159 4883
rect 12197 4878 12231 4883
rect 12269 4878 12303 4883
rect 12341 4878 12375 4883
rect 12413 4878 12447 4883
rect 12485 4878 12519 4883
rect 12557 4878 12591 4883
rect 12629 4878 12663 4883
rect 12701 4878 12735 4883
rect 12773 4878 12807 4883
rect 12845 4878 12879 4883
rect 12917 4878 12951 4883
rect 12989 4878 13023 4883
rect 13061 4878 13095 4883
rect 13133 4878 13167 4883
rect 13205 4878 13239 4883
rect 13277 4878 13311 4912
rect 13349 4883 13379 4912
rect 13379 4883 13383 4912
rect 13421 4883 13447 4912
rect 13447 4883 13455 4912
rect 13493 4883 13515 4912
rect 13515 4883 13527 4912
rect 13565 4883 13583 4912
rect 13583 4883 13599 4912
rect 13637 4883 13651 4912
rect 13651 4883 13671 4912
rect 13709 4883 13719 4912
rect 13719 4883 13743 4912
rect 13781 4883 13787 4912
rect 13787 4883 13815 4912
rect 13853 4883 13855 4912
rect 13855 4883 13887 4912
rect 13925 4883 13957 4912
rect 13957 4883 13959 4912
rect 13997 4883 14025 4912
rect 14025 4883 14031 4912
rect 14069 4883 14093 4912
rect 14093 4883 14103 4912
rect 14141 4883 14161 4912
rect 14161 4883 14175 4912
rect 14213 4883 14229 4912
rect 14229 4883 14247 4912
rect 14285 4883 14297 4912
rect 14297 4883 14319 4912
rect 14357 4883 14365 4912
rect 14365 4883 14391 4912
rect 14429 4883 14433 4912
rect 14433 4883 14463 4912
rect 13349 4878 13383 4883
rect 13421 4878 13455 4883
rect 13493 4878 13527 4883
rect 13565 4878 13599 4883
rect 13637 4878 13671 4883
rect 13709 4878 13743 4883
rect 13781 4878 13815 4883
rect 13853 4878 13887 4883
rect 13925 4878 13959 4883
rect 13997 4878 14031 4883
rect 14069 4878 14103 4883
rect 14141 4878 14175 4883
rect 14213 4878 14247 4883
rect 14285 4878 14319 4883
rect 14357 4878 14391 4883
rect 14429 4878 14463 4883
rect 14501 4878 14535 4912
rect 14573 4883 14603 4912
rect 14603 4883 14607 4912
rect 14645 4883 14671 4912
rect 14671 4883 14679 4912
rect 14717 4883 14739 4912
rect 14739 4883 14751 4912
rect 14789 4883 14807 4912
rect 14807 4883 14823 4912
rect 14861 4883 14875 4912
rect 14875 4883 14895 4912
rect 14933 4883 14943 4912
rect 14943 4883 14967 4912
rect 15005 4883 15011 4912
rect 15011 4883 15039 4912
rect 15077 4883 15079 4912
rect 15079 4883 15111 4912
rect 15149 4883 15181 4912
rect 15181 4883 15183 4912
rect 15221 4883 15249 4912
rect 15249 4883 15255 4912
rect 15293 4883 15317 4912
rect 15317 4883 15327 4912
rect 15365 4883 15385 4912
rect 15385 4883 15399 4912
rect 15437 4883 15453 4912
rect 15453 4883 15471 4912
rect 15509 4883 15521 4912
rect 15521 4883 15543 4912
rect 15581 4883 15589 4912
rect 15589 4883 15615 4912
rect 15653 4883 15657 4912
rect 15657 4883 15687 4912
rect 14573 4878 14607 4883
rect 14645 4878 14679 4883
rect 14717 4878 14751 4883
rect 14789 4878 14823 4883
rect 14861 4878 14895 4883
rect 14933 4878 14967 4883
rect 15005 4878 15039 4883
rect 15077 4878 15111 4883
rect 15149 4878 15183 4883
rect 15221 4878 15255 4883
rect 15293 4878 15327 4883
rect 15365 4878 15399 4883
rect 15437 4878 15471 4883
rect 15509 4878 15543 4883
rect 15581 4878 15615 4883
rect 15653 4878 15687 4883
rect 15725 4878 15759 4912
rect 15797 4883 15827 4912
rect 15827 4883 15831 4912
rect 15869 4883 15895 4912
rect 15895 4883 15903 4912
rect 15941 4883 15963 4912
rect 15963 4883 15975 4912
rect 16013 4883 16031 4912
rect 16031 4883 16047 4912
rect 16085 4883 16099 4912
rect 16099 4883 16119 4912
rect 16157 4883 16167 4912
rect 16167 4883 16191 4912
rect 16229 4883 16235 4912
rect 16235 4883 16263 4912
rect 16301 4883 16303 4912
rect 16303 4883 16335 4912
rect 16373 4883 16405 4912
rect 16405 4883 16407 4912
rect 16445 4883 16473 4912
rect 16473 4883 16479 4912
rect 16517 4883 16541 4912
rect 16541 4883 16551 4912
rect 16589 4883 16609 4912
rect 16609 4883 16623 4912
rect 16661 4883 16677 4912
rect 16677 4883 16695 4912
rect 16733 4883 16745 4912
rect 16745 4883 16767 4912
rect 16805 4883 16813 4912
rect 16813 4883 16839 4912
rect 16877 4883 16881 4912
rect 16881 4883 16911 4912
rect 15797 4878 15831 4883
rect 15869 4878 15903 4883
rect 15941 4878 15975 4883
rect 16013 4878 16047 4883
rect 16085 4878 16119 4883
rect 16157 4878 16191 4883
rect 16229 4878 16263 4883
rect 16301 4878 16335 4883
rect 16373 4878 16407 4883
rect 16445 4878 16479 4883
rect 16517 4878 16551 4883
rect 16589 4878 16623 4883
rect 16661 4878 16695 4883
rect 16733 4878 16767 4883
rect 16805 4878 16839 4883
rect 16877 4878 16911 4883
rect 16949 4878 16983 4912
rect 17021 4883 17051 4912
rect 17051 4883 17055 4912
rect 17093 4883 17119 4912
rect 17119 4883 17127 4912
rect 17165 4883 17187 4912
rect 17187 4883 17199 4912
rect 17237 4883 17255 4912
rect 17255 4883 17271 4912
rect 17309 4883 17323 4912
rect 17323 4883 17343 4912
rect 17381 4883 17391 4912
rect 17391 4883 17415 4912
rect 17453 4883 17459 4912
rect 17459 4883 17487 4912
rect 17525 4883 17527 4912
rect 17527 4883 17559 4912
rect 17597 4883 17629 4912
rect 17629 4883 17631 4912
rect 17669 4883 17697 4912
rect 17697 4883 17703 4912
rect 17741 4883 17765 4912
rect 17765 4883 17775 4912
rect 17813 4883 17833 4912
rect 17833 4883 17847 4912
rect 17885 4883 17901 4912
rect 17901 4883 17919 4912
rect 17957 4883 17969 4912
rect 17969 4883 17991 4912
rect 18029 4883 18037 4912
rect 18037 4883 18063 4912
rect 18101 4883 18105 4912
rect 18105 4883 18135 4912
rect 17021 4878 17055 4883
rect 17093 4878 17127 4883
rect 17165 4878 17199 4883
rect 17237 4878 17271 4883
rect 17309 4878 17343 4883
rect 17381 4878 17415 4883
rect 17453 4878 17487 4883
rect 17525 4878 17559 4883
rect 17597 4878 17631 4883
rect 17669 4878 17703 4883
rect 17741 4878 17775 4883
rect 17813 4878 17847 4883
rect 17885 4878 17919 4883
rect 17957 4878 17991 4883
rect 18029 4878 18063 4883
rect 18101 4878 18135 4883
rect 18173 4878 18207 4912
rect 18245 4883 18275 4912
rect 18275 4883 18279 4912
rect 18317 4883 18343 4912
rect 18343 4883 18351 4912
rect 18389 4883 18411 4912
rect 18411 4883 18423 4912
rect 18461 4883 18479 4912
rect 18479 4883 18495 4912
rect 18533 4883 18547 4912
rect 18547 4883 18567 4912
rect 18605 4883 18615 4912
rect 18615 4883 18639 4912
rect 18677 4883 18683 4912
rect 18683 4883 18711 4912
rect 18749 4883 18751 4912
rect 18751 4883 18783 4912
rect 18821 4883 18853 4912
rect 18853 4883 18855 4912
rect 18893 4883 18921 4912
rect 18921 4883 18927 4912
rect 18965 4883 18989 4912
rect 18989 4883 18999 4912
rect 19037 4883 19057 4912
rect 19057 4883 19071 4912
rect 19109 4883 19125 4912
rect 19125 4883 19143 4912
rect 19181 4883 19193 4912
rect 19193 4883 19215 4912
rect 19253 4883 19261 4912
rect 19261 4883 19287 4912
rect 19325 4883 19329 4912
rect 19329 4883 19359 4912
rect 18245 4878 18279 4883
rect 18317 4878 18351 4883
rect 18389 4878 18423 4883
rect 18461 4878 18495 4883
rect 18533 4878 18567 4883
rect 18605 4878 18639 4883
rect 18677 4878 18711 4883
rect 18749 4878 18783 4883
rect 18821 4878 18855 4883
rect 18893 4878 18927 4883
rect 18965 4878 18999 4883
rect 19037 4878 19071 4883
rect 19109 4878 19143 4883
rect 19181 4878 19215 4883
rect 19253 4878 19287 4883
rect 19325 4878 19359 4883
rect 19397 4878 19431 4912
rect 19469 4883 19499 4912
rect 19499 4883 19503 4912
rect 19541 4883 19567 4912
rect 19567 4883 19575 4912
rect 19613 4883 19635 4912
rect 19635 4883 19647 4912
rect 19685 4883 19703 4912
rect 19703 4883 19719 4912
rect 19757 4883 19771 4912
rect 19771 4883 19791 4912
rect 19829 4883 19839 4912
rect 19839 4883 19863 4912
rect 19901 4883 19907 4912
rect 19907 4883 19935 4912
rect 19469 4878 19503 4883
rect 19541 4878 19575 4883
rect 19613 4878 19647 4883
rect 19685 4878 19719 4883
rect 19757 4878 19791 4883
rect 19829 4878 19863 4883
rect 19901 4878 19935 4883
rect 8482 4814 8516 4838
rect 8482 4804 8516 4814
rect 8482 4745 8516 4764
rect 8482 4730 8516 4745
rect 8482 4676 8516 4690
rect 8482 4656 8516 4676
rect 8482 4607 8516 4616
rect 8482 4582 8516 4607
rect 8482 4538 8516 4542
rect 8482 4508 8516 4538
rect 8482 4434 8516 4468
rect 8482 4365 8516 4394
rect 8482 4360 8516 4365
rect 8482 4296 8516 4320
rect 8482 4286 8516 4296
rect 8482 4226 8516 4246
rect 8482 4212 8516 4226
rect 8482 4156 8516 4172
rect 8482 4138 8516 4156
rect 8482 4086 8516 4098
rect 8482 4064 8516 4086
rect 8482 4016 8516 4024
rect 8482 3990 8516 4016
rect 8482 3946 8516 3950
rect 8482 3916 8516 3946
rect 8482 3842 8516 3876
rect 8714 4792 8748 4808
rect 8714 4774 8748 4792
rect 8714 4724 8748 4736
rect 8714 4702 8748 4724
rect 8714 4656 8748 4664
rect 8714 4630 8748 4656
rect 8714 4588 8748 4592
rect 8714 4558 8748 4588
rect 8714 4486 8748 4520
rect 8714 4418 8748 4448
rect 8714 4414 8748 4418
rect 8714 4350 8748 4376
rect 8714 4342 8748 4350
rect 8714 4282 8748 4304
rect 8714 4270 8748 4282
rect 8714 4214 8748 4232
rect 8714 4198 8748 4214
rect 8714 4146 8748 4160
rect 8714 4126 8748 4146
rect 8714 4078 8748 4088
rect 8714 4054 8748 4078
rect 8714 4010 8748 4016
rect 8714 3982 8748 4010
rect 8714 3942 8748 3944
rect 8714 3910 8748 3942
rect 8714 3838 8748 3872
rect 8870 4792 8904 4808
rect 8870 4774 8904 4792
rect 8870 4724 8904 4736
rect 8870 4702 8904 4724
rect 8870 4656 8904 4664
rect 8870 4630 8904 4656
rect 8870 4588 8904 4592
rect 8870 4558 8904 4588
rect 8870 4486 8904 4520
rect 8870 4418 8904 4448
rect 8870 4414 8904 4418
rect 8870 4350 8904 4376
rect 8870 4342 8904 4350
rect 8870 4282 8904 4304
rect 8870 4270 8904 4282
rect 8870 4214 8904 4232
rect 8870 4198 8904 4214
rect 8870 4146 8904 4160
rect 8870 4126 8904 4146
rect 8870 4078 8904 4088
rect 8870 4054 8904 4078
rect 8870 4010 8904 4016
rect 8870 3982 8904 4010
rect 8870 3942 8904 3944
rect 8870 3910 8904 3942
rect 8870 3838 8904 3872
rect 9026 4792 9060 4808
rect 9026 4774 9060 4792
rect 9026 4724 9060 4736
rect 9026 4702 9060 4724
rect 9026 4656 9060 4664
rect 9026 4630 9060 4656
rect 9026 4588 9060 4592
rect 9026 4558 9060 4588
rect 9026 4486 9060 4520
rect 9026 4418 9060 4448
rect 9026 4414 9060 4418
rect 9026 4350 9060 4376
rect 9026 4342 9060 4350
rect 9026 4282 9060 4304
rect 9026 4270 9060 4282
rect 9026 4214 9060 4232
rect 9026 4198 9060 4214
rect 9026 4146 9060 4160
rect 9026 4126 9060 4146
rect 9026 4078 9060 4088
rect 9026 4054 9060 4078
rect 9026 4010 9060 4016
rect 9026 3982 9060 4010
rect 9026 3942 9060 3944
rect 9026 3910 9060 3942
rect 9026 3838 9060 3872
rect 9182 4792 9216 4808
rect 9182 4774 9216 4792
rect 9182 4724 9216 4736
rect 9182 4702 9216 4724
rect 9182 4656 9216 4664
rect 9182 4630 9216 4656
rect 9182 4588 9216 4592
rect 9182 4558 9216 4588
rect 9182 4486 9216 4520
rect 9182 4418 9216 4448
rect 9182 4414 9216 4418
rect 9182 4350 9216 4376
rect 9182 4342 9216 4350
rect 9182 4282 9216 4304
rect 9182 4270 9216 4282
rect 9182 4214 9216 4232
rect 9182 4198 9216 4214
rect 9182 4146 9216 4160
rect 9182 4126 9216 4146
rect 9182 4078 9216 4088
rect 9182 4054 9216 4078
rect 9182 4010 9216 4016
rect 9182 3982 9216 4010
rect 9182 3942 9216 3944
rect 9182 3910 9216 3942
rect 9182 3838 9216 3872
rect 9338 4792 9372 4808
rect 9338 4774 9372 4792
rect 9338 4724 9372 4736
rect 9338 4702 9372 4724
rect 9338 4656 9372 4664
rect 9338 4630 9372 4656
rect 9338 4588 9372 4592
rect 9338 4558 9372 4588
rect 9338 4486 9372 4520
rect 9338 4418 9372 4448
rect 9338 4414 9372 4418
rect 9338 4350 9372 4376
rect 9338 4342 9372 4350
rect 9338 4282 9372 4304
rect 9338 4270 9372 4282
rect 9338 4214 9372 4232
rect 9338 4198 9372 4214
rect 9338 4146 9372 4160
rect 9338 4126 9372 4146
rect 9338 4078 9372 4088
rect 9338 4054 9372 4078
rect 9338 4010 9372 4016
rect 9338 3982 9372 4010
rect 9338 3942 9372 3944
rect 9338 3910 9372 3942
rect 9338 3838 9372 3872
rect 9462 4792 9496 4808
rect 9462 4774 9496 4792
rect 9462 4724 9496 4736
rect 9462 4702 9496 4724
rect 9462 4656 9496 4664
rect 9462 4630 9496 4656
rect 9462 4588 9496 4592
rect 9462 4558 9496 4588
rect 9462 4486 9496 4520
rect 9462 4418 9496 4448
rect 9462 4414 9496 4418
rect 9462 4350 9496 4376
rect 9462 4342 9496 4350
rect 9462 4282 9496 4304
rect 9462 4270 9496 4282
rect 9462 4214 9496 4232
rect 9462 4198 9496 4214
rect 9462 4146 9496 4160
rect 9462 4126 9496 4146
rect 9462 4078 9496 4088
rect 9462 4054 9496 4078
rect 9462 4010 9496 4016
rect 9462 3982 9496 4010
rect 9462 3942 9496 3944
rect 9462 3910 9496 3942
rect 9462 3838 9496 3872
rect 9618 4792 9652 4808
rect 9618 4774 9652 4792
rect 9618 4724 9652 4736
rect 9618 4702 9652 4724
rect 9618 4656 9652 4664
rect 9618 4630 9652 4656
rect 9618 4588 9652 4592
rect 9618 4558 9652 4588
rect 9618 4486 9652 4520
rect 9618 4418 9652 4448
rect 9618 4414 9652 4418
rect 9618 4350 9652 4376
rect 9618 4342 9652 4350
rect 9618 4282 9652 4304
rect 9618 4270 9652 4282
rect 9618 4214 9652 4232
rect 9618 4198 9652 4214
rect 9618 4146 9652 4160
rect 9618 4126 9652 4146
rect 9618 4078 9652 4088
rect 9618 4054 9652 4078
rect 9618 4010 9652 4016
rect 9618 3982 9652 4010
rect 9618 3942 9652 3944
rect 9618 3910 9652 3942
rect 9618 3838 9652 3872
rect 9742 4792 9776 4808
rect 9742 4774 9776 4792
rect 9742 4724 9776 4736
rect 9742 4702 9776 4724
rect 9742 4656 9776 4664
rect 9742 4630 9776 4656
rect 9742 4588 9776 4592
rect 9742 4558 9776 4588
rect 9742 4486 9776 4520
rect 9742 4418 9776 4448
rect 9742 4414 9776 4418
rect 9742 4350 9776 4376
rect 9742 4342 9776 4350
rect 9742 4282 9776 4304
rect 9742 4270 9776 4282
rect 9742 4214 9776 4232
rect 9742 4198 9776 4214
rect 9742 4146 9776 4160
rect 9742 4126 9776 4146
rect 9742 4078 9776 4088
rect 9742 4054 9776 4078
rect 9742 4010 9776 4016
rect 9742 3982 9776 4010
rect 9742 3942 9776 3944
rect 9742 3910 9776 3942
rect 9742 3838 9776 3872
rect 9898 4792 9932 4808
rect 9898 4774 9932 4792
rect 9898 4724 9932 4736
rect 9898 4702 9932 4724
rect 9898 4656 9932 4664
rect 9898 4630 9932 4656
rect 9898 4588 9932 4592
rect 9898 4558 9932 4588
rect 9898 4486 9932 4520
rect 9898 4418 9932 4448
rect 9898 4414 9932 4418
rect 9898 4350 9932 4376
rect 9898 4342 9932 4350
rect 9898 4282 9932 4304
rect 9898 4270 9932 4282
rect 9898 4214 9932 4232
rect 9898 4198 9932 4214
rect 9898 4146 9932 4160
rect 9898 4126 9932 4146
rect 9898 4078 9932 4088
rect 9898 4054 9932 4078
rect 9898 4010 9932 4016
rect 9898 3982 9932 4010
rect 9898 3942 9932 3944
rect 9898 3910 9932 3942
rect 9898 3838 9932 3872
rect 10054 4792 10088 4808
rect 10054 4774 10088 4792
rect 10054 4724 10088 4736
rect 10054 4702 10088 4724
rect 10054 4656 10088 4664
rect 10054 4630 10088 4656
rect 10054 4588 10088 4592
rect 10054 4558 10088 4588
rect 10054 4486 10088 4520
rect 10054 4418 10088 4448
rect 10054 4414 10088 4418
rect 10054 4350 10088 4376
rect 10054 4342 10088 4350
rect 10054 4282 10088 4304
rect 10054 4270 10088 4282
rect 10054 4214 10088 4232
rect 10054 4198 10088 4214
rect 10054 4146 10088 4160
rect 10054 4126 10088 4146
rect 10054 4078 10088 4088
rect 10054 4054 10088 4078
rect 10054 4010 10088 4016
rect 10054 3982 10088 4010
rect 10054 3942 10088 3944
rect 10054 3910 10088 3942
rect 10054 3838 10088 3872
rect 10331 4792 10365 4808
rect 10331 4774 10365 4792
rect 10331 4724 10365 4736
rect 10331 4702 10365 4724
rect 10331 4656 10365 4664
rect 10331 4630 10365 4656
rect 10331 4588 10365 4592
rect 10331 4558 10365 4588
rect 10331 4486 10365 4520
rect 10331 4418 10365 4448
rect 10331 4414 10365 4418
rect 10331 4350 10365 4376
rect 10331 4342 10365 4350
rect 10331 4282 10365 4304
rect 10331 4270 10365 4282
rect 10331 4214 10365 4232
rect 10331 4198 10365 4214
rect 10331 4146 10365 4160
rect 10331 4126 10365 4146
rect 10331 4078 10365 4088
rect 10331 4054 10365 4078
rect 10331 4010 10365 4016
rect 10331 3982 10365 4010
rect 10331 3942 10365 3944
rect 10331 3910 10365 3942
rect 10331 3838 10365 3872
rect 10487 4792 10521 4808
rect 10487 4774 10521 4792
rect 10487 4724 10521 4736
rect 10487 4702 10521 4724
rect 10487 4656 10521 4664
rect 10487 4630 10521 4656
rect 10487 4588 10521 4592
rect 10487 4558 10521 4588
rect 10487 4486 10521 4520
rect 10487 4418 10521 4448
rect 10487 4414 10521 4418
rect 10487 4350 10521 4376
rect 10487 4342 10521 4350
rect 10487 4282 10521 4304
rect 10487 4270 10521 4282
rect 10487 4214 10521 4232
rect 10487 4198 10521 4214
rect 10487 4146 10521 4160
rect 10487 4126 10521 4146
rect 10487 4078 10521 4088
rect 10487 4054 10521 4078
rect 10487 4010 10521 4016
rect 10487 3982 10521 4010
rect 10487 3942 10521 3944
rect 10487 3910 10521 3942
rect 10487 3838 10521 3872
rect 10643 4792 10677 4808
rect 10643 4774 10677 4792
rect 10643 4724 10677 4736
rect 10643 4702 10677 4724
rect 10643 4656 10677 4664
rect 10643 4630 10677 4656
rect 10643 4588 10677 4592
rect 10643 4558 10677 4588
rect 10643 4486 10677 4520
rect 10643 4418 10677 4448
rect 10643 4414 10677 4418
rect 10643 4350 10677 4376
rect 10643 4342 10677 4350
rect 10643 4282 10677 4304
rect 10643 4270 10677 4282
rect 10643 4214 10677 4232
rect 10643 4198 10677 4214
rect 10643 4146 10677 4160
rect 10643 4126 10677 4146
rect 10643 4078 10677 4088
rect 10643 4054 10677 4078
rect 10643 4010 10677 4016
rect 10643 3982 10677 4010
rect 10643 3942 10677 3944
rect 10643 3910 10677 3942
rect 10643 3838 10677 3872
rect 10799 4792 10833 4808
rect 10799 4774 10833 4792
rect 10799 4724 10833 4736
rect 10799 4702 10833 4724
rect 10799 4656 10833 4664
rect 10799 4630 10833 4656
rect 10799 4588 10833 4592
rect 10799 4558 10833 4588
rect 10799 4486 10833 4520
rect 10799 4418 10833 4448
rect 10799 4414 10833 4418
rect 10799 4350 10833 4376
rect 10799 4342 10833 4350
rect 10799 4282 10833 4304
rect 10799 4270 10833 4282
rect 10799 4214 10833 4232
rect 10799 4198 10833 4214
rect 10799 4146 10833 4160
rect 10799 4126 10833 4146
rect 10799 4078 10833 4088
rect 10799 4054 10833 4078
rect 10799 4010 10833 4016
rect 10799 3982 10833 4010
rect 10799 3942 10833 3944
rect 10799 3910 10833 3942
rect 10799 3838 10833 3872
rect 10955 4792 10989 4808
rect 10955 4774 10989 4792
rect 10955 4724 10989 4736
rect 10955 4702 10989 4724
rect 10955 4656 10989 4664
rect 10955 4630 10989 4656
rect 10955 4588 10989 4592
rect 10955 4558 10989 4588
rect 10955 4486 10989 4520
rect 10955 4418 10989 4448
rect 10955 4414 10989 4418
rect 10955 4350 10989 4376
rect 10955 4342 10989 4350
rect 10955 4282 10989 4304
rect 10955 4270 10989 4282
rect 10955 4214 10989 4232
rect 10955 4198 10989 4214
rect 10955 4146 10989 4160
rect 10955 4126 10989 4146
rect 10955 4078 10989 4088
rect 10955 4054 10989 4078
rect 10955 4010 10989 4016
rect 10955 3982 10989 4010
rect 10955 3942 10989 3944
rect 10955 3910 10989 3942
rect 10955 3838 10989 3872
rect 11111 4792 11145 4808
rect 11111 4774 11145 4792
rect 11111 4724 11145 4736
rect 11111 4702 11145 4724
rect 11111 4656 11145 4664
rect 11111 4630 11145 4656
rect 11111 4588 11145 4592
rect 11111 4558 11145 4588
rect 11111 4486 11145 4520
rect 11111 4418 11145 4448
rect 11111 4414 11145 4418
rect 11111 4350 11145 4376
rect 11111 4342 11145 4350
rect 11111 4282 11145 4304
rect 11111 4270 11145 4282
rect 11111 4214 11145 4232
rect 11111 4198 11145 4214
rect 11111 4146 11145 4160
rect 11111 4126 11145 4146
rect 11111 4078 11145 4088
rect 11111 4054 11145 4078
rect 11111 4010 11145 4016
rect 11111 3982 11145 4010
rect 11111 3942 11145 3944
rect 11111 3910 11145 3942
rect 11111 3838 11145 3872
rect 11298 4806 11332 4840
rect 11298 4732 11332 4766
rect 11298 4658 11332 4692
rect 19973 4835 20007 4840
rect 19973 4806 19975 4835
rect 19975 4806 20007 4835
rect 19973 4733 20007 4767
rect 19973 4674 20007 4694
rect 19973 4660 19975 4674
rect 19975 4660 20007 4674
rect 11298 4584 11332 4618
rect 13493 4599 13527 4633
rect 13584 4599 13618 4633
rect 17403 4626 17437 4660
rect 11298 4510 11332 4544
rect 16721 4525 16755 4559
rect 16793 4525 16827 4559
rect 17403 4554 17437 4588
rect 17996 4626 18030 4660
rect 17684 4529 17718 4563
rect 17996 4554 18030 4588
rect 19973 4606 20007 4621
rect 19973 4587 19975 4606
rect 19975 4587 20007 4606
rect 11298 4436 11332 4470
rect 17684 4457 17718 4491
rect 19365 4530 19399 4564
rect 19365 4458 19399 4492
rect 19627 4530 19661 4564
rect 19627 4458 19661 4492
rect 11298 4362 11332 4396
rect 14725 4377 14759 4411
rect 14797 4377 14831 4411
rect 18469 4377 18503 4411
rect 18541 4377 18575 4411
rect 11298 4288 11332 4322
rect 11298 4214 11332 4248
rect 11298 4140 11332 4174
rect 11801 4277 11835 4311
rect 13933 4303 13967 4337
rect 14005 4303 14039 4337
rect 11801 4205 11835 4239
rect 13250 4220 13284 4254
rect 13322 4220 13356 4254
rect 11298 4066 11332 4100
rect 11580 4126 11614 4160
rect 12400 4123 12434 4157
rect 12472 4123 12506 4157
rect 15110 4229 15144 4263
rect 15182 4229 15216 4263
rect 16468 4231 16502 4265
rect 16540 4231 16574 4265
rect 17672 4231 17706 4265
rect 17744 4231 17778 4265
rect 15529 4155 15563 4189
rect 15601 4155 15635 4189
rect 19450 4371 19484 4405
rect 19043 4303 19077 4337
rect 19115 4303 19149 4337
rect 19450 4299 19484 4333
rect 11580 4054 11614 4088
rect 11298 3992 11332 4026
rect 13089 4080 13123 4114
rect 13161 4080 13195 4114
rect 12448 4024 12482 4058
rect 12520 4024 12554 4058
rect 11298 3918 11332 3952
rect 12739 4022 12773 4056
rect 14089 4080 14123 4114
rect 14161 4080 14195 4114
rect 14890 4080 14924 4114
rect 14962 4080 14996 4114
rect 15721 4080 15755 4114
rect 15794 4080 15828 4114
rect 15866 4080 15900 4114
rect 15938 4080 15972 4114
rect 16317 4087 16351 4121
rect 16389 4087 16423 4121
rect 16843 4081 16877 4115
rect 16943 4085 16977 4119
rect 17015 4085 17049 4119
rect 16843 4009 16877 4043
rect 12739 3950 12773 3984
rect 17779 4039 17813 4073
rect 17855 4039 17889 4073
rect 17931 4039 17965 4073
rect 18605 4065 18639 4099
rect 18677 4065 18711 4099
rect 18429 3969 18463 4003
rect 18501 3969 18535 4003
rect 19268 4056 19302 4090
rect 19973 4538 20007 4548
rect 19973 4514 19975 4538
rect 19975 4514 20007 4538
rect 19973 4470 20007 4475
rect 19973 4441 19975 4470
rect 19975 4441 20007 4470
rect 19973 4368 19975 4402
rect 19975 4368 20007 4402
rect 19973 4300 19975 4329
rect 19975 4300 20007 4329
rect 19973 4295 20007 4300
rect 19973 4232 19975 4256
rect 19975 4232 20007 4256
rect 19973 4222 20007 4232
rect 19729 4149 19763 4183
rect 19729 4077 19763 4111
rect 19973 4164 19975 4183
rect 19975 4164 20007 4183
rect 19973 4149 20007 4164
rect 19973 4096 19975 4110
rect 19975 4096 20007 4110
rect 19973 4076 20007 4096
rect 19268 3984 19302 4018
rect 19973 4028 19975 4037
rect 19975 4028 20007 4037
rect 19973 4003 20007 4028
rect 19973 3960 19975 3964
rect 19975 3960 20007 3964
rect 19973 3930 20007 3960
rect 11298 3844 11332 3878
rect 14298 3864 14332 3898
rect 14370 3864 14404 3898
rect 17116 3892 17150 3926
rect 8482 3772 8516 3802
rect 8482 3768 8516 3772
rect 17116 3820 17150 3854
rect 19973 3858 20007 3891
rect 19973 3857 19975 3858
rect 19975 3857 20007 3858
rect 11298 3770 11332 3804
rect 9812 3756 9846 3757
rect 8482 3702 8516 3728
rect 8482 3694 8516 3702
rect 8482 3632 8516 3654
rect 8482 3620 8516 3632
rect 8657 3722 8691 3756
rect 9223 3717 9257 3751
rect 9295 3722 9311 3751
rect 9311 3722 9329 3751
rect 9295 3717 9329 3722
rect 8657 3650 8691 3684
rect 9812 3723 9837 3756
rect 9837 3723 9846 3756
rect 9895 3756 9929 3757
rect 9977 3756 10011 3757
rect 9895 3723 9898 3756
rect 9898 3723 9929 3756
rect 9977 3723 9993 3756
rect 9993 3723 10011 3756
rect 10399 3722 10426 3756
rect 10426 3722 10433 3756
rect 10473 3722 10500 3756
rect 10500 3722 10507 3756
rect 10546 3722 10573 3756
rect 10573 3722 10580 3756
rect 10619 3722 10646 3756
rect 10646 3722 10653 3756
rect 10692 3722 10719 3756
rect 10719 3722 10726 3756
rect 10765 3722 10792 3756
rect 10792 3722 10799 3756
rect 10838 3722 10865 3756
rect 10865 3722 10872 3756
rect 10911 3722 10938 3756
rect 10938 3722 10945 3756
rect 10984 3722 11011 3756
rect 11011 3722 11018 3756
rect 11057 3722 11084 3756
rect 11084 3722 11091 3756
rect 11298 3696 11332 3730
rect 9465 3623 9499 3657
rect 9537 3634 9541 3657
rect 9541 3634 9571 3657
rect 9537 3623 9571 3634
rect 8482 3562 8516 3580
rect 8482 3546 8516 3562
rect 8482 3492 8516 3506
rect 8482 3472 8516 3492
rect 10636 3609 10640 3643
rect 10640 3609 10670 3643
rect 10778 3609 10808 3643
rect 10808 3609 10812 3643
rect 11298 3622 11332 3656
rect 19973 3790 20007 3818
rect 19973 3784 19975 3790
rect 19975 3784 20007 3790
rect 19973 3722 20007 3745
rect 19973 3711 19975 3722
rect 19975 3711 20007 3722
rect 19973 3654 20007 3672
rect 19973 3638 19975 3654
rect 19975 3638 20007 3654
rect 8889 3475 8905 3509
rect 8905 3475 8923 3509
rect 8961 3475 8973 3509
rect 8973 3475 8995 3509
rect 9033 3475 9041 3509
rect 9041 3475 9067 3509
rect 9105 3475 9109 3509
rect 9109 3475 9139 3509
rect 9177 3475 9211 3509
rect 9249 3475 9279 3509
rect 9279 3475 9283 3509
rect 9321 3475 9347 3509
rect 9347 3475 9355 3509
rect 9393 3475 9415 3509
rect 9415 3475 9427 3509
rect 9465 3475 9483 3509
rect 9483 3475 9499 3509
rect 9537 3475 9551 3509
rect 9551 3475 9571 3509
rect 9609 3475 9619 3509
rect 9619 3475 9643 3509
rect 9681 3475 9687 3509
rect 9687 3475 9715 3509
rect 9753 3475 9755 3509
rect 9755 3475 9787 3509
rect 9825 3475 9859 3509
rect 10891 3532 10925 3566
rect 10963 3532 10997 3566
rect 11298 3548 11332 3582
rect 8482 3422 8516 3432
rect 8482 3398 8516 3422
rect 8482 3352 8516 3358
rect 8482 3324 8516 3352
rect 9941 3448 9975 3455
rect 9941 3421 9975 3448
rect 11298 3470 11332 3504
rect 9941 3353 9975 3355
rect 8889 3319 8905 3353
rect 8905 3319 8923 3353
rect 8961 3319 8973 3353
rect 8973 3319 8995 3353
rect 9033 3319 9041 3353
rect 9041 3319 9067 3353
rect 9105 3319 9109 3353
rect 9109 3319 9139 3353
rect 9177 3319 9211 3353
rect 9249 3319 9279 3353
rect 9279 3319 9283 3353
rect 9321 3319 9347 3353
rect 9347 3319 9355 3353
rect 9393 3319 9415 3353
rect 9415 3319 9427 3353
rect 9465 3319 9483 3353
rect 9483 3319 9499 3353
rect 9537 3319 9551 3353
rect 9551 3319 9571 3353
rect 9609 3319 9619 3353
rect 9619 3319 9643 3353
rect 9681 3319 9687 3353
rect 9687 3319 9715 3353
rect 9753 3319 9755 3353
rect 9755 3319 9787 3353
rect 9825 3319 9859 3353
rect 9941 3321 9975 3353
rect 8482 3282 8516 3284
rect 8482 3250 8516 3282
rect 8482 3176 8516 3210
rect 9941 3224 9975 3254
rect 9941 3220 9975 3224
rect 10070 3335 10104 3337
rect 10186 3336 10220 3370
rect 10258 3336 10290 3370
rect 10290 3336 10292 3370
rect 10330 3336 10358 3370
rect 10358 3336 10364 3370
rect 10402 3336 10426 3370
rect 10426 3336 10436 3370
rect 10474 3336 10494 3370
rect 10494 3336 10508 3370
rect 10546 3336 10562 3370
rect 10562 3336 10580 3370
rect 10618 3336 10630 3370
rect 10630 3336 10652 3370
rect 10690 3336 10698 3370
rect 10698 3336 10724 3370
rect 10762 3336 10766 3370
rect 10766 3336 10796 3370
rect 10834 3336 10868 3370
rect 10906 3336 10936 3370
rect 10936 3336 10940 3370
rect 10978 3336 11004 3370
rect 11004 3336 11012 3370
rect 11050 3336 11072 3370
rect 11072 3336 11084 3370
rect 11122 3336 11140 3370
rect 11140 3336 11156 3370
rect 11298 3382 11332 3393
rect 19973 3586 20007 3599
rect 19973 3565 19975 3586
rect 19975 3565 20007 3586
rect 19973 3518 20007 3526
rect 19973 3492 19975 3518
rect 19975 3492 20007 3518
rect 19973 3450 20007 3454
rect 19973 3420 19975 3450
rect 19975 3420 20007 3450
rect 11298 3359 11322 3382
rect 11322 3359 11332 3382
rect 11565 3348 11594 3377
rect 11594 3348 11599 3377
rect 11638 3348 11662 3377
rect 11662 3348 11672 3377
rect 11711 3348 11730 3377
rect 11730 3348 11745 3377
rect 11784 3348 11798 3377
rect 11798 3348 11818 3377
rect 11857 3348 11866 3377
rect 11866 3348 11891 3377
rect 11930 3348 11934 3377
rect 11934 3348 11964 3377
rect 12003 3348 12036 3377
rect 12036 3348 12037 3377
rect 12076 3348 12104 3377
rect 12104 3348 12110 3377
rect 12149 3348 12172 3377
rect 12172 3348 12183 3377
rect 12222 3348 12240 3377
rect 12240 3348 12256 3377
rect 12295 3348 12308 3377
rect 12308 3348 12329 3377
rect 12368 3348 12376 3377
rect 12376 3348 12402 3377
rect 12441 3348 12444 3377
rect 12444 3348 12475 3377
rect 12514 3348 12546 3377
rect 12546 3348 12548 3377
rect 12587 3348 12614 3377
rect 12614 3348 12621 3377
rect 12660 3348 12682 3377
rect 12682 3348 12694 3377
rect 12733 3348 12750 3377
rect 12750 3348 12767 3377
rect 12806 3348 12818 3377
rect 12818 3348 12840 3377
rect 12879 3348 12886 3377
rect 12886 3348 12913 3377
rect 12952 3348 12954 3377
rect 12954 3348 12986 3377
rect 13025 3348 13056 3377
rect 13056 3348 13059 3377
rect 13098 3348 13124 3377
rect 13124 3348 13132 3377
rect 13171 3348 13192 3377
rect 13192 3348 13205 3377
rect 13244 3348 13260 3377
rect 13260 3348 13278 3377
rect 13317 3348 13328 3377
rect 13328 3348 13351 3377
rect 13390 3348 13396 3377
rect 13396 3348 13424 3377
rect 13463 3348 13464 3377
rect 13464 3348 13497 3377
rect 13536 3348 13566 3377
rect 13566 3348 13570 3377
rect 13609 3348 13634 3377
rect 13634 3348 13643 3377
rect 13682 3348 13702 3377
rect 13702 3348 13716 3377
rect 13755 3348 13770 3377
rect 13770 3348 13789 3377
rect 13828 3348 13838 3377
rect 13838 3348 13862 3377
rect 13901 3348 13906 3377
rect 13906 3348 13935 3377
rect 13974 3348 14008 3377
rect 14047 3348 14076 3377
rect 14076 3348 14081 3377
rect 14120 3348 14144 3377
rect 14144 3348 14154 3377
rect 14193 3348 14212 3377
rect 14212 3348 14227 3377
rect 14266 3348 14280 3377
rect 14280 3348 14300 3377
rect 14339 3348 14348 3377
rect 14348 3348 14373 3377
rect 14412 3348 14416 3377
rect 14416 3348 14446 3377
rect 14485 3348 14518 3377
rect 14518 3348 14519 3377
rect 14558 3348 14586 3377
rect 14586 3348 14592 3377
rect 14631 3348 14654 3377
rect 14654 3348 14665 3377
rect 14704 3348 14722 3377
rect 14722 3348 14738 3377
rect 14777 3348 14790 3377
rect 14790 3348 14811 3377
rect 14849 3348 14858 3377
rect 14858 3348 14883 3377
rect 14921 3348 14926 3377
rect 14926 3348 14955 3377
rect 14993 3348 14994 3377
rect 14994 3348 15027 3377
rect 15065 3348 15096 3377
rect 15096 3348 15099 3377
rect 15137 3348 15164 3377
rect 15164 3348 15171 3377
rect 15209 3348 15232 3377
rect 15232 3348 15243 3377
rect 15281 3348 15300 3377
rect 15300 3348 15315 3377
rect 15353 3348 15368 3377
rect 15368 3348 15387 3377
rect 15425 3348 15436 3377
rect 15436 3348 15459 3377
rect 15497 3348 15504 3377
rect 15504 3348 15531 3377
rect 15569 3348 15572 3377
rect 15572 3348 15603 3377
rect 15641 3348 15674 3377
rect 15674 3348 15675 3377
rect 15713 3348 15742 3377
rect 15742 3348 15747 3377
rect 15785 3348 15810 3377
rect 15810 3348 15819 3377
rect 15857 3348 15878 3377
rect 15878 3348 15891 3377
rect 15929 3348 15946 3377
rect 15946 3348 15963 3377
rect 16001 3348 16014 3377
rect 16014 3348 16035 3377
rect 16073 3348 16082 3377
rect 16082 3348 16107 3377
rect 16145 3348 16150 3377
rect 16150 3348 16179 3377
rect 16217 3348 16218 3377
rect 16218 3348 16251 3377
rect 16289 3348 16320 3377
rect 16320 3348 16323 3377
rect 16361 3348 16388 3377
rect 16388 3348 16395 3377
rect 16433 3348 16456 3377
rect 16456 3348 16467 3377
rect 16505 3348 16524 3377
rect 16524 3348 16539 3377
rect 16577 3348 16592 3377
rect 16592 3348 16611 3377
rect 16649 3348 16660 3377
rect 16660 3348 16683 3377
rect 16721 3348 16728 3377
rect 16728 3348 16755 3377
rect 16793 3348 16796 3377
rect 16796 3348 16827 3377
rect 16865 3348 16898 3377
rect 16898 3348 16899 3377
rect 16937 3348 16966 3377
rect 16966 3348 16971 3377
rect 17009 3348 17034 3377
rect 17034 3348 17043 3377
rect 17081 3348 17102 3377
rect 17102 3348 17115 3377
rect 17153 3348 17170 3377
rect 17170 3348 17187 3377
rect 17225 3348 17238 3377
rect 17238 3348 17259 3377
rect 17297 3348 17306 3377
rect 17306 3348 17331 3377
rect 17369 3348 17374 3377
rect 17374 3348 17403 3377
rect 17441 3348 17442 3377
rect 17442 3348 17475 3377
rect 17513 3348 17544 3377
rect 17544 3348 17547 3377
rect 17585 3348 17612 3377
rect 17612 3348 17619 3377
rect 17657 3348 17680 3377
rect 17680 3348 17691 3377
rect 17729 3348 17748 3377
rect 17748 3348 17763 3377
rect 17801 3348 17816 3377
rect 17816 3348 17835 3377
rect 17873 3348 17884 3377
rect 17884 3348 17907 3377
rect 17945 3348 17952 3377
rect 17952 3348 17979 3377
rect 18017 3348 18020 3377
rect 18020 3348 18051 3377
rect 18089 3348 18122 3377
rect 18122 3348 18123 3377
rect 18161 3348 18190 3377
rect 18190 3348 18195 3377
rect 18233 3348 18258 3377
rect 18258 3348 18267 3377
rect 18305 3348 18326 3377
rect 18326 3348 18339 3377
rect 18377 3348 18394 3377
rect 18394 3348 18411 3377
rect 18449 3348 18462 3377
rect 18462 3348 18483 3377
rect 18521 3348 18530 3377
rect 18530 3348 18555 3377
rect 18593 3348 18598 3377
rect 18598 3348 18627 3377
rect 18665 3348 18666 3377
rect 18666 3348 18699 3377
rect 18737 3348 18768 3377
rect 18768 3348 18771 3377
rect 18809 3348 18836 3377
rect 18836 3348 18843 3377
rect 18881 3348 18904 3377
rect 18904 3348 18915 3377
rect 18953 3348 18972 3377
rect 18972 3348 18987 3377
rect 19025 3348 19040 3377
rect 19040 3348 19059 3377
rect 19097 3348 19108 3377
rect 19108 3348 19131 3377
rect 19169 3348 19176 3377
rect 19176 3348 19203 3377
rect 19241 3348 19244 3377
rect 19244 3348 19275 3377
rect 19313 3348 19346 3377
rect 19346 3348 19347 3377
rect 19385 3348 19414 3377
rect 19414 3348 19419 3377
rect 19457 3348 19482 3377
rect 19482 3348 19491 3377
rect 19529 3348 19550 3377
rect 19550 3348 19563 3377
rect 19601 3348 19618 3377
rect 19618 3348 19635 3377
rect 19673 3348 19686 3377
rect 19686 3348 19707 3377
rect 19745 3348 19754 3377
rect 19754 3348 19779 3377
rect 19817 3348 19822 3377
rect 19822 3348 19851 3377
rect 19889 3348 19890 3377
rect 19890 3348 19923 3377
rect 10070 3303 10104 3335
rect 10070 3233 10104 3265
rect 10070 3231 10104 3233
rect 11565 3343 11599 3348
rect 11638 3343 11672 3348
rect 11711 3343 11745 3348
rect 11784 3343 11818 3348
rect 11857 3343 11891 3348
rect 11930 3343 11964 3348
rect 12003 3343 12037 3348
rect 12076 3343 12110 3348
rect 12149 3343 12183 3348
rect 12222 3343 12256 3348
rect 12295 3343 12329 3348
rect 12368 3343 12402 3348
rect 12441 3343 12475 3348
rect 12514 3343 12548 3348
rect 12587 3343 12621 3348
rect 12660 3343 12694 3348
rect 12733 3343 12767 3348
rect 12806 3343 12840 3348
rect 12879 3343 12913 3348
rect 12952 3343 12986 3348
rect 13025 3343 13059 3348
rect 13098 3343 13132 3348
rect 13171 3343 13205 3348
rect 13244 3343 13278 3348
rect 13317 3343 13351 3348
rect 13390 3343 13424 3348
rect 13463 3343 13497 3348
rect 13536 3343 13570 3348
rect 13609 3343 13643 3348
rect 13682 3343 13716 3348
rect 13755 3343 13789 3348
rect 13828 3343 13862 3348
rect 13901 3343 13935 3348
rect 13974 3343 14008 3348
rect 14047 3343 14081 3348
rect 14120 3343 14154 3348
rect 14193 3343 14227 3348
rect 14266 3343 14300 3348
rect 14339 3343 14373 3348
rect 14412 3343 14446 3348
rect 14485 3343 14519 3348
rect 14558 3343 14592 3348
rect 14631 3343 14665 3348
rect 14704 3343 14738 3348
rect 14777 3343 14811 3348
rect 14849 3343 14883 3348
rect 14921 3343 14955 3348
rect 14993 3343 15027 3348
rect 15065 3343 15099 3348
rect 15137 3343 15171 3348
rect 15209 3343 15243 3348
rect 15281 3343 15315 3348
rect 15353 3343 15387 3348
rect 15425 3343 15459 3348
rect 15497 3343 15531 3348
rect 15569 3343 15603 3348
rect 15641 3343 15675 3348
rect 15713 3343 15747 3348
rect 15785 3343 15819 3348
rect 15857 3343 15891 3348
rect 15929 3343 15963 3348
rect 16001 3343 16035 3348
rect 16073 3343 16107 3348
rect 16145 3343 16179 3348
rect 16217 3343 16251 3348
rect 16289 3343 16323 3348
rect 16361 3343 16395 3348
rect 16433 3343 16467 3348
rect 16505 3343 16539 3348
rect 16577 3343 16611 3348
rect 16649 3343 16683 3348
rect 16721 3343 16755 3348
rect 16793 3343 16827 3348
rect 16865 3343 16899 3348
rect 16937 3343 16971 3348
rect 17009 3343 17043 3348
rect 17081 3343 17115 3348
rect 17153 3343 17187 3348
rect 17225 3343 17259 3348
rect 17297 3343 17331 3348
rect 17369 3343 17403 3348
rect 17441 3343 17475 3348
rect 17513 3343 17547 3348
rect 17585 3343 17619 3348
rect 17657 3343 17691 3348
rect 17729 3343 17763 3348
rect 17801 3343 17835 3348
rect 17873 3343 17907 3348
rect 17945 3343 17979 3348
rect 18017 3343 18051 3348
rect 18089 3343 18123 3348
rect 18161 3343 18195 3348
rect 18233 3343 18267 3348
rect 18305 3343 18339 3348
rect 18377 3343 18411 3348
rect 18449 3343 18483 3348
rect 18521 3343 18555 3348
rect 18593 3343 18627 3348
rect 18665 3343 18699 3348
rect 18737 3343 18771 3348
rect 18809 3343 18843 3348
rect 18881 3343 18915 3348
rect 18953 3343 18987 3348
rect 19025 3343 19059 3348
rect 19097 3343 19131 3348
rect 19169 3343 19203 3348
rect 19241 3343 19275 3348
rect 19313 3343 19347 3348
rect 19385 3343 19419 3348
rect 19457 3343 19491 3348
rect 19529 3343 19563 3348
rect 19601 3343 19635 3348
rect 19673 3343 19707 3348
rect 19745 3343 19779 3348
rect 19817 3343 19851 3348
rect 19889 3343 19923 3348
rect 11298 3281 11332 3315
rect 8889 3163 8905 3197
rect 8905 3163 8923 3197
rect 8961 3163 8973 3197
rect 8973 3163 8995 3197
rect 9033 3163 9041 3197
rect 9041 3163 9067 3197
rect 9105 3163 9109 3197
rect 9109 3163 9139 3197
rect 9177 3163 9211 3197
rect 9249 3163 9279 3197
rect 9279 3163 9283 3197
rect 9321 3163 9347 3197
rect 9347 3163 9355 3197
rect 9393 3163 9415 3197
rect 9415 3163 9427 3197
rect 9465 3163 9483 3197
rect 9483 3163 9499 3197
rect 9537 3163 9551 3197
rect 9551 3163 9571 3197
rect 9609 3163 9619 3197
rect 9619 3163 9643 3197
rect 9681 3163 9687 3197
rect 9687 3163 9715 3197
rect 9753 3163 9755 3197
rect 9755 3163 9787 3197
rect 9825 3163 9859 3197
rect 10186 3180 10220 3214
rect 10258 3180 10290 3214
rect 10290 3180 10292 3214
rect 10330 3180 10358 3214
rect 10358 3180 10364 3214
rect 10402 3180 10426 3214
rect 10426 3180 10436 3214
rect 10474 3180 10494 3214
rect 10494 3180 10508 3214
rect 10546 3180 10562 3214
rect 10562 3180 10580 3214
rect 10618 3180 10630 3214
rect 10630 3180 10652 3214
rect 10690 3180 10698 3214
rect 10698 3180 10724 3214
rect 10762 3180 10766 3214
rect 10766 3180 10796 3214
rect 10834 3180 10868 3214
rect 10906 3180 10936 3214
rect 10936 3180 10940 3214
rect 10978 3180 11004 3214
rect 11004 3180 11012 3214
rect 11050 3180 11072 3214
rect 11072 3180 11084 3214
rect 11122 3180 11140 3214
rect 11140 3180 11156 3214
rect 11298 3203 11332 3237
rect 17954 3241 17988 3275
rect 3456 3077 3490 3094
rect 3528 3077 3562 3094
rect 3600 3077 3634 3094
rect 3672 3077 3706 3094
rect 3744 3077 3778 3094
rect 8482 3106 8516 3136
rect 8482 3102 8516 3106
rect 17104 3195 17117 3216
rect 17117 3195 17138 3216
rect 17189 3195 17219 3216
rect 17219 3195 17223 3216
rect 17273 3195 17287 3216
rect 17287 3195 17307 3216
rect 17357 3195 17389 3216
rect 17389 3195 17391 3216
rect 17441 3195 17457 3216
rect 17457 3195 17475 3216
rect 17525 3195 17559 3216
rect 17104 3182 17138 3195
rect 17189 3182 17223 3195
rect 17273 3182 17307 3195
rect 17357 3182 17391 3195
rect 17441 3182 17475 3195
rect 17525 3182 17559 3195
rect 11298 3125 11332 3159
rect 8482 3036 8516 3062
rect 8482 3028 8516 3036
rect 10362 3053 10396 3087
rect 10434 3053 10435 3087
rect 10435 3053 10468 3087
rect 10506 3053 10508 3087
rect 10508 3053 10540 3087
rect 10578 3053 10581 3087
rect 10581 3053 10612 3087
rect 10650 3053 10654 3087
rect 10654 3053 10684 3087
rect 10722 3053 10726 3087
rect 10726 3053 10756 3087
rect 10794 3053 10798 3087
rect 10798 3053 10828 3087
rect 10866 3053 10870 3087
rect 10870 3053 10900 3087
rect 10938 3053 10942 3087
rect 10942 3053 10972 3087
rect 11010 3053 11014 3087
rect 11014 3053 11044 3087
rect 11082 3053 11086 3087
rect 11086 3053 11116 3087
rect 11154 3053 11158 3087
rect 11158 3053 11188 3087
rect 11226 3053 11230 3087
rect 11230 3053 11260 3087
rect 17619 3168 17653 3202
rect 17619 3100 17653 3130
rect 17619 3096 17653 3100
rect 17207 3019 17219 3047
rect 17219 3019 17241 3047
rect 17291 3019 17321 3047
rect 17321 3019 17325 3047
rect 17374 3019 17389 3047
rect 17389 3019 17408 3047
rect 17457 3019 17491 3047
rect 17798 3148 17832 3178
rect 17798 3144 17832 3148
rect 17798 3080 17832 3106
rect 17798 3072 17832 3080
rect 18900 3271 18934 3305
rect 17954 3182 17988 3203
rect 17954 3169 17988 3182
rect 18110 3114 18144 3148
rect 18110 3046 18144 3076
rect 18110 3042 18144 3046
rect 18282 3114 18316 3148
rect 18282 3046 18316 3076
rect 18282 3042 18316 3046
rect 18438 3182 18472 3208
rect 18438 3174 18472 3182
rect 18438 3114 18472 3136
rect 18438 3102 18472 3114
rect 18438 3046 18472 3064
rect 18438 3030 18472 3046
rect 18594 3114 18628 3148
rect 18594 3046 18628 3076
rect 18594 3042 18628 3046
rect 18744 3114 18778 3148
rect 18744 3046 18778 3076
rect 18744 3042 18778 3046
rect 18900 3216 18934 3233
rect 18900 3199 18934 3216
rect 19056 3114 19090 3148
rect 19056 3046 19090 3076
rect 19056 3042 19090 3046
rect 20002 3182 20036 3216
rect 20002 3109 20036 3143
rect 20002 3036 20036 3070
rect 17207 3013 17241 3019
rect 17291 3013 17325 3019
rect 17374 3013 17408 3019
rect 17457 3013 17491 3019
rect 8482 2954 8516 2988
rect 8867 2968 8895 3002
rect 8895 2968 8901 3002
rect 8942 2968 8964 3002
rect 8964 2968 8976 3002
rect 9017 2968 9033 3002
rect 9033 2968 9051 3002
rect 9092 2968 9102 3002
rect 9102 2968 9126 3002
rect 9167 2968 9171 3002
rect 9171 2968 9201 3002
rect 9242 2968 9274 3002
rect 9274 2968 9276 3002
rect 9317 2968 9343 3002
rect 9343 2968 9351 3002
rect 9392 2968 9412 3002
rect 9412 2968 9426 3002
rect 9467 2968 9481 3002
rect 9481 2968 9501 3002
rect 9542 2968 9550 3002
rect 9550 2968 9576 3002
rect 9617 2968 9619 3002
rect 9619 2968 9651 3002
rect 9692 2968 9723 3002
rect 9723 2968 9726 3002
rect 9767 2968 9792 3002
rect 9792 2968 9801 3002
rect 9842 2968 9861 3002
rect 9861 2968 9876 3002
rect 9917 2968 9929 3002
rect 9929 2968 9951 3002
rect 9992 2968 9997 3002
rect 9997 2968 10026 3002
rect 10067 2968 10099 3002
rect 10099 2968 10101 3002
rect 10142 2968 10167 3002
rect 10167 2968 10176 3002
rect 10217 2968 10235 3002
rect 10235 2968 10251 3002
rect 10291 2968 10303 3002
rect 10303 2968 10325 3002
rect 17855 2942 17889 2976
rect 17954 2942 17988 2976
rect 18053 2942 18087 2976
rect 18339 2942 18373 2976
rect 18438 2942 18472 2976
rect 18537 2942 18571 2976
rect 18801 2942 18835 2976
rect 18900 2942 18934 2976
rect 18999 2942 19033 2976
rect 20002 2964 20036 2998
rect 8482 2880 8516 2914
rect 20002 2892 20036 2926
rect 8482 2806 8516 2840
rect 10488 2822 10522 2856
rect 10568 2855 10602 2856
rect 10647 2855 10681 2856
rect 10726 2855 10760 2856
rect 10805 2855 10839 2856
rect 10884 2855 10918 2856
rect 10963 2855 10997 2856
rect 11042 2855 11076 2856
rect 11121 2855 11155 2856
rect 11200 2855 11234 2856
rect 11279 2855 11313 2856
rect 10568 2822 10596 2855
rect 10596 2822 10602 2855
rect 10647 2822 10664 2855
rect 10664 2822 10681 2855
rect 10726 2822 10732 2855
rect 10732 2822 10760 2855
rect 10805 2822 10834 2855
rect 10834 2822 10839 2855
rect 10884 2822 10902 2855
rect 10902 2822 10918 2855
rect 10963 2822 10970 2855
rect 10970 2822 10997 2855
rect 11042 2822 11072 2855
rect 11072 2822 11076 2855
rect 11121 2822 11140 2855
rect 11140 2822 11155 2855
rect 11200 2822 11208 2855
rect 11208 2822 11234 2855
rect 11279 2822 11310 2855
rect 11310 2822 11313 2855
rect 12253 2821 12262 2849
rect 12262 2821 12287 2849
rect 12325 2821 12330 2849
rect 12330 2821 12359 2849
rect 12397 2821 12398 2849
rect 12398 2821 12431 2849
rect 12469 2821 12500 2849
rect 12500 2821 12503 2849
rect 12542 2821 12568 2849
rect 12568 2821 12576 2849
rect 12615 2821 12636 2849
rect 12636 2821 12649 2849
rect 12688 2821 12704 2849
rect 12704 2821 12722 2849
rect 12761 2821 12772 2849
rect 12772 2821 12795 2849
rect 12834 2821 12840 2849
rect 12840 2821 12868 2849
rect 12907 2821 12908 2849
rect 12908 2821 12941 2849
rect 12980 2821 13010 2849
rect 13010 2821 13014 2849
rect 13053 2821 13078 2849
rect 13078 2821 13087 2849
rect 13126 2821 13146 2849
rect 13146 2821 13160 2849
rect 13199 2821 13214 2849
rect 13214 2821 13233 2849
rect 13272 2821 13282 2849
rect 13282 2821 13306 2849
rect 13345 2821 13350 2849
rect 13350 2821 13379 2849
rect 13418 2821 13452 2849
rect 13491 2821 13520 2849
rect 13520 2821 13525 2849
rect 13564 2821 13588 2849
rect 13588 2821 13598 2849
rect 13637 2821 13656 2849
rect 13656 2821 13671 2849
rect 13710 2821 13724 2849
rect 13724 2821 13744 2849
rect 13783 2821 13792 2849
rect 13792 2821 13817 2849
rect 13856 2821 13860 2849
rect 13860 2821 13890 2849
rect 13929 2821 13962 2849
rect 13962 2821 13963 2849
rect 14002 2821 14030 2849
rect 14030 2821 14036 2849
rect 14075 2821 14098 2849
rect 14098 2821 14109 2849
rect 14148 2821 14166 2849
rect 14166 2821 14182 2849
rect 14221 2821 14234 2849
rect 14234 2821 14255 2849
rect 14294 2821 14302 2849
rect 14302 2821 14328 2849
rect 14367 2821 14370 2849
rect 14370 2821 14401 2849
rect 14440 2821 14472 2849
rect 14472 2821 14474 2849
rect 14513 2821 14540 2849
rect 14540 2821 14547 2849
rect 14586 2821 14608 2849
rect 14608 2821 14620 2849
rect 14659 2821 14676 2849
rect 14676 2821 14693 2849
rect 14732 2821 14744 2849
rect 14744 2821 14766 2849
rect 14805 2821 14812 2849
rect 14812 2821 14839 2849
rect 14878 2821 14880 2849
rect 14880 2821 14912 2849
rect 14951 2821 14982 2849
rect 14982 2821 14985 2849
rect 15024 2821 15050 2849
rect 15050 2821 15058 2849
rect 15097 2821 15118 2849
rect 15118 2821 15131 2849
rect 15170 2821 15186 2849
rect 15186 2821 15204 2849
rect 15243 2821 15254 2849
rect 15254 2821 15277 2849
rect 15316 2821 15322 2849
rect 15322 2821 15350 2849
rect 15389 2821 15390 2849
rect 15390 2821 15423 2849
rect 15462 2821 15492 2849
rect 15492 2821 15496 2849
rect 15535 2821 15560 2849
rect 15560 2821 15569 2849
rect 15608 2821 15628 2849
rect 15628 2821 15642 2849
rect 15681 2821 15696 2849
rect 15696 2821 15715 2849
rect 15754 2821 15764 2849
rect 15764 2821 15788 2849
rect 15827 2821 15832 2849
rect 15832 2821 15861 2849
rect 8482 2732 8516 2766
rect 8482 2657 8516 2691
rect 8482 2582 8516 2616
rect 582 2518 598 2552
rect 598 2518 616 2552
rect 660 2518 668 2552
rect 668 2518 694 2552
rect 738 2518 772 2552
rect 815 2518 842 2552
rect 842 2518 849 2552
rect 892 2518 912 2552
rect 912 2518 926 2552
rect 969 2518 982 2552
rect 982 2518 1003 2552
rect 1046 2518 1053 2552
rect 1053 2518 1080 2552
rect 1123 2518 1124 2552
rect 1124 2518 1157 2552
rect 1200 2518 1232 2552
rect 1232 2518 1234 2552
rect 1277 2518 1303 2552
rect 1303 2518 1311 2552
rect 1354 2518 1374 2552
rect 1374 2518 1388 2552
rect 1431 2518 1445 2552
rect 1445 2518 1465 2552
rect 1508 2518 1516 2552
rect 1516 2518 1542 2552
rect 2245 2465 2271 2499
rect 2271 2465 2279 2499
rect 2323 2465 2339 2499
rect 2339 2465 2357 2499
rect 2400 2465 2407 2499
rect 2407 2465 2434 2499
rect 2510 2465 2543 2499
rect 2543 2465 2544 2499
rect 2583 2465 2611 2499
rect 2611 2465 2617 2499
rect 2656 2465 2679 2499
rect 2679 2465 2690 2499
rect 2729 2465 2747 2499
rect 2747 2465 2763 2499
rect 2802 2465 2815 2499
rect 2815 2465 2836 2499
rect 2875 2465 2883 2499
rect 2883 2465 2909 2499
rect 2948 2465 2951 2499
rect 2951 2465 2982 2499
rect 3021 2465 3053 2499
rect 3053 2465 3055 2499
rect 3094 2465 3121 2499
rect 3121 2465 3128 2499
rect 3167 2465 3189 2499
rect 3189 2465 3201 2499
rect 3240 2465 3257 2499
rect 3257 2465 3274 2499
rect 3313 2465 3325 2499
rect 3325 2465 3347 2499
rect 3386 2465 3393 2499
rect 3393 2465 3420 2499
rect 3459 2465 3461 2499
rect 3461 2465 3493 2499
rect 3532 2465 3563 2499
rect 3563 2465 3566 2499
rect 3605 2465 3631 2499
rect 3631 2465 3639 2499
rect 3678 2465 3699 2499
rect 3699 2465 3712 2499
rect 3751 2465 3767 2499
rect 3767 2465 3785 2499
rect 3824 2465 3835 2499
rect 3835 2465 3858 2499
rect 3897 2465 3903 2499
rect 3903 2465 3931 2499
rect 3970 2465 3971 2499
rect 3971 2465 4004 2499
rect 4043 2465 4073 2499
rect 4073 2465 4077 2499
rect 4116 2465 4141 2499
rect 4141 2465 4150 2499
rect 4189 2465 4209 2499
rect 4209 2465 4223 2499
rect 4262 2465 4277 2499
rect 4277 2465 4296 2499
rect 4335 2465 4345 2499
rect 4345 2465 4369 2499
rect 4408 2465 4413 2499
rect 4413 2465 4442 2499
rect 4481 2465 4515 2499
rect 4554 2465 4583 2499
rect 4583 2465 4588 2499
rect 4627 2465 4651 2499
rect 4651 2465 4661 2499
rect 4700 2465 4719 2499
rect 4719 2465 4734 2499
rect 4773 2465 4787 2499
rect 4787 2465 4807 2499
rect 4846 2465 4855 2499
rect 4855 2465 4880 2499
rect 4919 2465 4923 2499
rect 4923 2465 4953 2499
rect 4992 2465 5025 2499
rect 5025 2465 5026 2499
rect 5065 2465 5093 2499
rect 5093 2465 5099 2499
rect 5138 2465 5161 2499
rect 5161 2465 5172 2499
rect 5211 2465 5229 2499
rect 5229 2465 5245 2499
rect 5284 2465 5297 2499
rect 5297 2465 5318 2499
rect 5357 2465 5365 2499
rect 5365 2465 5391 2499
rect 5430 2465 5433 2499
rect 5433 2465 5464 2499
rect 5503 2465 5535 2499
rect 5535 2465 5537 2499
rect 5576 2465 5603 2499
rect 5603 2465 5610 2499
rect 5649 2465 5671 2499
rect 5671 2465 5683 2499
rect 5722 2465 5739 2499
rect 5739 2465 5756 2499
rect 5795 2465 5807 2499
rect 5807 2465 5829 2499
rect 5868 2465 5875 2499
rect 5875 2465 5902 2499
rect 5941 2465 5943 2499
rect 5943 2465 5975 2499
rect 6014 2465 6045 2499
rect 6045 2465 6048 2499
rect 6087 2465 6113 2499
rect 6113 2465 6121 2499
rect 6160 2465 6181 2499
rect 6181 2465 6194 2499
rect 6233 2465 6249 2499
rect 6249 2465 6267 2499
rect 6306 2465 6317 2499
rect 6317 2465 6340 2499
rect 6379 2465 6385 2499
rect 6385 2465 6413 2499
rect 6452 2465 6453 2499
rect 6453 2465 6486 2499
rect 6525 2465 6555 2499
rect 6555 2465 6559 2499
rect 6598 2465 6623 2499
rect 6623 2465 6632 2499
rect 6671 2465 6691 2499
rect 6691 2465 6705 2499
rect 6744 2465 6759 2499
rect 6759 2465 6778 2499
rect 6816 2465 6827 2499
rect 6827 2465 6850 2499
rect 6888 2465 6895 2499
rect 6895 2465 6922 2499
rect 6960 2465 6963 2499
rect 6963 2465 6994 2499
rect 7032 2465 7065 2499
rect 7065 2465 7066 2499
rect 7104 2465 7133 2499
rect 7133 2465 7138 2499
rect 7176 2465 7201 2499
rect 7201 2465 7210 2499
rect 7248 2465 7269 2499
rect 7269 2465 7282 2499
rect 7320 2465 7337 2499
rect 7337 2465 7354 2499
rect 7392 2465 7405 2499
rect 7405 2465 7426 2499
rect 7464 2465 7473 2499
rect 7473 2465 7498 2499
rect 7536 2465 7541 2499
rect 7541 2465 7570 2499
rect 7608 2465 7609 2499
rect 7609 2465 7642 2499
rect 7680 2465 7711 2499
rect 7711 2465 7714 2499
rect 7752 2465 7779 2499
rect 7779 2465 7786 2499
rect 7824 2465 7847 2499
rect 7847 2465 7858 2499
rect 7896 2465 7915 2499
rect 7915 2465 7930 2499
rect 7968 2465 7983 2499
rect 7983 2465 8002 2499
rect 8040 2465 8051 2499
rect 8051 2465 8074 2499
rect 8112 2465 8119 2499
rect 8119 2465 8146 2499
rect 8184 2465 8187 2499
rect 8187 2465 8218 2499
rect 8256 2465 8289 2499
rect 8289 2465 8290 2499
rect 8328 2465 8357 2499
rect 8357 2465 8362 2499
rect 8400 2465 8425 2499
rect 8425 2465 8434 2499
rect 466 2407 500 2441
rect 570 2399 586 2433
rect 586 2399 604 2433
rect 642 2399 654 2433
rect 654 2399 676 2433
rect 714 2399 722 2433
rect 722 2399 748 2433
rect 786 2399 790 2433
rect 790 2399 820 2433
rect 858 2399 892 2433
rect 930 2399 960 2433
rect 960 2399 964 2433
rect 1002 2399 1028 2433
rect 1028 2399 1036 2433
rect 1074 2399 1096 2433
rect 1096 2399 1108 2433
rect 1146 2399 1164 2433
rect 1164 2399 1180 2433
rect 1218 2399 1232 2433
rect 1232 2399 1252 2433
rect 1290 2399 1300 2433
rect 1300 2399 1324 2433
rect 1362 2399 1368 2433
rect 1368 2399 1396 2433
rect 1434 2399 1436 2433
rect 1436 2399 1468 2433
rect 1506 2399 1540 2433
rect 466 2335 500 2369
rect 466 2263 500 2297
rect 1622 2347 1656 2380
rect 1622 2346 1656 2347
rect 1622 2279 1656 2308
rect 570 2243 586 2277
rect 586 2243 604 2277
rect 642 2243 654 2277
rect 654 2243 676 2277
rect 714 2243 722 2277
rect 722 2243 748 2277
rect 786 2243 790 2277
rect 790 2243 820 2277
rect 858 2243 892 2277
rect 930 2243 960 2277
rect 960 2243 964 2277
rect 1002 2243 1028 2277
rect 1028 2243 1036 2277
rect 1074 2243 1096 2277
rect 1096 2243 1108 2277
rect 1146 2243 1164 2277
rect 1164 2243 1180 2277
rect 1218 2243 1232 2277
rect 1232 2243 1252 2277
rect 1290 2243 1300 2277
rect 1300 2243 1324 2277
rect 1362 2243 1368 2277
rect 1368 2243 1396 2277
rect 1434 2243 1436 2277
rect 1436 2243 1468 2277
rect 1506 2243 1540 2277
rect 1622 2274 1656 2279
rect 2151 2397 2185 2402
rect 2151 2368 2185 2397
rect 2151 2295 2185 2329
rect 466 2191 500 2225
rect 2151 2227 2185 2256
rect 2151 2222 2185 2227
rect 2443 2219 2452 2231
rect 2452 2219 2477 2231
rect 2535 2219 2555 2231
rect 2555 2219 2569 2231
rect 2627 2219 2659 2231
rect 2659 2219 2661 2231
rect 3138 2219 3142 2231
rect 3142 2219 3172 2231
rect 3211 2219 3245 2231
rect 3284 2219 3314 2231
rect 3314 2219 3318 2231
rect 3357 2219 3383 2231
rect 3383 2219 3391 2231
rect 3430 2219 3452 2231
rect 3452 2219 3464 2231
rect 3503 2219 3521 2231
rect 3521 2219 3537 2231
rect 3576 2219 3590 2231
rect 3590 2219 3610 2231
rect 3649 2219 3659 2231
rect 3659 2219 3683 2231
rect 3722 2219 3728 2231
rect 3728 2219 3756 2231
rect 3795 2219 3796 2231
rect 3796 2219 3829 2231
rect 3868 2219 3898 2231
rect 3898 2219 3902 2231
rect 3941 2219 3966 2231
rect 3966 2219 3975 2231
rect 4014 2219 4034 2231
rect 4034 2219 4048 2231
rect 4087 2219 4102 2231
rect 4102 2219 4121 2231
rect 4160 2219 4170 2231
rect 4170 2219 4194 2231
rect 4233 2219 4238 2231
rect 4238 2219 4267 2231
rect 4306 2219 4340 2231
rect 4379 2219 4408 2231
rect 4408 2219 4413 2231
rect 4452 2219 4476 2231
rect 4476 2219 4486 2231
rect 4525 2219 4544 2231
rect 4544 2219 4559 2231
rect 4598 2219 4612 2231
rect 4612 2219 4632 2231
rect 4671 2219 4680 2231
rect 4680 2219 4705 2231
rect 4744 2219 4748 2231
rect 4748 2219 4778 2231
rect 4817 2219 4850 2231
rect 4850 2219 4851 2231
rect 4890 2219 4918 2231
rect 4918 2219 4924 2231
rect 4963 2219 4986 2231
rect 4986 2219 4997 2231
rect 5036 2219 5054 2231
rect 5054 2219 5070 2231
rect 5109 2219 5122 2231
rect 5122 2219 5143 2231
rect 5182 2219 5190 2231
rect 5190 2219 5216 2231
rect 5255 2219 5258 2231
rect 5258 2219 5289 2231
rect 5328 2219 5360 2231
rect 5360 2219 5362 2231
rect 5401 2219 5428 2231
rect 5428 2219 5435 2231
rect 5474 2219 5496 2231
rect 5496 2219 5508 2231
rect 5547 2219 5564 2231
rect 5564 2219 5581 2231
rect 5620 2219 5632 2231
rect 5632 2219 5654 2231
rect 5693 2219 5700 2231
rect 5700 2219 5727 2231
rect 5766 2219 5768 2231
rect 5768 2219 5800 2231
rect 5839 2219 5870 2231
rect 5870 2219 5873 2231
rect 5912 2219 5938 2231
rect 5938 2219 5946 2231
rect 5985 2219 6006 2231
rect 6006 2219 6019 2231
rect 6058 2219 6074 2231
rect 6074 2219 6092 2231
rect 6131 2219 6142 2231
rect 6142 2219 6165 2231
rect 6204 2219 6210 2231
rect 6210 2219 6238 2231
rect 6277 2219 6278 2231
rect 6278 2219 6311 2231
rect 6350 2219 6380 2231
rect 6380 2219 6384 2231
rect 6423 2219 6448 2231
rect 6448 2219 6457 2231
rect 6496 2219 6516 2231
rect 6516 2219 6530 2231
rect 6569 2219 6584 2231
rect 6584 2219 6603 2231
rect 6641 2219 6652 2231
rect 6652 2219 6675 2231
rect 6713 2219 6720 2231
rect 6720 2219 6747 2231
rect 6785 2219 6788 2231
rect 6788 2219 6819 2231
rect 6857 2219 6890 2231
rect 6890 2219 6891 2231
rect 6929 2219 6958 2231
rect 6958 2219 6963 2231
rect 2443 2197 2477 2219
rect 2535 2197 2569 2219
rect 2627 2197 2661 2219
rect 2790 2185 2824 2219
rect 2882 2185 2916 2219
rect 2974 2185 3008 2219
rect 3138 2197 3172 2219
rect 3211 2197 3245 2219
rect 3284 2197 3318 2219
rect 3357 2197 3391 2219
rect 3430 2197 3464 2219
rect 3503 2197 3537 2219
rect 3576 2197 3610 2219
rect 3649 2197 3683 2219
rect 3722 2197 3756 2219
rect 3795 2197 3829 2219
rect 3868 2197 3902 2219
rect 3941 2197 3975 2219
rect 4014 2197 4048 2219
rect 4087 2197 4121 2219
rect 4160 2197 4194 2219
rect 4233 2197 4267 2219
rect 4306 2197 4340 2219
rect 4379 2197 4413 2219
rect 4452 2197 4486 2219
rect 4525 2197 4559 2219
rect 4598 2197 4632 2219
rect 4671 2197 4705 2219
rect 4744 2197 4778 2219
rect 4817 2197 4851 2219
rect 4890 2197 4924 2219
rect 4963 2197 4997 2219
rect 5036 2197 5070 2219
rect 5109 2197 5143 2219
rect 5182 2197 5216 2219
rect 5255 2197 5289 2219
rect 5328 2197 5362 2219
rect 5401 2197 5435 2219
rect 5474 2197 5508 2219
rect 5547 2197 5581 2219
rect 5620 2197 5654 2219
rect 5693 2197 5727 2219
rect 5766 2197 5800 2219
rect 5839 2197 5873 2219
rect 5912 2197 5946 2219
rect 5985 2197 6019 2219
rect 6058 2197 6092 2219
rect 6131 2197 6165 2219
rect 6204 2197 6238 2219
rect 6277 2197 6311 2219
rect 6350 2197 6384 2219
rect 6423 2197 6457 2219
rect 6496 2197 6530 2219
rect 6569 2197 6603 2219
rect 6641 2197 6675 2219
rect 6713 2197 6747 2219
rect 6785 2197 6819 2219
rect 6857 2197 6891 2219
rect 6929 2197 6963 2219
rect 7667 2203 7685 2237
rect 7685 2203 7701 2237
rect 7744 2203 7753 2237
rect 7753 2203 7778 2237
rect 7821 2203 7855 2237
rect 7898 2203 7923 2237
rect 7923 2203 7932 2237
rect 7975 2203 7991 2237
rect 7991 2203 8009 2237
rect 8052 2203 8059 2237
rect 8059 2203 8086 2237
rect 8129 2203 8161 2237
rect 8161 2203 8163 2237
rect 8206 2203 8229 2237
rect 8229 2203 8240 2237
rect 8283 2203 8297 2237
rect 8297 2203 8317 2237
rect 8359 2203 8365 2237
rect 8365 2203 8393 2237
rect 8435 2203 8469 2237
rect 8613 2211 8647 2245
rect 466 2119 500 2153
rect 466 2047 500 2081
rect 466 1975 500 2009
rect 466 1903 500 1937
rect 574 2130 598 2162
rect 598 2130 608 2162
rect 648 2130 669 2162
rect 669 2130 682 2162
rect 722 2130 740 2162
rect 740 2130 756 2162
rect 796 2130 811 2162
rect 811 2130 830 2162
rect 870 2130 882 2162
rect 882 2130 904 2162
rect 944 2130 953 2162
rect 953 2130 978 2162
rect 1017 2130 1024 2162
rect 1024 2130 1051 2162
rect 1090 2130 1095 2162
rect 1095 2130 1124 2162
rect 1163 2130 1166 2162
rect 1166 2130 1197 2162
rect 1236 2130 1270 2162
rect 1309 2130 1340 2162
rect 1340 2130 1343 2162
rect 1382 2130 1410 2162
rect 1410 2130 1416 2162
rect 1455 2130 1480 2162
rect 1480 2130 1489 2162
rect 1528 2130 1550 2162
rect 1550 2130 1562 2162
rect 574 2128 608 2130
rect 648 2128 682 2130
rect 722 2128 756 2130
rect 796 2128 830 2130
rect 870 2128 904 2130
rect 944 2128 978 2130
rect 1017 2128 1051 2130
rect 1090 2128 1124 2130
rect 1163 2128 1197 2130
rect 1236 2128 1270 2130
rect 1309 2128 1343 2130
rect 1382 2128 1416 2130
rect 1455 2128 1489 2130
rect 1528 2128 1562 2130
rect 574 2028 608 2062
rect 648 2028 682 2062
rect 722 2028 756 2062
rect 796 2028 830 2062
rect 870 2028 904 2062
rect 944 2028 978 2062
rect 1017 2028 1051 2062
rect 1090 2028 1124 2062
rect 1163 2028 1197 2062
rect 1236 2028 1270 2062
rect 1309 2028 1343 2062
rect 1382 2028 1416 2062
rect 1455 2028 1489 2062
rect 1528 2028 1562 2062
rect 574 1960 608 1962
rect 648 1960 682 1962
rect 722 1960 756 1962
rect 796 1960 830 1962
rect 870 1960 904 1962
rect 944 1960 978 1962
rect 1017 1960 1051 1962
rect 1090 1960 1124 1962
rect 1163 1960 1197 1962
rect 1236 1960 1270 1962
rect 1309 1960 1343 1962
rect 1382 1960 1416 1962
rect 1455 1960 1489 1962
rect 1528 1960 1562 1962
rect 574 1928 598 1960
rect 598 1928 608 1960
rect 648 1928 669 1960
rect 669 1928 682 1960
rect 722 1928 740 1960
rect 740 1928 756 1960
rect 796 1928 811 1960
rect 811 1928 830 1960
rect 870 1928 882 1960
rect 882 1928 904 1960
rect 944 1928 953 1960
rect 953 1928 978 1960
rect 1017 1928 1024 1960
rect 1024 1928 1051 1960
rect 1090 1928 1095 1960
rect 1095 1928 1124 1960
rect 1163 1928 1166 1960
rect 1166 1928 1197 1960
rect 1236 1928 1270 1960
rect 1309 1928 1340 1960
rect 1340 1928 1343 1960
rect 1382 1928 1410 1960
rect 1410 1928 1416 1960
rect 1455 1928 1480 1960
rect 1480 1928 1489 1960
rect 1528 1928 1550 1960
rect 1550 1928 1562 1960
rect 2151 2159 2185 2182
rect 2151 2148 2185 2159
rect 8613 2158 8647 2173
rect 2151 2091 2185 2108
rect 2151 2074 2185 2091
rect 2420 2103 2436 2137
rect 2436 2103 2454 2137
rect 2492 2103 2504 2137
rect 2504 2103 2526 2137
rect 2564 2103 2572 2137
rect 2572 2103 2598 2137
rect 2636 2103 2640 2137
rect 2640 2103 2670 2137
rect 2708 2103 2742 2137
rect 2780 2103 2810 2137
rect 2810 2103 2814 2137
rect 2852 2103 2878 2137
rect 2878 2103 2886 2137
rect 2924 2103 2946 2137
rect 2946 2103 2958 2137
rect 2996 2103 3014 2137
rect 3014 2103 3030 2137
rect 3068 2103 3082 2137
rect 3082 2103 3102 2137
rect 3140 2103 3150 2137
rect 3150 2103 3174 2137
rect 3212 2103 3218 2137
rect 3218 2103 3246 2137
rect 3284 2103 3286 2137
rect 3286 2103 3318 2137
rect 3356 2103 3388 2137
rect 3388 2103 3390 2137
rect 3428 2103 3456 2137
rect 3456 2103 3462 2137
rect 3500 2103 3524 2137
rect 3524 2103 3534 2137
rect 3572 2103 3592 2137
rect 3592 2103 3606 2137
rect 3644 2103 3660 2137
rect 3660 2103 3678 2137
rect 3716 2103 3728 2137
rect 3728 2103 3750 2137
rect 3788 2103 3796 2137
rect 3796 2103 3822 2137
rect 3860 2103 3864 2137
rect 3864 2103 3894 2137
rect 3932 2103 3966 2137
rect 4004 2103 4034 2137
rect 4034 2103 4038 2137
rect 4076 2103 4102 2137
rect 4102 2103 4110 2137
rect 4148 2103 4170 2137
rect 4170 2103 4182 2137
rect 4220 2103 4238 2137
rect 4238 2103 4254 2137
rect 4292 2103 4306 2137
rect 4306 2103 4326 2137
rect 4364 2103 4374 2137
rect 4374 2103 4398 2137
rect 4688 2103 4712 2137
rect 4712 2103 4722 2137
rect 4760 2103 4780 2137
rect 4780 2103 4794 2137
rect 4832 2103 4848 2137
rect 4848 2103 4866 2137
rect 4904 2103 4916 2137
rect 4916 2103 4938 2137
rect 4976 2103 4984 2137
rect 4984 2103 5010 2137
rect 5048 2103 5052 2137
rect 5052 2103 5082 2137
rect 5120 2103 5154 2137
rect 5192 2103 5222 2137
rect 5222 2103 5226 2137
rect 5264 2103 5290 2137
rect 5290 2103 5298 2137
rect 5336 2103 5358 2137
rect 5358 2103 5370 2137
rect 5408 2103 5426 2137
rect 5426 2103 5442 2137
rect 5480 2103 5494 2137
rect 5494 2103 5514 2137
rect 5552 2103 5562 2137
rect 5562 2103 5586 2137
rect 5624 2103 5630 2137
rect 5630 2103 5658 2137
rect 5696 2103 5698 2137
rect 5698 2103 5730 2137
rect 5768 2103 5800 2137
rect 5800 2103 5802 2137
rect 5840 2103 5868 2137
rect 5868 2103 5874 2137
rect 5912 2103 5936 2137
rect 5936 2103 5946 2137
rect 5984 2103 6004 2137
rect 6004 2103 6018 2137
rect 6056 2103 6072 2137
rect 6072 2103 6090 2137
rect 6128 2103 6140 2137
rect 6140 2103 6162 2137
rect 6200 2103 6208 2137
rect 6208 2103 6234 2137
rect 6272 2103 6276 2137
rect 6276 2103 6306 2137
rect 6344 2103 6378 2137
rect 6416 2103 6446 2137
rect 6446 2103 6450 2137
rect 6488 2103 6514 2137
rect 6514 2103 6522 2137
rect 6560 2103 6582 2137
rect 6582 2103 6594 2137
rect 6632 2103 6650 2137
rect 6650 2103 6666 2137
rect 8613 2139 8639 2158
rect 8639 2139 8647 2158
rect 2151 2023 2185 2034
rect 2151 2000 2185 2023
rect 466 1831 500 1865
rect 2151 1955 2185 1960
rect 2151 1926 2185 1955
rect 4472 2076 4506 2082
rect 4472 2048 4506 2076
rect 4472 1974 4506 2005
rect 4472 1971 4506 1974
rect 4472 1906 4506 1928
rect 2151 1853 2185 1886
rect 2151 1852 2185 1853
rect 2420 1867 2436 1901
rect 2436 1867 2454 1901
rect 2492 1867 2504 1901
rect 2504 1867 2526 1901
rect 2564 1867 2572 1901
rect 2572 1867 2598 1901
rect 2636 1867 2640 1901
rect 2640 1867 2670 1901
rect 2708 1867 2742 1901
rect 2780 1867 2810 1901
rect 2810 1867 2814 1901
rect 2852 1867 2878 1901
rect 2878 1867 2886 1901
rect 2924 1867 2946 1901
rect 2946 1867 2958 1901
rect 2996 1867 3014 1901
rect 3014 1867 3030 1901
rect 3068 1867 3082 1901
rect 3082 1867 3102 1901
rect 3140 1867 3150 1901
rect 3150 1867 3174 1901
rect 3212 1867 3218 1901
rect 3218 1867 3246 1901
rect 3284 1867 3286 1901
rect 3286 1867 3318 1901
rect 3356 1867 3388 1901
rect 3388 1867 3390 1901
rect 3428 1867 3456 1901
rect 3456 1867 3462 1901
rect 3500 1867 3524 1901
rect 3524 1867 3534 1901
rect 3572 1867 3592 1901
rect 3592 1867 3606 1901
rect 3644 1867 3660 1901
rect 3660 1867 3678 1901
rect 3716 1867 3728 1901
rect 3728 1867 3750 1901
rect 3788 1867 3796 1901
rect 3796 1867 3822 1901
rect 3860 1867 3864 1901
rect 3864 1867 3894 1901
rect 3932 1867 3966 1901
rect 4004 1867 4034 1901
rect 4034 1867 4038 1901
rect 4076 1867 4102 1901
rect 4102 1867 4110 1901
rect 4148 1867 4170 1901
rect 4170 1867 4182 1901
rect 4220 1867 4238 1901
rect 4238 1867 4254 1901
rect 4292 1867 4306 1901
rect 4306 1867 4326 1901
rect 4364 1867 4374 1901
rect 4374 1867 4398 1901
rect 4472 1894 4506 1906
rect 570 1807 586 1841
rect 586 1807 604 1841
rect 642 1807 654 1841
rect 654 1807 676 1841
rect 714 1807 722 1841
rect 722 1807 748 1841
rect 786 1807 790 1841
rect 790 1807 820 1841
rect 858 1807 892 1841
rect 930 1807 960 1841
rect 960 1807 964 1841
rect 1002 1807 1028 1841
rect 1028 1807 1036 1841
rect 1074 1807 1096 1841
rect 1096 1807 1108 1841
rect 1146 1807 1164 1841
rect 1164 1807 1180 1841
rect 1218 1807 1232 1841
rect 1232 1807 1252 1841
rect 1290 1807 1300 1841
rect 1300 1807 1324 1841
rect 1362 1807 1368 1841
rect 1368 1807 1396 1841
rect 1434 1807 1436 1841
rect 1436 1807 1468 1841
rect 1506 1807 1540 1841
rect 466 1759 500 1793
rect 466 1687 500 1721
rect 1114 1730 1148 1764
rect 1186 1730 1220 1764
rect 570 1651 586 1685
rect 586 1651 604 1685
rect 642 1651 654 1685
rect 654 1651 676 1685
rect 714 1651 722 1685
rect 722 1651 748 1685
rect 786 1651 790 1685
rect 790 1651 820 1685
rect 858 1651 892 1685
rect 930 1651 960 1685
rect 960 1651 964 1685
rect 1002 1651 1028 1685
rect 1028 1651 1036 1685
rect 1074 1651 1096 1685
rect 1096 1651 1108 1685
rect 1146 1651 1164 1685
rect 1164 1651 1180 1685
rect 1218 1651 1232 1685
rect 1232 1651 1252 1685
rect 1290 1651 1300 1685
rect 1300 1651 1324 1685
rect 1362 1651 1368 1685
rect 1368 1651 1396 1685
rect 1434 1651 1436 1685
rect 1436 1651 1468 1685
rect 1506 1651 1540 1685
rect 466 1615 500 1649
rect 466 1543 500 1577
rect 1114 1573 1148 1607
rect 1186 1573 1220 1607
rect 2151 1785 2185 1812
rect 2151 1778 2185 1785
rect 2151 1717 2185 1738
rect 2151 1704 2185 1717
rect 2151 1649 2185 1664
rect 2151 1630 2185 1649
rect 4472 1838 4506 1851
rect 4472 1817 4506 1838
rect 4472 1770 4506 1774
rect 4472 1740 4506 1770
rect 4472 1668 4506 1697
rect 4580 2076 4614 2077
rect 4580 2043 4614 2076
rect 7499 2047 7515 2081
rect 7515 2047 7533 2081
rect 7571 2047 7583 2081
rect 7583 2047 7605 2081
rect 7643 2047 7651 2081
rect 7651 2047 7677 2081
rect 7715 2047 7719 2081
rect 7719 2047 7749 2081
rect 7787 2047 7821 2081
rect 7859 2047 7889 2081
rect 7889 2047 7893 2081
rect 7931 2047 7957 2081
rect 7957 2047 7965 2081
rect 8003 2047 8025 2081
rect 8025 2047 8037 2081
rect 8075 2047 8093 2081
rect 8093 2047 8109 2081
rect 8147 2047 8161 2081
rect 8161 2047 8181 2081
rect 8219 2047 8229 2081
rect 8229 2047 8253 2081
rect 8291 2047 8297 2081
rect 8297 2047 8325 2081
rect 8363 2047 8365 2081
rect 8365 2047 8397 2081
rect 8435 2047 8469 2081
rect 4580 1972 4614 1989
rect 4580 1955 4614 1972
rect 6829 1942 6863 1958
rect 6829 1924 6863 1942
rect 4580 1866 4614 1900
rect 4688 1867 4712 1901
rect 4712 1867 4722 1901
rect 4760 1867 4780 1901
rect 4780 1867 4794 1901
rect 4832 1867 4848 1901
rect 4848 1867 4866 1901
rect 4904 1867 4916 1901
rect 4916 1867 4938 1901
rect 4976 1867 4984 1901
rect 4984 1867 5010 1901
rect 5048 1867 5052 1901
rect 5052 1867 5082 1901
rect 5120 1867 5154 1901
rect 5192 1867 5222 1901
rect 5222 1867 5226 1901
rect 5264 1867 5290 1901
rect 5290 1867 5298 1901
rect 5336 1867 5358 1901
rect 5358 1867 5370 1901
rect 5408 1867 5426 1901
rect 5426 1867 5442 1901
rect 5480 1867 5494 1901
rect 5494 1867 5514 1901
rect 5552 1867 5562 1901
rect 5562 1867 5586 1901
rect 5624 1867 5630 1901
rect 5630 1867 5658 1901
rect 5696 1867 5698 1901
rect 5698 1867 5730 1901
rect 5768 1867 5800 1901
rect 5800 1867 5802 1901
rect 5840 1867 5868 1901
rect 5868 1867 5874 1901
rect 5912 1867 5936 1901
rect 5936 1867 5946 1901
rect 5984 1867 6004 1901
rect 6004 1867 6018 1901
rect 6056 1867 6072 1901
rect 6072 1867 6090 1901
rect 6128 1867 6140 1901
rect 6140 1867 6162 1901
rect 6200 1867 6208 1901
rect 6208 1867 6234 1901
rect 6272 1867 6276 1901
rect 6276 1867 6306 1901
rect 6344 1867 6378 1901
rect 6416 1867 6446 1901
rect 6446 1867 6450 1901
rect 6488 1867 6514 1901
rect 6514 1867 6522 1901
rect 6560 1867 6582 1901
rect 6582 1867 6594 1901
rect 6632 1867 6650 1901
rect 6650 1867 6666 1901
rect 6829 1852 6863 1886
rect 8485 1942 8519 1958
rect 8485 1924 8519 1942
rect 8485 1852 8519 1886
rect 9411 1967 9445 1987
rect 9411 1953 9445 1967
rect 9411 1899 9445 1908
rect 9411 1874 9445 1899
rect 6967 1822 7001 1823
rect 7043 1822 7077 1823
rect 7119 1822 7153 1823
rect 7195 1822 7229 1823
rect 7271 1822 7305 1823
rect 7347 1822 7381 1823
rect 7423 1822 7457 1823
rect 7499 1822 7533 1823
rect 7575 1822 7609 1823
rect 7651 1822 7685 1823
rect 7726 1822 7760 1823
rect 7801 1822 7835 1823
rect 7876 1822 7910 1823
rect 7951 1822 7985 1823
rect 8026 1822 8060 1823
rect 8101 1822 8135 1823
rect 8176 1822 8210 1823
rect 8251 1822 8285 1823
rect 8326 1822 8360 1823
rect 8401 1822 8435 1823
rect 4580 1796 4614 1811
rect 4580 1777 4614 1796
rect 6967 1789 6977 1822
rect 6977 1789 7001 1822
rect 7043 1789 7045 1822
rect 7045 1789 7077 1822
rect 7119 1789 7147 1822
rect 7147 1789 7153 1822
rect 7195 1789 7215 1822
rect 7215 1789 7229 1822
rect 7271 1789 7283 1822
rect 7283 1789 7305 1822
rect 7347 1789 7351 1822
rect 7351 1789 7381 1822
rect 7423 1789 7453 1822
rect 7453 1789 7457 1822
rect 7499 1789 7521 1822
rect 7521 1789 7533 1822
rect 7575 1789 7589 1822
rect 7589 1789 7609 1822
rect 7651 1789 7657 1822
rect 7657 1789 7685 1822
rect 7726 1789 7759 1822
rect 7759 1789 7760 1822
rect 7801 1789 7827 1822
rect 7827 1789 7835 1822
rect 7876 1789 7896 1822
rect 7896 1789 7910 1822
rect 7951 1789 7965 1822
rect 7965 1789 7985 1822
rect 8026 1789 8034 1822
rect 8034 1789 8060 1822
rect 8101 1789 8103 1822
rect 8103 1789 8135 1822
rect 8176 1789 8207 1822
rect 8207 1789 8210 1822
rect 8251 1789 8276 1822
rect 8276 1789 8285 1822
rect 8326 1789 8345 1822
rect 8345 1789 8360 1822
rect 8401 1789 8414 1822
rect 8414 1789 8435 1822
rect 9411 1797 9445 1829
rect 9411 1795 9445 1797
rect 4580 1692 4614 1722
rect 4580 1688 4614 1692
rect 6829 1724 6863 1758
rect 2420 1631 2436 1665
rect 2436 1631 2454 1665
rect 2492 1631 2504 1665
rect 2504 1631 2526 1665
rect 2564 1631 2572 1665
rect 2572 1631 2598 1665
rect 2636 1631 2640 1665
rect 2640 1631 2670 1665
rect 2708 1631 2742 1665
rect 2780 1631 2810 1665
rect 2810 1631 2814 1665
rect 2852 1631 2878 1665
rect 2878 1631 2886 1665
rect 2924 1631 2946 1665
rect 2946 1631 2958 1665
rect 2996 1631 3014 1665
rect 3014 1631 3030 1665
rect 3068 1631 3082 1665
rect 3082 1631 3102 1665
rect 3140 1631 3150 1665
rect 3150 1631 3174 1665
rect 3212 1631 3218 1665
rect 3218 1631 3246 1665
rect 3284 1631 3286 1665
rect 3286 1631 3318 1665
rect 3356 1631 3388 1665
rect 3388 1631 3390 1665
rect 3428 1631 3456 1665
rect 3456 1631 3462 1665
rect 3500 1631 3524 1665
rect 3524 1631 3534 1665
rect 3572 1631 3592 1665
rect 3592 1631 3606 1665
rect 3644 1631 3660 1665
rect 3660 1631 3678 1665
rect 3716 1631 3728 1665
rect 3728 1631 3750 1665
rect 3788 1631 3796 1665
rect 3796 1631 3822 1665
rect 3860 1631 3864 1665
rect 3864 1631 3894 1665
rect 3932 1631 3966 1665
rect 4004 1631 4034 1665
rect 4034 1631 4038 1665
rect 4076 1631 4102 1665
rect 4102 1631 4110 1665
rect 4148 1631 4170 1665
rect 4170 1631 4182 1665
rect 4220 1631 4238 1665
rect 4238 1631 4254 1665
rect 4292 1631 4306 1665
rect 4306 1631 4326 1665
rect 4364 1631 4374 1665
rect 4374 1631 4398 1665
rect 4472 1663 4506 1668
rect 6829 1668 6863 1686
rect 2151 1581 2185 1590
rect 2151 1556 2185 1581
rect 466 1471 500 1505
rect 570 1495 586 1529
rect 586 1495 604 1529
rect 642 1495 654 1529
rect 654 1495 676 1529
rect 714 1495 722 1529
rect 722 1495 748 1529
rect 786 1495 790 1529
rect 790 1495 820 1529
rect 858 1495 892 1529
rect 930 1495 960 1529
rect 960 1495 964 1529
rect 1002 1495 1028 1529
rect 1028 1495 1036 1529
rect 1074 1495 1096 1529
rect 1096 1495 1108 1529
rect 1146 1495 1164 1529
rect 1164 1495 1180 1529
rect 1218 1495 1232 1529
rect 1232 1495 1252 1529
rect 1290 1495 1300 1529
rect 1300 1495 1324 1529
rect 1362 1495 1368 1529
rect 1368 1495 1396 1529
rect 1434 1495 1436 1529
rect 1436 1495 1468 1529
rect 1506 1495 1540 1529
rect 466 1399 500 1433
rect 2151 1513 2185 1516
rect 2151 1482 2185 1513
rect 597 1367 598 1401
rect 598 1367 631 1401
rect 675 1367 702 1401
rect 702 1367 709 1401
rect 753 1367 772 1401
rect 772 1367 787 1401
rect 831 1367 842 1401
rect 842 1367 865 1401
rect 909 1367 912 1401
rect 912 1367 943 1401
rect 987 1367 1019 1401
rect 1019 1367 1021 1401
rect 1065 1367 1090 1401
rect 1090 1367 1099 1401
rect 1143 1367 1161 1401
rect 1161 1367 1177 1401
rect 1220 1367 1232 1401
rect 1232 1367 1254 1401
rect 1297 1367 1303 1401
rect 1303 1367 1331 1401
rect 1374 1367 1408 1401
rect 1451 1367 1479 1401
rect 1479 1367 1485 1401
rect 1528 1367 1550 1401
rect 1550 1367 1562 1401
rect 2151 1411 2185 1442
rect 2151 1408 2185 1411
rect 4688 1631 4712 1665
rect 4712 1631 4722 1665
rect 4760 1631 4780 1665
rect 4780 1631 4794 1665
rect 4832 1631 4848 1665
rect 4848 1631 4866 1665
rect 4904 1631 4916 1665
rect 4916 1631 4938 1665
rect 4976 1631 4984 1665
rect 4984 1631 5010 1665
rect 5048 1631 5052 1665
rect 5052 1631 5082 1665
rect 5120 1631 5154 1665
rect 5192 1631 5222 1665
rect 5222 1631 5226 1665
rect 5264 1631 5290 1665
rect 5290 1631 5298 1665
rect 5336 1631 5358 1665
rect 5358 1631 5370 1665
rect 5408 1631 5426 1665
rect 5426 1631 5442 1665
rect 5480 1631 5494 1665
rect 5494 1631 5514 1665
rect 5552 1631 5562 1665
rect 5562 1631 5586 1665
rect 5624 1631 5630 1665
rect 5630 1631 5658 1665
rect 5696 1631 5698 1665
rect 5698 1631 5730 1665
rect 5768 1631 5800 1665
rect 5800 1631 5802 1665
rect 5840 1631 5868 1665
rect 5868 1631 5874 1665
rect 5912 1631 5936 1665
rect 5936 1631 5946 1665
rect 5984 1631 6004 1665
rect 6004 1631 6018 1665
rect 6056 1631 6072 1665
rect 6072 1631 6090 1665
rect 6128 1631 6140 1665
rect 6140 1631 6162 1665
rect 6200 1631 6208 1665
rect 6208 1631 6234 1665
rect 6272 1631 6276 1665
rect 6276 1631 6306 1665
rect 6344 1631 6378 1665
rect 6416 1631 6446 1665
rect 6446 1631 6450 1665
rect 6488 1631 6514 1665
rect 6514 1631 6522 1665
rect 6560 1631 6582 1665
rect 6582 1631 6594 1665
rect 6632 1631 6650 1665
rect 6650 1631 6666 1665
rect 6829 1652 6863 1668
rect 8485 1724 8519 1758
rect 8485 1668 8519 1686
rect 8485 1652 8519 1668
rect 9411 1729 9445 1750
rect 9411 1716 9445 1729
rect 9411 1661 9445 1671
rect 9411 1637 9445 1661
rect 4472 1599 4506 1619
rect 4472 1585 4506 1599
rect 4472 1530 4506 1541
rect 4472 1507 4506 1530
rect 12253 2815 12287 2821
rect 12325 2815 12359 2821
rect 12397 2815 12431 2821
rect 12469 2815 12503 2821
rect 12542 2815 12576 2821
rect 12615 2815 12649 2821
rect 12688 2815 12722 2821
rect 12761 2815 12795 2821
rect 12834 2815 12868 2821
rect 12907 2815 12941 2821
rect 12980 2815 13014 2821
rect 13053 2815 13087 2821
rect 13126 2815 13160 2821
rect 13199 2815 13233 2821
rect 13272 2815 13306 2821
rect 13345 2815 13379 2821
rect 13418 2815 13452 2821
rect 13491 2815 13525 2821
rect 13564 2815 13598 2821
rect 13637 2815 13671 2821
rect 13710 2815 13744 2821
rect 13783 2815 13817 2821
rect 13856 2815 13890 2821
rect 13929 2815 13963 2821
rect 14002 2815 14036 2821
rect 14075 2815 14109 2821
rect 14148 2815 14182 2821
rect 14221 2815 14255 2821
rect 14294 2815 14328 2821
rect 14367 2815 14401 2821
rect 14440 2815 14474 2821
rect 14513 2815 14547 2821
rect 14586 2815 14620 2821
rect 14659 2815 14693 2821
rect 14732 2815 14766 2821
rect 14805 2815 14839 2821
rect 14878 2815 14912 2821
rect 14951 2815 14985 2821
rect 15024 2815 15058 2821
rect 15097 2815 15131 2821
rect 15170 2815 15204 2821
rect 15243 2815 15277 2821
rect 15316 2815 15350 2821
rect 15389 2815 15423 2821
rect 15462 2815 15496 2821
rect 15535 2815 15569 2821
rect 15608 2815 15642 2821
rect 15681 2815 15715 2821
rect 15754 2815 15788 2821
rect 15827 2815 15861 2821
rect 15900 2815 15934 2849
rect 15973 2821 16002 2849
rect 16002 2821 16007 2849
rect 16046 2821 16070 2849
rect 16070 2821 16080 2849
rect 16119 2821 16138 2849
rect 16138 2821 16153 2849
rect 16192 2821 16206 2849
rect 16206 2821 16226 2849
rect 16265 2821 16274 2849
rect 16274 2821 16299 2849
rect 16338 2821 16342 2849
rect 16342 2821 16372 2849
rect 18417 2849 18428 2883
rect 18428 2849 18451 2883
rect 18497 2849 18530 2883
rect 18530 2849 18531 2883
rect 18577 2849 18598 2883
rect 18598 2849 18611 2883
rect 18657 2849 18666 2883
rect 18666 2849 18691 2883
rect 18737 2849 18768 2883
rect 18768 2849 18771 2883
rect 18817 2849 18836 2883
rect 18836 2849 18851 2883
rect 18897 2849 18904 2883
rect 18904 2849 18931 2883
rect 18977 2849 19006 2883
rect 19006 2849 19011 2883
rect 19056 2849 19074 2883
rect 19074 2849 19090 2883
rect 15973 2815 16007 2821
rect 16046 2815 16080 2821
rect 16119 2815 16153 2821
rect 16192 2815 16226 2821
rect 16265 2815 16299 2821
rect 16338 2815 16372 2821
rect 20002 2820 20036 2854
rect 16410 2742 16444 2776
rect 17935 2768 17966 2778
rect 17966 2768 17969 2778
rect 18007 2768 18034 2778
rect 18034 2768 18041 2778
rect 17935 2744 17969 2768
rect 18007 2744 18041 2768
rect 20002 2748 20036 2782
rect 10613 2584 10647 2618
rect 10685 2584 10719 2618
rect 16410 2693 16444 2703
rect 16410 2669 16444 2693
rect 16410 2625 16444 2630
rect 16410 2596 16444 2625
rect 16410 2523 16444 2557
rect 16410 2455 16444 2484
rect 16410 2450 16444 2455
rect 16410 2387 16444 2411
rect 16410 2377 16444 2387
rect 16410 2319 16444 2338
rect 16410 2304 16444 2319
rect 16410 2251 16444 2265
rect 16410 2231 16444 2251
rect 10613 2188 10647 2213
rect 10613 2179 10634 2188
rect 10634 2179 10647 2188
rect 10685 2179 10719 2213
rect 16410 2183 16444 2192
rect 16410 2158 16444 2183
rect 16410 2115 16444 2119
rect 16410 2085 16444 2115
rect 10500 2013 10534 2047
rect 10573 2013 10590 2047
rect 10590 2013 10607 2047
rect 10646 2013 10658 2047
rect 10658 2013 10680 2047
rect 10719 2013 10726 2047
rect 10726 2013 10753 2047
rect 10792 2013 10794 2047
rect 10794 2013 10826 2047
rect 10865 2013 10896 2047
rect 10896 2013 10899 2047
rect 10938 2013 10964 2047
rect 10964 2013 10972 2047
rect 11010 2013 11032 2047
rect 11032 2013 11044 2047
rect 11082 2013 11100 2047
rect 11100 2013 11116 2047
rect 11154 2013 11168 2047
rect 11168 2013 11188 2047
rect 11226 2013 11236 2047
rect 11236 2013 11260 2047
rect 11298 2013 11304 2047
rect 11304 2013 11332 2047
rect 11370 2013 11372 2047
rect 11372 2013 11404 2047
rect 11442 2013 11474 2047
rect 11474 2013 11476 2047
rect 11514 2013 11542 2047
rect 11542 2013 11548 2047
rect 11586 2013 11610 2047
rect 11610 2013 11620 2047
rect 11658 2013 11678 2047
rect 11678 2013 11692 2047
rect 11730 2013 11746 2047
rect 11746 2013 11764 2047
rect 11802 2013 11814 2047
rect 11814 2013 11836 2047
rect 11874 2013 11882 2047
rect 11882 2013 11908 2047
rect 11946 2013 11950 2047
rect 11950 2013 11980 2047
rect 12018 2013 12052 2047
rect 12090 2013 12120 2047
rect 12120 2013 12124 2047
rect 12162 2013 12188 2047
rect 12188 2013 12196 2047
rect 12234 2013 12256 2047
rect 12256 2013 12268 2047
rect 12306 2013 12324 2047
rect 12324 2013 12340 2047
rect 12378 2013 12392 2047
rect 12392 2013 12412 2047
rect 12450 2013 12460 2047
rect 12460 2013 12484 2047
rect 12522 2013 12528 2047
rect 12528 2013 12556 2047
rect 12594 2013 12596 2047
rect 12596 2013 12628 2047
rect 12666 2013 12698 2047
rect 12698 2013 12700 2047
rect 12738 2013 12766 2047
rect 12766 2013 12772 2047
rect 12810 2013 12834 2047
rect 12834 2013 12844 2047
rect 12882 2013 12902 2047
rect 12902 2013 12916 2047
rect 12954 2013 12970 2047
rect 12970 2013 12988 2047
rect 13026 2013 13038 2047
rect 13038 2013 13060 2047
rect 13098 2013 13106 2047
rect 13106 2013 13132 2047
rect 13170 2013 13174 2047
rect 13174 2013 13204 2047
rect 13242 2013 13276 2047
rect 13314 2013 13344 2047
rect 13344 2013 13348 2047
rect 13386 2013 13412 2047
rect 13412 2013 13420 2047
rect 13458 2013 13480 2047
rect 13480 2013 13492 2047
rect 13530 2013 13548 2047
rect 13548 2013 13564 2047
rect 13602 2013 13616 2047
rect 13616 2013 13636 2047
rect 13674 2013 13684 2047
rect 13684 2013 13708 2047
rect 13746 2013 13752 2047
rect 13752 2013 13780 2047
rect 13818 2013 13820 2047
rect 13820 2013 13852 2047
rect 13890 2013 13922 2047
rect 13922 2013 13924 2047
rect 13962 2013 13990 2047
rect 13990 2013 13996 2047
rect 14034 2013 14058 2047
rect 14058 2013 14068 2047
rect 14106 2013 14126 2047
rect 14126 2013 14140 2047
rect 14178 2013 14194 2047
rect 14194 2013 14212 2047
rect 14250 2013 14262 2047
rect 14262 2013 14284 2047
rect 14322 2013 14330 2047
rect 14330 2013 14356 2047
rect 14394 2013 14398 2047
rect 14398 2013 14428 2047
rect 14466 2013 14500 2047
rect 14538 2013 14568 2047
rect 14568 2013 14572 2047
rect 14610 2013 14636 2047
rect 14636 2013 14644 2047
rect 14682 2013 14704 2047
rect 14704 2013 14716 2047
rect 14754 2013 14772 2047
rect 14772 2013 14788 2047
rect 14826 2013 14840 2047
rect 14840 2013 14860 2047
rect 14898 2013 14908 2047
rect 14908 2013 14932 2047
rect 14970 2013 14976 2047
rect 14976 2013 15004 2047
rect 15042 2013 15044 2047
rect 15044 2013 15076 2047
rect 15114 2013 15146 2047
rect 15146 2013 15148 2047
rect 15186 2013 15214 2047
rect 15214 2013 15220 2047
rect 15258 2013 15282 2047
rect 15282 2013 15292 2047
rect 15330 2013 15350 2047
rect 15350 2013 15364 2047
rect 15402 2013 15418 2047
rect 15418 2013 15436 2047
rect 15474 2013 15486 2047
rect 15486 2013 15508 2047
rect 15546 2013 15554 2047
rect 15554 2013 15580 2047
rect 15618 2013 15622 2047
rect 15622 2013 15652 2047
rect 15690 2013 15724 2047
rect 15762 2013 15792 2047
rect 15792 2013 15796 2047
rect 15834 2013 15860 2047
rect 15860 2013 15868 2047
rect 15906 2013 15928 2047
rect 15928 2013 15940 2047
rect 15978 2013 15996 2047
rect 15996 2013 16012 2047
rect 16050 2013 16064 2047
rect 16064 2013 16084 2047
rect 16122 2013 16132 2047
rect 16132 2013 16156 2047
rect 16194 2013 16200 2047
rect 16200 2013 16228 2047
rect 16266 2013 16268 2047
rect 16268 2013 16300 2047
rect 16338 2013 16370 2047
rect 16370 2013 16372 2047
rect 18430 2693 18462 2727
rect 18462 2693 18464 2727
rect 18509 2693 18530 2727
rect 18530 2693 18543 2727
rect 18588 2693 18598 2727
rect 18598 2693 18622 2727
rect 18666 2693 18700 2727
rect 18744 2693 18768 2727
rect 18768 2693 18778 2727
rect 18822 2693 18836 2727
rect 18836 2693 18856 2727
rect 18900 2693 18904 2727
rect 18904 2693 18934 2727
rect 18978 2693 19006 2727
rect 19006 2693 19012 2727
rect 19056 2693 19074 2727
rect 19074 2693 19090 2727
rect 20002 2676 20036 2710
rect 16601 2545 16635 2579
rect 16675 2545 16709 2579
rect 16749 2545 16783 2579
rect 16823 2545 16857 2579
rect 16897 2545 16931 2579
rect 16971 2545 17005 2579
rect 17045 2545 17079 2579
rect 17119 2545 17153 2579
rect 17192 2545 17226 2579
rect 17805 2572 17817 2606
rect 17817 2572 17839 2606
rect 17878 2572 17889 2606
rect 17889 2572 17912 2606
rect 17951 2572 17961 2606
rect 17961 2572 17985 2606
rect 18024 2572 18033 2606
rect 18033 2572 18058 2606
rect 18097 2572 18105 2606
rect 18105 2572 18131 2606
rect 18170 2572 18176 2606
rect 18176 2572 18204 2606
rect 18243 2572 18247 2606
rect 18247 2572 18277 2606
rect 18316 2572 18318 2606
rect 18318 2572 18350 2606
rect 18389 2572 18423 2606
rect 18462 2572 18494 2606
rect 18494 2572 18496 2606
rect 18535 2572 18565 2606
rect 18565 2572 18569 2606
rect 18608 2572 18636 2606
rect 18636 2572 18642 2606
rect 18680 2572 18707 2606
rect 18707 2572 18714 2606
rect 18752 2572 18778 2606
rect 18778 2572 18786 2606
rect 18824 2572 18849 2606
rect 18849 2572 18858 2606
rect 18896 2572 18920 2606
rect 18920 2572 18930 2606
rect 18968 2572 18991 2606
rect 18991 2572 19002 2606
rect 19040 2572 19062 2606
rect 19062 2572 19074 2606
rect 20002 2604 20036 2638
rect 16601 2473 16635 2507
rect 16675 2473 16709 2507
rect 16749 2473 16783 2507
rect 16823 2473 16857 2507
rect 16897 2473 16931 2507
rect 16971 2473 17005 2507
rect 17045 2473 17079 2507
rect 17119 2473 17153 2507
rect 17192 2473 17226 2507
rect 16601 2401 16635 2435
rect 16675 2401 16709 2435
rect 16749 2401 16783 2435
rect 16823 2401 16857 2435
rect 16897 2401 16931 2435
rect 16971 2401 17005 2435
rect 17045 2401 17079 2435
rect 17119 2401 17153 2435
rect 17192 2401 17226 2435
rect 20002 2532 20036 2566
rect 20002 2460 20036 2494
rect 16590 2329 16624 2363
rect 16662 2329 16696 2363
rect 16734 2329 16768 2363
rect 16806 2329 16840 2363
rect 20002 2388 20036 2422
rect 20002 2316 20036 2350
rect 16590 2242 16624 2276
rect 16662 2242 16696 2276
rect 16734 2242 16768 2276
rect 16806 2242 16840 2276
rect 16590 2154 16624 2188
rect 16662 2154 16696 2188
rect 16734 2154 16768 2188
rect 16806 2154 16840 2188
rect 16590 2070 16624 2100
rect 16662 2070 16696 2100
rect 16734 2070 16768 2100
rect 16806 2070 16840 2100
rect 16590 2066 16624 2070
rect 16662 2066 16696 2070
rect 16734 2066 16768 2070
rect 16806 2066 16840 2070
rect 16590 2001 16597 2012
rect 16597 2001 16624 2012
rect 16662 2001 16665 2012
rect 16665 2001 16696 2012
rect 16734 2001 16767 2012
rect 16767 2001 16768 2012
rect 16806 2001 16835 2012
rect 16835 2001 16840 2012
rect 16590 1978 16624 2001
rect 16662 1978 16696 2001
rect 16734 1978 16768 2001
rect 16806 1978 16840 2001
rect 9734 1898 9768 1918
rect 9808 1898 9842 1918
rect 9882 1898 9916 1918
rect 9956 1898 9990 1918
rect 10030 1898 10064 1918
rect 10104 1898 10138 1918
rect 10178 1898 10212 1918
rect 10252 1898 10286 1918
rect 10326 1898 10360 1918
rect 10400 1898 10434 1918
rect 10473 1898 10507 1918
rect 10546 1898 10580 1918
rect 10619 1898 10653 1918
rect 10692 1898 10726 1918
rect 10765 1898 10799 1918
rect 10838 1898 10872 1918
rect 10911 1898 10945 1918
rect 10984 1898 11018 1918
rect 11057 1898 11091 1918
rect 11130 1898 11164 1918
rect 11203 1898 11237 1918
rect 11276 1898 11310 1918
rect 11349 1898 11383 1918
rect 11422 1898 11456 1918
rect 11495 1898 11529 1918
rect 11568 1898 11602 1918
rect 11641 1898 11675 1918
rect 11714 1898 11748 1918
rect 11787 1898 11821 1918
rect 11860 1898 11894 1918
rect 11933 1898 11967 1918
rect 12006 1898 12040 1918
rect 12079 1898 12113 1918
rect 12152 1898 12186 1918
rect 12225 1898 12259 1918
rect 12298 1898 12332 1918
rect 12371 1898 12405 1918
rect 20002 2244 20036 2278
rect 20002 2172 20036 2206
rect 20002 2100 20036 2134
rect 20002 2028 20036 2062
rect 24045 1991 24079 2025
rect 24121 1991 24155 2025
rect 24197 1991 24231 2025
rect 24273 1991 24307 2025
rect 24349 1991 24383 2025
rect 24424 1991 24458 2025
rect 24499 1991 24533 2025
rect 24574 1991 24608 2025
rect 24649 1991 24683 2025
rect 20002 1956 20036 1990
rect 12756 1898 12790 1911
rect 12830 1898 12864 1911
rect 12904 1898 12938 1911
rect 12978 1898 13012 1911
rect 13052 1898 13086 1911
rect 13126 1898 13160 1911
rect 13200 1898 13234 1911
rect 13274 1898 13308 1911
rect 13348 1898 13382 1911
rect 13422 1898 13456 1911
rect 13496 1898 13530 1911
rect 13569 1898 13603 1911
rect 13642 1898 13676 1911
rect 13715 1898 13749 1911
rect 13788 1898 13822 1911
rect 13861 1898 13895 1911
rect 13934 1898 13968 1911
rect 14007 1898 14041 1911
rect 14080 1898 14114 1911
rect 14153 1898 14187 1911
rect 14226 1898 14260 1911
rect 14299 1898 14333 1911
rect 14372 1898 14406 1911
rect 14445 1898 14479 1911
rect 14518 1898 14552 1911
rect 14591 1898 14625 1911
rect 14664 1898 14698 1911
rect 14737 1898 14771 1911
rect 14810 1898 14844 1911
rect 14883 1898 14917 1911
rect 14956 1898 14990 1911
rect 15029 1898 15063 1911
rect 15102 1898 15136 1911
rect 15175 1898 15209 1911
rect 15248 1898 15282 1911
rect 15321 1898 15355 1911
rect 15394 1898 15428 1911
rect 15467 1898 15501 1911
rect 15540 1898 15574 1911
rect 15613 1898 15647 1911
rect 15686 1898 15720 1911
rect 15759 1898 15793 1911
rect 15832 1898 15866 1911
rect 15905 1898 15939 1911
rect 15978 1898 16012 1911
rect 16051 1898 16085 1911
rect 16124 1898 16158 1911
rect 16197 1898 16231 1911
rect 16270 1898 16304 1911
rect 16343 1898 16377 1911
rect 16416 1898 16450 1911
rect 16489 1898 16523 1911
rect 16562 1898 16563 1911
rect 16563 1898 16596 1911
rect 9734 1884 9750 1898
rect 9750 1884 9768 1898
rect 9808 1884 9819 1898
rect 9819 1884 9842 1898
rect 9882 1884 9888 1898
rect 9888 1884 9916 1898
rect 9956 1884 9957 1898
rect 9957 1884 9990 1898
rect 10030 1884 10060 1898
rect 10060 1884 10064 1898
rect 10104 1884 10129 1898
rect 10129 1884 10138 1898
rect 10178 1884 10198 1898
rect 10198 1884 10212 1898
rect 10252 1884 10267 1898
rect 10267 1884 10286 1898
rect 10326 1884 10336 1898
rect 10336 1884 10360 1898
rect 10400 1884 10405 1898
rect 10405 1884 10434 1898
rect 10473 1884 10474 1898
rect 10474 1884 10507 1898
rect 10546 1884 10578 1898
rect 10578 1884 10580 1898
rect 10619 1884 10647 1898
rect 10647 1884 10653 1898
rect 10692 1884 10716 1898
rect 10716 1884 10726 1898
rect 10765 1884 10785 1898
rect 10785 1884 10799 1898
rect 10838 1884 10854 1898
rect 10854 1884 10872 1898
rect 10911 1884 10923 1898
rect 10923 1884 10945 1898
rect 10984 1884 10992 1898
rect 10992 1884 11018 1898
rect 11057 1884 11061 1898
rect 11061 1884 11091 1898
rect 11130 1884 11164 1898
rect 11203 1884 11233 1898
rect 11233 1884 11237 1898
rect 11276 1884 11302 1898
rect 11302 1884 11310 1898
rect 11349 1884 11371 1898
rect 11371 1884 11383 1898
rect 11422 1884 11440 1898
rect 11440 1884 11456 1898
rect 11495 1884 11509 1898
rect 11509 1884 11529 1898
rect 11568 1884 11578 1898
rect 11578 1884 11602 1898
rect 11641 1884 11647 1898
rect 11647 1884 11675 1898
rect 11714 1884 11716 1898
rect 11716 1884 11748 1898
rect 11787 1884 11820 1898
rect 11820 1884 11821 1898
rect 11860 1884 11889 1898
rect 11889 1884 11894 1898
rect 11933 1884 11958 1898
rect 11958 1884 11967 1898
rect 12006 1884 12027 1898
rect 12027 1884 12040 1898
rect 12079 1884 12096 1898
rect 12096 1884 12113 1898
rect 12152 1884 12165 1898
rect 12165 1884 12186 1898
rect 12225 1884 12234 1898
rect 12234 1884 12259 1898
rect 12298 1884 12303 1898
rect 12303 1884 12332 1898
rect 12371 1884 12372 1898
rect 12372 1884 12405 1898
rect 12756 1877 12786 1898
rect 12786 1877 12790 1898
rect 12830 1877 12855 1898
rect 12855 1877 12864 1898
rect 12904 1877 12924 1898
rect 12924 1877 12938 1898
rect 12978 1877 12993 1898
rect 12993 1877 13012 1898
rect 13052 1877 13086 1898
rect 13126 1877 13160 1898
rect 13200 1877 13234 1898
rect 13274 1877 13308 1898
rect 13348 1877 13382 1898
rect 13422 1877 13456 1898
rect 13496 1877 13530 1898
rect 13569 1877 13603 1898
rect 13642 1877 13676 1898
rect 13715 1877 13749 1898
rect 13788 1877 13822 1898
rect 13861 1877 13895 1898
rect 13934 1877 13968 1898
rect 14007 1877 14041 1898
rect 14080 1877 14114 1898
rect 14153 1877 14187 1898
rect 14226 1877 14260 1898
rect 14299 1877 14333 1898
rect 14372 1877 14406 1898
rect 14445 1877 14479 1898
rect 14518 1877 14552 1898
rect 14591 1877 14625 1898
rect 14664 1877 14698 1898
rect 14737 1877 14771 1898
rect 14810 1877 14844 1898
rect 14883 1877 14917 1898
rect 14956 1877 14990 1898
rect 15029 1877 15063 1898
rect 15102 1877 15136 1898
rect 15175 1877 15209 1898
rect 15248 1877 15282 1898
rect 15321 1877 15355 1898
rect 15394 1877 15428 1898
rect 15467 1877 15501 1898
rect 15540 1877 15574 1898
rect 15613 1877 15647 1898
rect 15686 1877 15720 1898
rect 15759 1877 15793 1898
rect 15832 1877 15866 1898
rect 15905 1877 15939 1898
rect 15978 1877 16012 1898
rect 16051 1877 16085 1898
rect 16124 1877 16158 1898
rect 16197 1877 16231 1898
rect 16270 1877 16304 1898
rect 16343 1877 16377 1898
rect 16416 1877 16450 1898
rect 16489 1877 16523 1898
rect 16562 1877 16596 1898
rect 16635 1877 16669 1911
rect 16708 1877 16742 1911
rect 16847 1868 16881 1902
rect 16919 1868 16953 1902
rect 16991 1868 17025 1902
rect 17063 1868 17097 1902
rect 17135 1868 17169 1902
rect 17207 1868 17241 1902
rect 17279 1868 17313 1902
rect 17351 1868 17385 1902
rect 17423 1868 17457 1902
rect 17495 1868 17529 1902
rect 17567 1868 17601 1902
rect 17639 1868 17673 1902
rect 17711 1868 17745 1902
rect 17783 1868 17817 1902
rect 17855 1868 17889 1902
rect 17927 1868 17961 1902
rect 17999 1868 18033 1902
rect 18071 1868 18105 1902
rect 18143 1868 18177 1902
rect 18215 1868 18249 1902
rect 18287 1868 18321 1902
rect 18359 1868 18393 1902
rect 18431 1868 18465 1902
rect 18503 1868 18537 1902
rect 18575 1868 18609 1902
rect 18647 1868 18681 1902
rect 18719 1868 18753 1902
rect 18791 1868 18825 1902
rect 18863 1868 18897 1902
rect 18935 1868 18969 1902
rect 19007 1868 19011 1902
rect 19011 1868 19041 1902
rect 19079 1889 19113 1902
rect 19079 1868 19113 1889
rect 19151 1889 19152 1902
rect 19152 1889 19185 1902
rect 19151 1868 19185 1889
rect 9734 1830 9768 1836
rect 9808 1830 9842 1836
rect 9882 1830 9916 1836
rect 9956 1830 9990 1836
rect 10030 1830 10064 1836
rect 10104 1830 10138 1836
rect 10178 1830 10212 1836
rect 10252 1830 10286 1836
rect 10326 1830 10360 1836
rect 10400 1830 10434 1836
rect 10473 1830 10507 1836
rect 10546 1830 10580 1836
rect 10619 1830 10653 1836
rect 10692 1830 10726 1836
rect 10765 1830 10799 1836
rect 10838 1830 10872 1836
rect 10911 1830 10945 1836
rect 10984 1830 11018 1836
rect 11057 1830 11091 1836
rect 11130 1830 11164 1836
rect 11203 1830 11237 1836
rect 11276 1830 11310 1836
rect 11349 1830 11383 1836
rect 11422 1830 11456 1836
rect 11495 1830 11529 1836
rect 11568 1830 11602 1836
rect 11641 1830 11675 1836
rect 11714 1830 11748 1836
rect 11787 1830 11821 1836
rect 11860 1830 11894 1836
rect 11933 1830 11967 1836
rect 12006 1830 12040 1836
rect 12079 1830 12113 1836
rect 12152 1830 12186 1836
rect 12225 1830 12259 1836
rect 12298 1830 12332 1836
rect 12371 1830 12405 1836
rect 9734 1802 9750 1830
rect 9750 1802 9768 1830
rect 9808 1802 9819 1830
rect 9819 1802 9842 1830
rect 9882 1802 9888 1830
rect 9888 1802 9916 1830
rect 9956 1802 9957 1830
rect 9957 1802 9990 1830
rect 10030 1802 10060 1830
rect 10060 1802 10064 1830
rect 10104 1802 10129 1830
rect 10129 1802 10138 1830
rect 10178 1802 10198 1830
rect 10198 1802 10212 1830
rect 10252 1802 10267 1830
rect 10267 1802 10286 1830
rect 10326 1802 10336 1830
rect 10336 1802 10360 1830
rect 10400 1802 10405 1830
rect 10405 1802 10434 1830
rect 10473 1802 10474 1830
rect 10474 1802 10507 1830
rect 10546 1802 10578 1830
rect 10578 1802 10580 1830
rect 10619 1802 10647 1830
rect 10647 1802 10653 1830
rect 10692 1802 10716 1830
rect 10716 1802 10726 1830
rect 10765 1802 10785 1830
rect 10785 1802 10799 1830
rect 10838 1802 10854 1830
rect 10854 1802 10872 1830
rect 10911 1802 10923 1830
rect 10923 1802 10945 1830
rect 10984 1802 10992 1830
rect 10992 1802 11018 1830
rect 11057 1802 11061 1830
rect 11061 1802 11091 1830
rect 11130 1802 11164 1830
rect 11203 1802 11233 1830
rect 11233 1802 11237 1830
rect 11276 1802 11302 1830
rect 11302 1802 11310 1830
rect 11349 1802 11371 1830
rect 11371 1802 11383 1830
rect 11422 1802 11440 1830
rect 11440 1802 11456 1830
rect 11495 1802 11509 1830
rect 11509 1802 11529 1830
rect 11568 1802 11578 1830
rect 11578 1802 11602 1830
rect 11641 1802 11647 1830
rect 11647 1802 11675 1830
rect 11714 1802 11716 1830
rect 11716 1802 11748 1830
rect 11787 1802 11820 1830
rect 11820 1802 11821 1830
rect 11860 1802 11889 1830
rect 11889 1802 11894 1830
rect 11933 1802 11958 1830
rect 11958 1802 11967 1830
rect 12006 1802 12027 1830
rect 12027 1802 12040 1830
rect 12079 1802 12096 1830
rect 12096 1802 12113 1830
rect 12152 1802 12165 1830
rect 12165 1802 12186 1830
rect 12225 1802 12234 1830
rect 12234 1802 12259 1830
rect 12298 1802 12303 1830
rect 12303 1802 12332 1830
rect 12371 1802 12372 1830
rect 12372 1802 12405 1830
rect 16847 1782 16881 1816
rect 16919 1782 16953 1816
rect 16991 1782 17025 1816
rect 17063 1782 17097 1816
rect 17135 1782 17169 1816
rect 17207 1782 17241 1816
rect 17279 1782 17313 1816
rect 17351 1782 17385 1816
rect 17423 1782 17457 1816
rect 17495 1782 17529 1816
rect 17567 1782 17601 1816
rect 17639 1782 17673 1816
rect 17711 1782 17745 1816
rect 17783 1782 17817 1816
rect 17855 1782 17889 1816
rect 17927 1782 17961 1816
rect 17999 1782 18033 1816
rect 18071 1782 18105 1816
rect 18143 1782 18177 1816
rect 18215 1782 18249 1816
rect 18287 1782 18321 1816
rect 18359 1782 18393 1816
rect 18431 1782 18465 1816
rect 18503 1782 18537 1816
rect 18575 1782 18609 1816
rect 18647 1782 18681 1816
rect 18719 1782 18753 1816
rect 18791 1782 18825 1816
rect 18863 1782 18897 1816
rect 18935 1782 18969 1816
rect 19007 1782 19011 1816
rect 19011 1782 19041 1816
rect 19079 1815 19113 1816
rect 19079 1782 19113 1815
rect 19151 1815 19152 1816
rect 19152 1815 19185 1816
rect 19151 1782 19185 1815
rect 9734 1728 9750 1754
rect 9750 1728 9768 1754
rect 9808 1728 9819 1754
rect 9819 1728 9842 1754
rect 9882 1728 9888 1754
rect 9888 1728 9916 1754
rect 9956 1728 9957 1754
rect 9957 1728 9990 1754
rect 10030 1728 10060 1754
rect 10060 1728 10064 1754
rect 10104 1728 10129 1754
rect 10129 1728 10138 1754
rect 10178 1728 10198 1754
rect 10198 1728 10212 1754
rect 10252 1728 10267 1754
rect 10267 1728 10286 1754
rect 10326 1728 10336 1754
rect 10336 1728 10360 1754
rect 10400 1728 10405 1754
rect 10405 1728 10434 1754
rect 10473 1728 10474 1754
rect 10474 1728 10507 1754
rect 10546 1728 10578 1754
rect 10578 1728 10580 1754
rect 10619 1728 10647 1754
rect 10647 1728 10653 1754
rect 10692 1728 10716 1754
rect 10716 1728 10726 1754
rect 10765 1728 10785 1754
rect 10785 1728 10799 1754
rect 10838 1728 10854 1754
rect 10854 1728 10872 1754
rect 10911 1728 10923 1754
rect 10923 1728 10945 1754
rect 10984 1728 10992 1754
rect 10992 1728 11018 1754
rect 11057 1728 11061 1754
rect 11061 1728 11091 1754
rect 11130 1728 11164 1754
rect 11203 1728 11233 1754
rect 11233 1728 11237 1754
rect 11276 1728 11302 1754
rect 11302 1728 11310 1754
rect 11349 1728 11371 1754
rect 11371 1728 11383 1754
rect 11422 1728 11440 1754
rect 11440 1728 11456 1754
rect 11495 1728 11509 1754
rect 11509 1728 11529 1754
rect 11568 1728 11578 1754
rect 11578 1728 11602 1754
rect 11641 1728 11647 1754
rect 11647 1728 11675 1754
rect 11714 1728 11716 1754
rect 11716 1728 11748 1754
rect 11787 1728 11820 1754
rect 11820 1728 11821 1754
rect 11860 1728 11889 1754
rect 11889 1728 11894 1754
rect 11933 1728 11958 1754
rect 11958 1728 11967 1754
rect 12006 1728 12027 1754
rect 12027 1728 12040 1754
rect 12079 1728 12096 1754
rect 12096 1728 12113 1754
rect 12152 1728 12165 1754
rect 12165 1728 12186 1754
rect 12225 1728 12234 1754
rect 12234 1728 12259 1754
rect 12298 1728 12303 1754
rect 12303 1728 12332 1754
rect 12371 1728 12372 1754
rect 12372 1728 12405 1754
rect 9734 1720 9768 1728
rect 9808 1720 9842 1728
rect 9882 1720 9916 1728
rect 9956 1720 9990 1728
rect 10030 1720 10064 1728
rect 10104 1720 10138 1728
rect 10178 1720 10212 1728
rect 10252 1720 10286 1728
rect 10326 1720 10360 1728
rect 10400 1720 10434 1728
rect 10473 1720 10507 1728
rect 10546 1720 10580 1728
rect 10619 1720 10653 1728
rect 10692 1720 10726 1728
rect 10765 1720 10799 1728
rect 10838 1720 10872 1728
rect 10911 1720 10945 1728
rect 10984 1720 11018 1728
rect 11057 1720 11091 1728
rect 11130 1720 11164 1728
rect 11203 1720 11237 1728
rect 11276 1720 11310 1728
rect 11349 1720 11383 1728
rect 11422 1720 11456 1728
rect 11495 1720 11529 1728
rect 11568 1720 11602 1728
rect 11641 1720 11675 1728
rect 11714 1720 11748 1728
rect 11787 1720 11821 1728
rect 11860 1720 11894 1728
rect 11933 1720 11967 1728
rect 12006 1720 12040 1728
rect 12079 1720 12113 1728
rect 12152 1720 12186 1728
rect 12225 1720 12259 1728
rect 12298 1720 12332 1728
rect 12371 1720 12405 1728
rect 16847 1696 16881 1730
rect 16919 1696 16953 1730
rect 16991 1696 17025 1730
rect 17063 1696 17097 1730
rect 17135 1696 17169 1730
rect 17207 1696 17241 1730
rect 17279 1696 17313 1730
rect 17351 1696 17385 1730
rect 17423 1696 17457 1730
rect 17495 1696 17529 1730
rect 17567 1696 17601 1730
rect 17639 1696 17673 1730
rect 17711 1696 17745 1730
rect 17783 1696 17817 1730
rect 17855 1696 17889 1730
rect 17927 1696 17961 1730
rect 17999 1696 18033 1730
rect 18071 1696 18105 1730
rect 18143 1696 18177 1730
rect 18215 1696 18249 1730
rect 18287 1696 18321 1730
rect 18359 1696 18393 1730
rect 18431 1696 18465 1730
rect 18503 1696 18537 1730
rect 18575 1696 18609 1730
rect 18647 1696 18681 1730
rect 18719 1696 18753 1730
rect 18791 1696 18825 1730
rect 18863 1696 18897 1730
rect 18935 1696 18969 1730
rect 19007 1696 19011 1730
rect 19011 1696 19041 1730
rect 19079 1701 19113 1730
rect 19079 1696 19113 1701
rect 19151 1701 19185 1730
rect 19151 1696 19152 1701
rect 19152 1696 19185 1701
rect 9734 1660 9750 1672
rect 9750 1660 9768 1672
rect 9808 1660 9819 1672
rect 9819 1660 9842 1672
rect 9882 1660 9888 1672
rect 9888 1660 9916 1672
rect 9956 1660 9957 1672
rect 9957 1660 9990 1672
rect 10030 1660 10060 1672
rect 10060 1660 10064 1672
rect 10104 1660 10129 1672
rect 10129 1660 10138 1672
rect 10178 1660 10198 1672
rect 10198 1660 10212 1672
rect 10252 1660 10267 1672
rect 10267 1660 10286 1672
rect 10326 1660 10336 1672
rect 10336 1660 10360 1672
rect 10400 1660 10405 1672
rect 10405 1660 10434 1672
rect 10473 1660 10474 1672
rect 10474 1660 10507 1672
rect 10546 1660 10578 1672
rect 10578 1660 10580 1672
rect 10619 1660 10647 1672
rect 10647 1660 10653 1672
rect 10692 1660 10716 1672
rect 10716 1660 10726 1672
rect 10765 1660 10785 1672
rect 10785 1660 10799 1672
rect 10838 1660 10854 1672
rect 10854 1660 10872 1672
rect 10911 1660 10923 1672
rect 10923 1660 10945 1672
rect 10984 1660 10992 1672
rect 10992 1660 11018 1672
rect 11057 1660 11061 1672
rect 11061 1660 11091 1672
rect 11130 1660 11164 1672
rect 11203 1660 11233 1672
rect 11233 1660 11237 1672
rect 11276 1660 11302 1672
rect 11302 1660 11310 1672
rect 11349 1660 11371 1672
rect 11371 1660 11383 1672
rect 11422 1660 11440 1672
rect 11440 1660 11456 1672
rect 11495 1660 11509 1672
rect 11509 1660 11529 1672
rect 11568 1660 11578 1672
rect 11578 1660 11602 1672
rect 11641 1660 11647 1672
rect 11647 1660 11675 1672
rect 11714 1660 11716 1672
rect 11716 1660 11748 1672
rect 11787 1660 11820 1672
rect 11820 1660 11821 1672
rect 11860 1660 11889 1672
rect 11889 1660 11894 1672
rect 11933 1660 11958 1672
rect 11958 1660 11967 1672
rect 12006 1660 12027 1672
rect 12027 1660 12040 1672
rect 12079 1660 12096 1672
rect 12096 1660 12113 1672
rect 12152 1660 12165 1672
rect 12165 1660 12186 1672
rect 12225 1660 12234 1672
rect 12234 1660 12259 1672
rect 12298 1660 12303 1672
rect 12303 1660 12332 1672
rect 12371 1660 12372 1672
rect 12372 1660 12405 1672
rect 9734 1638 9768 1660
rect 9808 1638 9842 1660
rect 9882 1638 9916 1660
rect 9956 1638 9990 1660
rect 10030 1638 10064 1660
rect 10104 1638 10138 1660
rect 10178 1638 10212 1660
rect 10252 1638 10286 1660
rect 10326 1638 10360 1660
rect 10400 1638 10434 1660
rect 10473 1638 10507 1660
rect 10546 1638 10580 1660
rect 10619 1638 10653 1660
rect 10692 1638 10726 1660
rect 10765 1638 10799 1660
rect 10838 1638 10872 1660
rect 10911 1638 10945 1660
rect 10984 1638 11018 1660
rect 11057 1638 11091 1660
rect 11130 1638 11164 1660
rect 11203 1638 11237 1660
rect 11276 1638 11310 1660
rect 11349 1638 11383 1660
rect 11422 1638 11456 1660
rect 11495 1638 11529 1660
rect 11568 1638 11602 1660
rect 11641 1638 11675 1660
rect 11714 1638 11748 1660
rect 11787 1638 11821 1660
rect 11860 1638 11894 1660
rect 11933 1638 11967 1660
rect 12006 1638 12040 1660
rect 12079 1638 12113 1660
rect 12152 1638 12186 1660
rect 12225 1638 12259 1660
rect 12298 1638 12332 1660
rect 12371 1638 12405 1660
rect 16847 1610 16881 1644
rect 16919 1610 16953 1644
rect 16991 1610 17025 1644
rect 17063 1610 17097 1644
rect 17135 1610 17169 1644
rect 17207 1610 17241 1644
rect 17279 1610 17313 1644
rect 17351 1610 17385 1644
rect 17423 1610 17457 1644
rect 17495 1610 17529 1644
rect 17567 1610 17601 1644
rect 17639 1610 17673 1644
rect 17711 1610 17745 1644
rect 17783 1610 17817 1644
rect 17855 1610 17889 1644
rect 17927 1610 17961 1644
rect 17999 1610 18033 1644
rect 18071 1610 18105 1644
rect 18143 1610 18177 1644
rect 18215 1610 18249 1644
rect 18287 1610 18321 1644
rect 18359 1610 18393 1644
rect 18431 1610 18465 1644
rect 18503 1610 18537 1644
rect 18575 1610 18609 1644
rect 18647 1610 18681 1644
rect 18719 1610 18753 1644
rect 18791 1610 18825 1644
rect 18863 1610 18897 1644
rect 18935 1610 18969 1644
rect 19007 1610 19011 1644
rect 19011 1610 19041 1644
rect 19079 1627 19113 1644
rect 19079 1610 19113 1627
rect 19151 1627 19185 1644
rect 19151 1610 19152 1627
rect 19152 1610 19185 1627
rect 19973 1812 20007 1846
rect 25309 1794 25343 1828
rect 25381 1794 25415 1828
rect 19973 1734 20007 1768
rect 19973 1656 20007 1690
rect 9411 1559 9445 1592
rect 9411 1558 9445 1559
rect 9734 1556 9768 1590
rect 9808 1556 9842 1590
rect 9882 1556 9916 1590
rect 9956 1556 9990 1590
rect 10030 1556 10064 1590
rect 10104 1556 10138 1590
rect 10178 1556 10212 1590
rect 10252 1556 10286 1590
rect 10326 1556 10360 1590
rect 10400 1556 10434 1590
rect 10473 1556 10507 1590
rect 10546 1556 10580 1590
rect 10619 1556 10653 1590
rect 10692 1556 10726 1590
rect 10765 1556 10799 1590
rect 10838 1556 10872 1590
rect 10911 1556 10945 1590
rect 10984 1556 11018 1590
rect 11057 1556 11091 1590
rect 11130 1556 11164 1590
rect 11203 1556 11237 1590
rect 11276 1556 11310 1590
rect 11349 1556 11383 1590
rect 11422 1556 11456 1590
rect 11495 1556 11529 1590
rect 11568 1556 11602 1590
rect 11641 1556 11675 1590
rect 11714 1556 11748 1590
rect 11787 1556 11821 1590
rect 11860 1556 11894 1590
rect 11933 1556 11967 1590
rect 12006 1556 12040 1590
rect 12079 1556 12113 1590
rect 12152 1556 12186 1590
rect 12225 1556 12259 1590
rect 12298 1556 12332 1590
rect 12371 1556 12405 1590
rect 19973 1578 20007 1612
rect 2420 1395 2436 1429
rect 2436 1395 2454 1429
rect 2492 1395 2504 1429
rect 2504 1395 2526 1429
rect 2564 1395 2572 1429
rect 2572 1395 2598 1429
rect 2636 1395 2640 1429
rect 2640 1395 2670 1429
rect 2708 1395 2742 1429
rect 2780 1395 2810 1429
rect 2810 1395 2814 1429
rect 2852 1395 2878 1429
rect 2878 1395 2886 1429
rect 2924 1395 2946 1429
rect 2946 1395 2958 1429
rect 2996 1395 3014 1429
rect 3014 1395 3030 1429
rect 3068 1395 3082 1429
rect 3082 1395 3102 1429
rect 3140 1395 3150 1429
rect 3150 1395 3174 1429
rect 3212 1395 3218 1429
rect 3218 1395 3246 1429
rect 3284 1395 3286 1429
rect 3286 1395 3318 1429
rect 3356 1395 3388 1429
rect 3388 1395 3390 1429
rect 3428 1395 3456 1429
rect 3456 1395 3462 1429
rect 3500 1395 3524 1429
rect 3524 1395 3534 1429
rect 3572 1395 3592 1429
rect 3592 1395 3606 1429
rect 3644 1395 3660 1429
rect 3660 1395 3678 1429
rect 3716 1395 3728 1429
rect 3728 1395 3750 1429
rect 3788 1395 3796 1429
rect 3796 1395 3822 1429
rect 3860 1395 3864 1429
rect 3864 1395 3894 1429
rect 3932 1395 3966 1429
rect 4004 1395 4034 1429
rect 4034 1395 4038 1429
rect 4076 1395 4102 1429
rect 4102 1395 4110 1429
rect 4148 1395 4170 1429
rect 4170 1395 4182 1429
rect 4220 1395 4238 1429
rect 4238 1395 4254 1429
rect 4292 1395 4306 1429
rect 4306 1395 4326 1429
rect 4364 1395 4374 1429
rect 4374 1395 4398 1429
rect 7511 1439 7519 1473
rect 7519 1439 7545 1473
rect 7601 1439 7635 1473
rect 7691 1439 7716 1473
rect 7716 1439 7725 1473
rect 7781 1439 7793 1473
rect 7793 1439 7815 1473
rect 9411 1491 9445 1513
rect 9411 1479 9445 1491
rect 466 1327 500 1361
rect 466 1255 500 1289
rect 2151 1343 2185 1368
rect 2151 1334 2185 1343
rect 570 1245 586 1279
rect 586 1245 604 1279
rect 642 1245 654 1279
rect 654 1245 676 1279
rect 714 1245 722 1279
rect 722 1245 748 1279
rect 786 1245 790 1279
rect 790 1245 820 1279
rect 858 1245 892 1279
rect 930 1245 960 1279
rect 960 1245 964 1279
rect 1002 1245 1028 1279
rect 1028 1245 1036 1279
rect 1074 1245 1096 1279
rect 1096 1245 1108 1279
rect 1146 1245 1164 1279
rect 1164 1245 1180 1279
rect 1218 1245 1232 1279
rect 1232 1245 1252 1279
rect 1290 1245 1300 1279
rect 1300 1245 1324 1279
rect 1362 1245 1368 1279
rect 1368 1245 1396 1279
rect 1434 1245 1436 1279
rect 1436 1245 1468 1279
rect 1506 1245 1540 1279
rect 2151 1275 2185 1294
rect 2151 1260 2185 1275
rect 466 1183 500 1217
rect 466 1111 500 1145
rect 1622 1184 1656 1204
rect 1622 1170 1656 1184
rect 570 1089 586 1123
rect 586 1089 604 1123
rect 642 1089 654 1123
rect 654 1089 676 1123
rect 714 1089 722 1123
rect 722 1089 748 1123
rect 786 1089 790 1123
rect 790 1089 820 1123
rect 858 1089 892 1123
rect 930 1089 960 1123
rect 960 1089 964 1123
rect 1002 1089 1028 1123
rect 1028 1089 1036 1123
rect 1074 1089 1096 1123
rect 1096 1089 1108 1123
rect 1146 1089 1164 1123
rect 1164 1089 1180 1123
rect 1218 1089 1232 1123
rect 1232 1089 1252 1123
rect 1290 1089 1300 1123
rect 1300 1089 1324 1123
rect 1362 1089 1368 1123
rect 1368 1089 1396 1123
rect 1434 1089 1436 1123
rect 1436 1089 1468 1123
rect 1506 1089 1540 1123
rect 1622 1089 1656 1119
rect 466 1039 500 1073
rect 466 967 500 1001
rect 1622 1085 1656 1089
rect 1622 1028 1656 1033
rect 1622 999 1656 1028
rect 2151 1207 2185 1220
rect 2151 1186 2185 1207
rect 4688 1395 4712 1429
rect 4712 1395 4722 1429
rect 4760 1395 4780 1429
rect 4780 1395 4794 1429
rect 4832 1395 4848 1429
rect 4848 1395 4866 1429
rect 4904 1395 4916 1429
rect 4916 1395 4938 1429
rect 4976 1395 4984 1429
rect 4984 1395 5010 1429
rect 5048 1395 5052 1429
rect 5052 1395 5082 1429
rect 5120 1395 5154 1429
rect 5192 1395 5222 1429
rect 5222 1395 5226 1429
rect 5264 1395 5290 1429
rect 5290 1395 5298 1429
rect 5336 1395 5358 1429
rect 5358 1395 5370 1429
rect 5408 1395 5426 1429
rect 5426 1395 5442 1429
rect 5480 1395 5494 1429
rect 5494 1395 5514 1429
rect 5552 1395 5562 1429
rect 5562 1395 5586 1429
rect 5624 1395 5630 1429
rect 5630 1395 5658 1429
rect 5696 1395 5698 1429
rect 5698 1395 5730 1429
rect 5768 1395 5800 1429
rect 5800 1395 5802 1429
rect 5840 1395 5868 1429
rect 5868 1395 5874 1429
rect 5912 1395 5936 1429
rect 5936 1395 5946 1429
rect 5984 1395 6004 1429
rect 6004 1395 6018 1429
rect 6056 1395 6072 1429
rect 6072 1395 6090 1429
rect 6128 1395 6140 1429
rect 6140 1395 6162 1429
rect 6200 1395 6208 1429
rect 6208 1395 6234 1429
rect 6272 1395 6276 1429
rect 6276 1395 6306 1429
rect 6344 1395 6378 1429
rect 6416 1395 6446 1429
rect 6446 1395 6450 1429
rect 6488 1395 6514 1429
rect 6514 1395 6522 1429
rect 6560 1395 6582 1429
rect 6582 1395 6594 1429
rect 6632 1395 6650 1429
rect 6650 1395 6666 1429
rect 9411 1423 9445 1434
rect 9411 1400 9445 1423
rect 4486 1323 4520 1355
rect 4486 1321 4506 1323
rect 4506 1321 4520 1323
rect 4558 1334 4580 1355
rect 4580 1334 4592 1355
rect 4558 1321 4592 1334
rect 4486 1254 4520 1273
rect 4486 1239 4506 1254
rect 4506 1239 4520 1254
rect 4558 1254 4592 1273
rect 4558 1239 4580 1254
rect 4580 1239 4592 1254
rect 7424 1355 7458 1389
rect 7424 1295 7458 1317
rect 7424 1283 7458 1295
rect 7424 1227 7458 1245
rect 7424 1211 7458 1227
rect 2420 1159 2436 1193
rect 2436 1159 2454 1193
rect 2492 1159 2504 1193
rect 2504 1159 2526 1193
rect 2564 1159 2572 1193
rect 2572 1159 2598 1193
rect 2636 1159 2640 1193
rect 2640 1159 2670 1193
rect 2708 1159 2742 1193
rect 2780 1159 2810 1193
rect 2810 1159 2814 1193
rect 2852 1159 2878 1193
rect 2878 1159 2886 1193
rect 2924 1159 2946 1193
rect 2946 1159 2958 1193
rect 2996 1159 3014 1193
rect 3014 1159 3030 1193
rect 3068 1159 3082 1193
rect 3082 1159 3102 1193
rect 3140 1159 3150 1193
rect 3150 1159 3174 1193
rect 3212 1159 3218 1193
rect 3218 1159 3246 1193
rect 3284 1159 3286 1193
rect 3286 1159 3318 1193
rect 3356 1159 3388 1193
rect 3388 1159 3390 1193
rect 3428 1159 3456 1193
rect 3456 1159 3462 1193
rect 3500 1159 3524 1193
rect 3524 1159 3534 1193
rect 3572 1159 3592 1193
rect 3592 1159 3606 1193
rect 3644 1159 3660 1193
rect 3660 1159 3678 1193
rect 3716 1159 3728 1193
rect 3728 1159 3750 1193
rect 3788 1159 3796 1193
rect 3796 1159 3822 1193
rect 3860 1159 3864 1193
rect 3864 1159 3894 1193
rect 3932 1159 3966 1193
rect 4004 1159 4034 1193
rect 4034 1159 4038 1193
rect 4076 1159 4102 1193
rect 4102 1159 4110 1193
rect 4148 1159 4170 1193
rect 4170 1159 4182 1193
rect 4220 1159 4238 1193
rect 4238 1159 4254 1193
rect 4292 1159 4306 1193
rect 4306 1159 4326 1193
rect 4364 1159 4374 1193
rect 4374 1159 4398 1193
rect 4688 1159 4712 1193
rect 4712 1159 4722 1193
rect 4760 1159 4780 1193
rect 4780 1159 4794 1193
rect 4832 1159 4848 1193
rect 4848 1159 4866 1193
rect 4904 1159 4916 1193
rect 4916 1159 4938 1193
rect 4976 1159 4984 1193
rect 4984 1159 5010 1193
rect 5048 1159 5052 1193
rect 5052 1159 5082 1193
rect 5120 1159 5154 1193
rect 5192 1159 5222 1193
rect 5222 1159 5226 1193
rect 5264 1159 5290 1193
rect 5290 1159 5298 1193
rect 5336 1159 5358 1193
rect 5358 1159 5370 1193
rect 5408 1159 5426 1193
rect 5426 1159 5442 1193
rect 5480 1159 5494 1193
rect 5494 1159 5514 1193
rect 5552 1159 5562 1193
rect 5562 1159 5586 1193
rect 5624 1159 5630 1193
rect 5630 1159 5658 1193
rect 5696 1159 5698 1193
rect 5698 1159 5730 1193
rect 5768 1159 5800 1193
rect 5800 1159 5802 1193
rect 5840 1159 5868 1193
rect 5868 1159 5874 1193
rect 5912 1159 5936 1193
rect 5936 1159 5946 1193
rect 5984 1159 6004 1193
rect 6004 1159 6018 1193
rect 6056 1159 6072 1193
rect 6072 1159 6090 1193
rect 6128 1159 6140 1193
rect 6140 1159 6162 1193
rect 6200 1159 6208 1193
rect 6208 1159 6234 1193
rect 6272 1159 6276 1193
rect 6276 1159 6306 1193
rect 6344 1159 6378 1193
rect 6416 1159 6446 1193
rect 6446 1159 6450 1193
rect 6488 1159 6514 1193
rect 6514 1159 6522 1193
rect 6560 1159 6582 1193
rect 6582 1159 6594 1193
rect 6632 1159 6650 1193
rect 6650 1159 6666 1193
rect 7424 1159 7458 1173
rect 2151 1139 2185 1146
rect 2151 1112 2185 1139
rect 7424 1139 7458 1159
rect 2151 1071 2185 1072
rect 2151 1038 2185 1071
rect 2466 1064 2467 1098
rect 2467 1064 2500 1098
rect 2549 1064 2573 1098
rect 2573 1064 2583 1098
rect 2632 1064 2645 1098
rect 2645 1064 2666 1098
rect 2715 1064 2717 1098
rect 2717 1064 2749 1098
rect 2797 1064 2827 1098
rect 2827 1064 2831 1098
rect 2879 1064 2898 1098
rect 2898 1064 2913 1098
rect 2961 1064 2969 1098
rect 2969 1064 2995 1098
rect 3094 1064 3125 1098
rect 3125 1064 3128 1098
rect 3177 1064 3196 1098
rect 3196 1064 3211 1098
rect 3259 1064 3267 1098
rect 3267 1064 3293 1098
rect 3341 1064 3375 1098
rect 3423 1064 3449 1098
rect 3449 1064 3457 1098
rect 3505 1064 3521 1098
rect 3521 1064 3539 1098
rect 3587 1064 3593 1098
rect 3593 1064 3621 1098
rect 3842 1064 3873 1098
rect 3873 1064 3876 1098
rect 3933 1064 3934 1098
rect 3934 1064 3967 1098
rect 4023 1064 4029 1098
rect 4029 1064 4057 1098
rect 4147 1064 4151 1097
rect 4151 1064 4181 1097
rect 4252 1064 4280 1097
rect 4280 1064 4286 1097
rect 4357 1064 4375 1097
rect 4375 1064 4391 1097
rect 4147 1063 4181 1064
rect 4252 1063 4286 1064
rect 4357 1063 4391 1064
rect 570 933 586 967
rect 586 933 604 967
rect 642 933 654 967
rect 654 933 676 967
rect 714 933 722 967
rect 722 933 748 967
rect 786 933 790 967
rect 790 933 820 967
rect 858 933 892 967
rect 930 933 960 967
rect 960 933 964 967
rect 1002 933 1028 967
rect 1028 933 1036 967
rect 1074 933 1096 967
rect 1096 933 1108 967
rect 1146 933 1164 967
rect 1164 933 1180 967
rect 1218 933 1232 967
rect 1232 933 1252 967
rect 1290 933 1300 967
rect 1300 933 1324 967
rect 1362 933 1368 967
rect 1368 933 1396 967
rect 1434 933 1436 967
rect 1436 933 1468 967
rect 1506 933 1540 967
rect 2151 969 2185 998
rect 2151 964 2185 969
rect 4603 1064 4619 1097
rect 4619 1064 4637 1097
rect 4603 1063 4637 1064
rect 4677 1063 4711 1097
rect 4751 1063 4785 1097
rect 4825 1064 4843 1097
rect 4843 1064 4859 1097
rect 4825 1063 4859 1064
rect 5071 1064 5087 1097
rect 5087 1064 5105 1097
rect 5144 1064 5157 1097
rect 5157 1064 5178 1097
rect 5217 1064 5226 1097
rect 5226 1064 5251 1097
rect 5289 1064 5295 1097
rect 5295 1064 5323 1097
rect 5361 1064 5364 1097
rect 5364 1064 5395 1097
rect 5433 1064 5467 1097
rect 5730 1064 5763 1098
rect 5763 1064 5764 1098
rect 5807 1064 5824 1098
rect 5824 1064 5841 1098
rect 5884 1064 5918 1098
rect 6226 1064 6231 1098
rect 6231 1064 6260 1098
rect 6298 1064 6332 1098
rect 6442 1064 6461 1096
rect 6461 1064 6476 1096
rect 6516 1064 6544 1096
rect 6544 1064 6550 1096
rect 5071 1063 5105 1064
rect 5144 1063 5178 1064
rect 5217 1063 5251 1064
rect 5289 1063 5323 1064
rect 5361 1063 5395 1064
rect 5433 1063 5467 1064
rect 6442 1062 6476 1064
rect 6516 1062 6550 1064
rect 6590 1062 6624 1096
rect 6663 1062 6697 1096
rect 6736 1064 6743 1096
rect 6743 1064 6770 1096
rect 6925 1064 6947 1090
rect 6947 1064 6959 1090
rect 7424 1091 7458 1101
rect 7424 1067 7458 1091
rect 6736 1062 6770 1064
rect 6925 1056 6959 1064
rect 466 895 500 929
rect 466 823 500 857
rect 1427 855 1461 889
rect 1499 855 1533 889
rect 2151 901 2185 924
rect 2151 890 2185 901
rect 2151 833 2185 850
rect 2151 816 2185 833
rect 466 751 500 785
rect 570 777 586 811
rect 586 777 604 811
rect 642 777 654 811
rect 654 777 676 811
rect 714 777 722 811
rect 722 777 748 811
rect 786 777 790 811
rect 790 777 820 811
rect 858 777 892 811
rect 930 777 960 811
rect 960 777 964 811
rect 1002 777 1028 811
rect 1028 777 1036 811
rect 1074 777 1096 811
rect 1096 777 1108 811
rect 1146 777 1164 811
rect 1164 777 1180 811
rect 1218 777 1232 811
rect 1232 777 1252 811
rect 1290 777 1300 811
rect 1300 777 1324 811
rect 1362 777 1368 811
rect 1368 777 1396 811
rect 1434 777 1436 811
rect 1436 777 1468 811
rect 1506 777 1540 811
rect 466 679 500 713
rect 1622 716 1656 736
rect 1622 702 1656 716
rect 466 607 500 641
rect 570 621 586 655
rect 586 621 604 655
rect 642 621 654 655
rect 654 621 676 655
rect 714 621 722 655
rect 722 621 748 655
rect 786 621 790 655
rect 790 621 820 655
rect 858 621 892 655
rect 930 621 960 655
rect 960 621 964 655
rect 1002 621 1028 655
rect 1028 621 1036 655
rect 1074 621 1096 655
rect 1096 621 1108 655
rect 1146 621 1164 655
rect 1164 621 1180 655
rect 1218 621 1232 655
rect 1232 621 1252 655
rect 1290 621 1300 655
rect 1300 621 1324 655
rect 1362 621 1368 655
rect 1368 621 1396 655
rect 1434 621 1436 655
rect 1436 621 1468 655
rect 1506 621 1540 655
rect 1622 621 1656 640
rect 466 535 500 569
rect 1622 606 1656 621
rect 1622 526 1656 544
rect 1622 510 1656 526
rect 2151 765 2185 776
rect 2151 742 2185 765
rect 2151 697 2185 702
rect 2151 668 2185 697
rect 2151 595 2185 628
rect 2151 594 2185 595
rect 466 463 500 497
rect 570 465 586 499
rect 586 465 604 499
rect 642 465 654 499
rect 654 465 676 499
rect 714 465 722 499
rect 722 465 748 499
rect 786 465 790 499
rect 790 465 820 499
rect 858 465 892 499
rect 930 465 960 499
rect 960 465 964 499
rect 1002 465 1028 499
rect 1028 465 1036 499
rect 1074 465 1096 499
rect 1096 465 1108 499
rect 1146 465 1164 499
rect 1164 465 1180 499
rect 1218 465 1232 499
rect 1232 465 1252 499
rect 1290 465 1300 499
rect 1300 465 1324 499
rect 1362 465 1368 499
rect 1368 465 1396 499
rect 1434 465 1436 499
rect 1436 465 1468 499
rect 1506 465 1540 499
rect 2151 527 2185 554
rect 2151 520 2185 527
rect 466 391 500 425
rect 1427 387 1461 421
rect 1499 387 1533 421
rect 2151 459 2185 480
rect 2151 446 2185 459
rect 2151 391 2185 406
rect 2151 372 2185 391
rect 466 319 500 353
rect 570 309 586 343
rect 586 309 604 343
rect 642 309 654 343
rect 654 309 676 343
rect 714 309 722 343
rect 722 309 748 343
rect 786 309 790 343
rect 790 309 820 343
rect 858 309 892 343
rect 930 309 960 343
rect 960 309 964 343
rect 1002 309 1028 343
rect 1028 309 1036 343
rect 1074 309 1096 343
rect 1096 309 1108 343
rect 1146 309 1164 343
rect 1164 309 1180 343
rect 1218 309 1232 343
rect 1232 309 1252 343
rect 1290 309 1300 343
rect 1300 309 1324 343
rect 1362 309 1368 343
rect 1368 309 1396 343
rect 1434 309 1436 343
rect 1436 309 1468 343
rect 1506 309 1540 343
rect 466 247 500 281
rect 466 175 500 209
rect 1622 248 1656 268
rect 1622 234 1656 248
rect 570 153 586 187
rect 586 153 604 187
rect 642 153 654 187
rect 654 153 676 187
rect 714 153 722 187
rect 722 153 748 187
rect 786 153 790 187
rect 790 153 820 187
rect 858 153 892 187
rect 930 153 960 187
rect 960 153 964 187
rect 1002 153 1028 187
rect 1028 153 1036 187
rect 1074 153 1096 187
rect 1096 153 1108 187
rect 1146 153 1164 187
rect 1164 153 1180 187
rect 1218 153 1232 187
rect 1232 153 1252 187
rect 1290 153 1300 187
rect 1300 153 1324 187
rect 1362 153 1368 187
rect 1368 153 1396 187
rect 1434 153 1436 187
rect 1436 153 1468 187
rect 1506 153 1540 187
rect 1622 153 1656 172
rect 466 103 500 137
rect 466 31 500 65
rect 1622 138 1656 153
rect 1622 58 1656 76
rect 1622 42 1656 58
rect 2151 323 2185 332
rect 2151 298 2185 323
rect 2151 255 2185 258
rect 2151 224 2185 255
rect 2151 153 2185 184
rect 2151 150 2185 153
rect 2151 85 2185 110
rect 2151 76 2185 85
rect 570 -3 586 31
rect 586 -3 604 31
rect 642 -3 654 31
rect 654 -3 676 31
rect 714 -3 722 31
rect 722 -3 748 31
rect 786 -3 790 31
rect 790 -3 820 31
rect 858 -3 892 31
rect 930 -3 960 31
rect 960 -3 964 31
rect 1002 -3 1028 31
rect 1028 -3 1036 31
rect 1074 -3 1096 31
rect 1096 -3 1108 31
rect 1146 -3 1164 31
rect 1164 -3 1180 31
rect 1218 -3 1232 31
rect 1232 -3 1252 31
rect 1290 -3 1300 31
rect 1300 -3 1324 31
rect 1362 -3 1368 31
rect 1368 -3 1396 31
rect 1434 -3 1436 31
rect 1436 -3 1468 31
rect 1506 -3 1540 31
rect 2151 17 2185 36
rect 2151 2 2185 17
rect 2406 948 2440 982
rect 2406 878 2440 910
rect 2406 876 2440 878
rect 2406 810 2440 838
rect 2406 804 2440 810
rect 2406 742 2440 766
rect 2406 732 2440 742
rect 2406 674 2440 694
rect 2406 660 2440 674
rect 2406 606 2440 622
rect 2406 588 2440 606
rect 2406 538 2440 550
rect 2406 516 2440 538
rect 2406 470 2440 478
rect 2406 444 2440 470
rect 2406 402 2440 406
rect 2406 372 2440 402
rect 2406 300 2440 334
rect 2406 232 2440 262
rect 2406 228 2440 232
rect 2406 164 2440 190
rect 2406 156 2440 164
rect 2406 96 2440 118
rect 2406 84 2440 96
rect 2406 28 2440 46
rect 2406 12 2440 28
rect 2562 948 2596 982
rect 2562 878 2596 910
rect 2562 876 2596 878
rect 2562 810 2596 838
rect 2562 804 2596 810
rect 2562 742 2596 766
rect 2562 732 2596 742
rect 2562 674 2596 694
rect 2562 660 2596 674
rect 2562 606 2596 622
rect 2562 588 2596 606
rect 2562 538 2596 550
rect 2562 516 2596 538
rect 2562 470 2596 478
rect 2562 444 2596 470
rect 2562 402 2596 406
rect 2562 372 2596 402
rect 2562 300 2596 334
rect 2562 232 2596 262
rect 2562 228 2596 232
rect 2562 164 2596 190
rect 2562 156 2596 164
rect 2562 96 2596 118
rect 2562 84 2596 96
rect 2562 28 2596 46
rect 2562 12 2596 28
rect 2718 948 2752 982
rect 2718 878 2752 910
rect 2718 876 2752 878
rect 2718 810 2752 838
rect 2718 804 2752 810
rect 2718 742 2752 766
rect 2718 732 2752 742
rect 2718 674 2752 694
rect 2718 660 2752 674
rect 2718 606 2752 622
rect 2718 588 2752 606
rect 2718 538 2752 550
rect 2718 516 2752 538
rect 2718 470 2752 478
rect 2718 444 2752 470
rect 2718 402 2752 406
rect 2718 372 2752 402
rect 2718 300 2752 334
rect 2718 232 2752 262
rect 2718 228 2752 232
rect 2718 164 2752 190
rect 2718 156 2752 164
rect 2718 96 2752 118
rect 2718 84 2752 96
rect 2718 28 2752 46
rect 2718 12 2752 28
rect 2874 948 2908 982
rect 2874 878 2908 910
rect 2874 876 2908 878
rect 2874 810 2908 838
rect 2874 804 2908 810
rect 2874 742 2908 766
rect 2874 732 2908 742
rect 2874 674 2908 694
rect 2874 660 2908 674
rect 2874 606 2908 622
rect 2874 588 2908 606
rect 2874 538 2908 550
rect 2874 516 2908 538
rect 2874 470 2908 478
rect 2874 444 2908 470
rect 2874 402 2908 406
rect 2874 372 2908 402
rect 2874 300 2908 334
rect 2874 232 2908 262
rect 2874 228 2908 232
rect 2874 164 2908 190
rect 2874 156 2908 164
rect 2874 96 2908 118
rect 2874 84 2908 96
rect 2874 28 2908 46
rect 2874 12 2908 28
rect 3030 948 3064 982
rect 3030 878 3064 910
rect 3030 876 3064 878
rect 3030 810 3064 838
rect 3030 804 3064 810
rect 3030 742 3064 766
rect 3030 732 3064 742
rect 3030 674 3064 694
rect 3030 660 3064 674
rect 3030 606 3064 622
rect 3030 588 3064 606
rect 3030 538 3064 550
rect 3030 516 3064 538
rect 3030 470 3064 478
rect 3030 444 3064 470
rect 3030 402 3064 406
rect 3030 372 3064 402
rect 3030 300 3064 334
rect 3030 232 3064 262
rect 3030 228 3064 232
rect 3030 164 3064 190
rect 3030 156 3064 164
rect 3030 96 3064 118
rect 3030 84 3064 96
rect 3030 28 3064 46
rect 3030 12 3064 28
rect 3186 948 3220 982
rect 3186 878 3220 910
rect 3186 876 3220 878
rect 3186 810 3220 838
rect 3186 804 3220 810
rect 3186 742 3220 766
rect 3186 732 3220 742
rect 3186 674 3220 694
rect 3186 660 3220 674
rect 3186 606 3220 622
rect 3186 588 3220 606
rect 3186 538 3220 550
rect 3186 516 3220 538
rect 3186 470 3220 478
rect 3186 444 3220 470
rect 3186 402 3220 406
rect 3186 372 3220 402
rect 3186 300 3220 334
rect 3186 232 3220 262
rect 3186 228 3220 232
rect 3186 164 3220 190
rect 3186 156 3220 164
rect 3186 96 3220 118
rect 3186 84 3220 96
rect 3186 28 3220 46
rect 3186 12 3220 28
rect 3342 948 3376 982
rect 3342 878 3376 910
rect 3342 876 3376 878
rect 3342 810 3376 838
rect 3342 804 3376 810
rect 3342 742 3376 766
rect 3342 732 3376 742
rect 3342 674 3376 694
rect 3342 660 3376 674
rect 3342 606 3376 622
rect 3342 588 3376 606
rect 3342 538 3376 550
rect 3342 516 3376 538
rect 3342 470 3376 478
rect 3342 444 3376 470
rect 3342 402 3376 406
rect 3342 372 3376 402
rect 3342 300 3376 334
rect 3342 232 3376 262
rect 3342 228 3376 232
rect 3342 164 3376 190
rect 3342 156 3376 164
rect 3342 96 3376 118
rect 3342 84 3376 96
rect 3342 28 3376 46
rect 3342 12 3376 28
rect 3498 948 3532 982
rect 3498 878 3532 910
rect 3498 876 3532 878
rect 3498 810 3532 838
rect 3498 804 3532 810
rect 3498 742 3532 766
rect 3498 732 3532 742
rect 3498 674 3532 694
rect 3498 660 3532 674
rect 3498 606 3532 622
rect 3498 588 3532 606
rect 3498 538 3532 550
rect 3498 516 3532 538
rect 3498 470 3532 478
rect 3498 444 3532 470
rect 3498 402 3532 406
rect 3498 372 3532 402
rect 3498 300 3532 334
rect 3498 232 3532 262
rect 3498 228 3532 232
rect 3498 164 3532 190
rect 3498 156 3532 164
rect 3498 96 3532 118
rect 3498 84 3532 96
rect 3498 28 3532 46
rect 3498 12 3532 28
rect 3654 948 3688 982
rect 3654 878 3688 910
rect 3654 876 3688 878
rect 3654 810 3688 838
rect 3654 804 3688 810
rect 3654 742 3688 766
rect 3654 732 3688 742
rect 3654 674 3688 694
rect 3654 660 3688 674
rect 3654 606 3688 622
rect 3654 588 3688 606
rect 3654 538 3688 550
rect 3654 516 3688 538
rect 3654 470 3688 478
rect 3654 444 3688 470
rect 3654 402 3688 406
rect 3654 372 3688 402
rect 3654 300 3688 334
rect 3654 232 3688 262
rect 3654 228 3688 232
rect 3654 164 3688 190
rect 3654 156 3688 164
rect 3654 96 3688 118
rect 3654 84 3688 96
rect 3654 28 3688 46
rect 3654 12 3688 28
rect 3778 948 3812 982
rect 3778 878 3812 910
rect 3778 876 3812 878
rect 3778 810 3812 838
rect 3778 804 3812 810
rect 3778 742 3812 766
rect 3778 732 3812 742
rect 3778 674 3812 694
rect 3778 660 3812 674
rect 3778 606 3812 622
rect 3778 588 3812 606
rect 3778 538 3812 550
rect 3778 516 3812 538
rect 3778 470 3812 478
rect 3778 444 3812 470
rect 3778 402 3812 406
rect 3778 372 3812 402
rect 3778 300 3812 334
rect 3778 232 3812 262
rect 3778 228 3812 232
rect 3778 164 3812 190
rect 3778 156 3812 164
rect 3778 96 3812 118
rect 3778 84 3812 96
rect 3778 28 3812 46
rect 3778 12 3812 28
rect 3934 948 3968 982
rect 3934 878 3968 910
rect 3934 876 3968 878
rect 3934 810 3968 838
rect 3934 804 3968 810
rect 3934 742 3968 766
rect 3934 732 3968 742
rect 3934 674 3968 694
rect 3934 660 3968 674
rect 3934 606 3968 622
rect 3934 588 3968 606
rect 3934 538 3968 550
rect 3934 516 3968 538
rect 3934 470 3968 478
rect 3934 444 3968 470
rect 3934 402 3968 406
rect 3934 372 3968 402
rect 3934 300 3968 334
rect 3934 232 3968 262
rect 3934 228 3968 232
rect 3934 164 3968 190
rect 3934 156 3968 164
rect 3934 96 3968 118
rect 3934 84 3968 96
rect 3934 28 3968 46
rect 3934 12 3968 28
rect 4090 948 4124 982
rect 4090 878 4124 910
rect 4090 876 4124 878
rect 4090 810 4124 838
rect 4090 804 4124 810
rect 4090 742 4124 766
rect 4090 732 4124 742
rect 4090 674 4124 694
rect 4090 660 4124 674
rect 4090 606 4124 622
rect 4090 588 4124 606
rect 4090 538 4124 550
rect 4090 516 4124 538
rect 4090 470 4124 478
rect 4090 444 4124 470
rect 4090 402 4124 406
rect 4090 372 4124 402
rect 4090 300 4124 334
rect 4090 232 4124 262
rect 4090 228 4124 232
rect 4090 164 4124 190
rect 4090 156 4124 164
rect 4090 96 4124 118
rect 4090 84 4124 96
rect 4090 28 4124 46
rect 4090 12 4124 28
rect 4246 948 4280 982
rect 4246 878 4280 910
rect 4246 876 4280 878
rect 4246 810 4280 838
rect 4246 804 4280 810
rect 4246 742 4280 766
rect 4246 732 4280 742
rect 4246 674 4280 694
rect 4246 660 4280 674
rect 4246 606 4280 622
rect 4246 588 4280 606
rect 4246 538 4280 550
rect 4246 516 4280 538
rect 4246 470 4280 478
rect 4246 444 4280 470
rect 4246 402 4280 406
rect 4246 372 4280 402
rect 4246 300 4280 334
rect 4246 232 4280 262
rect 4246 228 4280 232
rect 4246 164 4280 190
rect 4246 156 4280 164
rect 4246 96 4280 118
rect 4246 84 4280 96
rect 4246 28 4280 46
rect 4246 12 4280 28
rect 4402 948 4436 982
rect 4558 948 4592 982
rect 4402 878 4436 910
rect 4402 876 4436 878
rect 4558 878 4592 910
rect 4558 876 4592 878
rect 4402 810 4436 838
rect 4402 804 4436 810
rect 4558 810 4592 838
rect 4558 804 4592 810
rect 4402 742 4436 766
rect 4402 732 4436 742
rect 4558 742 4592 766
rect 4558 732 4592 742
rect 4402 674 4436 694
rect 4402 660 4436 674
rect 4558 674 4592 694
rect 4558 660 4592 674
rect 4402 606 4436 622
rect 4402 588 4436 606
rect 4558 606 4592 622
rect 4558 588 4592 606
rect 4402 538 4436 550
rect 4402 516 4436 538
rect 4558 538 4592 550
rect 4558 516 4592 538
rect 4402 470 4436 478
rect 4402 444 4436 470
rect 4558 470 4592 478
rect 4558 444 4592 470
rect 4402 402 4436 406
rect 4402 372 4436 402
rect 4558 402 4592 406
rect 4558 372 4592 402
rect 4402 300 4436 334
rect 4558 300 4592 334
rect 4402 232 4436 262
rect 4402 228 4436 232
rect 4558 232 4592 262
rect 4558 228 4592 232
rect 4402 164 4436 190
rect 4402 156 4436 164
rect 4558 164 4592 190
rect 4558 156 4592 164
rect 4402 96 4436 118
rect 4402 84 4436 96
rect 4558 96 4592 118
rect 4558 84 4592 96
rect 4402 28 4436 46
rect 4402 12 4436 28
rect 4558 28 4592 46
rect 4558 12 4592 28
rect 4714 948 4748 982
rect 4714 878 4748 910
rect 4714 876 4748 878
rect 4714 810 4748 838
rect 4714 804 4748 810
rect 4714 742 4748 766
rect 4714 732 4748 742
rect 4714 674 4748 694
rect 4714 660 4748 674
rect 4714 606 4748 622
rect 4714 588 4748 606
rect 4714 538 4748 550
rect 4714 516 4748 538
rect 4714 470 4748 478
rect 4714 444 4748 470
rect 4714 402 4748 406
rect 4714 372 4748 402
rect 4714 300 4748 334
rect 4714 232 4748 262
rect 4714 228 4748 232
rect 4714 164 4748 190
rect 4714 156 4748 164
rect 4714 96 4748 118
rect 4714 84 4748 96
rect 4714 28 4748 46
rect 4714 12 4748 28
rect 4870 948 4904 982
rect 5026 948 5060 982
rect 4870 878 4904 910
rect 4870 876 4904 878
rect 5026 878 5060 910
rect 5026 876 5060 878
rect 4870 810 4904 838
rect 4870 804 4904 810
rect 5026 810 5060 838
rect 5026 804 5060 810
rect 4870 742 4904 766
rect 4870 732 4904 742
rect 5026 742 5060 766
rect 5026 732 5060 742
rect 4870 674 4904 694
rect 4870 660 4904 674
rect 5026 674 5060 694
rect 5026 660 5060 674
rect 4870 606 4904 622
rect 4870 588 4904 606
rect 5026 606 5060 622
rect 5026 588 5060 606
rect 4870 538 4904 550
rect 4870 516 4904 538
rect 5026 538 5060 550
rect 5026 516 5060 538
rect 4870 470 4904 478
rect 4870 444 4904 470
rect 5026 470 5060 478
rect 5026 444 5060 470
rect 4870 402 4904 406
rect 4870 372 4904 402
rect 5026 402 5060 406
rect 5026 372 5060 402
rect 4870 300 4904 334
rect 5026 300 5060 334
rect 4870 232 4904 262
rect 4870 228 4904 232
rect 5026 232 5060 262
rect 5026 228 5060 232
rect 4870 164 4904 190
rect 4870 156 4904 164
rect 5026 164 5060 190
rect 5026 156 5060 164
rect 4870 96 4904 118
rect 4870 84 4904 96
rect 5026 96 5060 118
rect 5026 84 5060 96
rect 4870 28 4904 46
rect 4870 12 4904 28
rect 5026 28 5060 46
rect 5026 12 5060 28
rect 5182 948 5216 982
rect 5182 878 5216 910
rect 5182 876 5216 878
rect 5182 810 5216 838
rect 5182 804 5216 810
rect 5182 742 5216 766
rect 5182 732 5216 742
rect 5182 674 5216 694
rect 5182 660 5216 674
rect 5182 606 5216 622
rect 5182 588 5216 606
rect 5182 538 5216 550
rect 5182 516 5216 538
rect 5182 470 5216 478
rect 5182 444 5216 470
rect 5182 402 5216 406
rect 5182 372 5216 402
rect 5182 300 5216 334
rect 5182 232 5216 262
rect 5182 228 5216 232
rect 5182 164 5216 190
rect 5182 156 5216 164
rect 5182 96 5216 118
rect 5182 84 5216 96
rect 5182 28 5216 46
rect 5182 12 5216 28
rect 5338 948 5372 982
rect 5338 878 5372 910
rect 5338 876 5372 878
rect 5338 810 5372 838
rect 5338 804 5372 810
rect 5338 742 5372 766
rect 5338 732 5372 742
rect 5338 674 5372 694
rect 5338 660 5372 674
rect 5338 606 5372 622
rect 5338 588 5372 606
rect 5338 538 5372 550
rect 5338 516 5372 538
rect 5338 470 5372 478
rect 5338 444 5372 470
rect 5338 402 5372 406
rect 5338 372 5372 402
rect 5338 300 5372 334
rect 5338 232 5372 262
rect 5338 228 5372 232
rect 5338 164 5372 190
rect 5338 156 5372 164
rect 5338 96 5372 118
rect 5338 84 5372 96
rect 5338 28 5372 46
rect 5338 12 5372 28
rect 5494 948 5528 982
rect 5494 878 5528 910
rect 5494 876 5528 878
rect 5494 810 5528 838
rect 5494 804 5528 810
rect 5494 742 5528 766
rect 5494 732 5528 742
rect 5494 674 5528 694
rect 5494 660 5528 674
rect 5494 606 5528 622
rect 5494 588 5528 606
rect 5494 538 5528 550
rect 5494 516 5528 538
rect 5494 470 5528 478
rect 5494 444 5528 470
rect 5494 402 5528 406
rect 5494 372 5528 402
rect 5494 300 5528 334
rect 5494 232 5528 262
rect 5494 228 5528 232
rect 5494 164 5528 190
rect 5494 156 5528 164
rect 5494 96 5528 118
rect 5494 84 5528 96
rect 5494 28 5528 46
rect 5494 12 5528 28
rect 5668 948 5702 982
rect 5668 878 5702 910
rect 5668 876 5702 878
rect 5668 810 5702 838
rect 5668 804 5702 810
rect 5668 742 5702 766
rect 5668 732 5702 742
rect 5668 674 5702 694
rect 5668 660 5702 674
rect 5668 606 5702 622
rect 5668 588 5702 606
rect 5668 538 5702 550
rect 5668 516 5702 538
rect 5668 470 5702 478
rect 5668 444 5702 470
rect 5668 402 5702 406
rect 5668 372 5702 402
rect 5668 300 5702 334
rect 5668 232 5702 262
rect 5668 228 5702 232
rect 5668 164 5702 190
rect 5668 156 5702 164
rect 5668 96 5702 118
rect 5668 84 5702 96
rect 5668 28 5702 46
rect 5668 12 5702 28
rect 5824 948 5858 982
rect 5824 878 5858 910
rect 5824 876 5858 878
rect 5824 810 5858 838
rect 5824 804 5858 810
rect 5824 742 5858 766
rect 5824 732 5858 742
rect 5824 674 5858 694
rect 5824 660 5858 674
rect 5824 606 5858 622
rect 5824 588 5858 606
rect 5824 538 5858 550
rect 5824 516 5858 538
rect 5824 470 5858 478
rect 5824 444 5858 470
rect 5824 402 5858 406
rect 5824 372 5858 402
rect 5824 300 5858 334
rect 5824 232 5858 262
rect 5824 228 5858 232
rect 5824 164 5858 190
rect 5824 156 5858 164
rect 5824 96 5858 118
rect 5824 84 5858 96
rect 5824 28 5858 46
rect 5824 12 5858 28
rect 5980 948 6014 982
rect 5980 878 6014 910
rect 5980 876 6014 878
rect 5980 810 6014 838
rect 5980 804 6014 810
rect 5980 742 6014 766
rect 5980 732 6014 742
rect 5980 674 6014 694
rect 5980 660 6014 674
rect 5980 606 6014 622
rect 5980 588 6014 606
rect 5980 538 6014 550
rect 5980 516 6014 538
rect 5980 470 6014 478
rect 5980 444 6014 470
rect 5980 402 6014 406
rect 5980 372 6014 402
rect 5980 300 6014 334
rect 5980 232 6014 262
rect 5980 228 6014 232
rect 5980 164 6014 190
rect 5980 156 6014 164
rect 5980 96 6014 118
rect 5980 84 6014 96
rect 5980 28 6014 46
rect 5980 12 6014 28
rect 6136 948 6170 982
rect 6136 878 6170 910
rect 6136 876 6170 878
rect 6136 810 6170 838
rect 6136 804 6170 810
rect 6136 742 6170 766
rect 6136 732 6170 742
rect 6136 674 6170 694
rect 6136 660 6170 674
rect 6136 606 6170 622
rect 6136 588 6170 606
rect 6136 538 6170 550
rect 6136 516 6170 538
rect 6136 470 6170 478
rect 6136 444 6170 470
rect 6136 402 6170 406
rect 6136 372 6170 402
rect 6136 300 6170 334
rect 6136 232 6170 262
rect 6136 228 6170 232
rect 6136 164 6170 190
rect 6136 156 6170 164
rect 6136 96 6170 118
rect 6136 84 6170 96
rect 6136 28 6170 46
rect 6136 12 6170 28
rect 6292 948 6326 982
rect 6292 878 6326 910
rect 6292 876 6326 878
rect 6292 810 6326 838
rect 6292 804 6326 810
rect 6292 742 6326 766
rect 6292 732 6326 742
rect 6292 674 6326 694
rect 6292 660 6326 674
rect 6292 606 6326 622
rect 6292 588 6326 606
rect 6292 538 6326 550
rect 6292 516 6326 538
rect 6292 470 6326 478
rect 6292 444 6326 470
rect 6292 402 6326 406
rect 6292 372 6326 402
rect 6292 300 6326 334
rect 6292 232 6326 262
rect 6292 228 6326 232
rect 6292 164 6326 190
rect 6292 156 6326 164
rect 6292 96 6326 118
rect 6292 84 6326 96
rect 6292 28 6326 46
rect 6292 12 6326 28
rect 6416 948 6450 982
rect 6416 878 6450 910
rect 6416 876 6450 878
rect 6416 810 6450 838
rect 6416 804 6450 810
rect 6416 742 6450 766
rect 6416 732 6450 742
rect 6416 674 6450 694
rect 6416 660 6450 674
rect 6416 606 6450 622
rect 6416 588 6450 606
rect 6416 538 6450 550
rect 6416 516 6450 538
rect 6416 470 6450 478
rect 6416 444 6450 470
rect 6416 402 6450 406
rect 6416 372 6450 402
rect 6416 300 6450 334
rect 6416 232 6450 262
rect 6416 228 6450 232
rect 6416 164 6450 190
rect 6416 156 6450 164
rect 6416 96 6450 118
rect 6416 84 6450 96
rect 6416 28 6450 46
rect 6416 12 6450 28
rect 6572 948 6606 982
rect 6572 878 6606 910
rect 6572 876 6606 878
rect 6572 810 6606 838
rect 6572 804 6606 810
rect 6572 742 6606 766
rect 6572 732 6606 742
rect 6572 674 6606 694
rect 6572 660 6606 674
rect 6572 606 6606 622
rect 6572 588 6606 606
rect 6572 538 6606 550
rect 6572 516 6606 538
rect 6572 470 6606 478
rect 6572 444 6606 470
rect 6572 402 6606 406
rect 6572 372 6606 402
rect 6572 300 6606 334
rect 6572 232 6606 262
rect 6572 228 6606 232
rect 6572 164 6606 190
rect 6572 156 6606 164
rect 6572 96 6606 118
rect 6572 84 6606 96
rect 6572 28 6606 46
rect 6572 12 6606 28
rect 6696 948 6730 982
rect 6696 878 6730 910
rect 6696 876 6730 878
rect 6696 810 6730 838
rect 6696 804 6730 810
rect 6696 742 6730 766
rect 6696 732 6730 742
rect 6696 674 6730 694
rect 6696 660 6730 674
rect 6696 606 6730 622
rect 6696 588 6730 606
rect 6696 538 6730 550
rect 6696 516 6730 538
rect 6696 470 6730 478
rect 6696 444 6730 470
rect 6696 402 6730 406
rect 6696 372 6730 402
rect 6696 300 6730 334
rect 6696 232 6730 262
rect 6696 228 6730 232
rect 6696 164 6730 190
rect 6696 156 6730 164
rect 6696 96 6730 118
rect 6696 84 6730 96
rect 6696 28 6730 46
rect 6696 12 6730 28
rect 6852 948 6886 982
rect 6925 980 6959 1014
rect 7424 1023 7458 1029
rect 7424 995 7458 1023
rect 6852 878 6886 910
rect 6852 876 6886 878
rect 6852 810 6886 838
rect 6852 804 6886 810
rect 6852 742 6886 766
rect 6852 732 6886 742
rect 6852 674 6886 694
rect 6852 660 6886 674
rect 6852 606 6886 622
rect 6852 588 6886 606
rect 6852 538 6886 550
rect 6852 516 6886 538
rect 6852 470 6886 478
rect 6852 444 6886 470
rect 6852 402 6886 406
rect 6852 372 6886 402
rect 6852 300 6886 334
rect 6852 232 6886 262
rect 6852 228 6886 232
rect 6852 164 6886 190
rect 6852 156 6886 164
rect 6852 96 6886 118
rect 6852 84 6886 96
rect 6852 28 6886 46
rect 6852 12 6886 28
rect 7008 948 7042 982
rect 7008 878 7042 910
rect 7008 876 7042 878
rect 7008 810 7042 838
rect 7008 804 7042 810
rect 7008 742 7042 766
rect 7008 732 7042 742
rect 7008 674 7042 694
rect 7008 660 7042 674
rect 7008 606 7042 622
rect 7008 588 7042 606
rect 7008 538 7042 550
rect 7008 516 7042 538
rect 7008 470 7042 478
rect 7008 444 7042 470
rect 7008 402 7042 406
rect 7008 372 7042 402
rect 7008 300 7042 334
rect 7008 232 7042 262
rect 7008 228 7042 232
rect 7008 164 7042 190
rect 7008 156 7042 164
rect 7008 96 7042 118
rect 7008 84 7042 96
rect 7008 28 7042 46
rect 7008 12 7042 28
rect 7424 955 7458 957
rect 7424 923 7458 955
rect 7424 853 7458 885
rect 7424 851 7458 853
rect 7424 785 7458 813
rect 7424 779 7458 785
rect 7424 717 7458 741
rect 7424 707 7458 717
rect 7424 649 7458 669
rect 7424 635 7458 649
rect 7424 581 7458 597
rect 7424 563 7458 581
rect 7424 513 7458 525
rect 7424 491 7458 513
rect 7424 445 7458 453
rect 7424 419 7458 445
rect 7424 377 7458 381
rect 7424 347 7458 377
rect 7424 275 7458 309
rect 7424 207 7458 237
rect 7424 203 7458 207
rect 7424 139 7458 165
rect 7424 131 7458 139
rect 7424 71 7458 93
rect 7424 59 7458 71
rect 466 -41 500 -7
rect 466 -113 500 -79
rect 1427 -81 1461 -47
rect 1499 -81 1533 -47
rect 7424 3 7458 21
rect 7424 -13 7458 3
rect 7510 1355 7544 1389
rect 7510 1295 7544 1317
rect 7510 1283 7544 1295
rect 7510 1227 7544 1245
rect 7510 1211 7544 1227
rect 7510 1159 7544 1173
rect 7510 1139 7544 1159
rect 7510 1091 7544 1101
rect 7510 1067 7544 1091
rect 7510 1023 7544 1029
rect 7510 995 7544 1023
rect 7510 955 7544 957
rect 7510 923 7544 955
rect 7510 853 7544 885
rect 7510 851 7544 853
rect 7510 785 7544 813
rect 7510 779 7544 785
rect 7510 717 7544 741
rect 7510 707 7544 717
rect 7510 649 7544 669
rect 7510 635 7544 649
rect 7510 581 7544 597
rect 7510 563 7544 581
rect 7510 513 7544 525
rect 7510 491 7544 513
rect 7510 445 7544 453
rect 7510 419 7544 445
rect 7510 377 7544 381
rect 7510 347 7544 377
rect 7510 275 7544 309
rect 7510 207 7544 237
rect 7510 203 7544 207
rect 7510 139 7544 165
rect 7510 131 7544 139
rect 7510 71 7544 93
rect 7510 59 7544 71
rect 7510 3 7544 21
rect 7510 -13 7544 3
rect 7596 1355 7630 1389
rect 7596 1295 7630 1317
rect 7596 1283 7630 1295
rect 7596 1227 7630 1245
rect 7596 1211 7630 1227
rect 7596 1159 7630 1173
rect 7596 1139 7630 1159
rect 7596 1091 7630 1101
rect 7596 1067 7630 1091
rect 7596 1023 7630 1029
rect 7596 995 7630 1023
rect 7596 955 7630 957
rect 7596 923 7630 955
rect 7596 853 7630 885
rect 7596 851 7630 853
rect 7596 785 7630 813
rect 7596 779 7630 785
rect 7596 717 7630 741
rect 7596 707 7630 717
rect 7596 649 7630 669
rect 7596 635 7630 649
rect 7596 581 7630 597
rect 7596 563 7630 581
rect 7596 513 7630 525
rect 7596 491 7630 513
rect 7596 445 7630 453
rect 7596 419 7630 445
rect 7596 377 7630 381
rect 7596 347 7630 377
rect 7596 275 7630 309
rect 7596 207 7630 237
rect 7596 203 7630 207
rect 7596 139 7630 165
rect 7596 131 7630 139
rect 7596 71 7630 93
rect 7596 59 7630 71
rect 7596 3 7630 21
rect 7596 -13 7630 3
rect 7682 1355 7716 1389
rect 7682 1295 7716 1317
rect 7682 1283 7716 1295
rect 7682 1227 7716 1245
rect 7682 1211 7716 1227
rect 7682 1159 7716 1173
rect 7682 1139 7716 1159
rect 7682 1091 7716 1101
rect 7682 1067 7716 1091
rect 7682 1023 7716 1029
rect 7682 995 7716 1023
rect 7682 955 7716 957
rect 7682 923 7716 955
rect 7682 853 7716 885
rect 7682 851 7716 853
rect 7682 785 7716 813
rect 7682 779 7716 785
rect 7682 717 7716 741
rect 7682 707 7716 717
rect 7682 649 7716 669
rect 7682 635 7716 649
rect 7682 581 7716 597
rect 7682 563 7716 581
rect 7682 513 7716 525
rect 7682 491 7716 513
rect 7682 445 7716 453
rect 7682 419 7716 445
rect 7682 377 7716 381
rect 7682 347 7716 377
rect 7682 275 7716 309
rect 7682 207 7716 237
rect 7682 203 7716 207
rect 7682 139 7716 165
rect 7682 131 7716 139
rect 7682 71 7716 93
rect 7682 59 7716 71
rect 7682 3 7716 21
rect 7682 -13 7716 3
rect 7768 1355 7802 1389
rect 7768 1295 7802 1317
rect 7768 1283 7802 1295
rect 7768 1227 7802 1245
rect 7768 1211 7802 1227
rect 7768 1159 7802 1173
rect 7768 1139 7802 1159
rect 7768 1091 7802 1101
rect 7768 1067 7802 1091
rect 7768 1023 7802 1029
rect 7768 995 7802 1023
rect 7768 955 7802 957
rect 7768 923 7802 955
rect 7768 853 7802 885
rect 7768 851 7802 853
rect 7768 785 7802 813
rect 7768 779 7802 785
rect 7768 717 7802 741
rect 7768 707 7802 717
rect 7768 649 7802 669
rect 7768 635 7802 649
rect 7768 581 7802 597
rect 7768 563 7802 581
rect 7768 513 7802 525
rect 7768 491 7802 513
rect 7768 445 7802 453
rect 7768 419 7802 445
rect 7768 377 7802 381
rect 7768 347 7802 377
rect 7768 275 7802 309
rect 7768 207 7802 237
rect 7768 203 7802 207
rect 7768 139 7802 165
rect 7768 131 7802 139
rect 7768 71 7802 93
rect 7768 59 7802 71
rect 7768 3 7802 21
rect 7768 -13 7802 3
rect 7854 1355 7888 1389
rect 7854 1295 7888 1317
rect 19973 1500 20007 1534
rect 25243 1496 25277 1530
rect 25315 1496 25349 1530
rect 19973 1422 20007 1456
rect 9483 1321 9513 1355
rect 9513 1321 9517 1355
rect 9556 1321 9581 1355
rect 9581 1321 9590 1355
rect 9629 1321 9649 1355
rect 9649 1321 9663 1355
rect 9702 1321 9717 1355
rect 9717 1321 9736 1355
rect 9775 1321 9785 1355
rect 9785 1321 9809 1355
rect 9848 1321 9853 1355
rect 9853 1321 9882 1355
rect 9921 1321 9955 1355
rect 9994 1321 10023 1355
rect 10023 1321 10028 1355
rect 10067 1321 10091 1355
rect 10091 1321 10101 1355
rect 10140 1321 10159 1355
rect 10159 1321 10174 1355
rect 10213 1321 10227 1355
rect 10227 1321 10247 1355
rect 10286 1321 10295 1355
rect 10295 1321 10320 1355
rect 10359 1321 10363 1355
rect 10363 1321 10393 1355
rect 10432 1321 10465 1355
rect 10465 1321 10466 1355
rect 10505 1321 10533 1355
rect 10533 1321 10539 1355
rect 10578 1321 10601 1355
rect 10601 1321 10612 1355
rect 10651 1321 10669 1355
rect 10669 1321 10685 1355
rect 10724 1321 10737 1355
rect 10737 1321 10758 1355
rect 10797 1321 10805 1355
rect 10805 1321 10831 1355
rect 10870 1321 10873 1355
rect 10873 1321 10904 1355
rect 10943 1321 10975 1355
rect 10975 1321 10977 1355
rect 11016 1321 11043 1355
rect 11043 1321 11050 1355
rect 11089 1321 11111 1355
rect 11111 1321 11123 1355
rect 11162 1321 11179 1355
rect 11179 1321 11196 1355
rect 11235 1321 11247 1355
rect 11247 1321 11269 1355
rect 11308 1321 11315 1355
rect 11315 1321 11342 1355
rect 11381 1321 11383 1355
rect 11383 1321 11415 1355
rect 11454 1321 11485 1355
rect 11485 1321 11488 1355
rect 11527 1321 11553 1355
rect 11553 1321 11561 1355
rect 11600 1321 11621 1355
rect 11621 1321 11634 1355
rect 11672 1321 11689 1355
rect 11689 1321 11706 1355
rect 11744 1321 11757 1355
rect 11757 1321 11778 1355
rect 11816 1321 11825 1355
rect 11825 1321 11850 1355
rect 11888 1321 11893 1355
rect 11893 1321 11922 1355
rect 11960 1321 11961 1355
rect 11961 1321 11994 1355
rect 12032 1321 12063 1355
rect 12063 1321 12066 1355
rect 12104 1321 12131 1355
rect 12131 1321 12138 1355
rect 12176 1321 12199 1355
rect 12199 1321 12210 1355
rect 12248 1321 12267 1355
rect 12267 1321 12282 1355
rect 12320 1321 12335 1355
rect 12335 1321 12354 1355
rect 13526 1321 13559 1355
rect 13559 1321 13560 1355
rect 13599 1321 13627 1355
rect 13627 1321 13633 1355
rect 13672 1321 13695 1355
rect 13695 1321 13706 1355
rect 13745 1321 13763 1355
rect 13763 1321 13779 1355
rect 13818 1321 13831 1355
rect 13831 1321 13852 1355
rect 13891 1321 13899 1355
rect 13899 1321 13925 1355
rect 13964 1321 13967 1355
rect 13967 1321 13998 1355
rect 14037 1321 14069 1355
rect 14069 1321 14071 1355
rect 14110 1321 14137 1355
rect 14137 1321 14144 1355
rect 14183 1321 14205 1355
rect 14205 1321 14217 1355
rect 14255 1321 14273 1355
rect 14273 1321 14289 1355
rect 14327 1321 14341 1355
rect 14341 1321 14361 1355
rect 14399 1321 14409 1355
rect 14409 1321 14433 1355
rect 14471 1321 14477 1355
rect 14477 1321 14505 1355
rect 14543 1321 14545 1355
rect 14545 1321 14577 1355
rect 14615 1321 14647 1355
rect 14647 1321 14649 1355
rect 14687 1321 14715 1355
rect 14715 1321 14721 1355
rect 14759 1321 14783 1355
rect 14783 1321 14793 1355
rect 14831 1321 14851 1355
rect 14851 1321 14865 1355
rect 14903 1321 14919 1355
rect 14919 1321 14937 1355
rect 14975 1321 14987 1355
rect 14987 1321 15009 1355
rect 15047 1321 15055 1355
rect 15055 1321 15081 1355
rect 15119 1321 15123 1355
rect 15123 1321 15153 1355
rect 15191 1321 15225 1355
rect 15263 1321 15293 1355
rect 15293 1321 15297 1355
rect 15335 1321 15361 1355
rect 15361 1321 15369 1355
rect 15407 1321 15429 1355
rect 15429 1321 15441 1355
rect 15479 1321 15497 1355
rect 15497 1321 15513 1355
rect 15551 1321 15565 1355
rect 15565 1321 15585 1355
rect 15623 1321 15633 1355
rect 15633 1321 15657 1355
rect 15695 1321 15701 1355
rect 15701 1321 15729 1355
rect 15767 1321 15769 1355
rect 15769 1321 15801 1355
rect 15839 1321 15871 1355
rect 15871 1321 15873 1355
rect 15911 1321 15939 1355
rect 15939 1321 15945 1355
rect 15983 1321 16007 1355
rect 16007 1321 16017 1355
rect 16055 1321 16075 1355
rect 16075 1321 16089 1355
rect 16127 1321 16143 1355
rect 16143 1321 16161 1355
rect 16199 1321 16211 1355
rect 16211 1321 16233 1355
rect 16271 1321 16279 1355
rect 16279 1321 16305 1355
rect 16343 1321 16347 1355
rect 16347 1321 16377 1355
rect 16415 1321 16449 1355
rect 16487 1321 16517 1355
rect 16517 1321 16521 1355
rect 16559 1321 16585 1355
rect 16585 1321 16593 1355
rect 16631 1321 16653 1355
rect 16653 1321 16665 1355
rect 16703 1321 16721 1355
rect 16721 1321 16737 1355
rect 16775 1321 16789 1355
rect 16789 1321 16809 1355
rect 16847 1321 16857 1355
rect 16857 1321 16881 1355
rect 16919 1321 16925 1355
rect 16925 1321 16953 1355
rect 16991 1321 16993 1355
rect 16993 1321 17025 1355
rect 17063 1321 17095 1355
rect 17095 1321 17097 1355
rect 17135 1321 17163 1355
rect 17163 1321 17169 1355
rect 17207 1321 17231 1355
rect 17231 1321 17241 1355
rect 17279 1321 17299 1355
rect 17299 1321 17313 1355
rect 17351 1321 17367 1355
rect 17367 1321 17385 1355
rect 17423 1321 17435 1355
rect 17435 1321 17457 1355
rect 17495 1321 17503 1355
rect 17503 1321 17529 1355
rect 17567 1321 17571 1355
rect 17571 1321 17601 1355
rect 17639 1321 17673 1355
rect 17711 1321 17741 1355
rect 17741 1321 17745 1355
rect 17783 1321 17809 1355
rect 17809 1321 17817 1355
rect 17855 1321 17877 1355
rect 17877 1321 17889 1355
rect 17927 1321 17945 1355
rect 17945 1321 17961 1355
rect 17999 1321 18013 1355
rect 18013 1321 18033 1355
rect 18071 1321 18081 1355
rect 18081 1321 18105 1355
rect 18143 1321 18149 1355
rect 18149 1321 18177 1355
rect 18215 1321 18217 1355
rect 18217 1321 18249 1355
rect 18287 1321 18319 1355
rect 18319 1321 18321 1355
rect 18359 1321 18387 1355
rect 18387 1321 18393 1355
rect 18431 1321 18455 1355
rect 18455 1321 18465 1355
rect 18503 1321 18523 1355
rect 18523 1321 18537 1355
rect 18575 1321 18591 1355
rect 18591 1321 18609 1355
rect 18647 1321 18659 1355
rect 18659 1321 18681 1355
rect 18719 1321 18727 1355
rect 18727 1321 18753 1355
rect 18791 1321 18795 1355
rect 18795 1321 18825 1355
rect 7854 1283 7888 1295
rect 7854 1227 7888 1245
rect 7854 1211 7888 1227
rect 7854 1159 7888 1173
rect 7854 1139 7888 1159
rect 18863 1248 18897 1250
rect 18863 1216 18897 1248
rect 19973 1344 20007 1378
rect 19973 1266 20007 1300
rect 20252 1428 20286 1433
rect 20252 1399 20286 1428
rect 20252 1310 20286 1325
rect 25243 1320 25277 1354
rect 25315 1320 25349 1354
rect 20252 1291 20286 1310
rect 19973 1188 20007 1222
rect 7854 1091 7888 1101
rect 7854 1067 7888 1091
rect 12868 1080 12902 1114
rect 15219 1101 15253 1135
rect 15411 1101 15445 1135
rect 15506 1101 15540 1135
rect 15644 1101 15678 1135
rect 15736 1101 15770 1135
rect 8352 1030 8386 1033
rect 8431 1030 8465 1033
rect 8510 1030 8544 1033
rect 8589 1030 8623 1033
rect 7854 1023 7888 1029
rect 7854 995 7888 1023
rect 8352 999 8379 1030
rect 8379 999 8386 1030
rect 8431 999 8450 1030
rect 8450 999 8465 1030
rect 8510 999 8521 1030
rect 8521 999 8544 1030
rect 8589 999 8593 1030
rect 8593 999 8623 1030
rect 8668 999 8702 1033
rect 8747 1030 8781 1033
rect 8825 1030 8859 1033
rect 12868 1030 12902 1042
rect 13072 1035 13088 1069
rect 13088 1035 13106 1069
rect 13144 1035 13156 1069
rect 13156 1035 13178 1069
rect 13216 1035 13224 1069
rect 13224 1035 13250 1069
rect 13288 1035 13292 1069
rect 13292 1035 13322 1069
rect 13360 1035 13394 1069
rect 13432 1035 13462 1069
rect 13462 1035 13466 1069
rect 13504 1035 13530 1069
rect 13530 1035 13538 1069
rect 13576 1035 13598 1069
rect 13598 1035 13610 1069
rect 13648 1035 13666 1069
rect 13666 1035 13682 1069
rect 13720 1035 13734 1069
rect 13734 1035 13754 1069
rect 13792 1035 13802 1069
rect 13802 1035 13826 1069
rect 13864 1035 13870 1069
rect 13870 1035 13898 1069
rect 13936 1035 13938 1069
rect 13938 1035 13970 1069
rect 14008 1035 14040 1069
rect 14040 1035 14042 1069
rect 14080 1035 14108 1069
rect 14108 1035 14114 1069
rect 14152 1035 14176 1069
rect 14176 1035 14186 1069
rect 14224 1035 14244 1069
rect 14244 1035 14258 1069
rect 14296 1035 14312 1069
rect 14312 1035 14330 1069
rect 14368 1035 14380 1069
rect 14380 1035 14402 1069
rect 14440 1035 14448 1069
rect 14448 1035 14474 1069
rect 14512 1035 14516 1069
rect 14516 1035 14546 1069
rect 14584 1035 14618 1069
rect 14656 1035 14686 1069
rect 14686 1035 14690 1069
rect 14728 1035 14754 1069
rect 14754 1035 14762 1069
rect 14800 1035 14822 1069
rect 14822 1035 14834 1069
rect 14872 1035 14890 1069
rect 14890 1035 14906 1069
rect 14944 1035 14958 1069
rect 14958 1035 14978 1069
rect 15016 1035 15026 1069
rect 15026 1035 15050 1069
rect 8747 999 8775 1030
rect 8775 999 8781 1030
rect 8825 999 8847 1030
rect 8847 999 8859 1030
rect 8967 996 8969 1030
rect 8969 996 9001 1030
rect 9041 996 9043 1030
rect 9043 996 9075 1030
rect 9115 996 9116 1030
rect 9116 996 9149 1030
rect 9189 996 9223 1030
rect 9263 996 9296 1030
rect 9296 996 9297 1030
rect 9337 996 9369 1030
rect 9369 996 9371 1030
rect 9411 996 9442 1030
rect 9442 996 9445 1030
rect 9485 996 9515 1030
rect 9515 996 9519 1030
rect 9558 996 9588 1030
rect 9588 996 9592 1030
rect 9631 996 9661 1030
rect 9661 996 9665 1030
rect 9745 996 9749 1030
rect 9749 996 9779 1030
rect 9819 996 9822 1030
rect 9822 996 9853 1030
rect 9893 996 9895 1030
rect 9895 996 9927 1030
rect 9967 996 9968 1030
rect 9968 996 10001 1030
rect 10041 996 10075 1030
rect 10116 996 10148 1030
rect 10148 996 10150 1030
rect 10191 996 10221 1030
rect 10221 996 10225 1030
rect 10266 996 10294 1030
rect 10294 996 10300 1030
rect 10341 996 10367 1030
rect 10367 996 10375 1030
rect 10416 996 10441 1030
rect 10441 996 10450 1030
rect 10604 977 10638 1011
rect 10805 996 10838 1030
rect 10838 996 10839 1030
rect 10877 996 10909 1030
rect 10909 996 10911 1030
rect 10949 996 10980 1030
rect 10980 996 10983 1030
rect 11021 996 11051 1030
rect 11051 996 11055 1030
rect 11093 996 11122 1030
rect 11122 996 11127 1030
rect 11165 996 11193 1030
rect 11193 996 11199 1030
rect 11237 996 11264 1030
rect 11264 996 11271 1030
rect 11309 996 11335 1030
rect 11335 996 11343 1030
rect 11381 996 11406 1030
rect 11406 996 11415 1030
rect 11453 996 11477 1030
rect 11477 996 11487 1030
rect 11525 996 11548 1030
rect 11548 996 11559 1030
rect 11597 996 11619 1030
rect 11619 996 11631 1030
rect 11669 996 11690 1030
rect 11690 996 11703 1030
rect 11741 996 11761 1030
rect 11761 996 11775 1030
rect 11813 996 11832 1030
rect 11832 996 11847 1030
rect 11885 996 11903 1030
rect 11903 996 11919 1030
rect 11957 996 11974 1030
rect 11974 996 11991 1030
rect 12029 996 12044 1030
rect 12044 996 12063 1030
rect 12101 996 12114 1030
rect 12114 996 12135 1030
rect 12173 996 12184 1030
rect 12184 996 12207 1030
rect 12245 996 12254 1030
rect 12254 996 12279 1030
rect 12868 1008 12878 1030
rect 12878 1008 12902 1030
rect 15122 1023 15156 1057
rect 7854 955 7888 957
rect 7854 923 7888 955
rect 7854 853 7888 885
rect 7854 851 7888 853
rect 7854 785 7888 813
rect 7854 779 7888 785
rect 7854 717 7888 741
rect 7854 707 7888 717
rect 7854 649 7888 669
rect 7854 635 7888 649
rect 7854 581 7888 597
rect 7854 563 7888 581
rect 7854 513 7888 525
rect 7854 491 7888 513
rect 7854 445 7888 453
rect 7854 419 7888 445
rect 7854 377 7888 381
rect 7854 347 7888 377
rect 7854 275 7888 309
rect 7854 207 7888 237
rect 7854 203 7888 207
rect 7854 139 7888 165
rect 7854 131 7888 139
rect 7854 71 7888 93
rect 7854 59 7888 71
rect 7854 3 7888 21
rect 7854 -13 7888 3
rect 10604 924 10638 936
rect 8177 908 8202 914
rect 8202 908 8211 914
rect 8177 880 8211 908
rect 8177 836 8202 838
rect 8202 836 8211 838
rect 8177 804 8211 836
rect 8177 728 8211 762
rect 8177 654 8211 686
rect 8177 652 8202 654
rect 8202 652 8211 654
rect 8177 582 8211 610
rect 8177 576 8202 582
rect 8202 576 8211 582
rect 8177 510 8211 533
rect 8177 499 8202 510
rect 8202 499 8211 510
rect 8177 438 8211 456
rect 8177 422 8202 438
rect 8202 422 8211 438
rect 8177 366 8211 379
rect 8177 345 8202 366
rect 8202 345 8211 366
rect 8177 294 8211 302
rect 8177 268 8202 294
rect 8202 268 8211 294
rect 8177 222 8211 225
rect 8177 191 8202 222
rect 8202 191 8211 222
rect 8177 116 8202 148
rect 8202 116 8211 148
rect 8177 114 8211 116
rect 8177 44 8202 71
rect 8202 44 8211 71
rect 8177 37 8211 44
rect 2151 -51 2185 -38
rect 2151 -72 2185 -51
rect 8177 -28 8202 -6
rect 8202 -28 8211 -6
rect 8177 -40 8211 -28
rect 8284 880 8318 914
rect 8284 810 8318 842
rect 8284 808 8318 810
rect 8284 742 8318 770
rect 8284 736 8318 742
rect 8284 674 8318 698
rect 8284 664 8318 674
rect 8284 606 8318 626
rect 8284 592 8318 606
rect 8284 538 8318 554
rect 8284 520 8318 538
rect 8284 470 8318 482
rect 8284 448 8318 470
rect 8284 402 8318 410
rect 8284 376 8318 402
rect 8284 334 8318 338
rect 8284 304 8318 334
rect 8284 232 8318 266
rect 8284 164 8318 194
rect 8284 160 8318 164
rect 8284 96 8318 122
rect 8284 88 8318 96
rect 8284 28 8318 50
rect 8284 16 8318 28
rect 8284 -40 8318 -22
rect 8284 -56 8318 -40
rect 8440 880 8474 914
rect 8440 810 8474 842
rect 8440 808 8474 810
rect 8440 742 8474 770
rect 8440 736 8474 742
rect 8440 674 8474 698
rect 8440 664 8474 674
rect 8440 606 8474 626
rect 8440 592 8474 606
rect 8440 538 8474 554
rect 8440 520 8474 538
rect 8440 470 8474 482
rect 8440 448 8474 470
rect 8440 402 8474 410
rect 8440 376 8474 402
rect 8440 334 8474 338
rect 8440 304 8474 334
rect 8440 232 8474 266
rect 8440 164 8474 194
rect 8440 160 8474 164
rect 8440 96 8474 122
rect 8440 88 8474 96
rect 8440 28 8474 50
rect 8440 16 8474 28
rect 8440 -40 8474 -22
rect 8440 -56 8474 -40
rect 8596 880 8630 914
rect 8596 810 8630 842
rect 8596 808 8630 810
rect 8596 742 8630 770
rect 8596 736 8630 742
rect 8596 674 8630 698
rect 8596 664 8630 674
rect 8596 606 8630 626
rect 8596 592 8630 606
rect 8596 538 8630 554
rect 8596 520 8630 538
rect 8596 470 8630 482
rect 8596 448 8630 470
rect 8596 402 8630 410
rect 8596 376 8630 402
rect 8596 334 8630 338
rect 8596 304 8630 334
rect 8596 232 8630 266
rect 8596 164 8630 194
rect 8596 160 8630 164
rect 8596 96 8630 122
rect 8596 88 8630 96
rect 8596 28 8630 50
rect 8596 16 8630 28
rect 8596 -40 8630 -22
rect 8596 -56 8630 -40
rect 8752 880 8786 914
rect 8752 810 8786 842
rect 8752 808 8786 810
rect 8752 742 8786 770
rect 8752 736 8786 742
rect 8752 674 8786 698
rect 8752 664 8786 674
rect 8752 606 8786 626
rect 8752 592 8786 606
rect 8752 538 8786 554
rect 8752 520 8786 538
rect 8752 470 8786 482
rect 8752 448 8786 470
rect 8752 402 8786 410
rect 8752 376 8786 402
rect 8752 334 8786 338
rect 8752 304 8786 334
rect 8752 232 8786 266
rect 8752 164 8786 194
rect 8752 160 8786 164
rect 8752 96 8786 122
rect 8752 88 8786 96
rect 8752 28 8786 50
rect 8752 16 8786 28
rect 8752 -40 8786 -22
rect 8752 -56 8786 -40
rect 8908 880 8942 914
rect 8908 810 8942 842
rect 8908 808 8942 810
rect 8908 742 8942 770
rect 8908 736 8942 742
rect 8908 674 8942 698
rect 8908 664 8942 674
rect 8908 606 8942 626
rect 8908 592 8942 606
rect 8908 538 8942 554
rect 8908 520 8942 538
rect 8908 470 8942 482
rect 8908 448 8942 470
rect 8908 402 8942 410
rect 8908 376 8942 402
rect 8908 334 8942 338
rect 8908 304 8942 334
rect 8908 232 8942 266
rect 8908 164 8942 194
rect 8908 160 8942 164
rect 8908 96 8942 122
rect 8908 88 8942 96
rect 8908 28 8942 50
rect 8908 16 8942 28
rect 8908 -40 8942 -22
rect 8908 -56 8942 -40
rect 9064 880 9098 914
rect 9064 810 9098 842
rect 9064 808 9098 810
rect 9064 742 9098 770
rect 9064 736 9098 742
rect 9064 674 9098 698
rect 9064 664 9098 674
rect 9064 606 9098 626
rect 9064 592 9098 606
rect 9064 538 9098 554
rect 9064 520 9098 538
rect 9064 470 9098 482
rect 9064 448 9098 470
rect 9064 402 9098 410
rect 9064 376 9098 402
rect 9064 334 9098 338
rect 9064 304 9098 334
rect 9064 232 9098 266
rect 9064 164 9098 194
rect 9064 160 9098 164
rect 9064 96 9098 122
rect 9064 88 9098 96
rect 9064 28 9098 50
rect 9064 16 9098 28
rect 9064 -40 9098 -22
rect 9064 -56 9098 -40
rect 9220 880 9254 914
rect 9220 810 9254 842
rect 9220 808 9254 810
rect 9220 742 9254 770
rect 9220 736 9254 742
rect 9220 674 9254 698
rect 9220 664 9254 674
rect 9220 606 9254 626
rect 9220 592 9254 606
rect 9220 538 9254 554
rect 9220 520 9254 538
rect 9220 470 9254 482
rect 9220 448 9254 470
rect 9220 402 9254 410
rect 9220 376 9254 402
rect 9220 334 9254 338
rect 9220 304 9254 334
rect 9220 232 9254 266
rect 9220 164 9254 194
rect 9220 160 9254 164
rect 9220 96 9254 122
rect 9220 88 9254 96
rect 9220 28 9254 50
rect 9220 16 9254 28
rect 9220 -40 9254 -22
rect 9220 -56 9254 -40
rect 9376 880 9410 914
rect 9376 810 9410 842
rect 9376 808 9410 810
rect 9376 742 9410 770
rect 9376 736 9410 742
rect 9376 674 9410 698
rect 9376 664 9410 674
rect 9376 606 9410 626
rect 9376 592 9410 606
rect 9376 538 9410 554
rect 9376 520 9410 538
rect 9376 470 9410 482
rect 9376 448 9410 470
rect 9376 402 9410 410
rect 9376 376 9410 402
rect 9376 334 9410 338
rect 9376 304 9410 334
rect 9376 232 9410 266
rect 9376 164 9410 194
rect 9376 160 9410 164
rect 9376 96 9410 122
rect 9376 88 9410 96
rect 9376 28 9410 50
rect 9376 16 9410 28
rect 9376 -40 9410 -22
rect 9376 -56 9410 -40
rect 9532 880 9566 914
rect 9532 810 9566 842
rect 9532 808 9566 810
rect 9532 742 9566 770
rect 9532 736 9566 742
rect 9532 674 9566 698
rect 9532 664 9566 674
rect 9532 606 9566 626
rect 9532 592 9566 606
rect 9532 538 9566 554
rect 9532 520 9566 538
rect 9532 470 9566 482
rect 9532 448 9566 470
rect 9532 402 9566 410
rect 9532 376 9566 402
rect 9532 334 9566 338
rect 9532 304 9566 334
rect 9532 232 9566 266
rect 9532 164 9566 194
rect 9532 160 9566 164
rect 9532 96 9566 122
rect 9532 88 9566 96
rect 9532 28 9566 50
rect 9532 16 9566 28
rect 9532 -40 9566 -22
rect 9532 -56 9566 -40
rect 9688 880 9722 914
rect 9688 810 9722 842
rect 9688 808 9722 810
rect 9688 742 9722 770
rect 9688 736 9722 742
rect 9688 674 9722 698
rect 9688 664 9722 674
rect 9688 606 9722 626
rect 9688 592 9722 606
rect 9688 538 9722 554
rect 9688 520 9722 538
rect 9688 470 9722 482
rect 9688 448 9722 470
rect 9688 402 9722 410
rect 9688 376 9722 402
rect 9688 334 9722 338
rect 9688 304 9722 334
rect 9688 232 9722 266
rect 9688 164 9722 194
rect 9688 160 9722 164
rect 9688 96 9722 122
rect 9688 88 9722 96
rect 9688 28 9722 50
rect 9688 16 9722 28
rect 9688 -40 9722 -22
rect 9688 -56 9722 -40
rect 9844 880 9878 914
rect 9844 810 9878 842
rect 9844 808 9878 810
rect 9844 742 9878 770
rect 9844 736 9878 742
rect 9844 674 9878 698
rect 9844 664 9878 674
rect 9844 606 9878 626
rect 9844 592 9878 606
rect 9844 538 9878 554
rect 9844 520 9878 538
rect 9844 470 9878 482
rect 9844 448 9878 470
rect 9844 402 9878 410
rect 9844 376 9878 402
rect 9844 334 9878 338
rect 9844 304 9878 334
rect 9844 232 9878 266
rect 9844 164 9878 194
rect 9844 160 9878 164
rect 9844 96 9878 122
rect 9844 88 9878 96
rect 9844 28 9878 50
rect 9844 16 9878 28
rect 9844 -40 9878 -22
rect 9844 -56 9878 -40
rect 10000 880 10034 914
rect 10000 810 10034 842
rect 10000 808 10034 810
rect 10000 742 10034 770
rect 10000 736 10034 742
rect 10000 674 10034 698
rect 10000 664 10034 674
rect 10000 606 10034 626
rect 10000 592 10034 606
rect 10000 538 10034 554
rect 10000 520 10034 538
rect 10000 470 10034 482
rect 10000 448 10034 470
rect 10000 402 10034 410
rect 10000 376 10034 402
rect 10000 334 10034 338
rect 10000 304 10034 334
rect 10000 232 10034 266
rect 10000 164 10034 194
rect 10000 160 10034 164
rect 10000 96 10034 122
rect 10000 88 10034 96
rect 10000 28 10034 50
rect 10000 16 10034 28
rect 10000 -40 10034 -22
rect 10000 -56 10034 -40
rect 10156 880 10190 914
rect 10156 810 10190 842
rect 10156 808 10190 810
rect 10156 742 10190 770
rect 10156 736 10190 742
rect 10156 674 10190 698
rect 10156 664 10190 674
rect 10156 606 10190 626
rect 10156 592 10190 606
rect 10156 538 10190 554
rect 10156 520 10190 538
rect 10156 470 10190 482
rect 10156 448 10190 470
rect 10156 402 10190 410
rect 10156 376 10190 402
rect 10156 334 10190 338
rect 10156 304 10190 334
rect 10156 232 10190 266
rect 10156 164 10190 194
rect 10156 160 10190 164
rect 10156 96 10190 122
rect 10156 88 10190 96
rect 10156 28 10190 50
rect 10156 16 10190 28
rect 10156 -40 10190 -22
rect 10156 -56 10190 -40
rect 10312 880 10346 914
rect 10312 810 10346 842
rect 10312 808 10346 810
rect 10312 742 10346 770
rect 10312 736 10346 742
rect 10312 674 10346 698
rect 10312 664 10346 674
rect 10312 606 10346 626
rect 10312 592 10346 606
rect 10312 538 10346 554
rect 10312 520 10346 538
rect 10312 470 10346 482
rect 10312 448 10346 470
rect 10312 402 10346 410
rect 10312 376 10346 402
rect 10312 334 10346 338
rect 10312 304 10346 334
rect 10312 232 10346 266
rect 10312 164 10346 194
rect 10312 160 10346 164
rect 10312 96 10346 122
rect 10312 88 10346 96
rect 10312 28 10346 50
rect 10312 16 10346 28
rect 10312 -40 10346 -22
rect 10312 -56 10346 -40
rect 10468 880 10502 914
rect 10468 810 10502 842
rect 10468 808 10502 810
rect 10468 742 10502 770
rect 10468 736 10502 742
rect 10468 674 10502 698
rect 10468 664 10502 674
rect 10468 606 10502 626
rect 10468 592 10502 606
rect 10468 538 10502 554
rect 10468 520 10502 538
rect 10468 470 10502 482
rect 10468 448 10502 470
rect 10468 402 10502 410
rect 10468 376 10502 402
rect 10468 334 10502 338
rect 10468 304 10502 334
rect 10468 232 10502 266
rect 10468 164 10502 194
rect 10468 160 10502 164
rect 10468 96 10502 122
rect 10468 88 10502 96
rect 10468 28 10502 50
rect 10468 16 10502 28
rect 10468 -40 10502 -22
rect 10468 -56 10502 -40
rect 10604 902 10638 924
rect 10604 854 10638 861
rect 10604 827 10638 854
rect 10604 784 10638 786
rect 10604 752 10638 784
rect 10604 680 10638 710
rect 10604 676 10638 680
rect 10604 610 10638 634
rect 10604 600 10638 610
rect 10604 540 10638 558
rect 10604 524 10638 540
rect 10604 469 10638 482
rect 10604 448 10638 469
rect 10604 398 10638 406
rect 10604 372 10638 398
rect 10604 327 10638 330
rect 10604 296 10638 327
rect 10604 220 10638 254
rect 10604 148 10638 178
rect 10604 144 10638 148
rect 10604 77 10638 102
rect 10604 68 10638 77
rect 10604 6 10638 26
rect 10604 -8 10638 6
rect 466 -185 500 -151
rect 570 -159 586 -125
rect 586 -159 604 -125
rect 642 -159 654 -125
rect 654 -159 676 -125
rect 714 -159 722 -125
rect 722 -159 748 -125
rect 786 -159 790 -125
rect 790 -159 820 -125
rect 858 -159 892 -125
rect 930 -159 960 -125
rect 960 -159 964 -125
rect 1002 -159 1028 -125
rect 1028 -159 1036 -125
rect 1074 -159 1096 -125
rect 1096 -159 1108 -125
rect 1146 -159 1164 -125
rect 1164 -159 1180 -125
rect 1218 -159 1232 -125
rect 1232 -159 1252 -125
rect 1290 -159 1300 -125
rect 1300 -159 1324 -125
rect 1362 -159 1368 -125
rect 1368 -159 1396 -125
rect 1434 -159 1436 -125
rect 1436 -159 1468 -125
rect 1506 -159 1540 -125
rect 2151 -119 2185 -112
rect 2151 -146 2185 -119
rect 2410 -92 2422 -58
rect 2422 -92 2444 -58
rect 2483 -92 2491 -58
rect 2491 -92 2517 -58
rect 2556 -92 2560 -58
rect 2560 -92 2590 -58
rect 2629 -92 2663 -58
rect 2702 -92 2732 -58
rect 2732 -92 2736 -58
rect 2775 -92 2801 -58
rect 2801 -92 2809 -58
rect 2848 -92 2870 -58
rect 2870 -92 2882 -58
rect 2921 -92 2939 -58
rect 2939 -92 2955 -58
rect 2994 -92 3008 -58
rect 3008 -92 3028 -58
rect 3067 -92 3077 -58
rect 3077 -92 3101 -58
rect 3140 -92 3146 -58
rect 3146 -92 3174 -58
rect 3213 -92 3215 -58
rect 3215 -92 3247 -58
rect 3286 -92 3319 -58
rect 3319 -92 3320 -58
rect 3359 -92 3388 -58
rect 3388 -92 3393 -58
rect 3432 -92 3457 -58
rect 3457 -92 3466 -58
rect 3505 -92 3526 -58
rect 3526 -92 3539 -58
rect 3578 -92 3595 -58
rect 3595 -92 3612 -58
rect 3651 -92 3664 -58
rect 3664 -92 3685 -58
rect 3724 -92 3733 -58
rect 3733 -92 3758 -58
rect 3797 -92 3802 -58
rect 3802 -92 3831 -58
rect 3870 -92 3871 -58
rect 3871 -92 3904 -58
rect 3943 -92 3974 -58
rect 3974 -92 3977 -58
rect 4016 -92 4042 -58
rect 4042 -92 4050 -58
rect 4089 -92 4110 -58
rect 4110 -92 4123 -58
rect 4161 -92 4178 -58
rect 4178 -92 4195 -58
rect 4233 -92 4246 -58
rect 4246 -92 4267 -58
rect 4305 -92 4314 -58
rect 4314 -92 4339 -58
rect 4377 -92 4382 -58
rect 4382 -92 4411 -58
rect 4449 -92 4450 -58
rect 4450 -92 4483 -58
rect 4521 -92 4552 -58
rect 4552 -92 4555 -58
rect 4593 -92 4620 -58
rect 4620 -92 4627 -58
rect 4665 -92 4688 -58
rect 4688 -92 4699 -58
rect 4737 -92 4756 -58
rect 4756 -92 4771 -58
rect 4809 -92 4824 -58
rect 4824 -92 4843 -58
rect 4881 -92 4892 -58
rect 4892 -92 4915 -58
rect 4953 -92 4960 -58
rect 4960 -92 4987 -58
rect 5025 -92 5028 -58
rect 5028 -92 5059 -58
rect 5097 -92 5130 -58
rect 5130 -92 5131 -58
rect 5169 -92 5198 -58
rect 5198 -92 5203 -58
rect 5241 -92 5266 -58
rect 5266 -92 5275 -58
rect 5313 -92 5334 -58
rect 5334 -92 5347 -58
rect 5385 -92 5402 -58
rect 5402 -92 5419 -58
rect 5457 -92 5470 -58
rect 5470 -92 5491 -58
rect 5529 -92 5538 -58
rect 5538 -92 5563 -58
rect 5601 -92 5606 -58
rect 5606 -92 5635 -58
rect 5686 -92 5708 -58
rect 5708 -92 5720 -58
rect 5760 -92 5776 -58
rect 5776 -92 5794 -58
rect 5834 -92 5844 -58
rect 5844 -92 5868 -58
rect 5908 -92 5912 -58
rect 5912 -92 5942 -58
rect 5982 -92 6014 -58
rect 6014 -92 6016 -58
rect 6056 -92 6082 -58
rect 6082 -92 6090 -58
rect 6129 -92 6150 -58
rect 6150 -92 6163 -58
rect 6202 -92 6218 -58
rect 6218 -92 6236 -58
rect 6275 -92 6286 -58
rect 6286 -92 6309 -58
rect 6348 -92 6354 -58
rect 6354 -92 6382 -58
rect 6421 -92 6422 -58
rect 6422 -92 6455 -58
rect 6494 -92 6524 -58
rect 6524 -92 6528 -58
rect 6567 -92 6592 -58
rect 6592 -92 6601 -58
rect 6640 -92 6660 -58
rect 6660 -92 6674 -58
rect 6713 -92 6728 -58
rect 6728 -92 6747 -58
rect 6786 -92 6796 -58
rect 6796 -92 6820 -58
rect 6859 -92 6864 -58
rect 6864 -92 6893 -58
rect 10604 -84 10638 -50
rect 10737 880 10771 914
rect 10737 810 10771 842
rect 10737 808 10771 810
rect 10737 742 10771 770
rect 10737 736 10771 742
rect 10737 674 10771 698
rect 10737 664 10771 674
rect 10737 606 10771 626
rect 10737 592 10771 606
rect 10737 538 10771 554
rect 10737 520 10771 538
rect 10737 470 10771 482
rect 10737 448 10771 470
rect 10737 402 10771 410
rect 10737 376 10771 402
rect 10737 334 10771 338
rect 10737 304 10771 334
rect 10737 232 10771 266
rect 10737 164 10771 194
rect 10737 160 10771 164
rect 10737 96 10771 122
rect 10737 88 10771 96
rect 10737 28 10771 50
rect 10737 16 10771 28
rect 10737 -40 10771 -22
rect 10737 -56 10771 -40
rect 11193 880 11227 914
rect 11193 810 11227 842
rect 11193 808 11227 810
rect 11193 742 11227 770
rect 11193 736 11227 742
rect 11193 674 11227 698
rect 11193 664 11227 674
rect 11193 606 11227 626
rect 11193 592 11227 606
rect 11193 538 11227 554
rect 11193 520 11227 538
rect 11193 470 11227 482
rect 11193 448 11227 470
rect 11193 402 11227 410
rect 11193 376 11227 402
rect 11193 334 11227 338
rect 11193 304 11227 334
rect 11193 232 11227 266
rect 11193 164 11227 194
rect 11193 160 11227 164
rect 11193 96 11227 122
rect 11193 88 11227 96
rect 11193 28 11227 50
rect 11193 16 11227 28
rect 11193 -40 11227 -22
rect 11193 -56 11227 -40
rect 11649 880 11683 914
rect 11649 810 11683 842
rect 11649 808 11683 810
rect 11649 742 11683 770
rect 11649 736 11683 742
rect 11649 674 11683 698
rect 11649 664 11683 674
rect 11649 606 11683 626
rect 11649 592 11683 606
rect 11649 538 11683 554
rect 11649 520 11683 538
rect 11649 470 11683 482
rect 11649 448 11683 470
rect 11649 402 11683 410
rect 11649 376 11683 402
rect 11649 334 11683 338
rect 11649 304 11683 334
rect 11649 232 11683 266
rect 11649 164 11683 194
rect 11649 160 11683 164
rect 11649 96 11683 122
rect 11649 88 11683 96
rect 11649 28 11683 50
rect 11649 16 11683 28
rect 11649 -40 11683 -22
rect 11649 -56 11683 -40
rect 12105 880 12139 914
rect 12105 810 12139 842
rect 12105 808 12139 810
rect 12105 742 12139 770
rect 12105 736 12139 742
rect 12105 674 12139 698
rect 12105 664 12139 674
rect 12105 606 12139 626
rect 12105 592 12139 606
rect 12105 538 12139 554
rect 12105 520 12139 538
rect 12105 470 12139 482
rect 12105 448 12139 470
rect 12105 402 12139 410
rect 12105 376 12139 402
rect 12105 334 12139 338
rect 12105 304 12139 334
rect 12105 232 12139 266
rect 12105 164 12139 194
rect 12105 160 12139 164
rect 12105 96 12139 122
rect 12105 88 12139 96
rect 12105 28 12139 50
rect 12105 16 12139 28
rect 12105 -40 12139 -22
rect 12105 -56 12139 -40
rect 12561 880 12595 914
rect 12561 810 12595 842
rect 12561 808 12595 810
rect 12561 742 12595 770
rect 12783 896 12817 927
rect 12783 893 12817 896
rect 12783 794 12817 805
rect 12783 771 12817 794
rect 12959 896 12993 927
rect 12959 893 12993 896
rect 15122 974 15124 979
rect 15124 974 15156 979
rect 15122 945 15156 974
rect 15122 872 15156 901
rect 15122 867 15124 872
rect 15124 867 15156 872
rect 12959 794 12993 805
rect 13072 799 13088 833
rect 13088 799 13106 833
rect 13144 799 13156 833
rect 13156 799 13178 833
rect 13216 799 13224 833
rect 13224 799 13250 833
rect 13288 799 13292 833
rect 13292 799 13322 833
rect 13360 799 13394 833
rect 13432 799 13462 833
rect 13462 799 13466 833
rect 13504 799 13530 833
rect 13530 799 13538 833
rect 13576 799 13598 833
rect 13598 799 13610 833
rect 13648 799 13666 833
rect 13666 799 13682 833
rect 13720 799 13734 833
rect 13734 799 13754 833
rect 13792 799 13802 833
rect 13802 799 13826 833
rect 13864 799 13870 833
rect 13870 799 13898 833
rect 13936 799 13938 833
rect 13938 799 13970 833
rect 14008 799 14040 833
rect 14040 799 14042 833
rect 14080 799 14108 833
rect 14108 799 14114 833
rect 14152 799 14176 833
rect 14176 799 14186 833
rect 14224 799 14244 833
rect 14244 799 14258 833
rect 14296 799 14312 833
rect 14312 799 14330 833
rect 14368 799 14380 833
rect 14380 799 14402 833
rect 14440 799 14448 833
rect 14448 799 14474 833
rect 14512 799 14516 833
rect 14516 799 14546 833
rect 14584 799 14618 833
rect 14656 799 14686 833
rect 14686 799 14690 833
rect 14728 799 14754 833
rect 14754 799 14762 833
rect 14800 799 14822 833
rect 14822 799 14834 833
rect 14872 799 14890 833
rect 14890 799 14906 833
rect 14944 799 14958 833
rect 14958 799 14978 833
rect 15016 799 15026 833
rect 15026 799 15050 833
rect 15223 1022 15257 1038
rect 15223 1004 15257 1022
rect 15223 954 15257 966
rect 15223 932 15257 954
rect 15223 886 15257 894
rect 15223 860 15257 886
rect 15317 1029 15351 1063
rect 15317 949 15351 983
rect 15317 869 15351 903
rect 12959 771 12993 794
rect 15122 804 15156 823
rect 15122 789 15124 804
rect 15124 789 15156 804
rect 15459 1022 15493 1038
rect 15459 1004 15493 1022
rect 15459 954 15493 966
rect 15459 932 15493 954
rect 15459 886 15493 894
rect 15459 860 15493 886
rect 15572 1024 15606 1058
rect 15572 947 15606 981
rect 15572 870 15606 904
rect 15317 789 15351 823
rect 15695 1022 15729 1038
rect 15695 1004 15729 1022
rect 15695 954 15729 966
rect 15695 932 15729 954
rect 15695 886 15729 894
rect 15695 860 15729 886
rect 15827 1029 15861 1063
rect 15827 954 15861 988
rect 15827 879 15861 913
rect 15572 792 15606 826
rect 15827 805 15861 839
rect 15931 1022 15965 1038
rect 15931 1004 15965 1022
rect 15931 954 15965 966
rect 15931 932 15965 954
rect 15931 886 15965 894
rect 15931 860 15965 886
rect 16049 1017 16083 1051
rect 16049 944 16083 978
rect 16049 871 16083 905
rect 16167 1022 16201 1038
rect 16167 1004 16201 1022
rect 16167 954 16201 966
rect 16167 932 16201 954
rect 16167 886 16201 894
rect 16167 860 16201 886
rect 16352 1061 16386 1073
rect 16352 1039 16386 1061
rect 16352 974 16386 999
rect 16352 965 16386 974
rect 16352 891 16386 925
rect 16049 798 16083 832
rect 16352 817 16386 851
rect 12561 736 12595 742
rect 12561 674 12595 698
rect 12561 664 12595 674
rect 15122 736 15156 745
rect 15572 744 15594 748
rect 15594 744 15606 748
rect 15827 744 15834 765
rect 15834 744 15861 765
rect 16049 744 16072 759
rect 16072 744 16083 759
rect 15122 711 15124 736
rect 15124 711 15156 736
rect 15317 709 15351 743
rect 12561 606 12595 626
rect 12561 592 12595 606
rect 12561 538 12595 554
rect 12561 520 12595 538
rect 12561 470 12595 482
rect 12561 448 12595 470
rect 12561 402 12595 410
rect 12561 376 12595 402
rect 12561 334 12595 338
rect 12561 304 12595 334
rect 12561 232 12595 266
rect 12561 164 12595 194
rect 12561 160 12595 164
rect 12561 96 12595 122
rect 12561 88 12595 96
rect 12561 28 12595 50
rect 12561 16 12595 28
rect 12561 -40 12595 -22
rect 12561 -56 12595 -40
rect 12678 620 12712 636
rect 12678 602 12712 620
rect 15122 634 15124 667
rect 15124 634 15156 667
rect 15122 633 15156 634
rect 13072 563 13088 597
rect 13088 563 13106 597
rect 13144 563 13156 597
rect 13156 563 13178 597
rect 13216 563 13224 597
rect 13224 563 13250 597
rect 13288 563 13292 597
rect 13292 563 13322 597
rect 13360 563 13394 597
rect 13432 563 13462 597
rect 13462 563 13466 597
rect 13504 563 13530 597
rect 13530 563 13538 597
rect 13576 563 13598 597
rect 13598 563 13610 597
rect 13648 563 13666 597
rect 13666 563 13682 597
rect 13720 563 13734 597
rect 13734 563 13754 597
rect 13792 563 13802 597
rect 13802 563 13826 597
rect 13864 563 13870 597
rect 13870 563 13898 597
rect 13936 563 13938 597
rect 13938 563 13970 597
rect 14008 563 14040 597
rect 14040 563 14042 597
rect 14080 563 14108 597
rect 14108 563 14114 597
rect 14152 563 14176 597
rect 14176 563 14186 597
rect 14224 563 14244 597
rect 14244 563 14258 597
rect 14296 563 14312 597
rect 14312 563 14330 597
rect 14368 563 14380 597
rect 14380 563 14402 597
rect 14440 563 14448 597
rect 14448 563 14474 597
rect 14512 563 14516 597
rect 14516 563 14546 597
rect 14584 563 14618 597
rect 14656 563 14686 597
rect 14686 563 14690 597
rect 14728 563 14754 597
rect 14754 563 14762 597
rect 14800 563 14822 597
rect 14822 563 14834 597
rect 14872 563 14890 597
rect 14890 563 14906 597
rect 14944 563 14958 597
rect 14958 563 14978 597
rect 15016 563 15026 597
rect 15026 563 15050 597
rect 12678 547 12712 560
rect 12678 526 12712 547
rect 15122 565 15124 589
rect 15124 565 15156 589
rect 15122 555 15156 565
rect 12678 474 12712 484
rect 12678 450 12712 474
rect 12678 401 12712 408
rect 12816 482 12850 516
rect 12889 482 12923 516
rect 12816 410 12850 444
rect 12889 410 12923 444
rect 12962 410 15084 516
rect 15122 496 15124 511
rect 15124 496 15156 511
rect 15122 477 15156 496
rect 15223 627 15257 653
rect 15223 619 15257 627
rect 15223 559 15257 581
rect 15223 547 15257 559
rect 15223 491 15257 509
rect 15223 475 15257 491
rect 15572 714 15606 744
rect 15317 629 15351 663
rect 15317 550 15351 584
rect 15122 427 15124 433
rect 15124 427 15156 433
rect 12678 374 12712 401
rect 15122 399 15156 427
rect 15317 471 15351 505
rect 15459 627 15493 653
rect 15459 619 15493 627
rect 15459 559 15493 581
rect 15459 547 15493 559
rect 15459 491 15493 509
rect 15459 475 15493 491
rect 15827 731 15861 744
rect 15572 636 15606 670
rect 15572 558 15606 592
rect 15572 480 15606 514
rect 15317 398 15351 426
rect 15695 627 15729 653
rect 15695 619 15729 627
rect 15695 559 15729 581
rect 15695 547 15729 559
rect 15695 491 15729 509
rect 15695 475 15729 491
rect 15827 657 15861 691
rect 16049 725 16083 744
rect 15827 583 15861 617
rect 15827 509 15861 543
rect 15572 402 15606 436
rect 15931 627 15965 653
rect 15931 619 15965 627
rect 15931 559 15965 581
rect 15931 547 15965 559
rect 15931 491 15965 509
rect 15931 475 15965 491
rect 16049 652 16083 686
rect 16352 766 16386 777
rect 16352 743 16386 766
rect 16049 579 16083 613
rect 16049 506 16083 540
rect 15827 435 15861 469
rect 16167 627 16201 653
rect 16167 619 16201 627
rect 16167 559 16201 581
rect 16167 547 16201 559
rect 16167 491 16201 509
rect 16167 475 16201 491
rect 16352 679 16386 703
rect 16352 669 16386 679
rect 16352 626 16386 629
rect 16352 595 16386 626
rect 16352 539 16386 555
rect 16352 521 16386 539
rect 16049 433 16083 467
rect 16352 452 16386 481
rect 16352 447 16386 452
rect 15317 392 15318 398
rect 15318 392 15351 398
rect 12678 328 12712 332
rect 12678 298 12712 328
rect 13072 327 13088 361
rect 13088 327 13106 361
rect 13144 327 13156 361
rect 13156 327 13178 361
rect 13216 327 13224 361
rect 13224 327 13250 361
rect 13288 327 13292 361
rect 13292 327 13322 361
rect 13360 327 13394 361
rect 13432 327 13462 361
rect 13462 327 13466 361
rect 13504 327 13530 361
rect 13530 327 13538 361
rect 13576 327 13598 361
rect 13598 327 13610 361
rect 13648 327 13666 361
rect 13666 327 13682 361
rect 13720 327 13734 361
rect 13734 327 13754 361
rect 13792 327 13802 361
rect 13802 327 13826 361
rect 13864 327 13870 361
rect 13870 327 13898 361
rect 13936 327 13938 361
rect 13938 327 13970 361
rect 14008 327 14040 361
rect 14040 327 14042 361
rect 14080 327 14108 361
rect 14108 327 14114 361
rect 14152 327 14176 361
rect 14176 327 14186 361
rect 14224 327 14244 361
rect 14244 327 14258 361
rect 14296 327 14312 361
rect 14312 327 14330 361
rect 14368 327 14380 361
rect 14380 327 14402 361
rect 14440 327 14448 361
rect 14448 327 14474 361
rect 14512 327 14516 361
rect 14516 327 14546 361
rect 14584 327 14618 361
rect 14656 327 14686 361
rect 14686 327 14690 361
rect 14728 327 14754 361
rect 14754 327 14762 361
rect 14800 327 14822 361
rect 14822 327 14834 361
rect 14872 327 14890 361
rect 14890 327 14906 361
rect 14944 327 14958 361
rect 14958 327 14978 361
rect 15016 327 15026 361
rect 15026 327 15050 361
rect 15899 364 15902 395
rect 15902 364 15933 395
rect 15974 364 16004 395
rect 16004 364 16008 395
rect 16352 373 16386 407
rect 12678 255 12712 256
rect 12678 222 12712 255
rect 15122 323 15156 354
rect 15122 320 15124 323
rect 15124 320 15156 323
rect 15899 361 15933 364
rect 15974 361 16008 364
rect 15572 324 15606 358
rect 15122 254 15156 275
rect 15122 241 15124 254
rect 15124 241 15156 254
rect 15223 282 15257 298
rect 15223 264 15257 282
rect 15223 214 15257 226
rect 12678 148 12712 180
rect 12678 146 12712 148
rect 15223 192 15257 214
rect 15223 146 15257 154
rect 12678 75 12712 104
rect 13072 91 13088 125
rect 13088 91 13106 125
rect 13144 91 13156 125
rect 13156 91 13178 125
rect 13216 91 13224 125
rect 13224 91 13250 125
rect 13288 91 13292 125
rect 13292 91 13322 125
rect 13360 91 13394 125
rect 13432 91 13462 125
rect 13462 91 13466 125
rect 13504 91 13530 125
rect 13530 91 13538 125
rect 13576 91 13598 125
rect 13598 91 13610 125
rect 13648 91 13666 125
rect 13666 91 13682 125
rect 13720 91 13734 125
rect 13734 91 13754 125
rect 13792 91 13802 125
rect 13802 91 13826 125
rect 13864 91 13870 125
rect 13870 91 13898 125
rect 13936 91 13938 125
rect 13938 91 13970 125
rect 14008 91 14040 125
rect 14040 91 14042 125
rect 14080 91 14108 125
rect 14108 91 14114 125
rect 14152 91 14176 125
rect 14176 91 14186 125
rect 14224 91 14244 125
rect 14244 91 14258 125
rect 14296 91 14312 125
rect 14312 91 14330 125
rect 14368 91 14380 125
rect 14380 91 14402 125
rect 14440 91 14448 125
rect 14448 91 14474 125
rect 14512 91 14516 125
rect 14516 91 14546 125
rect 14584 91 14618 125
rect 14656 91 14686 125
rect 14686 91 14690 125
rect 14728 91 14754 125
rect 14754 91 14762 125
rect 14800 91 14822 125
rect 14822 91 14834 125
rect 14872 91 14890 125
rect 14890 91 14906 125
rect 14944 91 14958 125
rect 14958 91 14978 125
rect 15016 91 15026 125
rect 15026 91 15050 125
rect 15223 120 15257 146
rect 15459 282 15493 298
rect 15459 264 15493 282
rect 15459 214 15493 226
rect 15459 192 15493 214
rect 16352 331 16386 333
rect 16352 299 16386 331
rect 18937 1110 18971 1144
rect 19011 1110 19045 1144
rect 19085 1110 19119 1144
rect 19159 1110 19193 1144
rect 19233 1110 19267 1144
rect 19307 1110 19341 1144
rect 19381 1110 19415 1144
rect 19455 1110 19489 1144
rect 19529 1110 19563 1144
rect 19603 1110 19637 1144
rect 19677 1110 19711 1144
rect 19751 1110 19785 1144
rect 19826 1110 19860 1144
rect 19901 1110 19935 1144
rect 18863 1044 18897 1072
rect 18863 1038 18897 1044
rect 18863 976 18897 995
rect 18863 961 18897 976
rect 18863 908 18897 918
rect 18863 884 18897 908
rect 18863 840 18897 842
rect 18863 808 18897 840
rect 18863 738 18897 766
rect 18863 732 18897 738
rect 18863 670 18897 690
rect 18863 656 18897 670
rect 18863 602 18897 614
rect 18863 580 18897 602
rect 18863 534 18897 538
rect 18863 504 18897 534
rect 18863 432 18897 462
rect 18863 428 18897 432
rect 18382 338 18416 341
rect 18454 338 18488 341
rect 18382 307 18414 338
rect 18414 307 18416 338
rect 18454 307 18482 338
rect 18482 307 18488 338
rect 18863 364 18897 386
rect 18863 352 18897 364
rect 15572 246 15606 280
rect 15572 168 15606 202
rect 15695 282 15729 298
rect 15695 264 15729 282
rect 15695 214 15729 226
rect 15911 225 15945 259
rect 15983 225 16013 259
rect 16013 225 16017 259
rect 16097 225 16101 259
rect 16101 225 16131 259
rect 16173 225 16203 259
rect 16203 225 16207 259
rect 16352 244 16386 259
rect 16352 225 16386 244
rect 18863 296 18897 310
rect 18863 276 18897 296
rect 15695 192 15729 214
rect 15459 146 15493 154
rect 15459 120 15493 146
rect 15695 146 15729 154
rect 15695 120 15729 146
rect 18647 223 18678 257
rect 18678 223 18681 257
rect 18719 223 18746 257
rect 18746 223 18753 257
rect 16352 157 16386 185
rect 16352 151 16386 157
rect 18863 228 18897 234
rect 18863 200 18897 228
rect 15884 109 15918 143
rect 12678 70 12712 75
rect 12678 2 12712 27
rect 12678 -7 12712 2
rect 15884 39 15918 71
rect 15884 37 15918 39
rect 15884 -29 15918 -1
rect 15884 -35 15918 -29
rect 13146 -37 13180 -36
rect 13219 -37 13253 -36
rect 13292 -37 13326 -36
rect 13365 -37 13399 -36
rect 13438 -37 13472 -36
rect 13511 -37 13545 -36
rect 13584 -37 13618 -36
rect 13657 -37 13691 -36
rect 13730 -37 13764 -36
rect 13803 -37 13837 -36
rect 13876 -37 13910 -36
rect 13949 -37 13983 -36
rect 14022 -37 14056 -36
rect 14095 -37 14129 -36
rect 14168 -37 14202 -36
rect 14241 -37 14275 -36
rect 14314 -37 14348 -36
rect 14387 -37 14421 -36
rect 14460 -37 14494 -36
rect 14533 -37 14567 -36
rect 14606 -37 14640 -36
rect 14679 -37 14713 -36
rect 14752 -37 14786 -36
rect 14825 -37 14859 -36
rect 14898 -37 14932 -36
rect 14971 -37 15005 -36
rect 15043 -37 15077 -36
rect 15115 -37 15149 -36
rect 15187 -37 15221 -36
rect 15259 -37 15293 -36
rect 15331 -37 15365 -36
rect 15403 -37 15437 -36
rect 15475 -37 15509 -36
rect 15547 -37 15581 -36
rect 15619 -37 15653 -36
rect 12678 -71 12712 -50
rect 13146 -70 13176 -37
rect 13176 -70 13180 -37
rect 13219 -70 13245 -37
rect 13245 -70 13253 -37
rect 13292 -70 13314 -37
rect 13314 -70 13326 -37
rect 13365 -70 13383 -37
rect 13383 -70 13399 -37
rect 13438 -70 13452 -37
rect 13452 -70 13472 -37
rect 13511 -70 13520 -37
rect 13520 -70 13545 -37
rect 13584 -70 13588 -37
rect 13588 -70 13618 -37
rect 13657 -70 13690 -37
rect 13690 -70 13691 -37
rect 13730 -70 13758 -37
rect 13758 -70 13764 -37
rect 13803 -70 13826 -37
rect 13826 -70 13837 -37
rect 13876 -70 13894 -37
rect 13894 -70 13910 -37
rect 13949 -70 13962 -37
rect 13962 -70 13983 -37
rect 14022 -70 14030 -37
rect 14030 -70 14056 -37
rect 14095 -70 14098 -37
rect 14098 -70 14129 -37
rect 14168 -70 14200 -37
rect 14200 -70 14202 -37
rect 14241 -70 14268 -37
rect 14268 -70 14275 -37
rect 14314 -70 14336 -37
rect 14336 -70 14348 -37
rect 14387 -70 14404 -37
rect 14404 -70 14421 -37
rect 14460 -70 14472 -37
rect 14472 -70 14494 -37
rect 14533 -70 14540 -37
rect 14540 -70 14567 -37
rect 14606 -70 14608 -37
rect 14608 -70 14640 -37
rect 14679 -70 14710 -37
rect 14710 -70 14713 -37
rect 14752 -70 14778 -37
rect 14778 -70 14786 -37
rect 14825 -70 14846 -37
rect 14846 -70 14859 -37
rect 14898 -70 14914 -37
rect 14914 -70 14932 -37
rect 14971 -70 14982 -37
rect 14982 -70 15005 -37
rect 15043 -70 15050 -37
rect 15050 -70 15077 -37
rect 15115 -70 15118 -37
rect 15118 -70 15149 -37
rect 15187 -70 15220 -37
rect 15220 -70 15221 -37
rect 15259 -70 15288 -37
rect 15288 -70 15293 -37
rect 15331 -70 15356 -37
rect 15356 -70 15365 -37
rect 15403 -70 15424 -37
rect 15424 -70 15437 -37
rect 15475 -70 15492 -37
rect 15492 -70 15509 -37
rect 15547 -70 15560 -37
rect 15560 -70 15581 -37
rect 15619 -70 15628 -37
rect 15628 -70 15653 -37
rect 15709 -71 15730 -69
rect 15730 -71 15743 -69
rect 12678 -84 12712 -71
rect 466 -257 500 -223
rect 1622 -220 1656 -200
rect 1622 -234 1656 -220
rect 466 -329 500 -295
rect 570 -315 586 -281
rect 586 -315 604 -281
rect 642 -315 654 -281
rect 654 -315 676 -281
rect 714 -315 722 -281
rect 722 -315 748 -281
rect 786 -315 790 -281
rect 790 -315 820 -281
rect 858 -315 892 -281
rect 930 -315 960 -281
rect 960 -315 964 -281
rect 1002 -315 1028 -281
rect 1028 -315 1036 -281
rect 1074 -315 1096 -281
rect 1096 -315 1108 -281
rect 1146 -315 1164 -281
rect 1164 -315 1180 -281
rect 1218 -315 1232 -281
rect 1232 -315 1252 -281
rect 1290 -315 1300 -281
rect 1300 -315 1324 -281
rect 1362 -315 1368 -281
rect 1368 -315 1396 -281
rect 1434 -315 1436 -281
rect 1436 -315 1468 -281
rect 1506 -315 1540 -281
rect 1622 -315 1656 -285
rect 466 -402 500 -368
rect 1622 -319 1656 -315
rect 1622 -376 1656 -371
rect 2151 -220 2185 -186
rect 2151 -268 2185 -260
rect 2151 -294 2185 -268
rect 15709 -103 15743 -71
rect 15781 -103 15815 -69
rect 15709 -176 15743 -142
rect 15781 -176 15815 -142
rect 15709 -249 15743 -215
rect 15781 -249 15815 -215
rect 15709 -322 15743 -288
rect 15781 -322 15815 -288
rect 2227 -360 2253 -332
rect 2253 -360 2261 -332
rect 2303 -360 2321 -332
rect 2321 -360 2337 -332
rect 2379 -360 2389 -332
rect 2389 -360 2413 -332
rect 2455 -360 2457 -332
rect 2457 -360 2489 -332
rect 2531 -360 2559 -332
rect 2559 -360 2565 -332
rect 2607 -360 2627 -332
rect 2627 -360 2641 -332
rect 2683 -360 2695 -332
rect 2695 -360 2717 -332
rect 2759 -360 2763 -332
rect 2763 -360 2793 -332
rect 2835 -360 2865 -332
rect 2865 -360 2869 -332
rect 2911 -360 2933 -332
rect 2933 -360 2945 -332
rect 2987 -360 3001 -332
rect 3001 -360 3021 -332
rect 3063 -360 3069 -332
rect 3069 -360 3097 -332
rect 3140 -360 3171 -332
rect 3171 -360 3174 -332
rect 3217 -360 3239 -332
rect 3239 -360 3251 -332
rect 3294 -360 3307 -332
rect 3307 -360 3328 -332
rect 2227 -366 2261 -360
rect 2303 -366 2337 -360
rect 2379 -366 2413 -360
rect 2455 -366 2489 -360
rect 2531 -366 2565 -360
rect 2607 -366 2641 -360
rect 2683 -366 2717 -360
rect 2759 -366 2793 -360
rect 2835 -366 2869 -360
rect 2911 -366 2945 -360
rect 2987 -366 3021 -360
rect 3063 -366 3097 -360
rect 3140 -366 3174 -360
rect 3217 -366 3251 -360
rect 3294 -366 3328 -360
rect 1622 -405 1656 -376
rect 466 -475 500 -441
rect 570 -471 586 -437
rect 586 -471 604 -437
rect 642 -471 654 -437
rect 654 -471 676 -437
rect 714 -471 722 -437
rect 722 -471 748 -437
rect 786 -471 790 -437
rect 790 -471 820 -437
rect 858 -471 892 -437
rect 930 -471 960 -437
rect 960 -471 964 -437
rect 1002 -471 1028 -437
rect 1028 -471 1036 -437
rect 1074 -471 1096 -437
rect 1096 -471 1108 -437
rect 1146 -471 1164 -437
rect 1164 -471 1180 -437
rect 1218 -471 1232 -437
rect 1232 -471 1252 -437
rect 1290 -471 1300 -437
rect 1300 -471 1324 -437
rect 1362 -471 1368 -437
rect 1368 -471 1396 -437
rect 1434 -471 1436 -437
rect 1436 -471 1468 -437
rect 1506 -471 1540 -437
rect 466 -548 500 -514
rect 1427 -549 1461 -515
rect 1499 -549 1533 -515
rect 1802 -565 1836 -531
rect 466 -621 500 -587
rect 570 -627 586 -593
rect 586 -627 604 -593
rect 642 -627 654 -593
rect 654 -627 676 -593
rect 714 -627 722 -593
rect 722 -627 748 -593
rect 786 -627 790 -593
rect 790 -627 820 -593
rect 858 -627 892 -593
rect 930 -627 960 -593
rect 960 -627 964 -593
rect 1002 -627 1028 -593
rect 1028 -627 1036 -593
rect 1074 -627 1096 -593
rect 1096 -627 1108 -593
rect 1146 -627 1164 -593
rect 1164 -627 1180 -593
rect 1218 -627 1232 -593
rect 1232 -627 1252 -593
rect 1290 -627 1300 -593
rect 1300 -627 1324 -593
rect 1362 -627 1368 -593
rect 1368 -627 1396 -593
rect 1434 -627 1436 -593
rect 1436 -627 1468 -593
rect 1506 -627 1540 -593
rect 1802 -637 1836 -603
rect 466 -694 500 -660
rect 466 -767 500 -733
rect 836 -783 858 -749
rect 858 -783 870 -749
rect 911 -783 926 -749
rect 926 -783 945 -749
rect 986 -783 994 -749
rect 994 -783 1020 -749
rect 1061 -783 1062 -749
rect 1062 -783 1095 -749
rect 1136 -783 1164 -749
rect 1164 -783 1170 -749
rect 1210 -783 1232 -749
rect 1232 -783 1244 -749
rect 1284 -783 1300 -749
rect 1300 -783 1318 -749
rect 1358 -783 1368 -749
rect 1368 -783 1392 -749
rect 1432 -783 1436 -749
rect 1436 -783 1466 -749
rect 1506 -783 1540 -749
rect 466 -840 500 -806
rect 466 -913 500 -879
rect 666 -917 668 -886
rect 668 -917 700 -886
rect 742 -917 772 -886
rect 772 -917 776 -886
rect 818 -917 842 -886
rect 842 -917 852 -886
rect 894 -917 912 -886
rect 912 -917 928 -886
rect 970 -917 982 -886
rect 982 -917 1004 -886
rect 1046 -917 1053 -886
rect 1053 -917 1080 -886
rect 1122 -917 1124 -886
rect 1124 -917 1156 -886
rect 666 -920 700 -917
rect 742 -920 776 -917
rect 818 -920 852 -917
rect 894 -920 928 -917
rect 970 -920 1004 -917
rect 1046 -920 1080 -917
rect 1122 -920 1156 -917
rect 1198 -920 1232 -886
rect 1274 -917 1303 -886
rect 1303 -917 1308 -886
rect 1350 -917 1374 -886
rect 1374 -917 1384 -886
rect 1426 -917 1445 -886
rect 1445 -917 1460 -886
rect 1502 -917 1516 -886
rect 1516 -917 1536 -886
rect 1274 -920 1308 -917
rect 1350 -920 1384 -917
rect 1426 -920 1460 -917
rect 1502 -920 1536 -917
rect 466 -986 500 -952
rect 466 -1059 500 -1025
rect 1103 -1068 1130 -1034
rect 1130 -1068 1137 -1034
rect 1183 -1068 1198 -1034
rect 1198 -1068 1217 -1034
rect 1263 -1068 1266 -1034
rect 1266 -1068 1297 -1034
rect 1343 -1068 1368 -1034
rect 1368 -1068 1377 -1034
rect 1423 -1068 1436 -1034
rect 1436 -1068 1457 -1034
rect 1503 -1068 1504 -1034
rect 1504 -1068 1537 -1034
rect 466 -1132 500 -1098
rect 466 -1205 500 -1171
rect 1622 -1129 1656 -1109
rect 1622 -1143 1656 -1129
rect 570 -1224 586 -1190
rect 586 -1224 604 -1190
rect 642 -1224 654 -1190
rect 654 -1224 676 -1190
rect 714 -1224 722 -1190
rect 722 -1224 748 -1190
rect 786 -1224 790 -1190
rect 790 -1224 820 -1190
rect 858 -1224 892 -1190
rect 930 -1224 960 -1190
rect 960 -1224 964 -1190
rect 1002 -1224 1028 -1190
rect 1028 -1224 1036 -1190
rect 1074 -1224 1096 -1190
rect 1096 -1224 1108 -1190
rect 1146 -1224 1164 -1190
rect 1164 -1224 1180 -1190
rect 1218 -1224 1232 -1190
rect 1232 -1224 1252 -1190
rect 1290 -1224 1300 -1190
rect 1300 -1224 1324 -1190
rect 1362 -1224 1368 -1190
rect 1368 -1224 1396 -1190
rect 1434 -1224 1436 -1190
rect 1436 -1224 1468 -1190
rect 1506 -1224 1540 -1190
rect 466 -1278 500 -1244
rect 466 -1351 500 -1317
rect 1622 -1265 1656 -1231
rect 15709 -395 15743 -361
rect 15781 -395 15815 -361
rect 15709 -468 15743 -434
rect 15781 -468 15815 -434
rect 15709 -541 15743 -507
rect 15781 -541 15815 -507
rect 15709 -614 15743 -580
rect 15781 -614 15815 -580
rect 15709 -687 15743 -653
rect 15781 -687 15815 -653
rect 15709 -761 15743 -727
rect 15781 -761 15815 -727
rect 15709 -835 15743 -801
rect 15781 -835 15815 -801
rect 15884 -97 15918 -73
rect 15884 -107 15918 -97
rect 15884 -165 15918 -145
rect 15884 -179 15918 -165
rect 15884 -233 15918 -217
rect 15884 -251 15918 -233
rect 15884 -301 15918 -289
rect 15884 -323 15918 -301
rect 15884 -369 15918 -361
rect 15884 -395 15918 -369
rect 15884 -437 15918 -433
rect 15884 -467 15918 -437
rect 15884 -539 15918 -505
rect 15884 -607 15918 -577
rect 15884 -611 15918 -607
rect 15884 -675 15918 -649
rect 15884 -683 15918 -675
rect 15884 -743 15918 -721
rect 15884 -755 15918 -743
rect 15884 -811 15918 -793
rect 15884 -827 15918 -811
rect 16040 109 16074 143
rect 16040 39 16074 71
rect 16040 37 16074 39
rect 16040 -29 16074 -1
rect 16040 -35 16074 -29
rect 16040 -97 16074 -73
rect 16040 -107 16074 -97
rect 16040 -165 16074 -145
rect 16040 -179 16074 -165
rect 16040 -233 16074 -217
rect 16040 -251 16074 -233
rect 16040 -301 16074 -289
rect 16040 -323 16074 -301
rect 16040 -369 16074 -361
rect 16040 -395 16074 -369
rect 16040 -437 16074 -433
rect 16040 -467 16074 -437
rect 16040 -539 16074 -505
rect 16040 -607 16074 -577
rect 16040 -611 16074 -607
rect 16040 -675 16074 -649
rect 16040 -683 16074 -675
rect 16040 -743 16074 -721
rect 16040 -755 16074 -743
rect 16040 -811 16074 -793
rect 16040 -827 16074 -811
rect 16196 109 16230 143
rect 16196 39 16230 71
rect 16196 37 16230 39
rect 16196 -29 16230 -1
rect 16196 -35 16230 -29
rect 16196 -97 16230 -73
rect 16196 -107 16230 -97
rect 16196 -165 16230 -145
rect 16196 -179 16230 -165
rect 16196 -233 16230 -217
rect 16196 -251 16230 -233
rect 16196 -301 16230 -289
rect 16196 -323 16230 -301
rect 16196 -369 16230 -361
rect 16196 -395 16230 -369
rect 16196 -437 16230 -433
rect 16196 -467 16230 -437
rect 16196 -539 16230 -505
rect 16196 -607 16230 -577
rect 16196 -611 16230 -607
rect 16196 -675 16230 -649
rect 16196 -683 16230 -675
rect 16196 -743 16230 -721
rect 16196 -755 16230 -743
rect 16196 -811 16230 -793
rect 16196 -827 16230 -811
rect 18482 148 18516 182
rect 18554 148 18584 182
rect 18584 148 18588 182
rect 16352 104 16386 111
rect 16352 77 16386 104
rect 18647 71 18678 105
rect 18678 71 18681 105
rect 18719 71 18746 105
rect 18746 71 18753 105
rect 16352 17 16386 37
rect 16352 3 16386 17
rect 18953 52 18987 86
rect 18482 -8 18516 26
rect 18554 -8 18584 26
rect 18584 -8 18588 26
rect 16352 -70 16386 -38
rect 16352 -72 16386 -70
rect 16352 -147 16386 -113
rect 16352 -191 16386 -188
rect 16352 -222 16386 -191
rect 16352 -279 16386 -263
rect 16352 -297 16386 -279
rect 16352 -367 16386 -338
rect 16352 -372 16386 -367
rect 16352 -421 16386 -413
rect 16352 -447 16386 -421
rect 16352 -509 16386 -488
rect 16352 -522 16386 -509
rect 16352 -597 16386 -563
rect 16352 -672 16386 -638
rect 16352 -719 16386 -713
rect 16352 -747 16386 -719
rect 16352 -807 16386 -788
rect 16352 -822 16386 -807
rect 16352 -895 16386 -863
rect 16352 -897 16386 -895
rect 15917 -937 15951 -935
rect 15917 -969 15932 -937
rect 15932 -969 15951 -937
rect 15990 -937 16024 -935
rect 16063 -937 16097 -935
rect 15990 -969 15991 -937
rect 15991 -969 16024 -937
rect 16063 -969 16084 -937
rect 16084 -969 16097 -937
rect 16136 -969 16170 -935
rect 16208 -937 16242 -935
rect 16280 -937 16314 -935
rect 16208 -969 16210 -937
rect 16210 -969 16242 -937
rect 16280 -969 16302 -937
rect 16302 -969 16314 -937
rect 18953 -22 18987 12
rect 18953 -96 18987 -62
rect 18953 -170 18987 -136
rect 18953 -244 18987 -210
rect 18953 -318 18987 -284
rect 18953 -392 18987 -358
rect 18953 -466 18987 -432
rect 18953 -540 18987 -506
rect 18953 -614 18987 -580
rect 18953 -687 18987 -653
rect 18953 -760 18987 -726
rect 18953 -833 18987 -799
rect 18953 -906 18987 -872
rect 18953 -979 18987 -945
rect 18953 -1052 18987 -1018
rect 18953 -1125 18987 -1091
rect 18953 -1198 18987 -1164
rect 17961 -1286 17995 -1252
rect 18037 -1286 18071 -1252
rect 18113 -1286 18147 -1252
rect 18189 -1286 18223 -1252
rect 18265 -1286 18299 -1252
rect 18341 -1286 18375 -1252
rect 18417 -1286 18451 -1252
rect 18953 -1271 18987 -1237
rect 570 -1380 586 -1346
rect 586 -1380 604 -1346
rect 642 -1380 654 -1346
rect 654 -1380 676 -1346
rect 714 -1380 722 -1346
rect 722 -1380 748 -1346
rect 786 -1380 790 -1346
rect 790 -1380 820 -1346
rect 858 -1380 892 -1346
rect 930 -1380 960 -1346
rect 960 -1380 964 -1346
rect 1002 -1380 1028 -1346
rect 1028 -1380 1036 -1346
rect 1074 -1380 1096 -1346
rect 1096 -1380 1108 -1346
rect 1146 -1380 1164 -1346
rect 1164 -1380 1180 -1346
rect 1218 -1380 1232 -1346
rect 1232 -1380 1252 -1346
rect 1290 -1380 1300 -1346
rect 1300 -1380 1324 -1346
rect 1362 -1380 1368 -1346
rect 1368 -1380 1396 -1346
rect 1434 -1380 1436 -1346
rect 1436 -1380 1468 -1346
rect 1506 -1380 1540 -1346
rect 17961 -1366 17995 -1332
rect 18037 -1366 18071 -1332
rect 18113 -1366 18147 -1332
rect 18189 -1366 18223 -1332
rect 18265 -1366 18299 -1332
rect 18341 -1366 18375 -1332
rect 18417 -1366 18451 -1332
rect 18953 -1344 18987 -1310
rect 466 -1424 500 -1390
rect 466 -1497 500 -1463
rect 17961 -1446 17995 -1412
rect 18037 -1446 18071 -1412
rect 18113 -1446 18147 -1412
rect 18189 -1446 18223 -1412
rect 18265 -1446 18299 -1412
rect 18341 -1446 18375 -1412
rect 18417 -1446 18451 -1412
rect 18953 -1417 18987 -1383
rect 570 -1536 586 -1502
rect 586 -1536 604 -1502
rect 642 -1536 654 -1502
rect 654 -1536 676 -1502
rect 714 -1536 722 -1502
rect 722 -1536 748 -1502
rect 786 -1536 790 -1502
rect 790 -1536 820 -1502
rect 858 -1536 892 -1502
rect 930 -1536 960 -1502
rect 960 -1536 964 -1502
rect 1002 -1536 1028 -1502
rect 1028 -1536 1036 -1502
rect 1074 -1536 1096 -1502
rect 1096 -1536 1108 -1502
rect 1146 -1536 1164 -1502
rect 1164 -1536 1180 -1502
rect 1218 -1536 1232 -1502
rect 1232 -1536 1252 -1502
rect 1290 -1536 1300 -1502
rect 1300 -1536 1324 -1502
rect 1362 -1536 1368 -1502
rect 1368 -1536 1396 -1502
rect 1434 -1536 1436 -1502
rect 1436 -1536 1468 -1502
rect 1506 -1536 1540 -1502
rect 1622 -1536 1656 -1507
rect 466 -1570 500 -1536
rect 466 -1643 500 -1609
rect 1622 -1541 1656 -1536
rect 1622 -1597 1656 -1592
rect 1622 -1626 1656 -1597
rect 466 -1716 500 -1682
rect 570 -1692 586 -1658
rect 586 -1692 604 -1658
rect 642 -1692 654 -1658
rect 654 -1692 676 -1658
rect 714 -1692 722 -1658
rect 722 -1692 748 -1658
rect 786 -1692 790 -1658
rect 790 -1692 820 -1658
rect 858 -1692 892 -1658
rect 930 -1692 960 -1658
rect 960 -1692 964 -1658
rect 1002 -1692 1028 -1658
rect 1028 -1692 1036 -1658
rect 1074 -1692 1096 -1658
rect 1096 -1692 1108 -1658
rect 1146 -1692 1164 -1658
rect 1164 -1692 1180 -1658
rect 1218 -1692 1232 -1658
rect 1232 -1692 1252 -1658
rect 1290 -1692 1300 -1658
rect 1300 -1692 1324 -1658
rect 1362 -1692 1368 -1658
rect 1368 -1692 1396 -1658
rect 1434 -1692 1436 -1658
rect 1436 -1692 1468 -1658
rect 1506 -1692 1540 -1658
rect 466 -1789 500 -1755
rect 1622 -1753 1656 -1733
rect 1622 -1767 1656 -1753
rect 466 -1862 500 -1828
rect 570 -1848 586 -1814
rect 586 -1848 604 -1814
rect 642 -1848 654 -1814
rect 654 -1848 676 -1814
rect 714 -1848 722 -1814
rect 722 -1848 748 -1814
rect 786 -1848 790 -1814
rect 790 -1848 820 -1814
rect 858 -1848 892 -1814
rect 930 -1848 960 -1814
rect 960 -1848 964 -1814
rect 1002 -1848 1028 -1814
rect 1028 -1848 1036 -1814
rect 1074 -1848 1096 -1814
rect 1096 -1848 1108 -1814
rect 1146 -1848 1164 -1814
rect 1164 -1848 1180 -1814
rect 1218 -1848 1232 -1814
rect 1232 -1848 1252 -1814
rect 1290 -1848 1300 -1814
rect 1300 -1848 1324 -1814
rect 1362 -1848 1368 -1814
rect 1368 -1848 1396 -1814
rect 1434 -1848 1436 -1814
rect 1436 -1848 1468 -1814
rect 1506 -1848 1540 -1814
rect 1622 -1848 1656 -1818
rect 466 -1935 500 -1901
rect 1622 -1852 1656 -1848
rect 1622 -1909 1656 -1904
rect 1622 -1938 1656 -1909
rect 466 -2008 500 -1974
rect 570 -2004 586 -1970
rect 586 -2004 604 -1970
rect 642 -2004 654 -1970
rect 654 -2004 676 -1970
rect 714 -2004 722 -1970
rect 722 -2004 748 -1970
rect 786 -2004 790 -1970
rect 790 -2004 820 -1970
rect 858 -2004 892 -1970
rect 930 -2004 960 -1970
rect 960 -2004 964 -1970
rect 1002 -2004 1028 -1970
rect 1028 -2004 1036 -1970
rect 1074 -2004 1096 -1970
rect 1096 -2004 1108 -1970
rect 1146 -2004 1164 -1970
rect 1164 -2004 1180 -1970
rect 1218 -2004 1232 -1970
rect 1232 -2004 1252 -1970
rect 1290 -2004 1300 -1970
rect 1300 -2004 1324 -1970
rect 1362 -2004 1368 -1970
rect 1368 -2004 1396 -1970
rect 1434 -2004 1436 -1970
rect 1436 -2004 1468 -1970
rect 1506 -2004 1540 -1970
rect 466 -2081 500 -2047
rect 466 -2154 500 -2120
rect 1622 -2065 1656 -2045
rect 1622 -2079 1656 -2065
rect 570 -2160 586 -2126
rect 586 -2160 604 -2126
rect 644 -2160 654 -2126
rect 654 -2160 678 -2126
rect 718 -2160 722 -2126
rect 722 -2160 752 -2126
rect 792 -2160 824 -2126
rect 824 -2160 826 -2126
rect 865 -2160 892 -2126
rect 892 -2160 899 -2126
rect 938 -2160 960 -2126
rect 960 -2160 972 -2126
rect 1011 -2160 1028 -2126
rect 1028 -2160 1045 -2126
rect 1622 -2160 1656 -2130
rect 1622 -2164 1656 -2160
rect 1622 -2221 1656 -2216
rect 1622 -2250 1656 -2221
rect 570 -2316 586 -2282
rect 586 -2316 604 -2282
rect 642 -2316 654 -2282
rect 654 -2316 676 -2282
rect 714 -2316 722 -2282
rect 722 -2316 748 -2282
rect 786 -2316 790 -2282
rect 790 -2316 820 -2282
rect 858 -2316 892 -2282
rect 930 -2316 960 -2282
rect 960 -2316 964 -2282
rect 1002 -2316 1028 -2282
rect 1028 -2316 1036 -2282
rect 1074 -2316 1096 -2282
rect 1096 -2316 1108 -2282
rect 1146 -2316 1164 -2282
rect 1164 -2316 1180 -2282
rect 1218 -2316 1232 -2282
rect 1232 -2316 1252 -2282
rect 1290 -2316 1300 -2282
rect 1300 -2316 1324 -2282
rect 1362 -2316 1368 -2282
rect 1368 -2316 1396 -2282
rect 1434 -2316 1436 -2282
rect 1436 -2316 1468 -2282
rect 1506 -2316 1540 -2282
rect 597 -2398 631 -2397
rect 675 -2398 709 -2397
rect 753 -2398 787 -2397
rect 831 -2398 865 -2397
rect 909 -2398 943 -2397
rect 987 -2398 1021 -2397
rect 1065 -2398 1099 -2397
rect 1143 -2398 1177 -2397
rect 1220 -2398 1254 -2397
rect 1297 -2398 1331 -2397
rect 1374 -2398 1408 -2397
rect 1451 -2398 1485 -2397
rect 1528 -2398 1562 -2397
rect 597 -2431 598 -2398
rect 598 -2431 631 -2398
rect 675 -2431 702 -2398
rect 702 -2431 709 -2398
rect 753 -2431 772 -2398
rect 772 -2431 787 -2398
rect 831 -2431 842 -2398
rect 842 -2431 865 -2398
rect 909 -2431 912 -2398
rect 912 -2431 943 -2398
rect 987 -2431 1019 -2398
rect 1019 -2431 1021 -2398
rect 1065 -2431 1090 -2398
rect 1090 -2431 1099 -2398
rect 1143 -2431 1161 -2398
rect 1161 -2431 1177 -2398
rect 1220 -2431 1232 -2398
rect 1232 -2431 1254 -2398
rect 1297 -2431 1303 -2398
rect 1303 -2431 1331 -2398
rect 1374 -2431 1408 -2398
rect 1451 -2431 1479 -2398
rect 1479 -2431 1485 -2398
rect 1528 -2431 1550 -2398
rect 1550 -2431 1562 -2398
rect 407 -3277 441 -3243
rect 700 -3265 733 -3231
rect 733 -3265 734 -3231
rect 777 -3265 801 -3231
rect 801 -3265 811 -3231
rect 407 -3333 440 -3316
rect 440 -3333 441 -3316
rect 407 -3350 441 -3333
rect 1039 -3275 1073 -3241
rect 1039 -3321 1073 -3313
rect 1039 -3347 1073 -3321
rect 407 -3401 440 -3389
rect 440 -3401 441 -3389
rect 407 -3423 441 -3401
rect 890 -3403 896 -3369
rect 896 -3403 924 -3369
rect 1039 -3389 1073 -3385
rect 407 -3469 440 -3462
rect 440 -3469 441 -3462
rect 407 -3496 441 -3469
rect 890 -3475 924 -3441
rect 1039 -3419 1073 -3389
rect 407 -3537 440 -3535
rect 440 -3537 441 -3535
rect 407 -3569 441 -3537
rect 407 -3639 441 -3608
rect 407 -3642 440 -3639
rect 440 -3642 441 -3639
rect 407 -3715 441 -3681
rect 407 -3780 440 -3754
rect 440 -3780 441 -3754
rect 407 -3788 441 -3780
rect 407 -3848 440 -3827
rect 440 -3848 441 -3827
rect 407 -3861 441 -3848
rect 407 -3916 440 -3900
rect 440 -3916 441 -3900
rect 407 -3934 441 -3916
rect 407 -3984 440 -3973
rect 440 -3984 441 -3973
rect 407 -4007 441 -3984
rect 407 -4052 440 -4046
rect 440 -4052 441 -4046
rect 407 -4080 441 -4052
rect 407 -4120 440 -4119
rect 440 -4120 441 -4119
rect 407 -4153 441 -4120
rect 407 -4222 441 -4192
rect 407 -4226 440 -4222
rect 440 -4226 441 -4222
rect 407 -4290 441 -4265
rect 407 -4299 440 -4290
rect 440 -4299 441 -4290
rect 407 -4358 441 -4338
rect 407 -4372 440 -4358
rect 440 -4372 441 -4358
rect 407 -4426 441 -4411
rect 407 -4445 440 -4426
rect 440 -4445 441 -4426
rect 407 -4494 441 -4484
rect 407 -4518 440 -4494
rect 440 -4518 441 -4494
rect 407 -4562 441 -4557
rect 407 -4591 440 -4562
rect 440 -4591 441 -4562
rect 407 -4664 440 -4630
rect 440 -4664 441 -4630
rect 407 -4732 440 -4703
rect 440 -4732 441 -4703
rect 407 -4737 441 -4732
rect 407 -4800 440 -4775
rect 440 -4800 441 -4775
rect 407 -4809 441 -4800
rect 407 -4868 440 -4847
rect 440 -4868 441 -4847
rect 407 -4881 441 -4868
rect 407 -4936 440 -4919
rect 440 -4936 441 -4919
rect 407 -4953 441 -4936
rect 407 -5004 440 -4991
rect 440 -5004 441 -4991
rect 407 -5025 441 -5004
rect 407 -5072 440 -5063
rect 440 -5072 441 -5063
rect 407 -5097 441 -5072
rect 407 -5140 440 -5135
rect 440 -5140 441 -5135
rect 407 -5169 441 -5140
rect 407 -5208 440 -5207
rect 440 -5208 441 -5207
rect 407 -5241 441 -5208
rect 407 -5310 441 -5279
rect 407 -5313 440 -5310
rect 440 -5313 441 -5310
rect 407 -5378 441 -5351
rect 407 -5385 440 -5378
rect 440 -5385 441 -5378
rect 407 -5446 441 -5423
rect 407 -5457 440 -5446
rect 440 -5457 441 -5446
rect 407 -5514 441 -5495
rect 407 -5529 440 -5514
rect 440 -5529 441 -5514
rect 407 -5582 441 -5567
rect 407 -5601 440 -5582
rect 440 -5601 441 -5582
rect 407 -5650 441 -5639
rect 407 -5673 440 -5650
rect 440 -5673 441 -5650
rect 407 -5718 441 -5711
rect 407 -5745 440 -5718
rect 440 -5745 441 -5718
rect 407 -5786 441 -5783
rect 407 -5817 440 -5786
rect 440 -5817 441 -5786
rect 407 -5888 440 -5855
rect 440 -5888 441 -5855
rect 407 -5889 441 -5888
rect 407 -5956 440 -5927
rect 440 -5956 441 -5927
rect 407 -5961 441 -5956
rect 407 -6024 440 -5999
rect 440 -6024 441 -5999
rect 407 -6033 441 -6024
rect 407 -6092 440 -6071
rect 440 -6092 441 -6071
rect 407 -6105 441 -6092
rect 407 -6160 440 -6143
rect 440 -6160 441 -6143
rect 407 -6177 441 -6160
rect 407 -6228 440 -6215
rect 440 -6228 441 -6215
rect 407 -6249 441 -6228
rect 407 -6296 440 -6287
rect 440 -6296 441 -6287
rect 407 -6321 441 -6296
rect 407 -6364 440 -6359
rect 440 -6364 441 -6359
rect 407 -6393 441 -6364
rect 407 -6432 440 -6431
rect 440 -6432 441 -6431
rect 407 -6465 441 -6432
rect 407 -6534 441 -6503
rect 407 -6537 440 -6534
rect 440 -6537 441 -6534
rect 407 -6602 441 -6575
rect 407 -6609 440 -6602
rect 440 -6609 441 -6602
rect 407 -6670 441 -6647
rect 407 -6681 440 -6670
rect 440 -6681 441 -6670
rect 407 -6738 441 -6719
rect 407 -6753 440 -6738
rect 440 -6753 441 -6738
rect 407 -6806 441 -6791
rect 407 -6825 440 -6806
rect 440 -6825 441 -6806
rect 407 -6874 441 -6863
rect 407 -6897 440 -6874
rect 440 -6897 441 -6874
rect 407 -6942 441 -6935
rect 407 -6969 440 -6942
rect 440 -6969 441 -6942
rect 407 -7010 441 -7007
rect 407 -7041 440 -7010
rect 440 -7041 441 -7010
rect 407 -7112 440 -7079
rect 440 -7112 441 -7079
rect 407 -7113 441 -7112
rect 407 -7180 440 -7151
rect 440 -7180 441 -7151
rect 407 -7185 441 -7180
rect 407 -7248 440 -7223
rect 440 -7248 441 -7223
rect 407 -7257 441 -7248
rect 407 -7316 440 -7295
rect 440 -7316 441 -7295
rect 407 -7329 441 -7316
rect 407 -7384 440 -7367
rect 440 -7384 441 -7367
rect 407 -7401 441 -7384
rect 407 -7452 440 -7439
rect 440 -7452 441 -7439
rect 407 -7473 441 -7452
rect 407 -7520 440 -7511
rect 440 -7520 441 -7511
rect 407 -7545 441 -7520
rect 407 -7588 440 -7583
rect 440 -7588 441 -7583
rect 407 -7617 441 -7588
rect 407 -7656 440 -7655
rect 440 -7656 441 -7655
rect 407 -7689 441 -7656
rect 407 -7758 441 -7727
rect 407 -7761 440 -7758
rect 440 -7761 441 -7758
rect 407 -7826 441 -7799
rect 407 -7833 440 -7826
rect 440 -7833 441 -7826
rect 407 -7894 441 -7871
rect 407 -7905 440 -7894
rect 440 -7905 441 -7894
rect 407 -7962 441 -7943
rect 407 -7977 440 -7962
rect 440 -7977 441 -7962
rect 407 -8030 441 -8015
rect 407 -8049 440 -8030
rect 440 -8049 441 -8030
rect 407 -8098 441 -8087
rect 407 -8121 440 -8098
rect 440 -8121 441 -8098
rect 407 -8166 441 -8159
rect 407 -8193 440 -8166
rect 440 -8193 441 -8166
rect 407 -8234 441 -8231
rect 407 -8265 440 -8234
rect 440 -8265 441 -8234
rect 407 -8336 440 -8303
rect 440 -8336 441 -8303
rect 407 -8337 441 -8336
rect 407 -8404 440 -8375
rect 440 -8404 441 -8375
rect 407 -8409 441 -8404
rect 407 -8472 440 -8447
rect 440 -8472 441 -8447
rect 407 -8481 441 -8472
rect 407 -8540 440 -8519
rect 440 -8540 441 -8519
rect 407 -8553 441 -8540
rect 407 -8608 440 -8591
rect 440 -8608 441 -8591
rect 407 -8625 441 -8608
rect 407 -8676 440 -8663
rect 440 -8676 441 -8663
rect 407 -8697 441 -8676
rect 407 -8744 440 -8735
rect 440 -8744 441 -8735
rect 407 -8769 441 -8744
rect 407 -8812 440 -8807
rect 440 -8812 441 -8807
rect 407 -8841 441 -8812
rect 407 -8880 440 -8879
rect 440 -8880 441 -8879
rect 407 -8913 441 -8880
rect 407 -8982 441 -8951
rect 407 -8985 440 -8982
rect 440 -8985 441 -8982
rect 407 -9050 441 -9023
rect 407 -9057 440 -9050
rect 440 -9057 441 -9050
rect 407 -9118 441 -9095
rect 407 -9129 440 -9118
rect 440 -9129 441 -9118
rect 407 -9186 441 -9167
rect 407 -9201 440 -9186
rect 440 -9201 441 -9186
rect 407 -9254 441 -9239
rect 407 -9273 440 -9254
rect 440 -9273 441 -9254
rect 407 -9322 441 -9311
rect 407 -9345 440 -9322
rect 440 -9345 441 -9322
rect 407 -9390 441 -9383
rect 407 -9417 440 -9390
rect 440 -9417 441 -9390
rect 407 -9458 441 -9455
rect 407 -9489 440 -9458
rect 440 -9489 441 -9458
rect 407 -9560 440 -9527
rect 440 -9560 441 -9527
rect 407 -9561 441 -9560
rect 407 -9628 440 -9599
rect 440 -9628 441 -9599
rect 407 -9633 441 -9628
rect 407 -9696 440 -9671
rect 440 -9696 441 -9671
rect 407 -9705 441 -9696
rect 407 -9764 440 -9743
rect 440 -9764 441 -9743
rect 407 -9777 441 -9764
rect 407 -9832 440 -9815
rect 440 -9832 441 -9815
rect 407 -9849 441 -9832
rect 407 -9900 440 -9887
rect 440 -9900 441 -9887
rect 407 -9921 441 -9900
rect 407 -9968 440 -9959
rect 440 -9968 441 -9959
rect 407 -9993 441 -9968
rect 407 -10036 440 -10031
rect 440 -10036 441 -10031
rect 407 -10065 441 -10036
rect 407 -10104 440 -10103
rect 440 -10104 441 -10103
rect 407 -10137 441 -10104
rect 407 -10206 441 -10175
rect 407 -10209 440 -10206
rect 440 -10209 441 -10206
rect 407 -10274 441 -10247
rect 407 -10281 440 -10274
rect 440 -10281 441 -10274
rect 407 -10342 441 -10319
rect 407 -10353 440 -10342
rect 440 -10353 441 -10342
rect 407 -10410 441 -10391
rect 407 -10425 440 -10410
rect 440 -10425 441 -10410
rect 407 -10478 441 -10463
rect 407 -10497 440 -10478
rect 440 -10497 441 -10478
rect 407 -10546 441 -10535
rect 407 -10569 440 -10546
rect 440 -10569 441 -10546
rect 407 -10614 441 -10607
rect 407 -10641 440 -10614
rect 440 -10641 441 -10614
rect 407 -10682 441 -10679
rect 407 -10713 440 -10682
rect 440 -10713 441 -10682
rect 407 -10784 440 -10751
rect 440 -10784 441 -10751
rect 407 -10785 441 -10784
rect 407 -10852 440 -10823
rect 440 -10852 441 -10823
rect 1039 -3491 1073 -3457
rect 1039 -3559 1073 -3529
rect 1039 -3563 1073 -3559
rect 1039 -3627 1073 -3601
rect 1039 -3635 1073 -3627
rect 1039 -3695 1073 -3673
rect 1039 -3707 1073 -3695
rect 1039 -3763 1073 -3745
rect 1039 -3779 1073 -3763
rect 1039 -3831 1073 -3817
rect 1039 -3851 1073 -3831
rect 1039 -3899 1073 -3889
rect 1039 -3923 1073 -3899
rect 1039 -3967 1073 -3961
rect 1039 -3995 1073 -3967
rect 1039 -4035 1073 -4033
rect 1039 -4067 1073 -4035
rect 1039 -4137 1073 -4105
rect 1039 -4139 1073 -4137
rect 1039 -4205 1073 -4177
rect 1039 -4211 1073 -4205
rect 1039 -4273 1073 -4249
rect 1039 -4283 1073 -4273
rect 1039 -4341 1073 -4321
rect 1039 -4355 1073 -4341
rect 1039 -4409 1073 -4393
rect 1039 -4427 1073 -4409
rect 1039 -4477 1073 -4465
rect 1039 -4499 1073 -4477
rect 1039 -4545 1073 -4537
rect 1039 -4571 1073 -4545
rect 1039 -4613 1073 -4609
rect 1039 -4643 1073 -4613
rect 1039 -4715 1073 -4681
rect 1039 -4783 1073 -4753
rect 1039 -4787 1073 -4783
rect 1039 -4851 1073 -4825
rect 1039 -4859 1073 -4851
rect 1039 -4919 1073 -4897
rect 1039 -4931 1073 -4919
rect 1039 -4987 1073 -4969
rect 1039 -5003 1073 -4987
rect 1039 -5055 1073 -5041
rect 1039 -5075 1073 -5055
rect 1039 -5123 1073 -5113
rect 1039 -5147 1073 -5123
rect 1039 -5191 1073 -5185
rect 1039 -5219 1073 -5191
rect 1039 -5259 1073 -5257
rect 1039 -5291 1073 -5259
rect 1039 -5361 1073 -5329
rect 1039 -5363 1073 -5361
rect 1039 -5429 1073 -5401
rect 1039 -5435 1073 -5429
rect 1039 -5497 1073 -5473
rect 1039 -5507 1073 -5497
rect 1039 -5565 1073 -5545
rect 1039 -5579 1073 -5565
rect 1039 -5633 1073 -5617
rect 1039 -5651 1073 -5633
rect 1039 -5701 1073 -5689
rect 1039 -5723 1073 -5701
rect 1039 -5769 1073 -5761
rect 1039 -5795 1073 -5769
rect 1039 -5837 1073 -5833
rect 1039 -5867 1073 -5837
rect 1039 -5939 1073 -5905
rect 1039 -6007 1073 -5977
rect 1039 -6011 1073 -6007
rect 1039 -6075 1073 -6049
rect 1039 -6083 1073 -6075
rect 1039 -6143 1073 -6121
rect 1039 -6155 1073 -6143
rect 1039 -6211 1073 -6193
rect 1039 -6227 1073 -6211
rect 1039 -6279 1073 -6265
rect 1039 -6299 1073 -6279
rect 1039 -6347 1073 -6337
rect 1039 -6371 1073 -6347
rect 1039 -6415 1073 -6409
rect 1039 -6443 1073 -6415
rect 1039 -6483 1073 -6481
rect 1039 -6515 1073 -6483
rect 1039 -6585 1073 -6553
rect 1039 -6587 1073 -6585
rect 1039 -6653 1073 -6625
rect 1039 -6659 1073 -6653
rect 1039 -6721 1073 -6697
rect 1039 -6731 1073 -6721
rect 1039 -6789 1073 -6769
rect 1039 -6803 1073 -6789
rect 1039 -6857 1073 -6841
rect 1039 -6875 1073 -6857
rect 1039 -6925 1073 -6913
rect 1039 -6947 1073 -6925
rect 1039 -6993 1073 -6985
rect 1039 -7019 1073 -6993
rect 1039 -7061 1073 -7057
rect 1039 -7091 1073 -7061
rect 1039 -7163 1073 -7129
rect 1039 -7231 1073 -7201
rect 1039 -7235 1073 -7231
rect 1039 -7299 1073 -7273
rect 1039 -7307 1073 -7299
rect 1039 -7367 1073 -7345
rect 1039 -7379 1073 -7367
rect 1039 -7435 1073 -7417
rect 1039 -7451 1073 -7435
rect 1039 -7503 1073 -7489
rect 1039 -7523 1073 -7503
rect 1039 -7571 1073 -7561
rect 1039 -7595 1073 -7571
rect 1039 -7639 1073 -7633
rect 1039 -7667 1073 -7639
rect 1039 -7707 1073 -7705
rect 1039 -7739 1073 -7707
rect 1039 -7809 1073 -7777
rect 1039 -7811 1073 -7809
rect 1039 -7877 1073 -7849
rect 1039 -7883 1073 -7877
rect 1039 -7945 1073 -7921
rect 1039 -7955 1073 -7945
rect 1039 -8013 1073 -7993
rect 1039 -8027 1073 -8013
rect 1039 -8081 1073 -8065
rect 1039 -8099 1073 -8081
rect 1039 -8149 1073 -8137
rect 1039 -8171 1073 -8149
rect 1039 -8217 1073 -8209
rect 1039 -8243 1073 -8217
rect 1039 -8285 1073 -8281
rect 1039 -8315 1073 -8285
rect 1039 -8387 1073 -8353
rect 1039 -8455 1073 -8425
rect 1039 -8459 1073 -8455
rect 1039 -8523 1073 -8497
rect 1039 -8531 1073 -8523
rect 1039 -8591 1073 -8569
rect 1039 -8603 1073 -8591
rect 1039 -8659 1073 -8641
rect 1039 -8675 1073 -8659
rect 1039 -8727 1073 -8713
rect 1039 -8747 1073 -8727
rect 1039 -8795 1073 -8785
rect 1039 -8819 1073 -8795
rect 1039 -8863 1073 -8857
rect 1039 -8891 1073 -8863
rect 1039 -8931 1073 -8929
rect 1039 -8963 1073 -8931
rect 1039 -9033 1073 -9001
rect 1039 -9035 1073 -9033
rect 1039 -9101 1073 -9073
rect 1039 -9107 1073 -9101
rect 1039 -9169 1073 -9145
rect 1039 -9179 1073 -9169
rect 1039 -9237 1073 -9217
rect 1039 -9251 1073 -9237
rect 1039 -9305 1073 -9289
rect 1039 -9323 1073 -9305
rect 1039 -9373 1073 -9361
rect 1039 -9395 1073 -9373
rect 1039 -9441 1073 -9433
rect 1039 -9467 1073 -9441
rect 1039 -9509 1073 -9506
rect 1039 -9540 1073 -9509
rect 1039 -9611 1073 -9579
rect 1039 -9613 1073 -9611
rect 1039 -9679 1073 -9652
rect 1039 -9686 1073 -9679
rect 1039 -9747 1073 -9725
rect 1039 -9759 1073 -9747
rect 1039 -9815 1073 -9798
rect 1039 -9832 1073 -9815
rect 1039 -9883 1073 -9871
rect 1039 -9905 1073 -9883
rect 1039 -9951 1073 -9944
rect 1039 -9978 1073 -9951
rect 1039 -10019 1073 -10017
rect 1039 -10051 1073 -10019
rect 1039 -10121 1073 -10090
rect 1039 -10124 1073 -10121
rect 1039 -10189 1073 -10163
rect 2624 -9658 2658 -9624
rect 2624 -9730 2658 -9698
rect 2624 -9732 2658 -9730
rect 2624 -9798 2658 -9772
rect 2624 -9806 2658 -9798
rect 2624 -9866 2658 -9846
rect 2624 -9880 2658 -9866
rect 2624 -9934 2658 -9920
rect 2624 -9954 2658 -9934
rect 2624 -10002 2658 -9994
rect 2624 -10028 2658 -10002
rect 2624 -10070 2658 -10068
rect 2624 -10102 2658 -10070
rect 2624 -10172 2658 -10142
rect 2624 -10176 2658 -10172
rect 2780 -9658 2814 -9624
rect 2780 -9730 2814 -9698
rect 2780 -9732 2814 -9730
rect 2780 -9798 2814 -9772
rect 2780 -9806 2814 -9798
rect 2780 -9866 2814 -9846
rect 2780 -9880 2814 -9866
rect 2780 -9934 2814 -9920
rect 2780 -9954 2814 -9934
rect 2780 -10002 2814 -9994
rect 2780 -10028 2814 -10002
rect 2780 -10070 2814 -10068
rect 2780 -10102 2814 -10070
rect 2780 -10172 2814 -10142
rect 2780 -10176 2814 -10172
rect 2936 -9658 2970 -9624
rect 2936 -9730 2970 -9698
rect 2936 -9732 2970 -9730
rect 2936 -9798 2970 -9772
rect 2936 -9806 2970 -9798
rect 2936 -9866 2970 -9846
rect 2936 -9880 2970 -9866
rect 2936 -9934 2970 -9920
rect 2936 -9954 2970 -9934
rect 2936 -10002 2970 -9994
rect 2936 -10028 2970 -10002
rect 2936 -10070 2970 -10068
rect 2936 -10102 2970 -10070
rect 2936 -10172 2970 -10142
rect 2936 -10176 2970 -10172
rect 1039 -10197 1073 -10189
rect 1039 -10257 1073 -10236
rect 1039 -10270 1073 -10257
rect 2681 -10266 2685 -10232
rect 2685 -10266 2715 -10232
rect 2780 -10266 2814 -10232
rect 2879 -10266 2909 -10232
rect 2909 -10266 2913 -10232
rect 1039 -10325 1073 -10309
rect 1039 -10343 1073 -10325
rect 1039 -10393 1073 -10382
rect 1039 -10416 1073 -10393
rect 1039 -10461 1073 -10455
rect 1039 -10489 1073 -10461
rect 1039 -10529 1073 -10528
rect 1039 -10562 1073 -10529
rect 1039 -10631 1073 -10601
rect 1039 -10635 1073 -10631
rect 1039 -10699 1073 -10674
rect 1039 -10708 1073 -10699
rect 1039 -10767 1073 -10747
rect 1039 -10781 1073 -10767
rect 1039 -10835 1073 -10820
rect 407 -10857 441 -10852
rect 407 -10920 440 -10895
rect 440 -10920 441 -10895
rect 407 -10929 441 -10920
rect 548 -10880 582 -10846
rect 548 -10922 582 -10918
rect 1039 -10854 1073 -10835
rect 1039 -10903 1073 -10893
rect 548 -10952 582 -10922
rect 1039 -10927 1073 -10903
rect 407 -10988 440 -10967
rect 440 -10988 441 -10967
rect 407 -11001 441 -10988
rect 407 -11073 441 -11039
rect 1039 -10971 1073 -10966
rect 1039 -11000 1073 -10971
rect 1039 -11073 1073 -11039
rect 479 -11145 513 -11111
rect 559 -11145 593 -11111
rect 639 -11145 673 -11111
rect 719 -11145 753 -11111
rect 799 -11145 833 -11111
rect 879 -11145 913 -11111
rect 959 -11145 993 -11111
rect 18762 -11638 18796 -11604
rect 18762 -11726 18796 -11692
rect 18874 -12831 18908 -12797
rect 18874 -12969 18908 -12940
rect 18874 -12974 18908 -12969
rect 3080 -17018 3114 -17011
rect 3179 -17018 3213 -17011
rect 3278 -17018 3312 -17011
rect 3080 -17045 3084 -17018
rect 3084 -17045 3114 -17018
rect 3179 -17045 3213 -17018
rect 3278 -17045 3308 -17018
rect 3308 -17045 3312 -17018
rect 3023 -17452 3057 -17428
rect 3023 -17462 3057 -17452
rect 3023 -17520 3057 -17501
rect 3023 -17535 3057 -17520
rect 3023 -17588 3057 -17575
rect 3023 -17609 3057 -17588
rect 3023 -17683 3057 -17649
rect 3179 -17452 3213 -17431
rect 3179 -17465 3213 -17452
rect 3179 -17520 3213 -17503
rect 3179 -17537 3213 -17520
rect 3179 -17588 3213 -17576
rect 3179 -17610 3213 -17588
rect 3179 -17683 3213 -17649
rect 3335 -17452 3369 -17428
rect 3335 -17462 3369 -17452
rect 3335 -17520 3369 -17501
rect 3335 -17535 3369 -17520
rect 3335 -17588 3369 -17575
rect 3335 -17609 3369 -17588
rect 3335 -17683 3369 -17649
rect 2637 -17867 2641 -17833
rect 2641 -17867 2671 -17833
rect 2737 -17867 2770 -17833
rect 2770 -17867 2771 -17833
rect 2836 -17867 2865 -17833
rect 2865 -17867 2870 -17833
rect 2580 -18121 2614 -18114
rect 2580 -18148 2614 -18121
rect 2580 -18223 2614 -18194
rect 2580 -18228 2614 -18223
rect 2580 -18291 2614 -18274
rect 2580 -18308 2614 -18291
rect 2580 -18359 2614 -18354
rect 2580 -18388 2614 -18359
rect 2580 -18461 2614 -18435
rect 2580 -18469 2614 -18461
rect 2580 -18529 2614 -18516
rect 2580 -18550 2614 -18529
rect 2580 -18631 2614 -18597
rect 2580 -18699 2614 -18678
rect 2580 -18712 2614 -18699
rect 2736 -18223 2770 -18214
rect 2736 -18248 2770 -18223
rect 2736 -18291 2770 -18287
rect 2736 -18321 2770 -18291
rect 2736 -18393 2770 -18360
rect 2736 -18394 2770 -18393
rect 2736 -18461 2770 -18433
rect 2736 -18467 2770 -18461
rect 2736 -18529 2770 -18506
rect 2736 -18540 2770 -18529
rect 2736 -18597 2770 -18579
rect 2736 -18613 2770 -18597
rect 2736 -18665 2770 -18652
rect 2736 -18686 2770 -18665
rect 2736 -18733 2770 -18725
rect 2736 -18759 2770 -18733
rect 2736 -18801 2770 -18799
rect 2736 -18833 2770 -18801
rect 2736 -18903 2770 -18873
rect 2736 -18907 2770 -18903
rect 2892 -18121 2926 -18114
rect 2892 -18148 2926 -18121
rect 2892 -18189 2926 -18187
rect 2892 -18221 2926 -18189
rect 2892 -18291 2926 -18260
rect 2892 -18294 2926 -18291
rect 2892 -18359 2926 -18333
rect 2892 -18367 2926 -18359
rect 2892 -18427 2926 -18406
rect 2892 -18440 2926 -18427
rect 2892 -18495 2926 -18479
rect 2892 -18513 2926 -18495
rect 2892 -18563 2926 -18552
rect 2892 -18586 2926 -18563
rect 2892 -18631 2926 -18625
rect 2892 -18659 2926 -18631
rect 2892 -18733 2926 -18699
rect 2892 -18801 2926 -18773
rect 2892 -18807 2926 -18801
<< metal1 >>
rect 454 4994 7878 5000
rect 506 4960 539 4994
rect 573 4960 611 4994
rect 645 4960 683 4994
rect 717 4960 755 4994
rect 789 4960 827 4994
rect 861 4960 899 4994
rect 933 4960 971 4994
rect 1005 4960 1043 4994
rect 1077 4960 1115 4994
rect 1149 4960 1187 4994
rect 1221 4960 1259 4994
rect 1293 4960 1331 4994
rect 1365 4960 1403 4994
rect 1437 4960 1475 4994
rect 1509 4960 1547 4994
rect 1581 4960 1619 4994
rect 1653 4960 1691 4994
rect 1725 4960 1763 4994
rect 1797 4960 1835 4994
rect 1869 4960 1907 4994
rect 1941 4960 1979 4994
rect 2013 4960 2051 4994
rect 2085 4960 2123 4994
rect 2157 4960 2195 4994
rect 2229 4960 2267 4994
rect 2301 4960 2339 4994
rect 2373 4960 2411 4994
rect 2445 4960 2483 4994
rect 2517 4960 2555 4994
rect 2589 4960 2627 4994
rect 2661 4960 2699 4994
rect 2733 4960 2771 4994
rect 2805 4960 2843 4994
rect 2877 4960 2915 4994
rect 2949 4960 2987 4994
rect 3021 4960 3059 4994
rect 3093 4960 3131 4994
rect 3165 4960 3203 4994
rect 3237 4960 3275 4994
rect 3309 4960 3347 4994
rect 3381 4960 3419 4994
rect 3453 4960 3491 4994
rect 3525 4960 3563 4994
rect 3597 4960 3635 4994
rect 3669 4960 3707 4994
rect 3741 4960 3779 4994
rect 3813 4960 3851 4994
rect 3885 4960 3923 4994
rect 3957 4960 3995 4994
rect 4029 4960 4067 4994
rect 4101 4960 4139 4994
rect 4173 4960 4211 4994
rect 4245 4960 4283 4994
rect 4317 4960 4355 4994
rect 4389 4960 4427 4994
rect 4461 4960 4499 4994
rect 4533 4960 4571 4994
rect 4605 4960 4643 4994
rect 4677 4960 4715 4994
rect 4749 4960 4787 4994
rect 4821 4960 4859 4994
rect 4893 4960 4931 4994
rect 4965 4960 5003 4994
rect 5037 4960 5075 4994
rect 5109 4960 5147 4994
rect 5181 4960 5219 4994
rect 5253 4960 5291 4994
rect 5325 4960 5363 4994
rect 5397 4960 5435 4994
rect 5469 4960 5507 4994
rect 5541 4960 5579 4994
rect 5613 4960 5651 4994
rect 5685 4960 5723 4994
rect 5757 4960 5795 4994
rect 5829 4960 5868 4994
rect 5902 4960 5941 4994
rect 5975 4960 6014 4994
rect 6048 4960 6087 4994
rect 6121 4960 6160 4994
rect 6194 4960 6233 4994
rect 6267 4960 6306 4994
rect 6340 4960 6379 4994
rect 6413 4960 6452 4994
rect 6486 4960 6525 4994
rect 6559 4960 6598 4994
rect 6632 4960 6671 4994
rect 6705 4960 6744 4994
rect 6778 4960 6817 4994
rect 6851 4960 6890 4994
rect 6924 4960 6963 4994
rect 6997 4960 7036 4994
rect 7070 4960 7109 4994
rect 7143 4960 7182 4994
rect 7216 4960 7255 4994
rect 7289 4960 7328 4994
rect 7362 4960 7401 4994
rect 7435 4960 7474 4994
rect 7508 4960 7547 4994
rect 7581 4960 7620 4994
rect 7654 4960 7693 4994
rect 7727 4960 7766 4994
rect 7800 4960 7878 4994
rect 506 4954 7878 4960
rect 506 4942 514 4954
rect 454 4922 514 4942
rect 454 4912 467 4922
rect 501 4920 514 4922
tri 514 4920 548 4954 nw
tri 6824 4920 6858 4954 ne
rect 6858 4920 7878 4954
rect 501 4917 511 4920
tri 511 4917 514 4920 nw
tri 6858 4917 6861 4920 ne
rect 6861 4917 7838 4920
rect 501 4912 507 4917
tri 507 4913 511 4917 nw
rect 506 4860 507 4912
rect 569 4865 575 4917
rect 627 4865 639 4917
rect 691 4911 697 4917
tri 697 4911 703 4917 sw
tri 6861 4911 6867 4917 ne
rect 6867 4911 7838 4917
rect 691 4904 6811 4911
tri 6811 4904 6818 4911 sw
tri 6867 4904 6874 4911 ne
rect 6874 4904 7838 4911
rect 691 4900 6818 4904
tri 6818 4900 6822 4904 sw
tri 6874 4900 6878 4904 ne
rect 6878 4900 7838 4904
rect 691 4886 6822 4900
tri 6822 4886 6836 4900 sw
tri 6878 4886 6892 4900 ne
rect 6892 4886 7838 4900
rect 7872 4886 7878 4920
rect 691 4878 6836 4886
tri 6836 4878 6844 4886 sw
tri 6892 4878 6900 4886 ne
rect 6900 4878 7878 4886
rect 691 4865 6844 4878
tri 6844 4865 6857 4878 sw
tri 6900 4865 6913 4878 ne
rect 6913 4865 7878 4878
rect 454 4847 507 4860
rect 454 4830 467 4847
rect 501 4830 507 4847
tri 5275 4846 5294 4865 ne
rect 5294 4846 5362 4865
tri 5362 4846 5381 4865 nw
tri 5787 4846 5806 4865 ne
rect 5806 4846 5874 4865
tri 5874 4846 5893 4865 nw
tri 6299 4846 6318 4865 ne
rect 6318 4846 6386 4865
tri 6386 4846 6405 4865 nw
tri 6792 4846 6811 4865 ne
rect 6811 4856 6857 4865
tri 6857 4856 6866 4865 sw
tri 6913 4860 6918 4865 ne
rect 6918 4860 7878 4865
tri 6918 4856 6922 4860 ne
rect 6922 4856 6964 4860
rect 6811 4846 6866 4856
tri 6866 4846 6876 4856 sw
tri 6922 4846 6932 4856 ne
rect 6932 4846 6964 4856
tri 5294 4835 5305 4846 ne
rect 506 4778 507 4830
rect 454 4772 507 4778
rect 454 4748 467 4772
rect 501 4748 507 4772
rect 506 4696 507 4748
rect 454 4666 467 4696
rect 501 4666 507 4696
rect 506 4614 507 4666
rect 454 4588 467 4614
rect 501 4588 507 4614
rect 647 4831 2023 4835
rect 647 4824 1210 4831
rect 647 4823 952 4824
rect 647 4789 663 4823
rect 697 4789 871 4823
rect 905 4789 952 4823
rect 647 4772 952 4789
rect 1004 4772 1044 4824
rect 1096 4772 1135 4824
rect 1187 4779 1210 4824
rect 1262 4779 1279 4831
rect 1331 4779 1348 4831
rect 1400 4779 1417 4831
rect 1469 4779 1486 4831
rect 1538 4779 1554 4831
rect 1606 4779 1622 4831
rect 1674 4779 1690 4831
rect 1742 4823 1758 4831
rect 1742 4779 1758 4789
rect 1810 4779 1826 4831
rect 1878 4779 1894 4831
rect 1946 4779 1962 4831
rect 2014 4823 2023 4831
rect 2017 4789 2023 4823
rect 2014 4779 2023 4789
rect 1187 4772 2023 4779
rect 647 4753 2023 4772
rect 647 4751 1210 4753
rect 647 4740 871 4751
rect 647 4706 663 4740
rect 697 4717 871 4740
rect 905 4744 1210 4751
rect 905 4717 952 4744
rect 697 4706 952 4717
rect 647 4692 952 4706
rect 1004 4692 1044 4744
rect 1096 4692 1135 4744
rect 1187 4701 1210 4744
rect 1262 4701 1279 4753
rect 1331 4701 1348 4753
rect 1400 4701 1417 4753
rect 1469 4701 1486 4753
rect 1538 4701 1554 4753
rect 1606 4701 1622 4753
rect 1674 4701 1690 4753
rect 1742 4751 1758 4753
rect 1742 4701 1758 4717
rect 1810 4701 1826 4753
rect 1878 4701 1894 4753
rect 1946 4701 1962 4753
rect 2014 4751 2023 4753
rect 2017 4717 2023 4751
rect 2014 4701 2023 4717
rect 1187 4697 2023 4701
rect 2233 4823 2279 4835
rect 2233 4789 2239 4823
rect 2273 4789 2279 4823
rect 2233 4751 2279 4789
rect 2233 4717 2239 4751
rect 2273 4717 2279 4751
rect 1187 4692 1726 4697
rect 647 4667 1726 4692
tri 1726 4667 1756 4697 nw
rect 647 4664 1723 4667
tri 1723 4664 1726 4667 nw
rect 647 4657 952 4664
rect 647 4623 663 4657
rect 697 4652 952 4657
rect 1004 4652 1044 4664
rect 1096 4652 1135 4664
rect 1187 4661 1720 4664
tri 1720 4661 1723 4664 nw
rect 1187 4652 1686 4661
rect 697 4623 928 4652
rect 647 4618 928 4623
rect 1004 4618 1006 4652
rect 1040 4618 1044 4652
rect 1118 4618 1135 4652
rect 1196 4618 1239 4652
rect 1273 4618 1316 4652
rect 1350 4618 1393 4652
rect 1427 4618 1470 4652
rect 1504 4618 1547 4652
rect 1581 4618 1624 4652
rect 1658 4627 1686 4652
tri 1686 4627 1720 4661 nw
rect 1658 4618 1677 4627
tri 1677 4618 1686 4627 nw
rect 647 4612 952 4618
rect 1004 4612 1044 4618
rect 1096 4612 1135 4618
rect 1187 4615 1674 4618
tri 1674 4615 1677 4618 nw
rect 2039 4615 2045 4667
rect 2097 4615 2118 4667
rect 2170 4615 2176 4667
rect 1187 4612 1670 4615
rect 647 4611 1670 4612
tri 1670 4611 1674 4615 nw
tri 2212 4590 2233 4611 se
rect 2233 4590 2279 4717
rect 2486 4823 2538 4835
rect 2486 4819 2495 4823
rect 2529 4819 2538 4823
rect 2486 4755 2538 4767
rect 2486 4697 2538 4703
rect 2745 4823 2791 4835
rect 2745 4789 2751 4823
rect 2785 4789 2791 4823
rect 2745 4751 2791 4789
rect 2745 4717 2751 4751
rect 2785 4717 2791 4751
rect 2330 4615 2336 4667
rect 2388 4615 2413 4667
rect 2465 4615 2490 4667
rect 2542 4615 2567 4667
rect 2619 4615 2644 4667
rect 2696 4615 2702 4667
tri 2279 4590 2300 4611 sw
tri 2724 4590 2745 4611 se
rect 2745 4590 2791 4717
rect 2998 4823 3050 4835
rect 2998 4819 3007 4823
rect 3041 4819 3050 4823
rect 2998 4755 3050 4767
rect 2998 4697 3050 4703
rect 3257 4823 3303 4835
rect 3257 4789 3263 4823
rect 3297 4789 3303 4823
rect 3257 4751 3303 4789
rect 3257 4717 3263 4751
rect 3297 4717 3303 4751
rect 3510 4823 3562 4835
rect 3510 4819 3519 4823
rect 3553 4819 3562 4823
rect 3510 4755 3562 4767
tri 3479 4717 3510 4748 se
rect 2825 4615 2831 4667
rect 2883 4615 2898 4667
rect 2950 4661 2965 4667
rect 3017 4661 3031 4667
rect 3083 4661 3097 4667
rect 2956 4627 2965 4661
rect 3083 4627 3091 4661
rect 2950 4615 2965 4627
rect 3017 4615 3031 4627
rect 3083 4615 3097 4627
rect 3149 4615 3163 4667
rect 3215 4615 3221 4667
tri 3240 4590 3257 4607 se
rect 3257 4590 3303 4717
tri 3464 4702 3479 4717 se
rect 3479 4703 3510 4717
rect 3479 4702 3562 4703
tri 3460 4698 3464 4702 se
rect 3464 4698 3562 4702
tri 3459 4697 3460 4698 se
rect 3460 4697 3562 4698
rect 3769 4823 3815 4835
rect 3769 4789 3775 4823
rect 3809 4789 3815 4823
rect 3769 4751 3815 4789
rect 3769 4717 3775 4751
rect 3809 4717 3815 4751
tri 3429 4667 3459 4697 se
rect 3459 4667 3511 4697
tri 3511 4667 3541 4697 nw
rect 3373 4661 3508 4667
tri 3508 4664 3511 4667 nw
rect 3373 4627 3385 4661
rect 3419 4627 3462 4661
rect 3496 4627 3508 4661
rect 3373 4621 3508 4627
rect 3564 4615 3570 4667
rect 3622 4615 3679 4667
rect 3731 4615 3737 4667
rect 454 4584 507 4588
rect 506 4532 507 4584
tri 2204 4582 2212 4590 se
rect 2212 4582 2300 4590
tri 2300 4582 2308 4590 sw
tri 2716 4582 2724 4590 se
rect 2724 4582 2791 4590
tri 3232 4582 3240 4590 se
rect 3240 4582 3303 4590
tri 2203 4581 2204 4582 se
rect 2204 4581 2308 4582
tri 2308 4581 2309 4582 sw
tri 2715 4581 2716 4582 se
rect 2716 4581 2791 4582
rect 454 4513 467 4532
rect 501 4513 507 4532
rect 787 4529 793 4581
rect 845 4529 857 4581
rect 909 4529 2791 4581
tri 3226 4576 3232 4582 se
rect 3232 4576 3303 4582
rect 3001 4530 3303 4576
rect 3769 4590 3815 4717
rect 4022 4823 4074 4835
rect 4022 4819 4031 4823
rect 4065 4819 4074 4823
rect 4022 4755 4074 4767
rect 4022 4697 4074 4703
rect 4281 4823 4327 4835
rect 4281 4789 4287 4823
rect 4321 4789 4327 4823
rect 4281 4751 4327 4789
rect 4281 4717 4287 4751
rect 4321 4717 4327 4751
rect 3846 4615 3852 4667
rect 3904 4615 3921 4667
rect 3973 4661 3990 4667
rect 4042 4661 4058 4667
rect 4110 4661 4126 4667
rect 3979 4627 3990 4661
rect 4110 4627 4119 4661
rect 3973 4615 3990 4627
rect 4042 4615 4058 4627
rect 4110 4615 4126 4627
rect 4178 4615 4194 4667
rect 4246 4615 4252 4667
rect 4281 4606 4327 4717
rect 4534 4823 4586 4835
rect 4534 4819 4543 4823
rect 4577 4819 4586 4823
rect 4534 4755 4586 4767
rect 4534 4697 4586 4703
rect 4793 4823 4839 4835
rect 4793 4789 4799 4823
rect 4833 4789 4839 4823
rect 4793 4751 4839 4789
rect 4793 4717 4799 4751
rect 4833 4717 4839 4751
rect 4359 4615 4365 4667
rect 4417 4615 4433 4667
rect 4485 4661 4501 4667
rect 4553 4661 4569 4667
rect 4621 4661 4636 4667
rect 4491 4627 4501 4661
rect 4621 4627 4629 4661
rect 4485 4615 4501 4627
rect 4553 4615 4569 4627
rect 4621 4615 4636 4627
rect 4688 4615 4703 4667
rect 4755 4615 4761 4667
tri 4327 4606 4328 4607 sw
tri 3815 4590 3829 4604 sw
tri 4267 4590 4281 4604 se
rect 4281 4590 4328 4606
tri 4328 4590 4344 4606 sw
tri 4777 4590 4793 4606 se
rect 4793 4590 4839 4717
rect 5046 4823 5098 4835
rect 5046 4819 5055 4823
rect 5089 4819 5098 4823
rect 5046 4755 5098 4767
rect 5305 4823 5351 4846
tri 5351 4835 5362 4846 nw
tri 5806 4835 5817 4846 ne
rect 5305 4789 5311 4823
rect 5345 4789 5351 4823
rect 5305 4751 5351 4789
rect 5305 4717 5311 4751
rect 5345 4717 5351 4751
rect 5305 4705 5351 4717
rect 5558 4823 5610 4835
rect 5558 4819 5567 4823
rect 5601 4819 5610 4823
rect 5558 4755 5610 4767
rect 5046 4697 5098 4703
rect 5817 4823 5863 4846
tri 5863 4835 5874 4846 nw
tri 6318 4835 6329 4846 ne
rect 5817 4789 5823 4823
rect 5857 4789 5863 4823
rect 5817 4751 5863 4789
rect 5817 4717 5823 4751
rect 5857 4717 5863 4751
rect 5817 4705 5863 4717
rect 6070 4823 6122 4835
rect 6070 4819 6079 4823
rect 6113 4819 6122 4823
rect 6070 4755 6122 4767
rect 5558 4697 5610 4703
rect 6329 4823 6375 4846
tri 6375 4835 6386 4846 nw
tri 6811 4839 6818 4846 ne
rect 6818 4839 6876 4846
tri 6818 4835 6822 4839 ne
rect 6822 4835 6876 4839
tri 6876 4835 6887 4846 sw
tri 6932 4835 6943 4846 ne
rect 6943 4835 6964 4846
rect 6329 4789 6335 4823
rect 6369 4789 6375 4823
rect 6329 4751 6375 4789
rect 6329 4717 6335 4751
rect 6369 4717 6375 4751
rect 6329 4705 6375 4717
rect 6582 4823 6634 4835
tri 6822 4825 6832 4835 ne
rect 6832 4825 6887 4835
tri 6832 4823 6834 4825 ne
rect 6834 4823 6887 4825
tri 6943 4823 6955 4835 ne
rect 6955 4823 6964 4835
rect 6582 4819 6591 4823
rect 6625 4819 6634 4823
tri 6834 4820 6837 4823 ne
rect 6837 4820 6847 4823
tri 6837 4816 6841 4820 ne
rect 6582 4755 6634 4767
rect 6070 4697 6122 4703
rect 6841 4789 6847 4820
rect 6881 4789 6887 4823
tri 6955 4820 6958 4823 ne
rect 6841 4751 6887 4789
rect 6841 4717 6847 4751
rect 6881 4717 6887 4751
rect 6841 4705 6887 4717
rect 6958 4808 6964 4823
rect 7016 4808 7029 4860
rect 7081 4808 7094 4860
rect 7146 4808 7158 4860
rect 7210 4808 7222 4860
rect 7274 4808 7286 4860
rect 7338 4808 7350 4860
rect 7402 4808 7414 4860
rect 7466 4808 7478 4860
rect 7530 4846 7878 4860
rect 7530 4825 7838 4846
rect 7530 4823 7712 4825
rect 7530 4808 7703 4823
rect 6958 4789 7703 4808
rect 6958 4773 7712 4789
rect 7764 4773 7820 4825
rect 7872 4773 7878 4846
rect 6958 4772 7878 4773
rect 6958 4751 7838 4772
rect 6958 4750 7703 4751
rect 6582 4697 6634 4703
rect 6958 4698 6964 4750
rect 7016 4698 7029 4750
rect 7081 4698 7094 4750
rect 7146 4698 7158 4750
rect 7210 4698 7222 4750
rect 7274 4698 7286 4750
rect 7338 4698 7350 4750
rect 7402 4698 7414 4750
rect 7466 4698 7478 4750
rect 7530 4717 7703 4750
rect 7737 4749 7838 4751
rect 7530 4698 7712 4717
rect 6958 4697 7712 4698
rect 7764 4697 7820 4749
rect 4869 4615 4875 4667
rect 4927 4615 4941 4667
rect 4993 4615 5007 4667
rect 5059 4661 5073 4667
rect 5125 4661 5139 4667
rect 5191 4661 5205 4667
rect 5257 4661 5271 4667
rect 5323 4661 5337 4667
rect 5389 4661 5403 4667
rect 5455 4661 5469 4667
rect 5063 4627 5073 4661
rect 5136 4627 5139 4661
rect 5389 4627 5394 4661
rect 5455 4627 5467 4661
rect 5059 4615 5073 4627
rect 5125 4615 5139 4627
rect 5191 4615 5205 4627
rect 5257 4615 5271 4627
rect 5323 4615 5337 4627
rect 5389 4615 5403 4627
rect 5455 4615 5469 4627
rect 5521 4615 5535 4667
rect 5587 4615 5601 4667
rect 5653 4615 5667 4667
rect 5719 4661 5732 4667
rect 5784 4661 5797 4667
rect 5849 4661 5862 4667
rect 5914 4661 5927 4667
rect 5979 4661 5992 4667
rect 6044 4661 6057 4667
rect 5720 4627 5732 4661
rect 5793 4627 5797 4661
rect 6044 4627 6051 4661
rect 5719 4615 5732 4627
rect 5784 4615 5797 4627
rect 5849 4615 5862 4627
rect 5914 4615 5927 4627
rect 5979 4615 5992 4627
rect 6044 4615 6057 4627
rect 6109 4615 6122 4667
rect 6174 4615 6187 4667
rect 6239 4615 6252 4667
rect 6304 4615 6317 4667
rect 6369 4661 6382 4667
rect 6434 4661 6447 4667
rect 6499 4661 6512 4667
rect 6377 4627 6382 4661
rect 6369 4615 6382 4627
rect 6434 4615 6447 4627
rect 6499 4615 6512 4627
rect 6564 4615 6577 4667
rect 6629 4615 6642 4667
rect 6694 4615 6707 4667
rect 6759 4615 6772 4667
rect 6824 4615 6830 4667
rect 6958 4664 7838 4697
rect 7872 4664 7878 4772
rect 6958 4652 7878 4664
rect 8473 4926 8482 4978
rect 8534 4926 8548 4978
rect 8600 4926 8614 4978
rect 8666 4926 8680 4978
rect 8732 4926 8746 4978
rect 8798 4926 8811 4978
rect 8863 4926 8876 4978
rect 8928 4926 8941 4978
rect 8993 4926 9006 4978
rect 9058 4926 9071 4978
rect 9123 4926 9136 4978
rect 9188 4926 9201 4978
rect 9253 4926 9266 4978
rect 9318 4926 9331 4978
rect 9383 4926 9396 4978
rect 9448 4926 9461 4978
rect 9513 4926 9526 4978
rect 9578 4926 9591 4978
rect 9643 4926 9656 4978
rect 9708 4926 9721 4978
rect 9773 4926 9786 4978
rect 9838 4926 9851 4978
rect 9903 4926 9916 4978
rect 9968 4926 9981 4978
rect 10033 4926 10046 4978
rect 10098 4926 10111 4978
rect 10163 4926 10176 4978
rect 10228 4926 10241 4978
rect 10293 4926 10306 4978
rect 10358 4926 10371 4978
rect 10423 4926 10436 4978
rect 10488 4926 10501 4978
rect 10553 4926 10566 4978
rect 10618 4926 10631 4978
rect 10683 4926 10696 4978
rect 10748 4926 10761 4978
rect 10813 4926 10826 4978
rect 10878 4926 10891 4978
rect 10943 4926 10956 4978
rect 11008 4926 11021 4978
rect 11073 4926 11086 4978
rect 11138 4926 11151 4978
rect 11203 4926 11216 4978
rect 11268 4926 11281 4978
rect 11333 4926 11346 4978
rect 11398 4926 11411 4978
rect 11463 4970 11655 4978
rect 11463 4926 11515 4970
rect 8473 4918 11515 4926
rect 11567 4918 11580 4970
rect 11632 4918 11644 4970
rect 11696 4918 11702 4970
rect 19023 4946 19109 4978
rect 19823 4976 20016 4978
rect 19755 4970 20016 4976
rect 18571 4918 19157 4946
rect 19807 4918 19819 4970
rect 19871 4918 19883 4970
rect 19935 4918 19947 4970
rect 19999 4918 20016 4970
rect 8473 4912 20016 4918
rect 8473 4908 8554 4912
rect 8588 4908 8627 4912
rect 8661 4908 8700 4912
rect 8734 4908 8773 4912
rect 8807 4908 8846 4912
rect 8880 4908 8919 4912
rect 8953 4908 8992 4912
rect 9026 4908 9065 4912
rect 9099 4908 9138 4912
rect 9172 4908 9211 4912
rect 9245 4908 9284 4912
rect 9318 4908 9357 4912
rect 9391 4908 9430 4912
rect 9464 4908 9503 4912
rect 9537 4908 9576 4912
rect 9610 4908 9649 4912
rect 9683 4908 9722 4912
rect 9756 4908 9795 4912
rect 9829 4908 9868 4912
rect 9902 4908 9941 4912
rect 9975 4908 10014 4912
rect 10048 4908 10087 4912
rect 10121 4908 10160 4912
rect 10194 4908 10233 4912
rect 10267 4908 10306 4912
rect 10340 4908 10379 4912
rect 10413 4908 10452 4912
rect 10486 4908 10525 4912
rect 10559 4908 10598 4912
rect 10632 4908 10671 4912
rect 10705 4908 10744 4912
rect 10778 4908 10817 4912
rect 10851 4908 10890 4912
rect 10924 4908 10963 4912
rect 10997 4908 11036 4912
rect 11070 4908 11109 4912
rect 11143 4908 11182 4912
rect 11216 4908 11255 4912
rect 11289 4908 11328 4912
rect 11362 4908 11401 4912
rect 11435 4908 11474 4912
rect 8473 4856 8482 4908
rect 8534 4856 8548 4908
rect 8600 4856 8614 4908
rect 8666 4856 8680 4908
rect 8734 4878 8746 4908
rect 8807 4878 8811 4908
rect 9058 4878 9065 4908
rect 8732 4856 8746 4878
rect 8798 4856 8811 4878
rect 8863 4856 8876 4878
rect 8928 4856 8941 4878
rect 8993 4856 9006 4878
rect 9058 4856 9071 4878
rect 9123 4856 9136 4908
rect 9188 4856 9201 4908
rect 9253 4856 9266 4908
rect 9318 4856 9331 4908
rect 9391 4878 9396 4908
rect 9643 4878 9649 4908
rect 9383 4856 9396 4878
rect 9448 4856 9461 4878
rect 9513 4856 9526 4878
rect 9578 4856 9591 4878
rect 9643 4856 9656 4878
rect 9708 4856 9721 4908
rect 9773 4856 9786 4908
rect 9838 4856 9851 4908
rect 9903 4856 9916 4908
rect 9975 4878 9981 4908
rect 10228 4878 10233 4908
rect 9968 4856 9981 4878
rect 10033 4856 10046 4878
rect 10098 4856 10111 4878
rect 10163 4856 10176 4878
rect 10228 4856 10241 4878
rect 10293 4856 10306 4908
rect 10358 4856 10371 4908
rect 10423 4856 10436 4908
rect 10488 4856 10501 4908
rect 10559 4878 10566 4908
rect 10813 4878 10817 4908
rect 10878 4878 10890 4908
rect 10553 4856 10566 4878
rect 10618 4856 10631 4878
rect 10683 4856 10696 4878
rect 10748 4856 10761 4878
rect 10813 4856 10826 4878
rect 10878 4856 10891 4878
rect 10943 4856 10956 4908
rect 11008 4856 11021 4908
rect 11073 4856 11086 4908
rect 11143 4878 11151 4908
rect 11398 4878 11401 4908
rect 11463 4878 11474 4908
rect 11508 4878 11547 4912
rect 11581 4878 11620 4912
rect 11654 4878 11693 4912
rect 11727 4878 11765 4912
rect 11799 4878 11837 4912
rect 11871 4878 11909 4912
rect 11943 4878 11981 4912
rect 12015 4878 12053 4912
rect 12087 4878 12125 4912
rect 12159 4878 12197 4912
rect 12231 4878 12269 4912
rect 12303 4878 12341 4912
rect 12375 4878 12413 4912
rect 12447 4878 12485 4912
rect 12519 4878 12557 4912
rect 12591 4878 12629 4912
rect 12663 4878 12701 4912
rect 12735 4878 12773 4912
rect 12807 4878 12845 4912
rect 12879 4878 12917 4912
rect 12951 4878 12989 4912
rect 13023 4878 13061 4912
rect 13095 4878 13133 4912
rect 13167 4878 13205 4912
rect 13239 4878 13277 4912
rect 13311 4878 13349 4912
rect 13383 4878 13421 4912
rect 13455 4878 13493 4912
rect 13527 4878 13565 4912
rect 13599 4878 13637 4912
rect 13671 4878 13709 4912
rect 13743 4878 13781 4912
rect 13815 4878 13853 4912
rect 13887 4878 13925 4912
rect 13959 4878 13997 4912
rect 14031 4878 14069 4912
rect 14103 4878 14141 4912
rect 14175 4878 14213 4912
rect 14247 4878 14285 4912
rect 14319 4878 14357 4912
rect 14391 4878 14429 4912
rect 14463 4878 14501 4912
rect 14535 4878 14573 4912
rect 14607 4878 14645 4912
rect 14679 4878 14717 4912
rect 14751 4878 14789 4912
rect 14823 4878 14861 4912
rect 14895 4878 14933 4912
rect 14967 4878 15005 4912
rect 15039 4878 15077 4912
rect 15111 4878 15149 4912
rect 15183 4878 15221 4912
rect 15255 4878 15293 4912
rect 15327 4878 15365 4912
rect 15399 4878 15437 4912
rect 15471 4878 15509 4912
rect 15543 4878 15581 4912
rect 15615 4878 15653 4912
rect 15687 4878 15725 4912
rect 15759 4878 15797 4912
rect 15831 4878 15869 4912
rect 15903 4878 15941 4912
rect 15975 4878 16013 4912
rect 16047 4878 16085 4912
rect 16119 4878 16157 4912
rect 16191 4878 16229 4912
rect 16263 4878 16301 4912
rect 16335 4878 16373 4912
rect 16407 4878 16445 4912
rect 16479 4878 16517 4912
rect 16551 4878 16589 4912
rect 16623 4878 16661 4912
rect 16695 4878 16733 4912
rect 16767 4878 16805 4912
rect 16839 4878 16877 4912
rect 16911 4878 16949 4912
rect 16983 4878 17021 4912
rect 17055 4878 17093 4912
rect 17127 4878 17165 4912
rect 17199 4878 17237 4912
rect 17271 4878 17309 4912
rect 17343 4878 17381 4912
rect 17415 4878 17453 4912
rect 17487 4878 17525 4912
rect 17559 4878 17597 4912
rect 17631 4878 17669 4912
rect 17703 4878 17741 4912
rect 17775 4878 17813 4912
rect 17847 4878 17885 4912
rect 17919 4878 17957 4912
rect 17991 4878 18029 4912
rect 18063 4878 18101 4912
rect 18135 4878 18173 4912
rect 18207 4878 18245 4912
rect 18279 4878 18317 4912
rect 18351 4878 18389 4912
rect 18423 4878 18461 4912
rect 18495 4878 18533 4912
rect 18567 4878 18605 4912
rect 18639 4878 18677 4912
rect 18711 4878 18749 4912
rect 18783 4878 18821 4912
rect 18855 4878 18893 4912
rect 18927 4878 18965 4912
rect 18999 4878 19037 4912
rect 19071 4878 19109 4912
rect 19143 4878 19181 4912
rect 19215 4878 19253 4912
rect 19287 4878 19325 4912
rect 19359 4878 19397 4912
rect 19431 4878 19469 4912
rect 19503 4878 19541 4912
rect 19575 4878 19613 4912
rect 19647 4878 19685 4912
rect 19719 4879 19757 4912
rect 19791 4879 19829 4912
rect 19863 4879 19901 4912
rect 19935 4879 20016 4912
rect 19719 4878 19755 4879
rect 11138 4856 11151 4878
rect 11203 4856 11216 4878
rect 11268 4856 11281 4878
rect 11333 4856 11346 4878
rect 11398 4856 11411 4878
rect 11463 4876 19755 4878
rect 11463 4856 11515 4876
rect 8473 4840 8534 4856
tri 8534 4840 8550 4856 nw
tri 8817 4840 8833 4856 ne
rect 8833 4840 8941 4856
tri 8941 4840 8957 4856 nw
tri 11260 4840 11276 4856 ne
rect 11276 4840 11393 4856
tri 11393 4840 11409 4856 nw
tri 11475 4840 11491 4856 ne
rect 11491 4840 11515 4856
rect 8473 4838 8525 4840
rect 8473 4806 8482 4838
rect 8516 4806 8525 4838
tri 8525 4831 8534 4840 nw
tri 8833 4831 8842 4840 ne
rect 8842 4831 8927 4840
tri 8842 4820 8853 4831 ne
rect 8853 4826 8927 4831
tri 8927 4826 8941 4840 nw
tri 11276 4826 11290 4840 ne
rect 8853 4820 8921 4826
tri 8921 4820 8927 4826 nw
rect 8473 4730 8482 4754
rect 8516 4730 8525 4754
rect 8473 4723 8525 4730
rect 8473 4665 8482 4671
tri 8473 4662 8476 4665 ne
rect 6958 4618 7066 4652
rect 7100 4618 7150 4652
rect 7184 4618 7235 4652
rect 7269 4618 7320 4652
rect 7354 4618 7405 4652
rect 7439 4618 7490 4652
rect 7524 4624 7878 4652
rect 8476 4656 8482 4665
rect 8516 4665 8525 4671
rect 8516 4664 8524 4665
tri 8524 4664 8525 4665 nw
rect 8708 4808 8754 4820
tri 8853 4812 8861 4820 ne
rect 8708 4774 8714 4808
rect 8748 4774 8754 4808
rect 8708 4736 8754 4774
rect 8708 4702 8714 4736
rect 8748 4702 8754 4736
rect 8708 4664 8754 4702
rect 8861 4808 8913 4820
tri 8913 4812 8921 4820 nw
rect 8861 4806 8870 4808
rect 8904 4806 8913 4808
rect 8861 4736 8913 4754
rect 8861 4723 8870 4736
rect 8904 4723 8913 4736
rect 8861 4665 8913 4671
tri 8861 4664 8862 4665 ne
rect 8862 4664 8912 4665
tri 8912 4664 8913 4665 nw
rect 9020 4808 9066 4820
rect 9020 4774 9026 4808
rect 9060 4774 9066 4808
rect 9020 4736 9066 4774
rect 9020 4702 9026 4736
rect 9060 4702 9066 4736
rect 9020 4664 9066 4702
rect 8516 4656 8522 4664
tri 8522 4662 8524 4664 nw
rect 7524 4618 7838 4624
rect 3769 4582 3829 4590
tri 3829 4582 3837 4590 sw
tri 4259 4582 4267 4590 se
rect 4267 4582 4344 4590
tri 4344 4582 4352 4590 sw
tri 4769 4582 4777 4590 se
rect 4777 4582 4839 4590
rect 3769 4576 3837 4582
tri 3837 4576 3843 4582 sw
tri 4253 4576 4259 4582 se
rect 4259 4576 4352 4582
tri 4352 4576 4358 4582 sw
tri 4763 4576 4769 4582 se
rect 4769 4576 4839 4582
rect 3769 4530 4839 4576
rect 6958 4590 7838 4618
rect 7872 4590 7878 4624
tri 8204 4620 8209 4625 se
rect 8209 4620 8215 4625
rect 6958 4550 7878 4590
rect 3001 4529 3073 4530
tri 3073 4529 3074 4530 nw
tri 3990 4529 3991 4530 ne
rect 3991 4529 4092 4530
rect 454 4502 507 4513
rect 506 4450 507 4502
rect 3001 4516 3060 4529
tri 3060 4516 3073 4529 nw
tri 3991 4516 4004 4529 ne
rect 4004 4516 4092 4529
tri 4092 4516 4106 4530 nw
tri 6944 4516 6958 4530 se
rect 6958 4516 7838 4550
rect 7872 4516 7878 4550
rect 3001 4508 3052 4516
tri 3052 4508 3060 4516 nw
tri 4004 4508 4012 4516 ne
rect 4012 4508 4084 4516
tri 4084 4508 4092 4516 nw
tri 6936 4508 6944 4516 se
rect 6944 4508 7878 4516
rect 3001 4505 3049 4508
tri 3049 4505 3052 4508 nw
tri 4012 4505 4015 4508 ne
rect 454 4438 467 4450
rect 501 4438 507 4450
rect 454 4420 507 4438
rect 506 4368 507 4420
rect 454 4363 467 4368
rect 501 4363 507 4368
rect 454 4338 507 4363
rect 506 4286 507 4338
rect 454 4256 507 4286
rect 641 4497 1670 4498
rect 641 4492 952 4497
rect 1004 4492 1044 4497
rect 1096 4492 1135 4497
rect 1187 4492 1670 4497
tri 1670 4492 1676 4498 sw
rect 641 4486 928 4492
rect 641 4452 660 4486
rect 694 4458 928 4486
rect 1004 4458 1006 4492
rect 1040 4458 1044 4492
rect 1118 4458 1135 4492
rect 1196 4458 1239 4492
rect 1273 4458 1316 4492
rect 1350 4458 1393 4492
rect 1427 4458 1470 4492
rect 1504 4458 1547 4492
rect 1581 4458 1624 4492
rect 1658 4486 1676 4492
tri 1676 4486 1682 4492 sw
rect 1658 4458 1682 4486
rect 694 4452 952 4458
rect 641 4445 952 4452
rect 1004 4445 1044 4458
rect 1096 4445 1135 4458
rect 1187 4452 1682 4458
tri 1682 4452 1716 4486 sw
rect 1187 4446 1716 4452
tri 1716 4446 1722 4452 sw
rect 1777 4446 1783 4498
rect 1835 4446 1850 4498
rect 1902 4446 1917 4498
rect 1969 4486 1983 4498
rect 2035 4486 2049 4498
rect 2101 4486 2115 4498
rect 2167 4486 2181 4498
rect 2233 4486 2247 4498
rect 1975 4452 1983 4486
rect 2167 4452 2169 4486
rect 2233 4452 2244 4486
rect 1969 4446 1983 4452
rect 2035 4446 2049 4452
rect 2101 4446 2115 4452
rect 2167 4446 2181 4452
rect 2233 4446 2247 4452
rect 2299 4446 2313 4498
rect 2365 4446 2379 4498
rect 2431 4446 2445 4498
rect 2497 4486 2511 4498
rect 2563 4486 2577 4498
rect 2629 4486 2643 4498
rect 2695 4486 2709 4498
rect 2761 4486 2775 4498
rect 2503 4452 2511 4486
rect 2761 4452 2769 4486
rect 2497 4446 2511 4452
rect 2563 4446 2577 4452
rect 2629 4446 2643 4452
rect 2695 4446 2709 4452
rect 2761 4446 2775 4452
rect 2827 4446 2841 4498
rect 2893 4446 2907 4498
rect 2959 4446 2965 4498
rect 1187 4445 1722 4446
rect 641 4441 1722 4445
tri 1722 4441 1727 4446 sw
rect 641 4434 1727 4441
tri 1727 4434 1734 4441 sw
rect 641 4417 1734 4434
rect 641 4404 952 4417
rect 641 4370 660 4404
rect 694 4393 952 4404
rect 694 4370 871 4393
rect 641 4359 871 4370
rect 905 4365 952 4393
rect 1004 4365 1044 4417
rect 1096 4365 1135 4417
rect 1187 4414 1734 4417
tri 1734 4414 1754 4434 sw
rect 1187 4413 1754 4414
tri 1754 4413 1755 4414 sw
rect 1187 4365 1665 4413
rect 905 4361 1665 4365
rect 1717 4393 1746 4413
rect 1717 4361 1727 4393
rect 1798 4361 1804 4413
rect 2230 4407 2282 4413
rect 905 4359 1727 4361
rect 1761 4359 1804 4361
rect 641 4337 1804 4359
rect 641 4321 952 4337
rect 641 4287 660 4321
rect 694 4287 871 4321
rect 905 4287 952 4321
rect 641 4285 952 4287
rect 1004 4285 1044 4337
rect 1096 4285 1135 4337
rect 1187 4285 1665 4337
rect 1717 4321 1746 4337
rect 1717 4287 1727 4321
rect 1717 4285 1746 4287
rect 1798 4285 1804 4337
rect 641 4275 1804 4285
rect 1977 4393 2023 4405
rect 1977 4359 1983 4393
rect 2017 4359 2023 4393
rect 1977 4321 2023 4359
rect 1977 4287 1983 4321
rect 2017 4287 2023 4321
rect 506 4204 507 4256
rect 454 4174 507 4204
tri 1969 4189 1977 4197 se
rect 1977 4189 2023 4287
rect 2742 4407 2794 4413
rect 2230 4343 2282 4355
rect 2230 4287 2239 4291
rect 2273 4287 2282 4291
rect 2230 4275 2282 4287
rect 2489 4393 2535 4405
rect 2489 4359 2495 4393
rect 2529 4359 2535 4393
rect 2489 4321 2535 4359
rect 2489 4287 2495 4321
rect 2529 4287 2535 4321
tri 2475 4198 2489 4212 se
rect 2489 4198 2535 4287
rect 2742 4343 2794 4355
rect 2742 4287 2751 4291
rect 2785 4287 2794 4291
rect 2742 4275 2794 4287
rect 3001 4393 3047 4505
tri 3047 4503 3049 4505 nw
rect 3083 4446 3089 4498
rect 3141 4446 3158 4498
rect 3210 4446 3227 4498
rect 3279 4486 3296 4498
rect 3348 4486 3365 4498
rect 3417 4486 3434 4498
rect 3486 4486 3502 4498
rect 3554 4486 3570 4498
rect 3285 4452 3296 4486
rect 3363 4452 3365 4486
rect 3554 4452 3563 4486
rect 3279 4446 3296 4452
rect 3348 4446 3365 4452
rect 3417 4446 3434 4452
rect 3486 4446 3502 4452
rect 3554 4446 3570 4452
rect 3622 4446 3638 4498
rect 3690 4446 3706 4498
rect 3758 4446 3764 4498
rect 3820 4486 3975 4492
rect 3820 4452 3832 4486
rect 3866 4452 3929 4486
rect 3963 4452 3975 4486
rect 3820 4446 3975 4452
tri 3861 4441 3866 4446 ne
rect 3866 4441 3962 4446
tri 3962 4441 3967 4446 nw
tri 3866 4434 3873 4441 ne
rect 3873 4434 3955 4441
tri 3955 4434 3962 4441 nw
tri 3873 4418 3889 4434 ne
rect 3001 4359 3007 4393
rect 3041 4359 3047 4393
rect 3001 4321 3047 4359
rect 3001 4287 3007 4321
rect 3041 4287 3047 4321
rect 3254 4407 3306 4413
rect 3766 4407 3818 4413
rect 3254 4343 3306 4355
rect 3254 4287 3263 4291
rect 3297 4287 3306 4291
rect 3001 4286 3047 4287
tri 3047 4286 3048 4287 sw
rect 3001 4275 3048 4286
tri 3048 4275 3059 4286 sw
rect 3254 4275 3306 4287
rect 3513 4393 3559 4405
rect 3513 4359 3519 4393
rect 3553 4359 3559 4393
rect 3513 4321 3559 4359
rect 3513 4287 3519 4321
rect 3553 4287 3559 4321
rect 3766 4343 3818 4355
rect 3766 4287 3775 4291
rect 3809 4287 3818 4291
rect 3513 4286 3559 4287
tri 3559 4286 3560 4287 sw
rect 3513 4285 3560 4286
tri 3560 4285 3561 4286 sw
rect 3513 4275 3561 4285
tri 3561 4275 3571 4285 sw
rect 3766 4275 3818 4287
rect 3889 4407 3941 4434
tri 3941 4420 3955 4434 nw
rect 3889 4343 3941 4355
rect 3889 4285 3941 4291
rect 4015 4393 4081 4508
tri 4081 4505 4084 4508 nw
tri 6933 4505 6936 4508 se
rect 6936 4505 7878 4508
tri 6927 4499 6933 4505 se
rect 6933 4499 7878 4505
rect 6668 4498 6801 4499
tri 6926 4498 6927 4499 se
rect 6927 4498 7878 4499
rect 4121 4446 4127 4498
rect 4179 4446 4218 4498
rect 4270 4446 4276 4498
rect 4332 4486 4497 4492
rect 4332 4452 4344 4486
rect 4378 4452 4451 4486
rect 4485 4452 4497 4486
rect 4332 4446 4497 4452
rect 4588 4446 4594 4498
rect 4646 4446 4659 4498
rect 4711 4446 4724 4498
rect 4776 4486 4789 4498
rect 4841 4486 4853 4498
rect 4905 4486 4917 4498
rect 4969 4486 4981 4498
rect 4784 4452 4789 4486
rect 4969 4452 4975 4486
rect 4776 4446 4789 4452
rect 4841 4446 4853 4452
rect 4905 4446 4917 4452
rect 4969 4446 4981 4452
rect 5033 4446 5045 4498
rect 5097 4446 5109 4498
rect 5161 4446 5173 4498
rect 5225 4486 5237 4498
rect 5289 4486 5301 4498
rect 5353 4486 5365 4498
rect 5417 4486 5429 4498
rect 5233 4452 5237 4486
rect 5417 4452 5421 4486
rect 5225 4446 5237 4452
rect 5289 4446 5301 4452
rect 5353 4446 5365 4452
rect 5417 4446 5429 4452
rect 5481 4446 5493 4498
rect 5545 4446 5557 4498
rect 5609 4446 5621 4498
rect 5673 4486 5685 4498
rect 5737 4486 5749 4498
rect 5801 4486 5813 4498
rect 5865 4486 5877 4498
rect 5929 4486 5941 4498
rect 5677 4452 5685 4486
rect 5929 4452 5939 4486
rect 5673 4446 5685 4452
rect 5737 4446 5749 4452
rect 5801 4446 5813 4452
rect 5865 4446 5877 4452
rect 5929 4446 5941 4452
rect 5993 4446 6005 4498
rect 6057 4446 6069 4498
rect 6121 4446 6133 4498
rect 6185 4486 6197 4498
rect 6249 4486 6261 4498
rect 6313 4486 6325 4498
rect 6377 4486 6389 4498
rect 6195 4452 6197 4486
rect 6377 4452 6383 4486
rect 6185 4446 6197 4452
rect 6249 4446 6261 4452
rect 6313 4446 6325 4452
rect 6377 4446 6389 4452
rect 6441 4446 6453 4498
rect 6505 4446 6517 4498
rect 6569 4446 6577 4498
rect 6668 4446 6674 4498
rect 6726 4446 6743 4498
rect 6795 4446 6801 4498
tri 6920 4492 6926 4498 se
rect 6926 4492 7878 4498
tri 6886 4458 6920 4492 se
rect 6920 4458 7066 4492
rect 7100 4458 7138 4492
rect 7172 4458 7210 4492
rect 7244 4458 7282 4492
rect 7316 4458 7355 4492
rect 7389 4458 7428 4492
rect 7462 4458 7501 4492
rect 7535 4458 7574 4492
rect 7608 4458 7647 4492
rect 7681 4475 7878 4492
rect 7681 4458 7838 4475
tri 6880 4452 6886 4458 se
rect 6886 4452 7838 4458
tri 4368 4441 4373 4446 ne
rect 4373 4441 4481 4446
tri 4481 4441 4486 4446 nw
tri 4373 4434 4380 4441 ne
rect 4380 4434 4474 4441
tri 4474 4434 4481 4441 nw
tri 4380 4414 4400 4434 ne
rect 4400 4414 4454 4434
tri 4454 4414 4474 4434 nw
tri 4400 4413 4401 4414 ne
rect 4015 4359 4031 4393
rect 4065 4359 4081 4393
rect 4015 4321 4081 4359
rect 4015 4287 4031 4321
rect 4065 4287 4081 4321
rect 4278 4407 4330 4413
rect 4278 4343 4330 4355
tri 4081 4287 4090 4296 sw
rect 4278 4287 4287 4291
rect 4321 4287 4330 4291
rect 4015 4286 4090 4287
tri 4090 4286 4091 4287 sw
rect 4015 4285 4091 4286
tri 4091 4285 4092 4286 sw
rect 4015 4275 4092 4285
tri 4092 4275 4102 4285 sw
rect 4278 4275 4330 4287
rect 4401 4407 4453 4414
tri 4453 4413 4454 4414 nw
rect 4790 4407 4842 4413
rect 4401 4343 4453 4355
rect 4401 4285 4453 4291
rect 4537 4393 4583 4405
rect 4537 4359 4543 4393
rect 4577 4359 4583 4393
rect 4537 4321 4583 4359
rect 4537 4287 4543 4321
rect 4577 4287 4583 4321
rect 5302 4407 5354 4413
rect 4790 4343 4842 4355
tri 4583 4287 4597 4301 sw
rect 5049 4393 5095 4405
rect 5049 4359 5055 4393
rect 5089 4359 5095 4393
rect 5049 4321 5095 4359
rect 4790 4287 4799 4291
rect 4833 4287 4842 4291
tri 5035 4287 5049 4301 se
rect 5049 4287 5055 4321
rect 5089 4287 5095 4321
rect 4537 4286 4597 4287
tri 4597 4286 4598 4287 sw
rect 4537 4275 4598 4286
tri 4598 4275 4609 4286 sw
rect 4790 4275 4842 4287
tri 5034 4286 5035 4287 se
rect 5035 4286 5095 4287
tri 5023 4275 5034 4286 se
rect 5034 4275 5095 4286
rect 5814 4407 5866 4413
rect 5302 4343 5354 4355
rect 5302 4287 5311 4291
rect 5345 4287 5354 4291
rect 5302 4275 5354 4287
rect 5561 4393 5607 4405
rect 5561 4359 5567 4393
rect 5601 4359 5607 4393
rect 5561 4321 5607 4359
rect 5561 4287 5567 4321
rect 5601 4287 5607 4321
rect 3001 4270 3059 4275
tri 3059 4270 3064 4275 sw
rect 3513 4270 3571 4275
tri 3571 4270 3576 4275 sw
rect 4015 4270 4102 4275
tri 4102 4270 4107 4275 sw
rect 4537 4270 4609 4275
tri 4609 4270 4614 4275 sw
tri 5018 4270 5023 4275 se
rect 5023 4270 5095 4275
rect 3001 4265 3064 4270
tri 3064 4265 3069 4270 sw
rect 3513 4265 3576 4270
tri 3576 4265 3581 4270 sw
rect 4015 4265 4107 4270
tri 4107 4265 4112 4270 sw
rect 4537 4265 4614 4270
tri 4614 4265 4619 4270 sw
tri 5013 4265 5018 4270 se
rect 5018 4265 5095 4270
rect 3001 4263 3069 4265
tri 3069 4263 3071 4265 sw
rect 3513 4263 3581 4265
tri 3581 4263 3583 4265 sw
rect 4015 4263 4112 4265
tri 4112 4263 4114 4265 sw
rect 4537 4263 4619 4265
tri 4619 4263 4621 4265 sw
tri 5011 4263 5013 4265 se
rect 5013 4263 5095 4265
rect 3001 4254 3071 4263
tri 3071 4254 3080 4263 sw
rect 3513 4254 3583 4263
tri 3583 4254 3592 4263 sw
rect 4015 4254 4114 4263
tri 4114 4254 4123 4263 sw
rect 4537 4254 4621 4263
tri 4621 4254 4630 4263 sw
tri 5002 4254 5011 4263 se
rect 5011 4254 5095 4263
rect 3001 4250 3080 4254
tri 3080 4250 3084 4254 sw
rect 3513 4250 3592 4254
tri 3592 4250 3596 4254 sw
rect 4015 4250 4123 4254
tri 4123 4250 4127 4254 sw
rect 4537 4250 4630 4254
tri 4630 4250 4634 4254 sw
tri 4998 4250 5002 4254 se
rect 5002 4250 5095 4254
rect 3001 4247 3084 4250
tri 3084 4247 3087 4250 sw
rect 3513 4247 3596 4250
tri 3596 4247 3599 4250 sw
rect 4015 4247 4127 4250
tri 4127 4247 4130 4250 sw
rect 4537 4247 4634 4250
tri 4634 4247 4637 4250 sw
tri 4995 4247 4998 4250 se
rect 4998 4247 5095 4250
tri 2535 4198 2549 4212 sw
tri 2474 4197 2475 4198 se
rect 2475 4197 2549 4198
tri 2023 4189 2031 4197 sw
tri 2466 4189 2474 4197 se
rect 2474 4195 2549 4197
tri 2549 4195 2552 4198 sw
rect 3001 4195 3007 4247
rect 3059 4195 3071 4247
rect 3123 4195 3129 4247
rect 3513 4195 3519 4247
rect 3571 4195 3583 4247
rect 3635 4195 3641 4247
rect 4015 4195 4365 4247
rect 4417 4195 4429 4247
rect 4481 4195 4487 4247
rect 4537 4195 4973 4247
rect 5025 4195 5037 4247
rect 5089 4195 5095 4247
tri 5559 4195 5561 4197 se
rect 5561 4195 5607 4287
rect 6326 4407 6378 4413
rect 5814 4343 5866 4355
rect 5814 4287 5823 4291
rect 5857 4287 5866 4291
rect 5814 4275 5866 4287
rect 6073 4393 6119 4405
rect 6073 4359 6079 4393
rect 6113 4359 6119 4393
rect 6073 4321 6119 4359
rect 6073 4287 6079 4321
rect 6113 4287 6119 4321
tri 6070 4198 6073 4201 se
rect 6073 4198 6119 4287
rect 6326 4343 6378 4355
rect 6326 4287 6335 4291
rect 6369 4287 6378 4291
rect 6326 4275 6378 4287
rect 6585 4393 6631 4405
rect 6585 4359 6591 4393
rect 6625 4359 6631 4393
rect 6585 4321 6631 4359
rect 6585 4287 6591 4321
rect 6625 4287 6631 4321
tri 6583 4204 6585 4206 se
rect 6585 4204 6631 4287
tri 6580 4201 6583 4204 se
rect 6583 4201 6631 4204
tri 6119 4198 6122 4201 sw
tri 6577 4198 6580 4201 se
rect 6580 4198 6631 4201
tri 6069 4197 6070 4198 se
rect 6070 4197 6122 4198
tri 5607 4195 5609 4197 sw
tri 6067 4195 6069 4197 se
rect 6069 4195 6122 4197
rect 2474 4189 2552 4195
tri 2552 4189 2558 4195 sw
tri 5553 4189 5559 4195 se
rect 5559 4189 5609 4195
tri 5609 4189 5615 4195 sw
tri 6061 4189 6067 4195 se
rect 6067 4189 6122 4195
tri 6122 4189 6131 4198 sw
tri 6568 4189 6577 4198 se
rect 6577 4189 6631 4198
tri 1955 4175 1969 4189 se
rect 1969 4175 2031 4189
tri 2031 4175 2045 4189 sw
tri 2452 4175 2466 4189 se
rect 2466 4175 2558 4189
tri 2558 4175 2572 4189 sw
tri 5539 4175 5553 4189 se
rect 5553 4175 5615 4189
tri 5615 4175 5629 4189 sw
tri 6047 4175 6061 4189 se
rect 6061 4175 6131 4189
tri 6131 4175 6145 4189 sw
tri 6554 4175 6568 4189 se
rect 6568 4175 6631 4189
rect 506 4122 507 4174
tri 1947 4167 1955 4175 se
rect 1955 4171 2045 4175
tri 2045 4171 2049 4175 sw
tri 2448 4171 2452 4175 se
rect 2452 4171 2572 4175
tri 2572 4171 2576 4175 sw
tri 5535 4171 5539 4175 se
rect 5539 4171 5629 4175
tri 5629 4171 5633 4175 sw
tri 6043 4171 6047 4175 se
rect 6047 4171 6145 4175
rect 1955 4167 2049 4171
tri 2049 4167 2053 4171 sw
tri 2444 4167 2448 4171 se
rect 2448 4167 2454 4171
rect 454 4097 507 4122
rect 454 4092 467 4097
rect 501 4092 507 4097
rect 506 4040 507 4092
rect 699 4161 2454 4167
rect 751 4119 2454 4161
rect 2506 4119 2518 4171
rect 2570 4167 2576 4171
tri 2576 4167 2580 4171 sw
tri 5531 4167 5535 4171 se
rect 5535 4167 5633 4171
tri 5633 4167 5637 4171 sw
tri 6039 4167 6043 4171 se
rect 6043 4167 6145 4171
tri 6145 4167 6153 4175 sw
tri 6546 4167 6554 4175 se
rect 6554 4167 6631 4175
rect 2570 4119 5908 4167
rect 751 4115 781 4119
tri 781 4115 785 4119 nw
tri 5898 4115 5902 4119 ne
rect 5902 4115 5908 4119
rect 5960 4115 5972 4167
rect 6024 4119 6631 4167
rect 6668 4250 6801 4446
tri 6869 4441 6880 4452 se
rect 6880 4441 7838 4452
rect 7872 4441 7878 4475
tri 6862 4434 6869 4441 se
rect 6869 4434 7878 4441
tri 6842 4414 6862 4434 se
rect 6862 4414 7878 4434
tri 6841 4413 6842 4414 se
rect 6842 4413 7878 4414
rect 6841 4359 6847 4413
rect 6899 4361 6953 4413
rect 7005 4361 7058 4413
rect 7110 4361 7163 4413
rect 7215 4361 7268 4413
rect 7320 4361 7373 4413
rect 7425 4361 7478 4413
rect 7530 4361 7597 4413
rect 7649 4393 7705 4413
rect 7757 4400 7878 4413
rect 7649 4361 7703 4393
rect 7757 4366 7838 4400
rect 7872 4366 7878 4400
rect 7757 4361 7878 4366
rect 6881 4359 7703 4361
rect 7737 4359 7878 4361
rect 6841 4337 7878 4359
rect 6841 4285 6847 4337
rect 6899 4285 6953 4337
rect 7005 4285 7058 4337
rect 7110 4285 7163 4337
rect 7215 4285 7268 4337
rect 7320 4285 7373 4337
rect 7425 4285 7478 4337
rect 7530 4285 7597 4337
rect 7649 4321 7705 4337
rect 7757 4325 7878 4337
rect 7649 4287 7703 4321
rect 7757 4291 7838 4325
rect 7872 4291 7878 4325
rect 7649 4285 7705 4287
rect 7757 4285 7878 4291
rect 6841 4275 7878 4285
tri 6920 4270 6925 4275 ne
rect 6925 4270 7878 4275
tri 6925 4265 6930 4270 ne
rect 6930 4265 7878 4270
tri 6930 4263 6932 4265 ne
rect 6932 4263 7878 4265
rect 8103 4614 8155 4620
tri 8202 4618 8204 4620 se
rect 8204 4618 8215 4620
tri 8200 4616 8202 4618 se
rect 8202 4616 8215 4618
tri 8199 4615 8200 4616 se
rect 8200 4615 8215 4616
tri 8195 4611 8199 4615 se
rect 8199 4611 8215 4615
rect 8103 4550 8155 4562
tri 7878 4263 7879 4264 sw
tri 6932 4254 6941 4263 ne
rect 6941 4254 7879 4263
tri 7879 4254 7888 4263 sw
tri 6941 4250 6945 4254 ne
rect 6945 4250 7888 4254
rect 6668 4198 6674 4250
rect 6726 4198 6743 4250
rect 6795 4198 6801 4250
tri 6945 4216 6979 4250 ne
rect 6979 4216 7838 4250
rect 7872 4248 7888 4250
tri 7888 4248 7894 4254 sw
rect 7872 4246 7894 4248
tri 7894 4246 7896 4248 sw
rect 7872 4232 7896 4246
tri 7896 4232 7910 4246 sw
rect 7872 4216 8059 4232
tri 6979 4215 6980 4216 ne
rect 6024 4115 6030 4119
tri 6030 4115 6034 4119 nw
rect 751 4114 780 4115
tri 780 4114 781 4115 nw
rect 751 4109 766 4114
rect 699 4100 766 4109
tri 766 4100 780 4114 nw
rect 699 4097 751 4100
rect 454 4022 507 4040
rect 454 4010 467 4022
rect 501 4010 507 4022
rect 506 3958 507 4010
rect 454 3947 507 3958
rect 454 3928 467 3947
rect 501 3928 507 3947
rect 617 4057 669 4063
tri 751 4085 766 4100 nw
rect 699 4039 751 4045
rect 1258 4027 1264 4079
rect 1316 4027 1328 4079
rect 1380 4027 3519 4079
rect 3571 4027 3583 4079
rect 3635 4027 4973 4079
rect 5025 4027 5037 4079
rect 5089 4027 5095 4079
rect 617 3993 669 4005
tri 669 3991 699 4021 sw
rect 669 3990 699 3991
tri 699 3990 700 3991 sw
rect 669 3987 700 3990
tri 700 3987 703 3990 sw
rect 669 3941 3007 3987
rect 617 3935 3007 3941
rect 3059 3935 3071 3987
rect 3123 3935 5607 3987
rect 506 3876 507 3928
tri 5532 3916 5551 3935 ne
rect 5551 3916 5607 3935
tri 5551 3910 5557 3916 ne
rect 5557 3910 5607 3916
tri 5557 3906 5561 3910 ne
rect 454 3872 507 3876
rect 454 3846 467 3872
rect 501 3846 507 3872
rect 506 3794 507 3846
rect 1977 3853 2454 3903
rect 1977 3851 2055 3853
tri 2055 3851 2057 3853 nw
tri 2446 3851 2448 3853 ne
rect 2448 3851 2454 3853
rect 2506 3851 2518 3903
rect 2570 3853 3047 3903
rect 2570 3851 2576 3853
tri 2576 3851 2578 3853 nw
tri 2973 3851 2975 3853 ne
rect 2975 3851 3047 3853
rect 1977 3841 2045 3851
tri 2045 3841 2055 3851 nw
tri 2448 3841 2458 3851 ne
rect 2458 3841 2566 3851
tri 2566 3841 2576 3851 nw
tri 2975 3841 2985 3851 ne
rect 2985 3841 3047 3851
rect 1977 3838 2042 3841
tri 2042 3838 2045 3841 nw
tri 2458 3838 2461 3841 ne
rect 2461 3838 2563 3841
tri 2563 3838 2566 3841 nw
tri 2985 3838 2988 3841 ne
rect 2988 3838 3047 3841
rect 1977 3825 2029 3838
tri 2029 3825 2042 3838 nw
tri 2461 3825 2474 3838 ne
rect 2474 3825 2550 3838
tri 2550 3825 2563 3838 nw
tri 2988 3825 3001 3838 ne
rect 454 3764 467 3794
rect 501 3764 507 3794
rect 506 3712 507 3764
rect 454 3688 467 3712
rect 501 3688 507 3712
rect 454 3681 507 3688
rect 506 3629 507 3681
rect 454 3613 467 3629
rect 501 3613 507 3629
rect 641 3815 1767 3825
rect 641 3813 952 3815
rect 641 3779 660 3813
rect 694 3779 871 3813
rect 905 3779 952 3813
rect 641 3763 952 3779
rect 1004 3763 1044 3815
rect 1096 3763 1135 3815
rect 1187 3763 1624 3815
rect 1676 3763 1709 3815
rect 1761 3763 1767 3815
rect 641 3741 1767 3763
rect 641 3731 871 3741
rect 641 3697 660 3731
rect 694 3707 871 3731
rect 905 3739 1727 3741
rect 905 3735 1624 3739
rect 905 3707 952 3735
rect 694 3697 952 3707
rect 641 3683 952 3697
rect 1004 3683 1044 3735
rect 1096 3683 1135 3735
rect 1187 3687 1624 3735
rect 1676 3687 1709 3739
rect 1761 3687 1767 3741
rect 1977 3820 2024 3825
tri 2024 3820 2029 3825 nw
rect 1977 3813 2023 3820
tri 2023 3819 2024 3820 nw
rect 1977 3779 1983 3813
rect 2017 3779 2023 3813
rect 1977 3741 2023 3779
rect 1977 3707 1983 3741
rect 2017 3707 2023 3741
rect 1977 3695 2023 3707
rect 2230 3813 2282 3825
tri 2474 3820 2479 3825 ne
rect 2479 3820 2545 3825
tri 2545 3820 2550 3825 nw
tri 2479 3818 2481 3820 ne
rect 2481 3818 2543 3820
tri 2543 3818 2545 3820 nw
tri 2481 3813 2486 3818 ne
rect 2486 3813 2538 3818
tri 2538 3813 2543 3818 nw
rect 2742 3813 2794 3825
rect 2230 3809 2239 3813
rect 2273 3809 2282 3813
tri 2486 3810 2489 3813 ne
rect 2230 3745 2282 3757
rect 2489 3779 2495 3813
rect 2529 3779 2535 3813
tri 2535 3810 2538 3813 nw
rect 2489 3741 2535 3779
rect 2489 3707 2495 3741
rect 2529 3707 2535 3741
rect 2489 3695 2535 3707
rect 2742 3809 2751 3813
rect 2785 3809 2794 3813
rect 2742 3745 2794 3757
rect 2230 3687 2282 3693
rect 3001 3813 3047 3838
rect 3513 3853 3519 3905
rect 3571 3853 3583 3905
rect 3635 3853 4071 3905
rect 3513 3851 3591 3853
tri 3591 3851 3593 3853 nw
tri 3991 3851 3993 3853 ne
rect 3993 3851 4071 3853
rect 3513 3845 3585 3851
tri 3585 3845 3591 3851 nw
tri 3993 3845 3999 3851 ne
rect 3999 3845 4071 3851
rect 4359 3853 4365 3905
rect 4417 3853 4429 3905
rect 4481 3853 4593 3905
rect 4966 3853 4973 3905
rect 5025 3853 5037 3905
rect 5089 3853 5095 3905
rect 4359 3845 4593 3853
rect 3513 3841 3581 3845
tri 3581 3841 3585 3845 nw
tri 3999 3841 4003 3845 ne
rect 4003 3841 4071 3845
tri 4501 3841 4505 3845 ne
rect 4505 3841 4593 3845
tri 5015 3841 5027 3853 ne
rect 5027 3841 5095 3853
rect 3513 3838 3578 3841
tri 3578 3838 3581 3841 nw
tri 4003 3838 4006 3841 ne
rect 4006 3838 4071 3841
tri 4505 3838 4508 3841 ne
rect 4508 3838 4593 3841
tri 5027 3838 5030 3841 ne
rect 5030 3838 5095 3841
rect 3513 3825 3565 3838
tri 3565 3825 3578 3838 nw
tri 4006 3825 4019 3838 ne
rect 4019 3825 4071 3838
tri 4508 3825 4521 3838 ne
rect 4521 3825 4593 3838
tri 5030 3825 5043 3838 ne
rect 5043 3825 5095 3838
rect 3001 3779 3007 3813
rect 3041 3779 3047 3813
rect 3001 3741 3047 3779
rect 3001 3707 3007 3741
rect 3041 3707 3047 3741
rect 3001 3695 3047 3707
rect 3254 3813 3307 3825
rect 3254 3809 3263 3813
rect 3297 3809 3307 3813
rect 3306 3757 3307 3809
rect 3254 3745 3307 3757
rect 2742 3687 2794 3693
rect 3306 3693 3307 3745
rect 3513 3820 3560 3825
tri 3560 3820 3565 3825 nw
rect 3513 3813 3559 3820
tri 3559 3819 3560 3820 nw
rect 3513 3779 3519 3813
rect 3553 3779 3559 3813
rect 3513 3741 3559 3779
rect 3513 3707 3519 3741
rect 3553 3707 3559 3741
rect 3513 3695 3559 3707
rect 3765 3813 3818 3825
tri 4019 3820 4024 3825 ne
rect 4024 3820 4071 3825
tri 4024 3819 4025 3820 ne
rect 3765 3809 3775 3813
rect 3809 3809 3818 3813
rect 3765 3757 3766 3809
rect 3765 3745 3818 3757
rect 3254 3687 3307 3693
rect 3765 3693 3766 3745
rect 4025 3813 4071 3820
rect 4025 3779 4031 3813
rect 4065 3779 4071 3813
rect 4025 3741 4071 3779
rect 4025 3707 4031 3741
rect 4065 3707 4071 3741
rect 4025 3695 4071 3707
rect 4145 3809 4197 3815
rect 4145 3745 4197 3757
rect 3765 3687 3818 3693
rect 1187 3684 1764 3687
tri 1764 3684 1767 3687 nw
rect 1187 3683 1734 3684
rect 641 3655 1734 3683
rect 641 3648 952 3655
rect 454 3598 507 3613
rect 506 3546 507 3598
rect 454 3538 467 3546
rect 501 3538 507 3546
rect 454 3515 507 3538
rect 506 3463 507 3515
rect 535 3617 587 3623
rect 641 3614 660 3648
rect 694 3642 952 3648
rect 1004 3642 1044 3655
rect 1096 3642 1135 3655
rect 1187 3654 1734 3655
tri 1734 3654 1764 3684 nw
tri 4115 3654 4145 3684 se
rect 4145 3654 4197 3693
rect 4278 3813 4331 3825
tri 4521 3820 4526 3825 ne
rect 4526 3820 4593 3825
tri 4526 3819 4527 3820 ne
rect 4278 3809 4287 3813
rect 4321 3809 4331 3813
rect 4330 3757 4331 3809
rect 4278 3745 4331 3757
rect 4330 3693 4331 3745
rect 4278 3687 4331 3693
rect 4527 3813 4593 3820
rect 4527 3779 4543 3813
rect 4577 3779 4593 3813
rect 4527 3741 4593 3779
rect 4527 3707 4543 3741
rect 4577 3707 4593 3741
tri 4197 3654 4227 3684 sw
rect 1187 3650 1730 3654
tri 1730 3650 1734 3654 nw
rect 1187 3648 1728 3650
tri 1728 3648 1730 3650 nw
rect 1187 3645 1725 3648
tri 1725 3645 1728 3648 nw
rect 1187 3642 1691 3645
rect 694 3614 928 3642
rect 641 3608 928 3614
rect 1004 3608 1006 3642
rect 1040 3608 1044 3642
rect 1118 3608 1135 3642
rect 1196 3608 1239 3642
rect 1273 3608 1316 3642
rect 1350 3608 1393 3642
rect 1427 3608 1470 3642
rect 1504 3608 1547 3642
rect 1581 3608 1624 3642
rect 1658 3611 1691 3642
tri 1691 3611 1725 3645 nw
rect 1658 3608 1688 3611
tri 1688 3608 1691 3611 nw
rect 641 3603 952 3608
rect 1004 3603 1044 3608
rect 1096 3603 1135 3608
rect 1187 3603 1682 3608
rect 641 3602 1682 3603
tri 1682 3602 1688 3608 nw
rect 2545 3601 2553 3653
rect 2605 3601 2618 3653
rect 2670 3601 2682 3653
rect 2734 3645 2746 3653
rect 2798 3645 2810 3653
rect 2862 3645 2874 3653
rect 2926 3645 2938 3653
rect 2743 3611 2746 3645
rect 2926 3611 2936 3645
rect 2734 3601 2746 3611
rect 2798 3601 2810 3611
rect 2862 3601 2874 3611
rect 2926 3601 2938 3611
rect 2990 3601 3002 3653
rect 3054 3601 3066 3653
rect 3118 3645 3130 3653
rect 3182 3645 3194 3653
rect 3246 3645 3258 3653
rect 3310 3645 3322 3653
rect 3120 3611 3130 3645
rect 3310 3611 3311 3645
rect 3118 3601 3130 3611
rect 3182 3601 3194 3611
rect 3246 3601 3258 3611
rect 3310 3601 3322 3611
rect 3374 3601 3386 3653
rect 3438 3601 3450 3653
rect 3502 3601 3514 3653
rect 3566 3645 3578 3653
rect 3630 3645 3642 3653
rect 3694 3645 3706 3653
rect 3758 3645 3770 3653
rect 3570 3611 3578 3645
rect 3758 3611 3761 3645
rect 3566 3601 3578 3611
rect 3630 3601 3642 3611
rect 3694 3601 3706 3611
rect 3758 3601 3770 3611
rect 3822 3601 3834 3653
rect 3886 3601 3898 3653
rect 3950 3601 3962 3653
rect 4014 3645 4032 3653
rect 4020 3611 4032 3645
rect 4014 3601 4032 3611
rect 4076 3648 4241 3654
rect 4076 3614 4088 3648
rect 4122 3614 4195 3648
rect 4229 3614 4241 3648
rect 4076 3608 4241 3614
rect 4320 3645 4338 3653
rect 4320 3611 4332 3645
rect 4320 3601 4338 3611
rect 4390 3601 4433 3653
rect 4485 3601 4491 3653
tri 587 3599 589 3601 sw
rect 587 3592 589 3599
tri 589 3592 596 3599 sw
rect 587 3582 596 3592
tri 596 3582 606 3592 sw
tri 4517 3582 4527 3592 se
rect 4527 3582 4593 3707
rect 4657 3809 4709 3815
rect 4657 3745 4709 3757
rect 4657 3682 4709 3693
rect 4790 3813 4842 3825
tri 5043 3820 5048 3825 ne
rect 5048 3820 5095 3825
tri 5048 3819 5049 3820 ne
rect 4790 3809 4799 3813
rect 4833 3809 4842 3813
rect 4790 3745 4842 3757
rect 5049 3813 5095 3820
rect 5049 3779 5055 3813
rect 5089 3779 5095 3813
rect 5049 3741 5095 3779
rect 5049 3707 5055 3741
rect 5089 3707 5095 3741
rect 5049 3695 5095 3707
rect 5302 3813 5354 3825
rect 5302 3809 5311 3813
rect 5345 3809 5354 3813
rect 5302 3745 5354 3757
rect 4790 3687 4842 3693
rect 5561 3813 5607 3910
rect 5902 3853 5908 3905
rect 5960 3853 5972 3905
rect 6024 3853 6631 3905
tri 6039 3841 6051 3853 ne
rect 6051 3841 6141 3853
tri 6141 3841 6153 3853 nw
tri 6551 3841 6563 3853 ne
rect 6563 3841 6631 3853
tri 6051 3838 6054 3841 ne
rect 6054 3838 6138 3841
tri 6138 3838 6141 3841 nw
tri 6563 3838 6566 3841 ne
rect 6566 3838 6631 3841
tri 6054 3825 6067 3838 ne
rect 6067 3825 6125 3838
tri 6125 3825 6138 3838 nw
tri 6566 3825 6579 3838 ne
rect 6579 3825 6631 3838
rect 5561 3779 5567 3813
rect 5601 3779 5607 3813
rect 5561 3741 5607 3779
rect 5561 3707 5567 3741
rect 5601 3707 5607 3741
rect 5561 3695 5607 3707
rect 5814 3813 5866 3825
tri 6067 3820 6072 3825 ne
rect 6072 3820 6120 3825
tri 6120 3820 6125 3825 nw
tri 6072 3819 6073 3820 ne
rect 5814 3809 5823 3813
rect 5857 3809 5866 3813
rect 5814 3745 5866 3757
rect 5302 3687 5354 3693
rect 6073 3813 6119 3820
tri 6119 3819 6120 3820 nw
rect 6073 3779 6079 3813
rect 6113 3779 6119 3813
rect 6073 3741 6119 3779
rect 6073 3707 6079 3741
rect 6113 3707 6119 3741
rect 6073 3695 6119 3707
rect 6326 3813 6378 3825
tri 6579 3820 6584 3825 ne
rect 6584 3820 6631 3825
tri 6584 3819 6585 3820 ne
rect 6326 3809 6335 3813
rect 6369 3809 6378 3813
rect 6326 3745 6378 3757
rect 5814 3687 5866 3693
rect 6585 3813 6631 3820
rect 6585 3779 6591 3813
rect 6625 3779 6631 3813
rect 6585 3741 6631 3779
rect 6585 3707 6591 3741
rect 6625 3707 6631 3741
rect 6585 3695 6631 3707
rect 6326 3687 6378 3693
tri 4709 3682 4711 3684 sw
tri 4629 3654 4657 3682 se
rect 4657 3654 4711 3682
tri 4711 3654 4739 3682 sw
rect 4629 3648 4788 3654
rect 6668 3653 6801 4198
rect 6980 4204 8059 4216
rect 6980 4198 7905 4204
tri 7905 4198 7911 4204 nw
tri 8004 4198 8010 4204 ne
rect 8010 4198 8059 4204
rect 6980 4189 7896 4198
tri 7896 4189 7905 4198 nw
tri 8010 4189 8019 4198 ne
rect 8019 4189 8059 4198
rect 6980 4177 7884 4189
tri 7884 4177 7896 4189 nw
tri 8019 4177 8031 4189 ne
rect 6980 4175 7881 4177
rect 6980 4170 7838 4175
rect 7872 4174 7881 4175
tri 7881 4174 7884 4177 nw
rect 7872 4172 7879 4174
tri 7879 4172 7881 4174 nw
rect 7872 4170 7878 4172
tri 7878 4171 7879 4172 nw
rect 6980 4118 7826 4170
rect 6980 4106 7878 4118
rect 6980 4054 7826 4106
rect 6980 4025 7878 4054
rect 6980 3991 7838 4025
rect 7872 3991 7878 4025
rect 6980 3950 7878 3991
rect 6980 3916 7838 3950
rect 7872 3916 7878 3950
rect 6980 3875 7878 3916
tri 6947 3841 6980 3874 se
rect 6980 3841 7838 3875
rect 7872 3841 7878 3875
tri 6944 3838 6947 3841 se
rect 6947 3838 7878 3841
tri 6931 3825 6944 3838 se
rect 6944 3825 7878 3838
rect 6841 3815 7878 3825
rect 6841 3763 6847 3815
rect 6899 3763 6954 3815
rect 7006 3763 7061 3815
rect 7113 3763 7168 3815
rect 7220 3763 7275 3815
rect 7327 3763 7382 3815
rect 7434 3813 7878 3815
rect 7434 3779 7703 3813
rect 7737 3800 7878 3813
rect 7737 3779 7838 3800
rect 7434 3766 7838 3779
rect 7872 3766 7878 3800
rect 7434 3763 7878 3766
rect 6841 3741 7878 3763
rect 6841 3687 6847 3741
rect 6881 3739 7703 3741
rect 6899 3687 6954 3739
rect 7006 3687 7061 3739
rect 7113 3687 7168 3739
rect 7220 3687 7275 3739
rect 7327 3687 7382 3739
rect 7434 3707 7703 3739
rect 7737 3725 7878 3741
rect 7737 3707 7838 3725
rect 7434 3691 7838 3707
rect 7872 3691 7878 3725
rect 7434 3687 7878 3691
tri 6940 3684 6943 3687 ne
rect 6943 3684 7878 3687
tri 6943 3654 6973 3684 ne
rect 6973 3654 7878 3684
rect 4629 3614 4641 3648
rect 4675 3614 4742 3648
rect 4776 3614 4788 3648
rect 4629 3608 4788 3614
rect 4832 3645 4850 3653
rect 4902 3645 4921 3653
rect 4973 3645 4992 3653
rect 5044 3645 5062 3653
rect 4832 3611 4844 3645
rect 4902 3611 4916 3645
rect 4973 3611 4988 3645
rect 5044 3611 5060 3645
rect 4832 3601 4850 3611
rect 4902 3601 4921 3611
rect 4973 3601 4992 3611
rect 5044 3601 5062 3611
rect 5114 3601 5132 3653
rect 5184 3601 5202 3653
rect 5254 3601 5272 3653
rect 5324 3601 5342 3653
rect 5394 3601 5412 3653
rect 5464 3601 5482 3653
rect 5534 3601 5552 3653
rect 5604 3601 5649 3653
rect 5701 3601 5715 3653
rect 5767 3601 5780 3653
rect 5832 3645 5845 3653
rect 5897 3645 5910 3653
rect 5962 3645 5975 3653
rect 6027 3645 6040 3653
rect 6092 3645 6105 3653
rect 5837 3611 5845 3645
rect 6092 3611 6099 3645
rect 5832 3601 5845 3611
rect 5897 3601 5910 3611
rect 5962 3601 5975 3611
rect 6027 3601 6040 3611
rect 6092 3601 6105 3611
rect 6157 3601 6170 3653
rect 6222 3601 6235 3653
rect 6287 3601 6293 3653
rect 6404 3601 6410 3653
rect 6462 3601 6523 3653
rect 6575 3601 6581 3653
rect 6668 3601 6674 3653
rect 6726 3601 6743 3653
rect 6795 3601 6801 3653
tri 6973 3650 6977 3654 ne
rect 6977 3650 7878 3654
tri 6977 3648 6979 3650 ne
rect 6979 3648 7838 3650
tri 6979 3647 6980 3648 ne
tri 4593 3582 4603 3592 sw
rect 587 3580 606 3582
tri 606 3580 608 3582 sw
tri 4515 3580 4517 3582 se
rect 4517 3580 4603 3582
tri 4603 3580 4605 3582 sw
rect 587 3575 608 3580
tri 608 3575 613 3580 sw
tri 4510 3575 4515 3580 se
rect 4515 3575 4605 3580
tri 4605 3575 4610 3580 sw
rect 587 3567 613 3575
tri 613 3567 621 3575 sw
tri 4502 3567 4510 3575 se
rect 4510 3567 4610 3575
tri 4610 3567 4618 3575 sw
rect 587 3565 4839 3567
rect 535 3553 4839 3565
rect 587 3521 4839 3553
rect 587 3509 601 3521
tri 601 3509 613 3521 nw
tri 3739 3509 3751 3521 ne
rect 3751 3509 3833 3521
tri 3833 3509 3845 3521 nw
tri 4251 3509 4263 3521 ne
rect 4263 3509 4345 3521
tri 4345 3509 4357 3521 nw
tri 4763 3509 4775 3521 ne
rect 4775 3509 4839 3521
rect 587 3506 598 3509
tri 598 3506 601 3509 nw
tri 3751 3506 3754 3509 ne
rect 3754 3506 3830 3509
tri 3830 3506 3833 3509 nw
tri 4263 3506 4266 3509 ne
rect 4266 3506 4342 3509
tri 4342 3506 4345 3509 nw
tri 4775 3506 4778 3509 ne
rect 4778 3506 4839 3509
rect 587 3501 592 3506
rect 535 3500 592 3501
tri 592 3500 598 3506 nw
tri 3754 3500 3760 3506 ne
rect 3760 3500 3824 3506
tri 3824 3500 3830 3506 nw
tri 4266 3500 4272 3506 ne
rect 4272 3500 4336 3506
tri 4336 3500 4342 3506 nw
tri 4778 3500 4784 3506 ne
rect 4784 3500 4839 3506
rect 535 3495 587 3500
tri 587 3495 592 3500 nw
tri 3760 3495 3765 3500 ne
rect 3765 3495 3815 3500
tri 3765 3491 3769 3495 ne
rect 946 3488 952 3489
rect 454 3432 507 3463
rect 506 3380 507 3432
rect 454 3350 507 3380
rect 454 3349 467 3350
rect 501 3349 507 3350
rect 506 3297 507 3349
rect 454 3276 507 3297
rect 454 3266 467 3276
rect 501 3266 507 3276
rect 506 3214 507 3266
rect 641 3482 952 3488
rect 1004 3482 1044 3489
rect 1096 3482 1135 3489
rect 1187 3488 1193 3489
rect 1187 3482 1670 3488
rect 641 3476 928 3482
rect 641 3442 660 3476
rect 694 3448 928 3476
rect 1004 3448 1006 3482
rect 1040 3448 1044 3482
rect 1118 3448 1135 3482
rect 1196 3448 1239 3482
rect 1273 3448 1316 3482
rect 1350 3448 1393 3482
rect 1427 3448 1470 3482
rect 1504 3448 1547 3482
rect 1581 3448 1624 3482
rect 1658 3448 1670 3482
rect 694 3442 952 3448
rect 641 3437 952 3442
rect 1004 3437 1044 3448
rect 1096 3437 1135 3448
rect 1187 3437 1670 3448
rect 641 3425 1670 3437
rect 1772 3433 1778 3485
rect 1830 3433 1844 3485
rect 1896 3433 1910 3485
rect 1962 3476 1976 3485
rect 2028 3476 2042 3485
rect 2094 3476 2108 3485
rect 2160 3476 2174 3485
rect 2226 3476 2240 3485
rect 2292 3476 2306 3485
rect 2358 3476 2372 3485
rect 1966 3442 1976 3476
rect 2039 3442 2042 3476
rect 2292 3442 2297 3476
rect 2358 3442 2370 3476
rect 1962 3433 1976 3442
rect 2028 3433 2042 3442
rect 2094 3433 2108 3442
rect 2160 3433 2174 3442
rect 2226 3433 2240 3442
rect 2292 3433 2306 3442
rect 2358 3433 2372 3442
rect 2424 3433 2437 3485
rect 2489 3433 2502 3485
rect 2554 3433 2567 3485
rect 2619 3476 2632 3485
rect 2684 3476 2697 3485
rect 2749 3476 2762 3485
rect 2814 3476 2827 3485
rect 2879 3476 2892 3485
rect 2944 3476 2957 3485
rect 2623 3442 2632 3476
rect 2696 3442 2697 3476
rect 2879 3442 2881 3476
rect 2944 3442 2954 3476
rect 2619 3433 2632 3442
rect 2684 3433 2697 3442
rect 2749 3433 2762 3442
rect 2814 3433 2827 3442
rect 2879 3433 2892 3442
rect 2944 3433 2957 3442
rect 3009 3433 3022 3485
rect 3074 3433 3087 3485
rect 3139 3433 3152 3485
rect 3204 3476 3217 3485
rect 3269 3476 3282 3485
rect 3334 3476 3347 3485
rect 3399 3476 3412 3485
rect 3464 3476 3477 3485
rect 3529 3476 3542 3485
rect 3207 3442 3217 3476
rect 3280 3442 3282 3476
rect 3464 3442 3465 3476
rect 3529 3442 3538 3476
rect 3204 3433 3217 3442
rect 3269 3433 3282 3442
rect 3334 3433 3347 3442
rect 3399 3433 3412 3442
rect 3464 3433 3477 3442
rect 3529 3433 3542 3442
rect 3594 3433 3607 3485
rect 3659 3433 3672 3485
rect 3724 3433 3730 3485
rect 641 3394 952 3425
rect 641 3360 660 3394
rect 694 3383 952 3394
rect 694 3360 871 3383
rect 641 3349 871 3360
rect 905 3373 952 3383
rect 1004 3373 1044 3425
rect 1096 3373 1135 3425
rect 1187 3403 1670 3425
rect 1187 3373 1581 3403
rect 905 3349 935 3373
tri 935 3349 959 3373 nw
tri 1230 3349 1254 3373 ne
rect 1254 3351 1581 3373
rect 1633 3351 1670 3403
rect 1974 3397 2026 3403
rect 1254 3349 1670 3351
rect 641 3311 912 3349
tri 912 3326 935 3349 nw
tri 1254 3340 1263 3349 ne
rect 1263 3327 1670 3349
rect 641 3277 660 3311
rect 694 3277 871 3311
rect 905 3277 912 3311
rect 641 3265 912 3277
rect 1263 3275 1581 3327
rect 1633 3275 1670 3327
rect 1263 3265 1670 3275
rect 1721 3383 1767 3395
rect 1721 3349 1727 3383
rect 1761 3349 1767 3383
rect 1721 3311 1767 3349
rect 1721 3277 1727 3311
rect 1761 3277 1767 3311
tri 1697 3241 1721 3265 se
rect 1721 3241 1767 3277
rect 2486 3397 2538 3403
rect 1974 3333 2026 3345
rect 1974 3277 1983 3281
rect 2017 3277 2026 3281
rect 1974 3265 2026 3277
rect 2233 3383 2279 3395
rect 2233 3349 2239 3383
rect 2273 3349 2279 3383
rect 2233 3311 2279 3349
rect 2233 3277 2239 3311
rect 2273 3277 2279 3311
tri 1767 3241 1791 3265 sw
tri 2209 3241 2233 3265 se
rect 2233 3241 2279 3277
rect 2998 3397 3050 3403
rect 2486 3333 2538 3345
rect 2486 3277 2495 3281
rect 2529 3277 2538 3281
rect 2486 3265 2538 3277
rect 2745 3383 2791 3395
rect 2745 3349 2751 3383
rect 2785 3349 2791 3383
rect 2745 3311 2791 3349
rect 2745 3277 2751 3311
rect 2785 3277 2791 3311
tri 2279 3241 2303 3265 sw
tri 2721 3241 2745 3265 se
rect 2745 3241 2791 3277
rect 3510 3397 3562 3403
rect 2998 3333 3050 3345
rect 2998 3277 3007 3281
rect 3041 3277 3050 3281
rect 2998 3265 3050 3277
rect 3257 3383 3303 3395
rect 3257 3349 3263 3383
rect 3297 3349 3303 3383
rect 3257 3311 3303 3349
rect 3257 3277 3263 3311
rect 3297 3277 3303 3311
tri 2791 3241 2815 3265 sw
tri 3233 3241 3257 3265 se
rect 3257 3241 3303 3277
rect 3510 3333 3562 3345
rect 3510 3277 3519 3281
rect 3553 3277 3562 3281
rect 3510 3265 3562 3277
rect 3769 3383 3815 3495
tri 3815 3491 3824 3500 nw
tri 4272 3491 4281 3500 ne
rect 3849 3433 3855 3485
rect 3907 3433 3922 3485
rect 3974 3476 3989 3485
rect 4041 3476 4056 3485
rect 4108 3476 4123 3485
rect 3980 3442 3989 3476
rect 4108 3442 4116 3476
rect 3974 3433 3989 3442
rect 4041 3433 4056 3442
rect 4108 3433 4123 3442
rect 4175 3433 4189 3485
rect 4241 3433 4247 3485
rect 3769 3349 3775 3383
rect 3809 3349 3815 3383
rect 3769 3311 3815 3349
rect 3769 3277 3775 3311
rect 3809 3277 3815 3311
rect 3769 3265 3815 3277
rect 4022 3397 4074 3403
rect 4022 3333 4074 3345
rect 4022 3277 4031 3281
rect 4065 3277 4074 3281
rect 4022 3265 4074 3277
rect 4281 3383 4327 3500
tri 4327 3491 4336 3500 nw
tri 4784 3491 4793 3500 ne
rect 4361 3433 4367 3485
rect 4419 3433 4434 3485
rect 4486 3476 4501 3485
rect 4553 3476 4568 3485
rect 4620 3476 4635 3485
rect 4492 3442 4501 3476
rect 4620 3442 4628 3476
rect 4486 3433 4501 3442
rect 4553 3433 4568 3442
rect 4620 3433 4635 3442
rect 4687 3433 4701 3485
rect 4753 3433 4759 3485
rect 4281 3349 4287 3383
rect 4321 3349 4327 3383
rect 4281 3311 4327 3349
rect 4281 3277 4287 3311
rect 4321 3277 4327 3311
rect 4281 3265 4327 3277
rect 4534 3397 4586 3403
rect 4534 3333 4586 3345
rect 4534 3277 4543 3281
rect 4577 3277 4586 3281
rect 4534 3265 4586 3277
rect 4793 3383 4839 3500
rect 6668 3485 6801 3601
rect 6980 3642 7838 3648
rect 6980 3608 6992 3642
rect 7026 3608 7064 3642
rect 7098 3608 7136 3642
rect 7170 3608 7208 3642
rect 7242 3608 7280 3642
rect 7314 3608 7353 3642
rect 7387 3608 7426 3642
rect 7460 3608 7499 3642
rect 7533 3616 7838 3642
rect 7872 3616 7878 3650
rect 7533 3608 7878 3616
rect 6980 3575 7878 3608
rect 6980 3541 7838 3575
rect 7872 3541 7878 3575
rect 6980 3500 7878 3541
rect 4873 3433 4879 3485
rect 4931 3433 4986 3485
rect 5038 3433 5044 3485
rect 5100 3476 5556 3482
rect 5100 3442 5112 3476
rect 5146 3442 5192 3476
rect 5226 3442 5272 3476
rect 5306 3442 5352 3476
rect 5386 3442 5431 3476
rect 5465 3442 5510 3476
rect 5544 3442 5556 3476
rect 5100 3436 5556 3442
tri 5097 3433 5100 3436 se
rect 5100 3433 5178 3436
tri 5096 3432 5097 3433 se
rect 5097 3432 5178 3433
tri 5178 3432 5182 3436 nw
tri 5275 3432 5279 3436 ne
rect 5279 3432 5376 3436
tri 5376 3432 5380 3436 nw
tri 5474 3432 5478 3436 ne
rect 5478 3433 5556 3436
tri 5556 3433 5559 3436 sw
rect 5612 3433 5618 3485
rect 5670 3433 5684 3485
rect 5736 3433 5750 3485
rect 5802 3476 5816 3485
rect 5868 3476 5882 3485
rect 5934 3476 5948 3485
rect 6000 3476 6014 3485
rect 5810 3442 5816 3476
rect 6000 3442 6004 3476
rect 5802 3433 5816 3442
rect 5868 3433 5882 3442
rect 5934 3433 5948 3442
rect 6000 3433 6014 3442
rect 6066 3433 6079 3485
rect 6131 3433 6144 3485
rect 6196 3433 6209 3485
rect 6261 3476 6274 3485
rect 6326 3476 6339 3485
rect 6391 3476 6404 3485
rect 6456 3476 6469 3485
rect 6266 3442 6274 3476
rect 6456 3442 6459 3476
rect 6261 3433 6274 3442
rect 6326 3433 6339 3442
rect 6391 3433 6404 3442
rect 6456 3433 6469 3442
rect 6521 3433 6534 3485
rect 6586 3433 6592 3485
rect 6668 3433 6674 3485
rect 6726 3433 6743 3485
rect 6795 3433 6801 3485
tri 6974 3482 6980 3488 se
rect 6980 3482 7838 3500
tri 6940 3448 6974 3482 se
rect 6974 3448 6992 3482
rect 7026 3448 7064 3482
rect 7098 3448 7136 3482
rect 7170 3448 7208 3482
rect 7242 3448 7280 3482
rect 7314 3448 7353 3482
rect 7387 3448 7426 3482
rect 7460 3448 7499 3482
rect 7533 3466 7838 3482
rect 7872 3466 7878 3500
rect 7533 3448 7878 3466
tri 6934 3442 6940 3448 se
rect 6940 3442 7878 3448
tri 6925 3433 6934 3442 se
rect 6934 3433 7878 3442
rect 5478 3432 5559 3433
tri 5559 3432 5560 3433 sw
tri 6924 3432 6925 3433 se
rect 6925 3432 7878 3433
tri 5089 3425 5096 3432 se
rect 5096 3425 5171 3432
tri 5171 3425 5178 3432 nw
tri 5279 3425 5286 3432 ne
rect 5286 3425 5369 3432
tri 5369 3425 5376 3432 nw
tri 5478 3425 5485 3432 ne
rect 5485 3425 5560 3432
tri 5560 3425 5567 3432 sw
tri 6917 3425 6924 3432 se
rect 6924 3425 7878 3432
tri 5067 3403 5089 3425 se
rect 5089 3403 5149 3425
tri 5149 3403 5171 3425 nw
tri 5286 3409 5302 3425 ne
rect 4793 3349 4799 3383
rect 4833 3349 4839 3383
rect 4793 3311 4839 3349
rect 4793 3277 4799 3311
rect 4833 3277 4839 3311
rect 4793 3265 4839 3277
rect 5046 3397 5137 3403
rect 5098 3391 5137 3397
tri 5137 3391 5149 3403 nw
rect 5302 3397 5354 3425
tri 5354 3410 5369 3425 nw
tri 5485 3410 5500 3425 ne
rect 5500 3410 5567 3425
tri 5500 3403 5507 3410 ne
rect 5507 3403 5567 3410
tri 5567 3403 5589 3425 sw
tri 6895 3403 6917 3425 se
rect 6917 3403 7838 3425
rect 5098 3383 5129 3391
tri 5129 3383 5137 3391 nw
tri 5507 3391 5519 3403 ne
rect 5519 3397 5610 3403
rect 5519 3391 5558 3397
tri 5519 3383 5527 3391 ne
rect 5527 3383 5558 3391
rect 6070 3397 6122 3403
tri 5098 3352 5129 3383 nw
rect 5046 3333 5098 3345
rect 5046 3277 5055 3281
rect 5089 3277 5098 3281
rect 5046 3265 5098 3277
tri 5527 3352 5558 3383 ne
rect 5302 3333 5354 3345
rect 5302 3277 5311 3281
rect 5345 3277 5354 3281
rect 5302 3275 5354 3277
rect 5558 3333 5610 3345
rect 5558 3277 5567 3281
rect 5601 3277 5610 3281
rect 5305 3265 5351 3275
rect 5558 3265 5610 3277
rect 5817 3383 5863 3395
rect 5817 3349 5823 3383
rect 5857 3349 5863 3383
rect 5817 3311 5863 3349
rect 5817 3277 5823 3311
rect 5857 3277 5863 3311
tri 3303 3241 3327 3265 sw
tri 5793 3241 5817 3265 se
rect 5817 3241 5863 3277
rect 6582 3397 6634 3403
rect 6070 3333 6122 3345
rect 6070 3277 6079 3281
rect 6113 3277 6122 3281
rect 6070 3265 6122 3277
rect 6329 3383 6375 3395
rect 6329 3349 6335 3383
rect 6369 3349 6375 3383
rect 6329 3311 6375 3349
rect 6329 3277 6335 3311
rect 6369 3277 6375 3311
tri 5863 3241 5887 3265 sw
tri 6305 3241 6329 3265 se
rect 6329 3241 6375 3277
tri 6887 3395 6895 3403 se
rect 6895 3395 6986 3403
rect 6582 3333 6634 3345
rect 6841 3383 6986 3395
rect 6841 3349 6847 3383
rect 6881 3351 6986 3383
rect 7038 3351 7085 3403
rect 7137 3351 7184 3403
rect 7236 3351 7283 3403
rect 7335 3351 7382 3403
rect 7434 3383 7712 3403
rect 7434 3351 7703 3383
rect 7764 3351 7820 3403
rect 7872 3351 7878 3425
rect 6881 3349 7703 3351
rect 7737 3350 7878 3351
rect 7737 3349 7838 3350
rect 6841 3327 7838 3349
rect 6841 3311 6986 3327
rect 6582 3277 6591 3281
rect 6625 3277 6634 3281
tri 6836 3277 6841 3282 se
rect 6841 3277 6847 3311
rect 6881 3277 6986 3311
rect 6582 3265 6634 3277
tri 6834 3275 6836 3277 se
rect 6836 3275 6986 3277
rect 7038 3275 7085 3327
rect 7137 3275 7184 3327
rect 7236 3275 7283 3327
rect 7335 3275 7382 3327
rect 7434 3311 7712 3327
rect 7434 3277 7703 3311
rect 7434 3275 7712 3277
rect 7764 3275 7820 3327
tri 6824 3265 6834 3275 se
rect 6834 3265 7838 3275
tri 6375 3241 6399 3265 sw
tri 6800 3241 6824 3265 se
rect 6824 3241 7838 3265
rect 7872 3241 7878 3350
tri 1691 3235 1697 3241 se
rect 1697 3235 1791 3241
tri 1791 3235 1797 3241 sw
tri 2203 3235 2209 3241 se
rect 2209 3235 2303 3241
tri 2303 3235 2309 3241 sw
tri 2715 3235 2721 3241 se
rect 2721 3235 2815 3241
tri 2815 3235 2821 3241 sw
tri 3227 3235 3233 3241 se
rect 3233 3235 3327 3241
tri 3327 3235 3333 3241 sw
tri 5787 3235 5793 3241 se
rect 5793 3235 5887 3241
tri 5887 3235 5893 3241 sw
tri 6299 3235 6305 3241 se
rect 6305 3235 6399 3241
tri 6399 3235 6405 3241 sw
tri 6794 3235 6800 3241 se
rect 6800 3235 7878 3241
rect 454 3202 507 3214
rect 454 3183 467 3202
rect 501 3183 507 3202
rect 506 3166 507 3183
rect 781 3229 3333 3235
rect 833 3203 3333 3229
tri 3562 3220 3577 3235 se
rect 3577 3220 5863 3235
tri 3556 3214 3562 3220 se
rect 3562 3214 5863 3220
tri 3555 3213 3556 3214 se
rect 3556 3213 5863 3214
rect 6283 3213 6289 3235
tri 3552 3210 3555 3213 se
rect 3555 3210 6289 3213
tri 3545 3203 3552 3210 se
rect 3552 3203 6289 3210
rect 833 3200 864 3203
tri 864 3200 867 3203 nw
tri 3542 3200 3545 3203 se
rect 3545 3200 3603 3203
tri 3603 3200 3606 3203 nw
tri 5797 3200 5800 3203 ne
rect 5800 3200 5880 3203
tri 5880 3200 5883 3203 nw
tri 6263 3200 6266 3203 ne
rect 6266 3200 6289 3203
rect 833 3183 847 3200
tri 847 3183 864 3200 nw
tri 3525 3183 3542 3200 se
rect 3542 3183 3586 3200
tri 3586 3183 3603 3200 nw
tri 5800 3183 5817 3200 ne
rect 5817 3183 5863 3200
tri 5863 3183 5880 3200 nw
tri 6266 3183 6283 3200 ne
rect 6283 3183 6289 3200
rect 6341 3183 6353 3235
rect 6405 3183 6411 3235
tri 6779 3220 6794 3235 se
rect 6794 3220 7878 3235
tri 6773 3214 6779 3220 se
rect 6779 3214 7878 3220
tri 6769 3210 6773 3214 se
rect 6773 3210 7878 3214
tri 6759 3200 6769 3210 se
rect 6769 3200 7878 3210
tri 6742 3183 6759 3200 se
rect 6759 3183 7838 3200
rect 833 3177 839 3183
rect 781 3175 839 3177
tri 839 3175 847 3183 nw
tri 3517 3175 3525 3183 se
rect 3525 3175 3578 3183
tri 3578 3175 3586 3183 nw
tri 6734 3175 6742 3183 se
rect 6742 3175 7838 3183
tri 507 3166 509 3168 sw
rect 506 3163 509 3166
tri 509 3163 512 3166 sw
rect 781 3165 833 3175
tri 833 3169 839 3175 nw
tri 880 3169 886 3175 se
rect 886 3169 3569 3175
tri 877 3166 880 3169 se
rect 880 3166 3569 3169
tri 3569 3166 3578 3175 nw
tri 6725 3166 6734 3175 se
rect 6734 3166 7838 3175
rect 7872 3166 7878 3200
rect 506 3159 512 3163
tri 512 3159 516 3163 sw
rect 506 3136 516 3159
tri 516 3136 539 3159 sw
rect 506 3134 539 3136
tri 539 3134 541 3136 sw
rect 506 3131 543 3134
rect 454 3128 543 3131
rect 454 3100 482 3128
rect 516 3094 543 3128
tri 874 3163 877 3166 se
rect 877 3163 3566 3166
tri 3566 3163 3569 3166 nw
tri 6722 3163 6725 3166 se
rect 6725 3163 7878 3166
tri 870 3159 874 3163 se
rect 874 3159 3562 3163
tri 3562 3159 3566 3163 nw
tri 6718 3159 6722 3163 se
rect 6722 3159 7878 3163
rect 781 3107 833 3113
tri 863 3152 870 3159 se
rect 870 3152 3555 3159
tri 3555 3152 3562 3159 nw
tri 6711 3152 6718 3159 se
rect 6718 3152 7878 3159
rect 863 3149 3552 3152
tri 3552 3149 3555 3152 nw
tri 6708 3149 6711 3152 se
rect 6711 3149 7878 3152
rect 863 3145 3548 3149
tri 3548 3145 3552 3149 nw
tri 6704 3145 6708 3149 se
rect 6708 3145 7878 3149
rect 863 3143 940 3145
rect 506 3088 543 3094
rect 915 3136 940 3143
tri 940 3136 949 3145 nw
tri 6695 3136 6704 3145 se
rect 6704 3136 7878 3145
rect 915 3134 938 3136
tri 938 3134 940 3136 nw
tri 6693 3134 6695 3136 se
rect 6695 3134 7878 3136
rect 915 3128 932 3134
tri 932 3128 938 3134 nw
tri 3804 3128 3810 3134 se
rect 3810 3128 5035 3134
rect 5087 3128 5102 3134
rect 5154 3128 5169 3134
rect 5221 3128 5236 3134
rect 5288 3128 5303 3134
rect 5355 3128 5371 3134
rect 5423 3128 7878 3134
rect 915 3117 921 3128
tri 921 3117 932 3128 nw
tri 3793 3117 3804 3128 se
rect 3804 3117 3888 3128
tri 915 3111 921 3117 nw
tri 1059 3111 1065 3117 se
rect 1065 3111 1582 3117
tri 1055 3107 1059 3111 se
rect 1059 3107 1077 3111
rect 506 3077 529 3088
tri 529 3077 540 3088 nw
rect 863 3079 915 3091
rect 506 3062 514 3077
tri 514 3062 529 3077 nw
tri 506 3054 514 3062 nw
rect 454 3002 506 3048
rect 863 3021 915 3027
tri 1039 3091 1055 3107 se
rect 1055 3091 1077 3107
rect 1039 3077 1077 3091
rect 1111 3077 1150 3111
rect 1184 3077 1223 3111
rect 1257 3077 1296 3111
rect 1330 3077 1368 3111
rect 1402 3077 1440 3111
rect 1474 3077 1512 3111
rect 1546 3077 1582 3111
rect 1039 3071 1582 3077
rect 1039 3065 1096 3071
tri 1096 3065 1102 3071 nw
tri 1570 3065 1576 3071 ne
rect 1576 3065 1582 3071
rect 1634 3065 1646 3117
rect 1698 3111 1964 3117
rect 2016 3111 2028 3117
rect 2080 3111 3888 3117
rect 1698 3077 1728 3111
rect 1762 3077 1800 3111
rect 1834 3077 1872 3111
rect 1906 3077 1944 3111
rect 2080 3077 2088 3111
rect 2122 3077 2160 3111
rect 2194 3077 2232 3111
rect 2266 3077 2304 3111
rect 2338 3077 2376 3111
rect 2410 3077 2448 3111
rect 2482 3077 2520 3111
rect 2554 3077 2592 3111
rect 2626 3077 2664 3111
rect 2698 3077 2736 3111
rect 2770 3077 2808 3111
rect 2842 3077 2880 3111
rect 2914 3077 2952 3111
rect 2986 3077 3024 3111
rect 3058 3077 3096 3111
rect 3130 3077 3168 3111
rect 3202 3077 3240 3111
rect 3274 3077 3312 3111
rect 3346 3077 3384 3111
rect 3418 3077 3456 3111
rect 3490 3077 3528 3111
rect 3562 3077 3600 3111
rect 3634 3077 3672 3111
rect 3706 3077 3744 3111
rect 3778 3094 3888 3111
rect 3922 3094 3962 3128
rect 3996 3094 4036 3128
rect 4070 3094 4110 3128
rect 4144 3094 4184 3128
rect 4218 3094 4258 3128
rect 4292 3094 4332 3128
rect 4366 3094 4406 3128
rect 4440 3094 4480 3128
rect 4514 3094 4553 3128
rect 4587 3094 4626 3128
rect 4660 3094 4699 3128
rect 4733 3094 4772 3128
rect 4806 3094 4845 3128
rect 4879 3094 4918 3128
rect 4952 3094 4991 3128
rect 5025 3094 5035 3128
rect 5098 3094 5102 3128
rect 5355 3094 5356 3128
rect 5423 3094 5429 3128
rect 5463 3094 5502 3128
rect 5536 3094 5575 3128
rect 5609 3094 5648 3128
rect 5682 3094 5721 3128
rect 5755 3094 5794 3128
rect 5828 3094 5867 3128
rect 5901 3094 5940 3128
rect 5974 3094 6013 3128
rect 6047 3094 6086 3128
rect 6120 3094 6159 3128
rect 6193 3094 6232 3128
rect 6266 3094 6305 3128
rect 6339 3094 6378 3128
rect 6412 3094 6451 3128
rect 6485 3094 6524 3128
rect 6558 3094 6597 3128
rect 6631 3094 6670 3128
rect 6704 3094 6743 3128
rect 6777 3094 6816 3128
rect 6850 3094 6889 3128
rect 6923 3094 6962 3128
rect 6996 3094 7035 3128
rect 7069 3094 7108 3128
rect 7142 3094 7181 3128
rect 7215 3094 7254 3128
rect 7288 3094 7327 3128
rect 7361 3094 7400 3128
rect 7434 3094 7473 3128
rect 7507 3094 7546 3128
rect 7580 3094 7619 3128
rect 7653 3094 7692 3128
rect 7726 3094 7765 3128
rect 7799 3094 7878 3128
rect 3778 3088 5035 3094
rect 3778 3087 3872 3088
tri 3872 3087 3873 3088 nw
tri 5023 3087 5024 3088 ne
rect 5024 3087 5035 3088
rect 3778 3077 3856 3087
rect 1698 3071 1964 3077
rect 1698 3065 1704 3071
tri 1704 3065 1710 3071 nw
tri 1953 3066 1958 3071 ne
rect 1958 3065 1964 3071
rect 2016 3065 2028 3077
rect 2080 3071 3856 3077
tri 3856 3071 3872 3087 nw
tri 5024 3082 5029 3087 ne
rect 5029 3082 5035 3087
rect 5087 3082 5102 3094
rect 5154 3082 5169 3094
rect 5221 3082 5236 3094
rect 5288 3082 5303 3094
rect 5355 3082 5371 3094
rect 5423 3088 7878 3094
rect 7936 4144 7988 4150
rect 7936 4080 7988 4092
rect 5423 3087 5436 3088
tri 5436 3087 5437 3088 nw
rect 5423 3082 5431 3087
tri 5431 3082 5436 3087 nw
rect 2080 3065 2086 3071
tri 2086 3065 2092 3071 nw
rect 1039 3062 1093 3065
tri 1093 3062 1096 3065 nw
tri 1591 3062 1594 3065 ne
rect 1594 3062 1676 3065
tri 1676 3062 1679 3065 nw
tri 7934 3062 7936 3064 se
rect 7936 3062 7988 4028
tri 8020 4078 8031 4089 se
rect 8031 4078 8059 4189
tri 8059 4078 8072 4091 sw
rect 8020 4072 8072 4078
rect 8020 4008 8072 4020
rect 8020 3950 8072 3956
tri 8020 3939 8031 3950 ne
tri 1038 3013 1039 3014 se
rect 1039 3013 1077 3062
tri 1077 3046 1093 3062 nw
tri 1594 3046 1610 3062 ne
rect 1610 3046 1651 3062
tri 1610 3037 1619 3046 ne
rect 1619 3037 1651 3046
tri 1651 3037 1676 3062 nw
tri 7913 3041 7934 3062 se
rect 7934 3041 7988 3062
tri 506 3002 517 3013 sw
tri 1027 3002 1038 3013 se
rect 1038 3002 1077 3013
rect 454 2993 517 3002
tri 517 2993 526 3002 sw
tri 1018 2993 1027 3002 se
rect 1027 2993 1077 3002
rect 454 2947 1077 2993
rect 1619 2986 1647 3037
tri 1647 3033 1651 3037 nw
rect 1745 2989 1751 3041
rect 1803 2989 1815 3041
rect 1867 3035 1913 3041
tri 1913 3035 1919 3041 sw
tri 2122 3035 2128 3041 se
rect 2128 3035 5166 3041
rect 1867 2989 5166 3035
rect 5218 2989 5230 3041
rect 5282 3030 6520 3041
tri 6520 3030 6531 3041 sw
tri 7902 3030 7913 3041 se
rect 7913 3030 7988 3041
rect 5282 3015 7988 3030
rect 5282 3013 7986 3015
tri 7986 3013 7988 3015 nw
rect 5282 3002 7975 3013
tri 7975 3002 7986 3013 nw
rect 5282 2989 7962 3002
tri 7962 2989 7975 3002 nw
tri 1647 2986 1649 2988 sw
rect 1619 2985 1649 2986
tri 1649 2985 1650 2986 sw
tri 8030 2985 8031 2986 se
rect 8031 2985 8059 3950
tri 8059 3937 8072 3950 nw
rect 1116 2975 1232 2981
rect 1017 2895 1069 2901
tri 1232 2954 1244 2966 sw
rect 1619 2961 1650 2985
tri 1650 2961 1674 2985 sw
tri 8006 2961 8030 2985 se
rect 8030 2966 8059 2985
rect 8030 2961 8054 2966
tri 8054 2961 8059 2966 nw
rect 1619 2954 8047 2961
tri 8047 2954 8054 2961 nw
rect 1232 2942 1244 2954
tri 1244 2942 1256 2954 sw
rect 1619 2942 8035 2954
tri 8035 2942 8047 2954 nw
rect 1232 2933 1256 2942
tri 1256 2933 1265 2942 sw
rect 1619 2933 8026 2942
tri 8026 2933 8035 2942 nw
tri 8097 2933 8103 2939 se
rect 8103 2933 8155 4498
rect 1232 2926 1265 2933
tri 1265 2926 1272 2933 sw
tri 8090 2926 8097 2933 se
rect 8097 2926 8155 2933
rect 1232 2914 1272 2926
tri 1272 2914 1284 2926 sw
tri 8078 2914 8090 2926 se
rect 8090 2914 8155 2926
rect 1232 2905 1284 2914
tri 1284 2905 1293 2914 sw
tri 8069 2905 8078 2914 se
rect 8078 2905 8155 2914
rect 1232 2886 8155 2905
rect 1232 2880 8149 2886
tri 8149 2880 8155 2886 nw
tri 8183 4599 8195 4611 se
rect 8195 4599 8215 4611
rect 8183 4573 8215 4599
rect 8267 4573 8279 4625
rect 8331 4573 8337 4625
rect 8476 4616 8522 4656
rect 8476 4582 8482 4616
rect 8516 4582 8522 4616
rect 8183 4558 8254 4573
tri 8254 4558 8269 4573 nw
rect 8183 4544 8240 4558
tri 8240 4544 8254 4558 nw
rect 8183 4542 8238 4544
tri 8238 4542 8240 4544 nw
rect 8476 4542 8522 4582
rect 1232 2859 8128 2880
tri 8128 2859 8149 2880 nw
tri 1069 2856 1072 2859 sw
rect 1116 2856 8125 2859
tri 8125 2856 8128 2859 nw
tri 8180 2856 8183 2859 se
rect 8183 2856 8235 4542
tri 8235 4539 8238 4542 nw
rect 8476 4508 8482 4542
rect 8516 4508 8522 4542
rect 8476 4468 8522 4508
rect 1069 2853 1072 2856
tri 1072 2853 1075 2856 sw
rect 1116 2853 8122 2856
tri 8122 2853 8125 2856 nw
tri 8177 2853 8180 2856 se
rect 8180 2853 8235 2856
rect 1069 2843 1075 2853
rect 1017 2840 1075 2843
tri 1075 2840 1088 2853 sw
tri 8164 2840 8177 2853 se
rect 8177 2840 8235 2853
rect 1017 2831 1088 2840
rect 1069 2825 1088 2831
tri 1088 2825 1103 2840 sw
tri 8149 2825 8164 2840 se
rect 8164 2825 8235 2840
rect 1069 2805 8235 2825
rect 1069 2782 8212 2805
tri 8212 2782 8235 2805 nw
rect 8263 4412 8269 4464
rect 8321 4412 8333 4464
rect 8385 4412 8391 4464
rect 8476 4434 8482 4468
rect 8516 4434 8522 4468
rect 8263 4411 8348 4412
tri 8348 4411 8349 4412 nw
rect 8263 4396 8333 4411
tri 8333 4396 8348 4411 nw
rect 8263 4394 8331 4396
tri 8331 4394 8333 4396 nw
rect 8476 4394 8522 4434
rect 1069 2779 8209 2782
tri 8209 2779 8212 2782 nw
rect 1017 2778 8208 2779
tri 8208 2778 8209 2779 nw
tri 8262 2778 8263 2779 se
rect 8263 2778 8315 4394
tri 8315 4378 8331 4394 nw
rect 8476 4360 8482 4394
rect 8516 4360 8522 4394
rect 8476 4320 8522 4360
rect 8476 4286 8482 4320
rect 8516 4286 8522 4320
rect 8476 4246 8522 4286
rect 8476 4212 8482 4246
rect 8516 4212 8522 4246
rect 8476 4172 8522 4212
rect 8476 4138 8482 4172
rect 8516 4138 8522 4172
rect 8476 4098 8522 4138
rect 8476 4064 8482 4098
rect 8516 4064 8522 4098
rect 8476 4024 8522 4064
rect 1017 2776 8206 2778
tri 8206 2776 8208 2778 nw
tri 8260 2776 8262 2778 se
rect 8262 2776 8315 2778
rect 1017 2773 8203 2776
tri 8203 2773 8206 2776 nw
tri 8257 2773 8260 2776 se
rect 8260 2773 8315 2776
tri 8250 2766 8257 2773 se
rect 8257 2766 8315 2773
tri 8229 2745 8250 2766 se
rect 8250 2745 8315 2766
rect 863 2739 8315 2745
rect 915 2736 8315 2739
rect 915 2732 8311 2736
tri 8311 2732 8315 2736 nw
rect 8348 4001 8400 4007
rect 8348 3937 8400 3949
rect 915 2727 8306 2732
tri 8306 2727 8311 2732 nw
rect 8348 2729 8400 3885
rect 8476 3990 8482 4024
rect 8516 3990 8522 4024
rect 8476 3950 8522 3990
rect 8708 4630 8714 4664
rect 8748 4630 8754 4664
tri 8862 4662 8864 4664 ne
rect 8708 4592 8754 4630
rect 8708 4558 8714 4592
rect 8748 4558 8754 4592
rect 8708 4520 8754 4558
rect 8708 4486 8714 4520
rect 8748 4486 8754 4520
rect 8708 4448 8754 4486
rect 8708 4414 8714 4448
rect 8748 4414 8754 4448
rect 8708 4376 8754 4414
rect 8708 4342 8714 4376
rect 8748 4342 8754 4376
rect 8708 4304 8754 4342
rect 8708 4270 8714 4304
rect 8748 4270 8754 4304
rect 8708 4232 8754 4270
rect 8708 4198 8714 4232
rect 8748 4198 8754 4232
rect 8708 4160 8754 4198
rect 8708 4126 8714 4160
rect 8748 4126 8754 4160
rect 8708 4088 8754 4126
rect 8708 4054 8714 4088
rect 8748 4054 8754 4088
rect 8708 4016 8754 4054
rect 8708 3982 8714 4016
rect 8748 3982 8754 4016
tri 8697 3961 8708 3972 se
rect 8708 3961 8754 3982
rect 8864 4630 8870 4664
rect 8904 4630 8910 4664
tri 8910 4662 8912 4664 nw
rect 8864 4592 8910 4630
rect 8864 4558 8870 4592
rect 8904 4558 8910 4592
rect 8864 4520 8910 4558
rect 8864 4486 8870 4520
rect 8904 4486 8910 4520
rect 8864 4448 8910 4486
rect 8864 4414 8870 4448
rect 8904 4414 8910 4448
rect 8864 4376 8910 4414
rect 8864 4342 8870 4376
rect 8904 4342 8910 4376
rect 8864 4304 8910 4342
rect 8864 4270 8870 4304
rect 8904 4270 8910 4304
rect 8864 4232 8910 4270
rect 8864 4198 8870 4232
rect 8904 4198 8910 4232
rect 8864 4160 8910 4198
rect 8864 4126 8870 4160
rect 8904 4126 8910 4160
rect 8864 4088 8910 4126
rect 8864 4054 8870 4088
rect 8904 4054 8910 4088
rect 8864 4016 8910 4054
rect 8864 3982 8870 4016
rect 8904 3982 8910 4016
tri 8688 3952 8697 3961 se
rect 8697 3952 8754 3961
tri 8754 3952 8763 3961 sw
rect 8476 3916 8482 3950
rect 8516 3916 8522 3950
tri 8680 3944 8688 3952 se
rect 8688 3947 8763 3952
tri 8763 3947 8768 3952 sw
rect 8688 3944 8768 3947
tri 8768 3944 8771 3947 sw
rect 8864 3944 8910 3982
rect 9020 4630 9026 4664
rect 9060 4630 9066 4664
rect 9020 4592 9066 4630
rect 9020 4558 9026 4592
rect 9060 4558 9066 4592
rect 9020 4520 9066 4558
rect 9020 4486 9026 4520
rect 9060 4486 9066 4520
rect 9020 4448 9066 4486
rect 9020 4414 9026 4448
rect 9060 4414 9066 4448
rect 9020 4376 9066 4414
rect 9020 4342 9026 4376
rect 9060 4342 9066 4376
rect 9020 4304 9066 4342
rect 9020 4270 9026 4304
rect 9060 4270 9066 4304
rect 9020 4232 9066 4270
rect 9020 4198 9026 4232
rect 9060 4198 9066 4232
rect 9020 4160 9066 4198
rect 9020 4126 9026 4160
rect 9060 4126 9066 4160
rect 9020 4088 9066 4126
rect 9020 4054 9026 4088
rect 9060 4054 9066 4088
rect 9020 4016 9066 4054
rect 9020 3982 9026 4016
rect 9060 3982 9066 4016
tri 9000 3952 9020 3972 se
rect 9020 3952 9066 3982
rect 9176 4808 9222 4820
rect 9176 4774 9182 4808
rect 9216 4774 9222 4808
rect 9176 4736 9222 4774
rect 9176 4702 9182 4736
rect 9216 4702 9222 4736
rect 9176 4664 9222 4702
rect 9176 4630 9182 4664
rect 9216 4630 9222 4664
rect 9176 4592 9222 4630
rect 9176 4558 9182 4592
rect 9216 4558 9222 4592
rect 9176 4520 9222 4558
rect 9176 4486 9182 4520
rect 9216 4486 9222 4520
rect 9176 4448 9222 4486
rect 9176 4414 9182 4448
rect 9216 4414 9222 4448
rect 9176 4376 9222 4414
rect 9176 4342 9182 4376
rect 9216 4342 9222 4376
rect 9176 4304 9222 4342
rect 9176 4270 9182 4304
rect 9216 4270 9222 4304
rect 9176 4232 9222 4270
rect 9176 4198 9182 4232
rect 9216 4198 9222 4232
rect 9176 4160 9222 4198
rect 9176 4126 9182 4160
rect 9216 4126 9222 4160
rect 9176 4088 9222 4126
rect 9176 4054 9182 4088
rect 9216 4054 9222 4088
rect 9176 4016 9222 4054
rect 9176 3982 9182 4016
rect 9216 3982 9222 4016
tri 9066 3952 9086 3972 sw
tri 8995 3947 9000 3952 se
rect 9000 3947 9086 3952
tri 9086 3947 9091 3952 sw
tri 8992 3944 8995 3947 se
rect 8995 3944 9091 3947
tri 9091 3944 9094 3947 sw
rect 9176 3944 9222 3982
rect 9332 4808 9378 4820
rect 9332 4774 9338 4808
rect 9372 4774 9378 4808
rect 9332 4736 9378 4774
rect 9332 4702 9338 4736
rect 9372 4702 9378 4736
rect 9332 4664 9378 4702
rect 9332 4630 9338 4664
rect 9372 4630 9378 4664
rect 9332 4592 9378 4630
rect 9332 4558 9338 4592
rect 9372 4558 9378 4592
rect 9332 4520 9378 4558
rect 9332 4486 9338 4520
rect 9372 4486 9378 4520
rect 9332 4448 9378 4486
rect 9332 4414 9338 4448
rect 9372 4414 9378 4448
rect 9332 4376 9378 4414
rect 9332 4342 9338 4376
rect 9372 4342 9378 4376
rect 9332 4304 9378 4342
rect 9332 4270 9338 4304
rect 9372 4270 9378 4304
rect 9332 4232 9378 4270
rect 9332 4198 9338 4232
rect 9372 4198 9378 4232
rect 9332 4160 9378 4198
rect 9332 4126 9338 4160
rect 9372 4126 9378 4160
rect 9332 4088 9378 4126
rect 9332 4054 9338 4088
rect 9372 4054 9378 4088
rect 9332 4016 9378 4054
rect 9332 3982 9338 4016
rect 9372 3982 9378 4016
rect 9456 4808 9502 4820
rect 9456 4774 9462 4808
rect 9496 4774 9502 4808
rect 9456 4736 9502 4774
rect 9456 4702 9462 4736
rect 9496 4702 9502 4736
rect 9456 4664 9502 4702
rect 9609 4808 9661 4820
rect 9609 4806 9618 4808
rect 9652 4806 9661 4808
rect 9609 4736 9661 4754
rect 9609 4723 9618 4736
rect 9652 4723 9661 4736
rect 9609 4665 9661 4671
tri 9609 4664 9610 4665 ne
rect 9610 4664 9660 4665
tri 9660 4664 9661 4665 nw
rect 9736 4808 9782 4820
rect 9736 4774 9742 4808
rect 9776 4774 9782 4808
rect 9736 4736 9782 4774
rect 9736 4702 9742 4736
rect 9776 4702 9782 4736
rect 9736 4664 9782 4702
rect 9889 4808 9941 4820
rect 9889 4806 9898 4808
rect 9932 4806 9941 4808
rect 9889 4736 9941 4754
rect 9889 4723 9898 4736
rect 9932 4723 9941 4736
rect 9889 4665 9941 4671
tri 9889 4664 9890 4665 ne
rect 9890 4664 9940 4665
tri 9940 4664 9941 4665 nw
rect 10048 4808 10094 4820
rect 10048 4774 10054 4808
rect 10088 4774 10094 4808
rect 10048 4736 10094 4774
rect 10048 4702 10054 4736
rect 10088 4702 10094 4736
rect 10048 4664 10094 4702
rect 10322 4808 10374 4820
rect 10322 4806 10331 4808
rect 10365 4806 10374 4808
rect 10322 4736 10374 4754
rect 10322 4723 10331 4736
rect 10365 4723 10374 4736
rect 10322 4665 10374 4671
tri 10322 4664 10323 4665 ne
rect 10323 4664 10373 4665
tri 10373 4664 10374 4665 nw
rect 10481 4808 10527 4820
rect 10481 4774 10487 4808
rect 10521 4774 10527 4808
rect 10481 4736 10527 4774
rect 10481 4702 10487 4736
rect 10521 4702 10527 4736
rect 10481 4664 10527 4702
rect 10634 4808 10686 4820
rect 10634 4806 10643 4808
rect 10677 4806 10686 4808
rect 10634 4736 10686 4754
rect 10634 4723 10643 4736
rect 10677 4723 10686 4736
rect 10634 4665 10686 4671
tri 10634 4664 10635 4665 ne
rect 10635 4664 10685 4665
tri 10685 4664 10686 4665 nw
rect 10793 4808 10839 4820
rect 10793 4774 10799 4808
rect 10833 4774 10839 4808
rect 10793 4736 10839 4774
rect 10793 4702 10799 4736
rect 10833 4702 10839 4736
rect 10793 4664 10839 4702
rect 10946 4808 10998 4820
rect 10946 4806 10955 4808
rect 10989 4806 10998 4808
rect 10946 4736 10998 4754
rect 10946 4723 10955 4736
rect 10989 4723 10998 4736
rect 10946 4665 10998 4671
tri 10946 4664 10947 4665 ne
rect 10947 4664 10997 4665
tri 10997 4664 10998 4665 nw
rect 11105 4808 11151 4820
rect 11105 4774 11111 4808
rect 11145 4774 11151 4808
rect 11105 4736 11151 4774
rect 11105 4702 11111 4736
rect 11145 4702 11151 4736
rect 11105 4664 11151 4702
rect 9456 4630 9462 4664
rect 9496 4630 9502 4664
tri 9610 4662 9612 4664 ne
rect 9456 4592 9502 4630
rect 9456 4558 9462 4592
rect 9496 4558 9502 4592
rect 9456 4520 9502 4558
rect 9456 4486 9462 4520
rect 9496 4486 9502 4520
rect 9456 4448 9502 4486
rect 9456 4414 9462 4448
rect 9496 4414 9502 4448
rect 9456 4376 9502 4414
rect 9456 4342 9462 4376
rect 9496 4342 9502 4376
rect 9456 4304 9502 4342
rect 9456 4270 9462 4304
rect 9496 4270 9502 4304
rect 9456 4232 9502 4270
rect 9456 4198 9462 4232
rect 9496 4198 9502 4232
rect 9456 4160 9502 4198
rect 9456 4126 9462 4160
rect 9496 4126 9502 4160
rect 9456 4088 9502 4126
rect 9456 4054 9462 4088
rect 9496 4054 9502 4088
rect 9456 4026 9502 4054
rect 9612 4630 9618 4664
rect 9652 4630 9658 4664
tri 9658 4662 9660 4664 nw
rect 9612 4592 9658 4630
rect 9612 4558 9618 4592
rect 9652 4558 9658 4592
rect 9612 4520 9658 4558
rect 9612 4486 9618 4520
rect 9652 4486 9658 4520
rect 9612 4448 9658 4486
rect 9612 4414 9618 4448
rect 9652 4414 9658 4448
rect 9612 4376 9658 4414
rect 9612 4342 9618 4376
rect 9652 4342 9658 4376
rect 9736 4630 9742 4664
rect 9776 4630 9782 4664
tri 9890 4662 9892 4664 ne
rect 9736 4592 9782 4630
rect 9736 4558 9742 4592
rect 9776 4558 9782 4592
rect 9736 4520 9782 4558
rect 9736 4486 9742 4520
rect 9776 4486 9782 4520
rect 9736 4448 9782 4486
rect 9736 4414 9742 4448
rect 9776 4414 9782 4448
rect 9736 4376 9782 4414
tri 9726 4342 9736 4352 se
rect 9736 4342 9742 4376
rect 9776 4343 9782 4376
rect 9892 4630 9898 4664
rect 9932 4630 9938 4664
tri 9938 4662 9940 4664 nw
rect 9892 4592 9938 4630
rect 9892 4558 9898 4592
rect 9932 4558 9938 4592
rect 9892 4520 9938 4558
rect 9892 4486 9898 4520
rect 9932 4486 9938 4520
rect 9892 4448 9938 4486
rect 9892 4414 9898 4448
rect 9932 4414 9938 4448
rect 9892 4376 9938 4414
rect 10048 4630 10054 4664
rect 10088 4630 10094 4664
tri 10323 4662 10325 4664 ne
rect 10048 4592 10094 4630
rect 10048 4558 10054 4592
rect 10088 4558 10094 4592
rect 10048 4520 10094 4558
rect 10048 4486 10054 4520
rect 10088 4486 10094 4520
rect 10048 4448 10094 4486
rect 10048 4414 10054 4448
rect 10088 4414 10094 4448
rect 10048 4380 10094 4414
rect 10325 4630 10331 4664
rect 10365 4630 10371 4664
tri 10371 4662 10373 4664 nw
rect 10325 4592 10371 4630
rect 10325 4558 10331 4592
rect 10365 4558 10371 4592
rect 10325 4520 10371 4558
rect 10325 4486 10331 4520
rect 10365 4486 10371 4520
rect 10325 4448 10371 4486
rect 10325 4414 10331 4448
rect 10365 4414 10371 4448
tri 9782 4343 9795 4356 sw
rect 9776 4342 9795 4343
tri 9795 4342 9796 4343 sw
rect 9892 4342 9898 4376
rect 9932 4342 9938 4376
rect 9612 4304 9658 4342
tri 9721 4337 9726 4342 se
rect 9726 4337 9796 4342
tri 9796 4337 9801 4342 sw
rect 9612 4270 9618 4304
rect 9652 4270 9658 4304
rect 9612 4232 9658 4270
tri 9706 4322 9721 4337 se
rect 9721 4323 9801 4337
tri 9801 4323 9815 4337 sw
rect 9721 4322 9815 4323
tri 9815 4322 9816 4323 sw
rect 9706 4270 9712 4322
rect 9764 4304 9776 4322
rect 9828 4270 9834 4322
rect 9892 4304 9938 4342
rect 9892 4270 9898 4304
rect 9932 4270 9938 4304
tri 9706 4265 9711 4270 ne
rect 9711 4265 9811 4270
tri 9811 4265 9816 4270 nw
tri 9711 4263 9713 4265 ne
rect 9713 4263 9809 4265
tri 9809 4263 9811 4265 nw
tri 9713 4254 9722 4263 ne
rect 9722 4254 9800 4263
tri 9800 4254 9809 4263 nw
tri 9722 4248 9728 4254 ne
rect 9728 4252 9798 4254
tri 9798 4252 9800 4254 nw
rect 9728 4248 9794 4252
tri 9794 4248 9798 4252 nw
tri 9728 4240 9736 4248 ne
rect 9612 4198 9618 4232
rect 9652 4198 9658 4232
rect 9612 4160 9658 4198
rect 9612 4126 9618 4160
rect 9652 4126 9658 4160
rect 9612 4088 9658 4126
rect 9612 4054 9618 4088
rect 9652 4054 9658 4088
tri 9502 4026 9517 4041 sw
rect 9456 4016 9517 4026
tri 9517 4016 9527 4026 sw
rect 9612 4016 9658 4054
tri 9312 3952 9332 3972 se
rect 9332 3952 9378 3982
tri 9448 4007 9456 4015 se
rect 9456 4007 9462 4016
rect 9496 4007 9527 4016
tri 9527 4007 9536 4016 sw
tri 9378 3952 9398 3972 sw
rect 9448 3955 9454 4007
rect 9506 3955 9518 4007
rect 9570 3955 9576 4007
rect 9612 3982 9618 4016
rect 9652 3982 9658 4016
tri 9448 3952 9451 3955 ne
rect 9451 3952 9533 3955
tri 9533 3952 9536 3955 nw
tri 9307 3947 9312 3952 se
rect 9312 3947 9398 3952
tri 9398 3947 9403 3952 sw
tri 9451 3947 9456 3952 ne
tri 9304 3944 9307 3947 se
rect 9307 3944 9403 3947
tri 9403 3944 9406 3947 sw
rect 9456 3944 9525 3952
tri 9525 3944 9533 3952 nw
rect 9612 3944 9658 3982
tri 8674 3938 8680 3944 se
rect 8680 3938 8714 3944
rect 8748 3938 8771 3944
tri 8771 3938 8777 3944 sw
rect 8476 3876 8522 3916
rect 8649 3886 8655 3938
rect 8707 3910 8714 3938
rect 8707 3886 8719 3910
rect 8771 3886 8777 3938
tri 8674 3878 8682 3886 ne
rect 8682 3879 8770 3886
tri 8770 3879 8777 3886 nw
rect 8864 3910 8870 3944
rect 8904 3910 8910 3944
tri 8986 3938 8992 3944 se
rect 8992 3938 9026 3944
rect 9060 3938 9094 3944
tri 9094 3938 9100 3944 sw
rect 8682 3878 8769 3879
tri 8769 3878 8770 3879 nw
rect 8476 3842 8482 3876
rect 8516 3842 8522 3876
tri 8682 3872 8688 3878 ne
rect 8688 3872 8763 3878
tri 8763 3872 8769 3878 nw
rect 8864 3872 8910 3910
rect 8972 3886 8978 3938
rect 9030 3886 9042 3910
rect 9094 3886 9100 3938
tri 8986 3879 8993 3886 ne
rect 8993 3879 9093 3886
tri 9093 3879 9100 3886 nw
rect 9176 3910 9182 3944
rect 9216 3910 9222 3944
tri 9298 3938 9304 3944 se
rect 9304 3938 9338 3944
rect 9372 3938 9406 3944
tri 9406 3938 9412 3944 sw
tri 8993 3878 8994 3879 ne
rect 8994 3878 9092 3879
tri 9092 3878 9093 3879 nw
tri 9175 3878 9176 3879 se
rect 9176 3878 9222 3910
rect 9290 3886 9296 3938
rect 9348 3886 9360 3910
rect 9412 3886 9418 3938
rect 9456 3910 9462 3944
rect 9496 3938 9519 3944
tri 9519 3938 9525 3944 nw
rect 9496 3910 9502 3938
tri 9502 3921 9519 3938 nw
tri 9298 3878 9306 3886 ne
rect 9306 3878 9404 3886
tri 9404 3878 9412 3886 nw
tri 8994 3872 9000 3878 ne
rect 9000 3872 9086 3878
tri 9086 3872 9092 3878 nw
tri 9169 3872 9175 3878 se
rect 9175 3872 9222 3878
tri 9306 3872 9312 3878 ne
rect 9312 3872 9398 3878
tri 9398 3872 9404 3878 nw
rect 9456 3872 9502 3910
tri 8688 3863 8697 3872 ne
rect 8697 3863 8714 3872
tri 8697 3852 8708 3863 ne
rect 8476 3802 8522 3842
rect 8708 3838 8714 3863
rect 8748 3838 8754 3872
tri 8754 3863 8763 3872 nw
rect 8708 3826 8754 3838
rect 8864 3838 8870 3872
rect 8904 3838 8910 3872
tri 9000 3852 9020 3872 ne
rect 8864 3826 8910 3838
rect 9020 3838 9026 3872
rect 9060 3838 9066 3872
tri 9066 3852 9086 3872 nw
tri 9149 3852 9169 3872 se
rect 9169 3852 9182 3872
tri 9135 3838 9149 3852 se
rect 9149 3838 9182 3852
rect 9216 3838 9222 3872
tri 9312 3852 9332 3872 ne
rect 9020 3826 9066 3838
tri 9123 3826 9135 3838 se
rect 9135 3826 9222 3838
rect 9332 3838 9338 3872
rect 9372 3838 9378 3872
tri 9378 3852 9398 3872 nw
rect 9332 3826 9378 3838
rect 9456 3838 9462 3872
rect 9496 3838 9502 3872
rect 9456 3826 9502 3838
rect 9612 3910 9618 3944
rect 9652 3910 9658 3944
rect 9612 3872 9658 3910
rect 9612 3838 9618 3872
rect 9652 3838 9658 3872
rect 9612 3826 9658 3838
rect 9736 4232 9782 4248
tri 9782 4236 9794 4248 nw
rect 9736 4198 9742 4232
rect 9776 4198 9782 4232
rect 9736 4160 9782 4198
rect 9736 4126 9742 4160
rect 9776 4126 9782 4160
rect 9736 4088 9782 4126
rect 9736 4054 9742 4088
rect 9776 4054 9782 4088
rect 9736 4016 9782 4054
rect 9736 3982 9742 4016
rect 9776 3982 9782 4016
rect 9736 3944 9782 3982
rect 9736 3910 9742 3944
rect 9776 3910 9782 3944
rect 9736 3872 9782 3910
rect 9736 3838 9742 3872
rect 9776 3838 9782 3872
rect 9736 3826 9782 3838
rect 9892 4232 9938 4270
rect 10045 4376 10097 4380
rect 10045 4374 10054 4376
rect 10088 4374 10097 4376
rect 10045 4310 10097 4322
rect 10045 4252 10097 4258
rect 10325 4376 10371 4414
rect 10325 4342 10331 4376
rect 10365 4342 10371 4376
rect 10325 4304 10371 4342
rect 10325 4270 10331 4304
rect 10365 4270 10371 4304
rect 9892 4198 9898 4232
rect 9932 4198 9938 4232
rect 9892 4160 9938 4198
rect 9892 4126 9898 4160
rect 9932 4126 9938 4160
rect 9892 4088 9938 4126
rect 9892 4054 9898 4088
rect 9932 4054 9938 4088
rect 9892 4016 9938 4054
rect 9892 3982 9898 4016
rect 9932 3982 9938 4016
rect 9892 3944 9938 3982
rect 9892 3910 9898 3944
rect 9932 3910 9938 3944
rect 9892 3872 9938 3910
rect 9892 3838 9898 3872
rect 9932 3838 9938 3872
rect 9892 3826 9938 3838
rect 10048 4232 10094 4252
rect 10048 4198 10054 4232
rect 10088 4198 10094 4232
rect 10325 4232 10371 4270
tri 10094 4198 10106 4210 sw
rect 10325 4198 10331 4232
rect 10365 4198 10371 4232
rect 10048 4189 10106 4198
tri 10106 4189 10115 4198 sw
rect 10048 4185 10115 4189
tri 10115 4185 10119 4189 sw
rect 10048 4182 10119 4185
tri 10119 4182 10122 4185 sw
rect 10048 4179 10122 4182
tri 10122 4179 10125 4182 sw
rect 10048 4174 10125 4179
tri 10125 4174 10130 4179 sw
rect 10048 4160 10130 4174
rect 10048 4126 10054 4160
rect 10088 4126 10130 4160
rect 10048 4088 10130 4126
rect 10048 4054 10054 4088
rect 10088 4054 10130 4088
rect 10048 4016 10130 4054
rect 10048 3982 10054 4016
rect 10088 3982 10130 4016
rect 10048 3944 10130 3982
rect 10048 3910 10054 3944
rect 10088 3910 10130 3944
rect 10048 3878 10130 3910
rect 10325 4160 10371 4198
rect 10481 4630 10487 4664
rect 10521 4630 10527 4664
tri 10635 4662 10637 4664 ne
rect 10481 4592 10527 4630
rect 10481 4558 10487 4592
rect 10521 4558 10527 4592
rect 10481 4520 10527 4558
rect 10481 4486 10487 4520
rect 10521 4486 10527 4520
rect 10481 4448 10527 4486
rect 10481 4414 10487 4448
rect 10521 4414 10527 4448
rect 10481 4376 10527 4414
rect 10481 4342 10487 4376
rect 10521 4342 10527 4376
rect 10481 4304 10527 4342
rect 10481 4270 10487 4304
rect 10521 4270 10527 4304
rect 10481 4232 10527 4270
rect 10481 4198 10487 4232
rect 10521 4198 10527 4232
rect 10325 4126 10331 4160
rect 10365 4126 10371 4160
rect 10325 4088 10371 4126
rect 10325 4054 10331 4088
rect 10365 4054 10371 4088
rect 10325 4016 10371 4054
tri 10478 4176 10481 4179 se
rect 10481 4176 10527 4198
rect 10637 4630 10643 4664
rect 10677 4630 10683 4664
tri 10683 4662 10685 4664 nw
rect 10637 4592 10683 4630
rect 10637 4558 10643 4592
rect 10677 4558 10683 4592
rect 10637 4520 10683 4558
rect 10637 4486 10643 4520
rect 10677 4486 10683 4520
rect 10637 4448 10683 4486
rect 10637 4414 10643 4448
rect 10677 4414 10683 4448
rect 10637 4376 10683 4414
rect 10637 4342 10643 4376
rect 10677 4342 10683 4376
rect 10637 4304 10683 4342
rect 10637 4270 10643 4304
rect 10677 4270 10683 4304
rect 10637 4232 10683 4270
rect 10637 4198 10643 4232
rect 10677 4198 10683 4232
tri 10527 4176 10530 4179 sw
rect 10478 4170 10530 4176
rect 10478 4104 10530 4118
rect 10478 4046 10530 4052
tri 10478 4043 10481 4046 ne
rect 10325 3982 10331 4016
rect 10365 3982 10371 4016
rect 10325 3944 10371 3982
rect 10325 3910 10331 3944
rect 10365 3910 10371 3944
tri 10130 3878 10132 3880 sw
rect 10048 3872 10132 3878
tri 10132 3872 10138 3878 sw
rect 10325 3872 10371 3910
rect 10048 3838 10054 3872
rect 10088 3855 10138 3872
tri 10138 3855 10155 3872 sw
rect 10088 3838 10155 3855
tri 10155 3838 10172 3855 sw
rect 10325 3838 10331 3872
rect 10365 3838 10371 3872
rect 10048 3826 10172 3838
tri 9117 3820 9123 3826 se
rect 9123 3825 9222 3826
rect 9123 3820 9217 3825
tri 9217 3820 9222 3825 nw
tri 10086 3820 10092 3826 ne
rect 10092 3820 10172 3826
tri 10172 3820 10190 3838 sw
rect 10325 3826 10371 3838
rect 10481 4016 10527 4046
tri 10527 4043 10530 4046 nw
rect 10637 4160 10683 4198
rect 10793 4630 10799 4664
rect 10833 4630 10839 4664
tri 10947 4662 10949 4664 ne
rect 10793 4592 10839 4630
rect 10793 4558 10799 4592
rect 10833 4558 10839 4592
rect 10793 4520 10839 4558
rect 10793 4486 10799 4520
rect 10833 4486 10839 4520
rect 10793 4448 10839 4486
rect 10793 4414 10799 4448
rect 10833 4414 10839 4448
rect 10793 4376 10839 4414
rect 10793 4342 10799 4376
rect 10833 4342 10839 4376
rect 10793 4304 10839 4342
rect 10793 4270 10799 4304
rect 10833 4270 10839 4304
rect 10793 4232 10839 4270
rect 10793 4198 10799 4232
rect 10833 4198 10839 4232
tri 10790 4179 10793 4182 se
rect 10793 4179 10839 4198
rect 10949 4630 10955 4664
rect 10989 4630 10995 4664
tri 10995 4662 10997 4664 nw
rect 10949 4592 10995 4630
rect 10949 4558 10955 4592
rect 10989 4558 10995 4592
rect 10949 4520 10995 4558
rect 10949 4486 10955 4520
rect 10989 4486 10995 4520
rect 10949 4448 10995 4486
rect 10949 4414 10955 4448
rect 10989 4414 10995 4448
rect 10949 4376 10995 4414
rect 10949 4342 10955 4376
rect 10989 4342 10995 4376
rect 10949 4304 10995 4342
rect 10949 4270 10955 4304
rect 10989 4270 10995 4304
rect 10949 4232 10995 4270
rect 10949 4198 10955 4232
rect 10989 4198 10995 4232
rect 10637 4126 10643 4160
rect 10677 4126 10683 4160
rect 10637 4088 10683 4126
rect 10637 4054 10643 4088
rect 10677 4054 10683 4088
rect 10481 3982 10487 4016
rect 10521 3982 10527 4016
rect 10481 3944 10527 3982
rect 10481 3910 10487 3944
rect 10521 3910 10527 3944
rect 10481 3872 10527 3910
rect 10481 3838 10487 3872
rect 10521 3838 10527 3872
rect 10481 3826 10527 3838
rect 10637 4016 10683 4054
tri 10787 4176 10790 4179 se
rect 10790 4176 10839 4179
rect 10787 4170 10839 4176
rect 10787 4104 10839 4118
rect 10787 4046 10839 4052
tri 10787 4043 10790 4046 ne
rect 10790 4043 10839 4046
tri 10790 4040 10793 4043 ne
rect 10637 3982 10643 4016
rect 10677 3982 10683 4016
rect 10637 3944 10683 3982
rect 10637 3910 10643 3944
rect 10677 3910 10683 3944
rect 10637 3872 10683 3910
rect 10637 3838 10643 3872
rect 10677 3838 10683 3872
rect 10637 3826 10683 3838
rect 10793 4016 10839 4043
rect 10793 3982 10799 4016
rect 10833 3982 10839 4016
rect 10793 3944 10839 3982
rect 10793 3910 10799 3944
rect 10833 3910 10839 3944
rect 10793 3872 10839 3910
rect 10793 3838 10799 3872
rect 10833 3838 10839 3872
rect 10793 3826 10839 3838
rect 10867 4179 10919 4185
rect 10867 4113 10919 4127
rect 10867 4055 10919 4061
rect 10949 4160 10995 4198
rect 10949 4126 10955 4160
rect 10989 4126 10995 4160
rect 10949 4088 10995 4126
tri 9115 3818 9117 3820 se
rect 9117 3818 9215 3820
tri 9215 3818 9217 3820 nw
tri 10092 3818 10094 3820 ne
rect 10094 3818 10190 3820
tri 10190 3818 10192 3820 sw
tri 9101 3804 9115 3818 se
rect 9115 3804 9201 3818
tri 9201 3804 9215 3818 nw
tri 10094 3804 10108 3818 ne
rect 10108 3804 10192 3818
tri 10192 3804 10206 3818 sw
rect 8476 3768 8482 3802
rect 8516 3768 8522 3802
tri 9076 3779 9101 3804 se
rect 9101 3779 9176 3804
tri 9176 3779 9201 3804 nw
tri 10108 3779 10133 3804 ne
rect 10133 3790 10206 3804
tri 10206 3790 10220 3804 sw
rect 10133 3779 10220 3790
tri 9067 3770 9076 3779 se
rect 9076 3770 9167 3779
tri 9167 3770 9176 3779 nw
tri 10133 3770 10142 3779 ne
rect 10142 3770 10220 3779
tri 10220 3770 10240 3790 sw
tri 10847 3770 10867 3790 se
rect 10867 3770 10918 4055
rect 10949 4054 10955 4088
rect 10989 4054 10995 4088
rect 10949 4016 10995 4054
rect 10949 3982 10955 4016
rect 10989 3982 10995 4016
rect 10949 3944 10995 3982
rect 10949 3910 10955 3944
rect 10989 3910 10995 3944
rect 11105 4630 11111 4664
rect 11145 4630 11151 4664
rect 11105 4592 11151 4630
rect 11105 4558 11111 4592
rect 11145 4558 11151 4592
rect 11105 4520 11151 4558
rect 11105 4486 11111 4520
rect 11145 4486 11151 4520
rect 11105 4448 11151 4486
rect 11105 4414 11111 4448
rect 11145 4414 11151 4448
rect 11105 4376 11151 4414
rect 11105 4342 11111 4376
rect 11145 4342 11151 4376
rect 11105 4304 11151 4342
rect 11105 4270 11111 4304
rect 11145 4270 11151 4304
rect 11105 4232 11151 4270
rect 11105 4198 11111 4232
rect 11145 4198 11151 4232
rect 11105 4160 11151 4198
rect 11105 4126 11111 4160
rect 11145 4126 11151 4160
rect 11105 4088 11151 4126
rect 11105 4054 11111 4088
rect 11145 4054 11151 4088
rect 11105 4016 11151 4054
rect 11105 3982 11111 4016
rect 11145 3982 11151 4016
rect 11105 3944 11151 3982
rect 10949 3872 10995 3910
rect 10949 3838 10955 3872
rect 10989 3838 10995 3872
rect 10949 3826 10995 3838
tri 11103 3927 11105 3929 se
rect 11105 3927 11111 3944
rect 11103 3921 11111 3927
rect 11145 3929 11151 3944
rect 11184 4809 11236 4815
rect 11184 4723 11236 4757
tri 11151 3929 11153 3931 sw
rect 11145 3927 11153 3929
tri 11153 3927 11155 3929 sw
rect 11145 3921 11155 3927
rect 11103 3855 11111 3869
rect 11145 3855 11155 3869
rect 11103 3797 11155 3803
tri 10918 3770 10938 3790 sw
tri 9065 3768 9067 3770 se
rect 9067 3768 9165 3770
tri 9165 3768 9167 3770 nw
tri 10142 3768 10144 3770 ne
rect 10144 3768 10240 3770
tri 10240 3768 10242 3770 sw
tri 10845 3768 10847 3770 se
rect 10847 3768 10938 3770
rect 8476 3728 8522 3768
rect 8476 3694 8482 3728
rect 8516 3694 8522 3728
rect 8476 3654 8522 3694
rect 8476 3620 8482 3654
rect 8516 3620 8522 3654
rect 8476 3580 8522 3620
rect 8476 3546 8482 3580
rect 8516 3546 8522 3580
rect 8476 3506 8522 3546
rect 8646 3756 8698 3768
rect 8646 3722 8657 3756
rect 8691 3722 8698 3756
rect 8646 3684 8698 3722
rect 8646 3667 8657 3684
rect 8691 3667 8698 3684
rect 9065 3763 9160 3768
tri 9160 3763 9165 3768 nw
tri 10144 3763 10149 3768 ne
rect 10149 3763 10242 3768
tri 10242 3763 10247 3768 sw
tri 10840 3763 10845 3768 se
rect 10845 3763 10938 3768
tri 10938 3763 10945 3770 sw
rect 9065 3757 9154 3763
tri 9154 3757 9160 3763 nw
rect 9211 3757 9683 3763
tri 9683 3757 9689 3763 sw
rect 9800 3757 10023 3763
tri 10149 3757 10155 3763 ne
rect 10155 3762 10247 3763
tri 10247 3762 10248 3763 sw
tri 10839 3762 10840 3763 se
rect 10840 3762 10945 3763
tri 10945 3762 10946 3763 sw
rect 10155 3757 10248 3762
tri 10248 3757 10253 3762 sw
rect 9065 3751 9148 3757
tri 9148 3751 9154 3757 nw
rect 9211 3751 9689 3757
rect 9065 3669 9141 3751
tri 9141 3744 9148 3751 nw
rect 9211 3717 9223 3751
rect 9257 3717 9295 3751
rect 9329 3723 9689 3751
tri 9689 3723 9723 3757 sw
rect 9800 3723 9812 3757
rect 9846 3723 9895 3757
rect 9929 3723 9977 3757
rect 10011 3723 10023 3757
tri 10155 3756 10156 3757 ne
rect 10156 3756 10253 3757
tri 10253 3756 10254 3757 sw
rect 10387 3756 11103 3762
tri 10156 3735 10177 3756 ne
rect 10177 3735 10254 3756
tri 10254 3735 10275 3756 sw
rect 9329 3722 9723 3723
tri 9723 3722 9724 3723 sw
rect 9800 3722 10023 3723
tri 10023 3722 10036 3735 sw
tri 10177 3722 10190 3735 ne
rect 10190 3722 10275 3735
tri 10275 3722 10288 3735 sw
rect 10387 3722 10399 3756
rect 10433 3722 10473 3756
rect 10507 3722 10546 3756
rect 10580 3722 10619 3756
rect 10653 3722 10692 3756
rect 10726 3722 10765 3756
rect 10799 3722 10838 3756
rect 10872 3722 10911 3756
rect 10945 3722 10984 3756
rect 11018 3722 11057 3756
rect 11091 3722 11103 3756
rect 9329 3717 9724 3722
tri 9724 3717 9729 3722 sw
rect 9800 3717 10036 3722
tri 10036 3717 10041 3722 sw
tri 10190 3717 10195 3722 ne
rect 10195 3717 10288 3722
tri 10288 3717 10293 3722 sw
rect 9211 3711 9729 3717
tri 9729 3711 9735 3717 sw
tri 9966 3711 9972 3717 ne
rect 9972 3716 10041 3717
tri 10041 3716 10042 3717 sw
tri 10195 3716 10196 3717 ne
rect 10196 3716 10293 3717
tri 10293 3716 10294 3717 sw
rect 10387 3716 11103 3722
rect 9972 3711 10042 3716
tri 10042 3711 10047 3716 sw
tri 10196 3711 10201 3716 ne
rect 10201 3711 10294 3716
tri 10294 3711 10299 3716 sw
tri 9607 3696 9622 3711 ne
rect 9622 3696 9735 3711
tri 9735 3696 9750 3711 sw
tri 9972 3696 9987 3711 ne
rect 9987 3696 10047 3711
tri 10047 3696 10062 3711 sw
tri 10201 3696 10216 3711 ne
rect 10216 3696 10299 3711
tri 10299 3696 10314 3711 sw
tri 9622 3676 9642 3696 ne
rect 9642 3676 9750 3696
tri 9750 3676 9770 3696 sw
rect 9642 3669 9770 3676
tri 9987 3672 10011 3696 ne
rect 10011 3672 10062 3696
tri 10062 3672 10086 3696 sw
tri 10216 3672 10240 3696 ne
rect 10240 3672 10314 3696
tri 10314 3672 10338 3696 sw
tri 10011 3669 10014 3672 ne
rect 10014 3669 10086 3672
tri 10086 3669 10089 3672 sw
tri 10240 3669 10243 3672 ne
rect 10243 3669 10338 3672
tri 10338 3669 10341 3672 sw
rect 9013 3617 9019 3669
rect 9071 3617 9083 3669
rect 9135 3617 9141 3669
rect 9186 3617 9192 3669
rect 9244 3617 9256 3669
rect 9308 3657 9583 3669
rect 9308 3623 9465 3657
rect 9499 3623 9537 3657
rect 9571 3623 9583 3657
rect 9308 3617 9583 3623
rect 9642 3617 9648 3669
rect 9700 3617 9712 3669
rect 9764 3617 9770 3669
tri 10014 3664 10019 3669 ne
rect 10019 3664 10089 3669
tri 10089 3664 10094 3669 sw
tri 10243 3664 10248 3669 ne
rect 10248 3664 10341 3669
tri 10341 3664 10346 3669 sw
tri 10019 3660 10023 3664 ne
rect 10023 3660 10077 3664
tri 10023 3656 10027 3660 ne
rect 10027 3656 10077 3660
tri 10027 3643 10040 3656 ne
rect 10040 3643 10077 3656
tri 10040 3617 10066 3643 ne
rect 10066 3617 10077 3643
rect 8646 3603 8698 3615
tri 10066 3612 10071 3617 ne
rect 10071 3612 10077 3617
rect 10129 3612 10141 3664
rect 10193 3612 10199 3664
tri 10248 3659 10253 3664 ne
rect 10253 3659 10346 3664
tri 10346 3659 10351 3664 sw
tri 10253 3656 10256 3659 ne
rect 10256 3656 10824 3659
tri 10256 3649 10263 3656 ne
rect 10263 3649 10824 3656
tri 10263 3643 10269 3649 ne
rect 10269 3643 10824 3649
tri 10269 3612 10300 3643 ne
rect 10300 3612 10636 3643
tri 10300 3609 10303 3612 ne
rect 10303 3609 10636 3612
rect 10670 3609 10778 3643
rect 10812 3609 10824 3643
tri 10303 3603 10309 3609 ne
rect 10309 3603 10824 3609
tri 11180 3599 11184 3603 se
rect 11184 3599 11236 4671
tri 11164 3583 11180 3599 se
rect 11180 3583 11236 3599
tri 8841 3582 8842 3583 se
rect 8842 3582 10211 3583
tri 10211 3582 10212 3583 sw
tri 11163 3582 11164 3583 se
rect 11164 3582 11236 3583
tri 8825 3566 8841 3582 se
rect 8841 3572 10212 3582
tri 10212 3572 10222 3582 sw
tri 11153 3572 11163 3582 se
rect 11163 3572 11236 3582
rect 8841 3566 10222 3572
tri 10222 3566 10228 3572 sw
rect 10879 3566 11236 3572
tri 8815 3556 8825 3566 se
rect 8825 3556 10228 3566
tri 10228 3556 10238 3566 sw
rect 8646 3545 8698 3551
tri 8804 3545 8815 3556 se
rect 8815 3547 10723 3556
rect 8815 3545 8842 3547
tri 8792 3533 8804 3545 se
rect 8804 3533 8842 3545
tri 8842 3533 8856 3547 nw
tri 10161 3533 10175 3547 ne
rect 10175 3533 10723 3547
tri 8791 3532 8792 3533 se
rect 8792 3532 8841 3533
tri 8841 3532 8842 3533 nw
tri 10175 3532 10176 3533 ne
rect 10176 3532 10723 3533
tri 8785 3526 8791 3532 se
rect 8791 3526 8835 3532
tri 8835 3526 8841 3532 nw
tri 10176 3526 10182 3532 ne
rect 10182 3526 10723 3532
tri 8777 3518 8785 3526 se
rect 8785 3518 8827 3526
tri 8827 3518 8835 3526 nw
tri 10182 3518 10190 3526 ne
rect 10190 3518 10723 3526
tri 8768 3509 8777 3518 se
rect 8777 3509 8818 3518
tri 8818 3509 8827 3518 nw
tri 9722 3515 9725 3518 se
rect 9725 3515 9731 3518
rect 8877 3509 9731 3515
rect 9783 3509 9799 3518
rect 9851 3515 9857 3518
tri 9857 3515 9860 3518 sw
tri 10190 3515 10193 3518 ne
rect 10193 3515 10723 3518
rect 9851 3509 9871 3515
rect 8476 3472 8482 3506
rect 8516 3472 8522 3506
tri 8742 3483 8768 3509 se
rect 8768 3483 8792 3509
tri 8792 3483 8818 3509 nw
tri 8734 3475 8742 3483 se
rect 8742 3475 8784 3483
tri 8784 3475 8792 3483 nw
rect 8877 3475 8889 3509
rect 8923 3475 8961 3509
rect 8995 3475 9033 3509
rect 9067 3475 9105 3509
rect 9139 3475 9177 3509
rect 9211 3475 9249 3509
rect 9283 3475 9321 3509
rect 9355 3475 9393 3509
rect 9427 3475 9465 3509
rect 9499 3475 9537 3509
rect 9571 3475 9609 3509
rect 9643 3475 9681 3509
rect 9715 3475 9731 3509
rect 9787 3475 9799 3509
rect 9859 3475 9871 3509
tri 10193 3504 10204 3515 ne
rect 10204 3504 10723 3515
rect 10775 3504 10787 3556
rect 10839 3504 10845 3556
rect 10879 3532 10891 3566
rect 10925 3532 10963 3566
rect 10997 3532 11236 3566
rect 10879 3526 11236 3532
rect 11290 4807 11298 4840
rect 11332 4807 11379 4840
tri 11379 4826 11393 4840 nw
tri 11491 4826 11505 4840 ne
rect 11505 4826 11515 4840
tri 11505 4822 11509 4826 ne
rect 11509 4824 11515 4826
rect 11567 4824 11580 4876
rect 11632 4824 11644 4876
rect 11696 4872 19755 4876
rect 11696 4824 11702 4872
rect 11342 4755 11379 4807
rect 11290 4732 11298 4755
rect 11332 4732 11379 4755
rect 11290 4721 11379 4732
rect 11509 4782 11702 4824
rect 11509 4730 11515 4782
rect 11567 4730 11580 4782
rect 11632 4730 11644 4782
rect 11696 4730 11702 4782
rect 18571 4744 19157 4872
rect 19807 4827 19819 4879
rect 19871 4827 19883 4879
rect 19935 4827 19947 4879
rect 19999 4840 20016 4879
rect 19755 4806 19973 4827
rect 20007 4806 20016 4840
rect 19755 4788 20016 4806
rect 11342 4669 11379 4721
rect 19023 4720 19109 4744
rect 19807 4736 19819 4788
rect 19871 4736 19883 4788
rect 19935 4736 19947 4788
rect 19999 4767 20016 4788
rect 19755 4733 19973 4736
rect 20007 4733 20016 4767
rect 19755 4730 20016 4733
rect 19823 4720 20016 4730
tri 19930 4694 19956 4720 ne
rect 19956 4694 20016 4720
tri 19956 4686 19964 4694 ne
rect 19964 4686 19973 4694
rect 20007 4686 20016 4694
rect 11290 4658 11298 4669
rect 11332 4658 11379 4669
tri 17385 4660 17397 4672 se
rect 17397 4660 17443 4672
rect 11290 4618 11379 4658
tri 17381 4656 17385 4660 se
rect 17385 4656 17403 4660
rect 11290 4584 11298 4618
rect 11332 4584 11379 4618
rect 11665 4593 11671 4645
rect 11723 4593 11735 4645
rect 11787 4642 11793 4645
tri 11793 4642 11796 4645 sw
rect 11787 4639 11796 4642
tri 11796 4639 11799 4642 sw
tri 17048 4639 17051 4642 se
rect 17051 4639 17057 4642
rect 11787 4633 17057 4639
rect 11787 4599 13493 4633
rect 13527 4599 13584 4633
rect 13618 4599 17057 4633
rect 11787 4598 17057 4599
rect 11787 4593 14415 4598
tri 14415 4593 14420 4598 nw
tri 14596 4593 14601 4598 ne
rect 14601 4593 17057 4598
tri 17048 4590 17051 4593 ne
rect 17051 4590 17057 4593
rect 17109 4590 17121 4642
rect 17173 4590 17179 4642
rect 17397 4626 17403 4656
rect 17437 4626 17443 4660
rect 17397 4604 17443 4626
rect 17523 4620 17529 4672
rect 17581 4620 17593 4672
rect 17645 4660 18036 4672
rect 17645 4626 17996 4660
rect 18030 4626 18036 4660
rect 17645 4620 18036 4626
tri 17362 4593 17373 4604 ne
rect 17373 4593 17443 4604
tri 17373 4590 17376 4593 ne
rect 17376 4590 17443 4593
tri 17376 4588 17378 4590 ne
rect 17378 4588 17443 4590
tri 17890 4588 17922 4620 ne
rect 17922 4588 18036 4620
rect 11290 4544 11379 4584
tri 17378 4569 17397 4588 ne
rect 14437 4565 14443 4568
tri 11472 4559 11478 4565 se
rect 11478 4559 14443 4565
rect 11290 4510 11298 4544
rect 11332 4510 11379 4544
rect 11290 4470 11379 4510
rect 11290 4436 11298 4470
rect 11332 4436 11379 4470
rect 11290 4396 11379 4436
rect 11290 4362 11298 4396
rect 11332 4362 11379 4396
rect 11290 4322 11379 4362
rect 11290 4288 11298 4322
rect 11332 4288 11379 4322
rect 11290 4248 11379 4288
rect 11290 4214 11298 4248
rect 11332 4214 11379 4248
rect 11290 4174 11379 4214
rect 11290 4140 11298 4174
rect 11332 4140 11379 4174
rect 11290 4100 11379 4140
rect 11290 4066 11298 4100
rect 11332 4066 11379 4100
rect 11290 4026 11379 4066
rect 11290 3992 11298 4026
rect 11332 3992 11379 4026
rect 11290 3952 11379 3992
rect 11290 3918 11298 3952
rect 11332 3918 11379 3952
rect 11290 3878 11379 3918
rect 11290 3844 11298 3878
rect 11332 3844 11379 3878
rect 11290 3804 11379 3844
rect 11290 3770 11298 3804
rect 11332 3770 11379 3804
rect 11290 3730 11379 3770
tri 11444 4531 11472 4559 se
rect 11472 4531 14443 4559
rect 11444 4519 14443 4531
rect 11444 4516 11526 4519
tri 11526 4516 11529 4519 nw
rect 14437 4516 14443 4519
rect 14495 4516 14507 4568
rect 14559 4565 14565 4568
rect 14559 4559 16839 4565
rect 14559 4525 16721 4559
rect 16755 4525 16793 4559
rect 16827 4525 16839 4559
rect 17397 4554 17403 4588
rect 17437 4554 17443 4588
tri 17922 4586 17924 4588 ne
rect 17924 4586 17996 4588
rect 17397 4542 17443 4554
rect 17678 4563 17724 4575
rect 17678 4529 17684 4563
rect 17718 4529 17724 4563
rect 17990 4554 17996 4586
rect 18030 4554 18036 4588
rect 17990 4542 18036 4554
tri 18392 4624 18421 4653 se
rect 18421 4624 18726 4653
rect 18392 4614 18726 4624
rect 18392 4601 18452 4614
tri 18452 4601 18465 4614 nw
tri 18707 4601 18720 4614 ne
rect 18720 4601 18726 4614
rect 18778 4601 18790 4653
rect 18842 4601 18848 4653
rect 19964 4621 20016 4634
rect 18392 4587 18438 4601
tri 18438 4587 18452 4601 nw
rect 14559 4519 16839 4525
tri 17672 4519 17678 4525 se
rect 17678 4519 17724 4529
rect 14559 4516 14565 4519
tri 17669 4516 17672 4519 se
rect 17672 4516 17724 4519
rect 11444 4514 11524 4516
tri 11524 4514 11526 4516 nw
tri 17667 4514 17669 4516 se
rect 17669 4514 17724 4516
rect 11444 4492 11502 4514
tri 11502 4492 11524 4514 nw
tri 17645 4492 17667 4514 se
rect 17667 4492 17724 4514
tri 17724 4492 17727 4495 sw
rect 11444 4491 11501 4492
tri 11501 4491 11502 4492 nw
tri 17644 4491 17645 4492 se
rect 17645 4491 17727 4492
tri 17727 4491 17728 4492 sw
rect 11290 3696 11298 3730
rect 11332 3696 11379 3730
rect 11290 3656 11379 3696
rect 11290 3622 11298 3656
rect 11332 3622 11379 3656
rect 11290 3582 11379 3622
rect 11290 3548 11298 3582
rect 11332 3548 11379 3582
rect 11290 3504 11379 3548
rect 8476 3432 8522 3472
tri 8729 3470 8734 3475 se
rect 8734 3470 8779 3475
tri 8779 3470 8784 3475 nw
tri 8725 3466 8729 3470 se
rect 8729 3466 8775 3470
tri 8775 3466 8779 3470 nw
rect 8877 3469 9731 3475
tri 9722 3466 9725 3469 ne
rect 9725 3466 9731 3469
rect 9783 3466 9799 3475
rect 9851 3469 9871 3475
rect 11290 3470 11298 3504
rect 11332 3470 11379 3504
rect 9851 3467 9858 3469
tri 9858 3467 9860 3469 nw
rect 9851 3466 9857 3467
tri 9857 3466 9858 3467 nw
tri 9934 3466 9935 3467 se
rect 9935 3466 9981 3467
tri 8714 3455 8725 3466 se
rect 8725 3455 8764 3466
tri 8764 3455 8775 3466 nw
tri 9923 3455 9934 3466 se
rect 9934 3464 9981 3466
tri 9981 3464 9984 3467 sw
rect 9934 3455 11097 3464
tri 8700 3441 8714 3455 se
rect 8714 3441 8750 3455
tri 8750 3441 8764 3455 nw
tri 9909 3441 9923 3455 se
rect 9923 3441 9941 3455
tri 8696 3437 8700 3441 se
rect 8700 3437 8746 3441
tri 8746 3437 8750 3441 nw
tri 9340 3437 9344 3441 se
rect 9344 3437 9350 3441
tri 8692 3433 8696 3437 se
rect 8696 3433 8742 3437
tri 8742 3433 8746 3437 nw
tri 8787 3433 8791 3437 se
rect 8791 3433 9350 3437
rect 8476 3398 8482 3432
rect 8516 3398 8522 3432
tri 8680 3421 8692 3433 se
rect 8692 3432 8741 3433
tri 8741 3432 8742 3433 nw
tri 8786 3432 8787 3433 se
rect 8787 3432 9350 3433
rect 8692 3421 8730 3432
tri 8730 3421 8741 3432 nw
tri 8775 3421 8786 3432 se
rect 8786 3421 9350 3432
tri 8679 3420 8680 3421 se
rect 8680 3420 8729 3421
tri 8729 3420 8730 3421 nw
tri 8774 3420 8775 3421 se
rect 8775 3420 9350 3421
tri 8660 3401 8679 3420 se
rect 8679 3401 8710 3420
tri 8710 3401 8729 3420 nw
tri 8755 3401 8774 3420 se
rect 8774 3401 9350 3420
rect 8476 3358 8522 3398
tri 8652 3393 8660 3401 se
rect 8660 3393 8702 3401
tri 8702 3393 8710 3401 nw
tri 8747 3393 8755 3401 se
rect 8755 3393 8797 3401
tri 8797 3393 8805 3401 nw
tri 9332 3393 9340 3401 ne
rect 9340 3393 9350 3401
tri 8648 3389 8652 3393 se
rect 8652 3389 8698 3393
tri 8698 3389 8702 3393 nw
tri 8743 3389 8747 3393 se
rect 8747 3389 8793 3393
tri 8793 3389 8797 3393 nw
tri 9340 3389 9344 3393 ne
rect 9344 3389 9350 3393
rect 9402 3389 9414 3441
rect 9466 3437 9472 3441
tri 9472 3437 9476 3441 sw
tri 9905 3437 9909 3441 se
rect 9909 3437 9941 3441
rect 9466 3421 9941 3437
rect 9975 3421 11097 3455
rect 9466 3412 11097 3421
rect 11149 3412 11161 3464
rect 11213 3412 11219 3464
tri 11279 3420 11290 3431 se
rect 11290 3420 11379 3470
tri 11271 3412 11279 3420 se
rect 11279 3412 11379 3420
rect 9466 3401 10044 3412
tri 10044 3401 10055 3412 nw
tri 11260 3401 11271 3412 se
rect 11271 3401 11379 3412
rect 9466 3393 9478 3401
tri 9478 3393 9486 3401 nw
tri 9905 3393 9913 3401 ne
rect 9913 3393 10036 3401
tri 10036 3393 10044 3401 nw
tri 11252 3393 11260 3401 se
rect 11260 3393 11379 3401
rect 9466 3389 9474 3393
tri 9474 3389 9478 3393 nw
tri 9913 3389 9917 3393 ne
rect 9917 3389 10019 3393
tri 8642 3383 8648 3389 se
rect 8648 3387 8696 3389
tri 8696 3387 8698 3389 nw
tri 8741 3387 8743 3389 se
rect 8743 3387 8791 3389
tri 8791 3387 8793 3389 nw
tri 9917 3387 9919 3389 ne
rect 9919 3387 10019 3389
rect 8648 3383 8692 3387
tri 8692 3383 8696 3387 nw
tri 8737 3383 8741 3387 se
rect 8741 3383 8774 3387
tri 8629 3370 8642 3383 se
rect 8642 3382 8691 3383
tri 8691 3382 8692 3383 nw
tri 8736 3382 8737 3383 se
rect 8737 3382 8774 3383
rect 8642 3370 8679 3382
tri 8679 3370 8691 3382 nw
tri 8724 3370 8736 3382 se
rect 8736 3370 8774 3382
tri 8774 3370 8791 3387 nw
tri 9919 3371 9935 3387 ne
rect 9935 3376 10019 3387
tri 10019 3376 10036 3393 nw
tri 11235 3376 11252 3393 se
rect 11252 3376 11298 3393
rect 9935 3370 10013 3376
tri 10013 3370 10019 3376 nw
rect 10174 3370 11298 3376
rect 8476 3324 8482 3358
rect 8516 3324 8522 3358
tri 8614 3355 8629 3370 se
rect 8629 3355 8664 3370
tri 8664 3355 8679 3370 nw
tri 8709 3355 8724 3370 se
rect 8724 3359 8763 3370
tri 8763 3359 8774 3370 nw
rect 8724 3355 8759 3359
tri 8759 3355 8763 3359 nw
tri 8808 3355 8812 3359 se
rect 8812 3355 9871 3359
tri 8612 3353 8614 3355 se
rect 8614 3353 8662 3355
tri 8662 3353 8664 3355 nw
tri 8707 3353 8709 3355 se
rect 8709 3353 8757 3355
tri 8757 3353 8759 3355 nw
tri 8806 3353 8808 3355 se
rect 8808 3353 9871 3355
tri 8596 3337 8612 3353 se
rect 8612 3337 8646 3353
tri 8646 3337 8662 3353 nw
tri 8691 3337 8707 3353 se
rect 8707 3342 8746 3353
tri 8746 3342 8757 3353 nw
tri 8795 3342 8806 3353 se
rect 8806 3342 8889 3353
rect 8707 3337 8741 3342
tri 8741 3337 8746 3342 nw
tri 8790 3337 8795 3342 se
rect 8795 3337 8889 3342
tri 8592 3333 8596 3337 se
rect 8596 3333 8642 3337
tri 8642 3333 8646 3337 nw
tri 8687 3333 8691 3337 se
rect 8691 3333 8723 3337
rect 8476 3284 8522 3324
tri 8578 3319 8592 3333 se
rect 8592 3332 8641 3333
tri 8641 3332 8642 3333 nw
tri 8686 3332 8687 3333 se
rect 8687 3332 8723 3333
rect 8592 3319 8628 3332
tri 8628 3319 8641 3332 nw
tri 8673 3319 8686 3332 se
rect 8686 3319 8723 3332
tri 8723 3319 8741 3337 nw
tri 8772 3319 8790 3337 se
rect 8790 3319 8889 3337
rect 8923 3319 8961 3353
rect 8995 3319 9033 3353
rect 9067 3319 9105 3353
rect 9139 3319 9177 3353
rect 9211 3319 9249 3353
rect 9283 3319 9321 3353
rect 9355 3319 9393 3353
rect 9427 3319 9465 3353
rect 9499 3319 9537 3353
rect 9571 3319 9609 3353
rect 9643 3319 9681 3353
rect 9715 3319 9753 3353
rect 9787 3319 9825 3353
rect 9859 3319 9871 3353
tri 8562 3303 8578 3319 se
rect 8578 3303 8612 3319
tri 8612 3303 8628 3319 nw
tri 8657 3303 8673 3319 se
rect 8673 3303 8707 3319
tri 8707 3303 8723 3319 nw
tri 8756 3303 8772 3319 se
rect 8772 3313 9871 3319
rect 9935 3355 9992 3370
rect 9935 3321 9941 3355
rect 9975 3349 9992 3355
tri 9992 3349 10013 3370 nw
rect 9975 3321 9981 3349
tri 9981 3338 9992 3349 nw
rect 8772 3303 8822 3313
tri 8822 3303 8832 3313 nw
rect 8476 3250 8482 3284
rect 8516 3250 8522 3284
rect 8476 3210 8522 3250
rect 8476 3176 8482 3210
rect 8516 3176 8522 3210
rect 8476 3136 8522 3176
rect 8476 3102 8482 3136
rect 8516 3102 8522 3136
rect 8476 3062 8522 3102
rect 8476 3028 8482 3062
rect 8516 3028 8522 3062
tri 8470 3014 8476 3020 se
rect 8476 3014 8522 3028
rect 8470 3008 8522 3014
rect 8470 2954 8482 2956
rect 8516 2954 8522 2956
rect 8470 2944 8522 2954
rect 8470 2886 8482 2892
tri 8470 2880 8476 2886 ne
rect 8476 2880 8482 2886
rect 8516 2880 8522 2892
rect 915 2703 8282 2727
tri 8282 2703 8306 2727 nw
rect 915 2693 8272 2703
tri 8272 2693 8282 2703 nw
rect 915 2691 953 2693
tri 953 2691 955 2693 nw
rect 915 2687 927 2691
rect 863 2675 927 2687
rect 915 2665 927 2675
tri 927 2665 953 2691 nw
rect 8348 2665 8400 2677
rect 915 2657 919 2665
tri 919 2657 927 2665 nw
tri 2022 2657 2030 2665 se
rect 2030 2657 8093 2665
tri 915 2653 919 2657 nw
tri 2018 2653 2022 2657 se
rect 2022 2653 8093 2657
tri 2017 2652 2018 2653 se
rect 2018 2652 8093 2653
rect 863 2617 915 2623
rect 1734 2646 1786 2652
rect 1734 2582 1786 2594
rect 454 2552 1554 2558
rect 454 2518 582 2552
rect 616 2518 660 2552
rect 694 2518 738 2552
rect 772 2518 815 2552
rect 849 2518 892 2552
rect 926 2518 969 2552
rect 1003 2518 1046 2552
rect 1080 2518 1123 2552
rect 1157 2518 1200 2552
rect 1234 2518 1277 2552
rect 1311 2518 1354 2552
rect 1388 2518 1431 2552
rect 1465 2518 1508 2552
rect 1542 2518 1554 2552
rect 454 2512 1554 2518
rect 454 2507 563 2512
tri 563 2507 568 2512 nw
rect 454 2499 555 2507
tri 555 2499 563 2507 nw
rect 454 2465 521 2499
tri 521 2465 555 2499 nw
rect 454 2450 506 2465
tri 506 2450 521 2465 nw
rect 1334 2439 1386 2442
rect 454 2370 506 2398
rect 558 2436 1552 2439
rect 558 2433 1334 2436
rect 1386 2433 1552 2436
rect 558 2399 570 2433
rect 604 2399 642 2433
rect 676 2399 714 2433
rect 748 2399 786 2433
rect 820 2399 858 2433
rect 892 2399 930 2433
rect 964 2399 1002 2433
rect 1036 2399 1074 2433
rect 1108 2399 1146 2433
rect 1180 2399 1218 2433
rect 1252 2399 1290 2433
rect 1324 2399 1334 2433
rect 1396 2399 1434 2433
rect 1468 2399 1506 2433
rect 1540 2399 1552 2433
rect 558 2393 1334 2399
rect 454 2297 506 2318
rect 1386 2393 1552 2399
rect 1334 2372 1386 2384
rect 1616 2380 1662 2392
rect 1334 2314 1386 2320
rect 1487 2358 1539 2364
tri 1483 2314 1487 2318 se
tri 1477 2308 1483 2314 se
rect 1483 2308 1487 2314
rect 454 2290 466 2297
rect 500 2290 506 2297
tri 1452 2283 1477 2308 se
rect 1477 2306 1487 2308
rect 1616 2346 1622 2380
rect 1656 2346 1662 2380
tri 1539 2308 1549 2318 sw
rect 1616 2308 1662 2346
rect 1539 2306 1549 2308
rect 1477 2294 1549 2306
rect 1477 2283 1487 2294
rect 454 2225 506 2238
rect 558 2277 1487 2283
rect 1539 2283 1549 2294
tri 1549 2283 1574 2308 sw
rect 1539 2281 1574 2283
tri 1574 2281 1576 2283 sw
rect 1539 2277 1576 2281
rect 558 2243 570 2277
rect 604 2243 642 2277
rect 676 2243 714 2277
rect 748 2243 786 2277
rect 820 2243 858 2277
rect 892 2243 930 2277
rect 964 2243 1002 2277
rect 1036 2243 1074 2277
rect 1108 2243 1146 2277
rect 1180 2243 1218 2277
rect 1252 2243 1290 2277
rect 1324 2243 1362 2277
rect 1396 2243 1434 2277
rect 1468 2243 1487 2277
rect 1540 2244 1576 2277
rect 1540 2243 1568 2244
rect 558 2242 1487 2243
rect 1539 2242 1568 2243
rect 558 2237 1568 2242
tri 1452 2236 1453 2237 ne
rect 1453 2236 1568 2237
tri 1568 2236 1576 2244 nw
rect 1616 2274 1622 2308
rect 1656 2280 1662 2308
tri 1662 2280 1668 2286 sw
rect 1656 2274 1668 2280
tri 1453 2234 1455 2236 ne
rect 1455 2234 1566 2236
tri 1566 2234 1568 2236 nw
rect 454 2210 466 2225
rect 500 2222 506 2225
tri 506 2222 509 2225 sw
rect 500 2210 509 2222
rect 506 2197 509 2210
tri 509 2197 534 2222 sw
rect 1616 2210 1668 2222
rect 506 2185 534 2197
tri 534 2185 546 2197 sw
rect 506 2182 546 2185
tri 546 2182 549 2185 sw
rect 506 2169 549 2182
tri 549 2169 562 2182 sw
rect 506 2162 1574 2169
rect 506 2158 574 2162
rect 454 2153 574 2158
rect 454 2130 466 2153
rect 500 2130 574 2153
rect 506 2128 574 2130
rect 608 2128 648 2162
rect 682 2128 722 2162
rect 756 2128 796 2162
rect 830 2128 870 2162
rect 904 2128 944 2162
rect 978 2128 1017 2162
rect 1051 2128 1090 2162
rect 1124 2128 1163 2162
rect 1197 2128 1236 2162
rect 1270 2128 1309 2162
rect 1343 2128 1382 2162
rect 1416 2128 1455 2162
rect 1489 2128 1528 2162
rect 1562 2128 1574 2162
rect 1616 2152 1668 2158
tri 1730 2152 1734 2156 se
rect 1734 2152 1786 2530
tri 1726 2148 1730 2152 se
rect 1730 2148 1786 2152
tri 1717 2139 1726 2148 se
rect 1726 2139 1786 2148
tri 1715 2137 1717 2139 se
rect 1717 2137 1786 2139
rect 506 2078 1574 2128
tri 1700 2122 1715 2137 se
rect 1715 2122 1786 2137
rect 454 2050 466 2078
rect 500 2062 1574 2078
rect 1658 2070 1664 2122
rect 1716 2070 1728 2122
rect 1780 2070 1786 2122
rect 500 2050 574 2062
rect 506 2028 574 2050
rect 608 2028 648 2062
rect 682 2028 722 2062
rect 756 2028 796 2062
rect 830 2028 870 2062
rect 904 2028 944 2062
rect 978 2028 1017 2062
rect 1051 2028 1090 2062
rect 1124 2028 1163 2062
rect 1197 2028 1236 2062
rect 1270 2028 1309 2062
rect 1343 2028 1382 2062
rect 1416 2028 1455 2062
rect 1489 2028 1528 2062
rect 1562 2028 1574 2062
tri 1700 2048 1722 2070 ne
rect 1722 2048 1786 2070
tri 1722 2043 1727 2048 ne
rect 1727 2043 1786 2048
tri 1727 2036 1734 2043 ne
rect 506 1998 1574 2028
rect 454 1975 466 1998
rect 500 1975 1574 1998
rect 454 1970 1574 1975
rect 506 1962 1574 1970
rect 506 1928 574 1962
rect 608 1928 648 1962
rect 682 1928 722 1962
rect 756 1928 796 1962
rect 830 1928 870 1962
rect 904 1928 944 1962
rect 978 1928 1017 1962
rect 1051 1928 1090 1962
rect 1124 1928 1163 1962
rect 1197 1928 1236 1962
rect 1270 1928 1309 1962
rect 1343 1928 1382 1962
rect 1416 1928 1455 1962
rect 1489 1928 1528 1962
rect 1562 1928 1574 1962
rect 506 1921 1574 1928
rect 506 1918 542 1921
rect 454 1903 466 1918
rect 500 1903 542 1918
rect 454 1901 542 1903
tri 542 1901 562 1921 nw
rect 454 1890 527 1901
rect 506 1886 527 1890
tri 527 1886 542 1901 nw
tri 506 1865 527 1886 nw
tri 1274 1847 1277 1850 se
rect 1277 1847 1283 1850
rect 454 1831 466 1838
rect 500 1831 506 1838
rect 454 1810 506 1831
rect 558 1841 1283 1847
rect 558 1807 570 1841
rect 604 1807 642 1841
rect 676 1807 714 1841
rect 748 1807 786 1841
rect 820 1807 858 1841
rect 892 1807 930 1841
rect 964 1807 1002 1841
rect 1036 1807 1074 1841
rect 1108 1807 1146 1841
rect 1180 1807 1218 1841
rect 1252 1807 1283 1841
rect 558 1801 1283 1807
tri 1274 1798 1277 1801 ne
rect 1277 1798 1283 1801
rect 1335 1798 1347 1850
rect 1399 1847 1405 1850
tri 1405 1847 1408 1850 sw
rect 1399 1841 1552 1847
rect 1399 1807 1434 1841
rect 1468 1807 1506 1841
rect 1540 1807 1552 1841
rect 1399 1801 1552 1807
rect 1399 1798 1405 1801
tri 1405 1798 1408 1801 nw
rect 454 1730 506 1758
rect 1102 1721 1108 1773
rect 1160 1721 1174 1773
rect 1226 1721 1232 1773
rect 1610 1729 1662 1735
tri 1606 1721 1610 1725 se
tri 1589 1704 1606 1721 se
rect 1606 1704 1610 1721
tri 1582 1697 1589 1704 se
rect 1589 1697 1610 1704
tri 1576 1691 1582 1697 se
rect 1582 1691 1610 1697
rect 454 1650 506 1678
rect 558 1685 1610 1691
rect 558 1651 570 1685
rect 604 1651 642 1685
rect 676 1651 714 1685
rect 748 1651 786 1685
rect 820 1651 858 1685
rect 892 1651 930 1685
rect 964 1651 1002 1685
rect 1036 1651 1074 1685
rect 1108 1651 1146 1685
rect 1180 1651 1218 1685
rect 1252 1651 1290 1685
rect 1324 1651 1362 1685
rect 1396 1651 1434 1685
rect 1468 1651 1506 1685
rect 1540 1677 1610 1685
rect 1540 1665 1662 1677
rect 1540 1651 1610 1665
rect 558 1645 1610 1651
tri 1576 1630 1591 1645 ne
rect 1591 1630 1610 1645
tri 1591 1619 1602 1630 ne
rect 1602 1619 1610 1630
tri 1602 1615 1606 1619 ne
rect 1606 1615 1610 1619
rect 454 1577 506 1598
rect 454 1570 466 1577
rect 500 1570 506 1577
rect 1102 1563 1108 1615
rect 1160 1563 1174 1615
rect 1226 1563 1232 1615
tri 1606 1611 1610 1615 ne
rect 1610 1607 1662 1613
tri 1274 1535 1277 1538 se
rect 1277 1535 1283 1538
rect 454 1505 506 1518
rect 454 1490 466 1505
rect 500 1490 506 1505
rect 558 1529 1283 1535
rect 558 1495 570 1529
rect 604 1495 642 1529
rect 676 1495 714 1529
rect 748 1495 786 1529
rect 820 1495 858 1529
rect 892 1495 930 1529
rect 964 1495 1002 1529
rect 1036 1495 1074 1529
rect 1108 1495 1146 1529
rect 1180 1495 1218 1529
rect 1252 1495 1283 1529
rect 558 1489 1283 1495
tri 1274 1486 1277 1489 ne
rect 1277 1486 1283 1489
rect 1335 1486 1347 1538
rect 1399 1535 1405 1538
tri 1405 1535 1408 1538 sw
rect 1399 1529 1552 1535
rect 1399 1495 1434 1529
rect 1468 1495 1506 1529
rect 1540 1495 1552 1529
rect 1399 1489 1552 1495
rect 1399 1486 1405 1489
tri 1405 1486 1408 1489 nw
rect 454 1433 506 1438
rect 454 1410 466 1433
rect 500 1410 506 1433
rect 1734 1456 1786 2043
tri 506 1408 530 1432 sw
rect 506 1407 530 1408
tri 530 1407 531 1408 sw
rect 506 1401 1574 1407
rect 506 1367 597 1401
rect 631 1367 675 1401
rect 709 1367 753 1401
rect 787 1367 831 1401
rect 865 1367 909 1401
rect 943 1367 987 1401
rect 1021 1367 1065 1401
rect 1099 1367 1143 1401
rect 1177 1367 1220 1401
rect 1254 1367 1297 1401
rect 1331 1367 1374 1401
rect 1408 1367 1451 1401
rect 1485 1367 1528 1401
rect 1562 1367 1574 1401
rect 506 1361 1574 1367
rect 1734 1377 1786 1404
rect 454 1330 466 1358
rect 500 1330 506 1358
tri 506 1336 531 1361 nw
rect 1734 1319 1786 1325
rect 1821 2646 1873 2652
rect 1821 2582 1873 2594
rect 1821 2274 1873 2530
rect 1821 2210 1873 2222
tri 1810 1294 1821 1305 se
rect 1821 1294 1873 2158
tri 1807 1291 1810 1294 se
rect 1810 1291 1873 1294
tri 1250 1285 1256 1291 se
rect 1256 1285 1262 1291
rect 454 1255 466 1278
rect 500 1255 506 1278
rect 454 1250 506 1255
rect 558 1279 1262 1285
rect 1314 1279 1326 1291
rect 1378 1285 1384 1291
tri 1384 1285 1390 1291 sw
tri 1801 1285 1807 1291 se
rect 1807 1285 1873 1291
rect 1378 1279 1552 1285
rect 558 1245 570 1279
rect 604 1245 642 1279
rect 676 1245 714 1279
rect 748 1245 786 1279
rect 820 1245 858 1279
rect 892 1245 930 1279
rect 964 1245 1002 1279
rect 1036 1245 1074 1279
rect 1108 1245 1146 1279
rect 1180 1245 1218 1279
rect 1252 1245 1262 1279
rect 1324 1245 1326 1279
rect 1396 1245 1434 1279
rect 1468 1245 1506 1279
rect 1540 1245 1552 1279
tri 1781 1265 1801 1285 se
rect 1801 1282 1873 1285
rect 1801 1265 1856 1282
tri 1856 1265 1873 1282 nw
rect 1901 2646 1953 2652
tri 2003 2638 2017 2652 se
rect 2017 2638 8093 2652
tri 1995 2630 2003 2638 se
rect 2003 2630 8093 2638
rect 1901 2582 1953 2594
rect 1901 1729 1953 2530
rect 1901 1660 1953 1677
rect 1901 1591 1953 1608
rect 1901 1522 1953 1539
rect 1901 1452 1953 1470
tri 1776 1260 1781 1265 se
rect 1781 1260 1851 1265
tri 1851 1260 1856 1265 nw
tri 1896 1260 1901 1265 se
rect 1901 1260 1953 1400
rect 558 1239 1262 1245
rect 1314 1239 1326 1245
rect 1378 1239 1552 1245
tri 1755 1239 1776 1260 se
rect 1776 1239 1835 1260
tri 1835 1244 1851 1260 nw
tri 1880 1244 1896 1260 se
rect 1896 1253 1953 1260
rect 1896 1244 1939 1253
tri 1875 1239 1880 1244 se
rect 1880 1239 1939 1244
tri 1939 1239 1953 1253 nw
tri 1983 2618 1995 2630 se
rect 1995 2618 8093 2630
rect 1983 2613 8093 2618
rect 8145 2613 8157 2665
rect 8209 2613 8215 2665
rect 1983 2585 2041 2613
tri 2041 2585 2069 2613 nw
tri 8322 2585 8348 2611 se
rect 8348 2585 8400 2613
rect 1983 2584 2040 2585
tri 2040 2584 2041 2585 nw
tri 2110 2584 2111 2585 se
rect 2111 2584 6269 2585
rect 1983 2582 2038 2584
tri 2038 2582 2040 2584 nw
tri 2108 2582 2110 2584 se
rect 2110 2582 6269 2584
tri 1736 1220 1755 1239 se
rect 1755 1220 1835 1239
tri 1732 1216 1736 1220 se
rect 1736 1216 1835 1220
rect 454 1183 466 1198
rect 500 1183 506 1198
rect 454 1170 506 1183
rect 1616 1204 1835 1216
rect 781 1167 833 1173
tri 777 1159 781 1163 se
tri 764 1146 777 1159 se
rect 777 1146 781 1159
tri 747 1129 764 1146 se
rect 764 1129 781 1146
rect 454 1111 466 1118
rect 500 1111 506 1118
rect 454 1090 506 1111
rect 558 1123 781 1129
rect 1616 1170 1622 1204
rect 1656 1170 1835 1204
tri 833 1159 837 1163 sw
rect 833 1146 837 1159
tri 837 1146 850 1159 sw
rect 833 1129 850 1146
tri 850 1129 867 1146 sw
rect 833 1123 1552 1129
rect 558 1089 570 1123
rect 604 1089 642 1123
rect 676 1089 714 1123
rect 748 1115 781 1123
rect 833 1115 858 1123
rect 748 1097 786 1115
rect 820 1097 858 1115
rect 748 1089 781 1097
rect 833 1089 858 1097
rect 892 1089 930 1123
rect 964 1089 1002 1123
rect 1036 1089 1074 1123
rect 1108 1089 1146 1123
rect 1180 1089 1218 1123
rect 1252 1089 1290 1123
rect 1324 1089 1362 1123
rect 1396 1089 1434 1123
rect 1468 1089 1506 1123
rect 1540 1089 1552 1123
rect 558 1083 781 1089
tri 747 1072 758 1083 ne
rect 758 1072 781 1083
tri 758 1049 781 1072 ne
rect 833 1083 1552 1089
rect 1616 1119 1835 1170
rect 1616 1085 1622 1119
rect 1656 1085 1835 1119
rect 833 1072 856 1083
tri 856 1072 867 1083 nw
tri 833 1049 856 1072 nw
rect 781 1039 833 1045
rect 454 1010 506 1038
rect 1616 1033 1835 1085
rect 1616 999 1622 1033
rect 1656 999 1835 1033
tri 1253 973 1256 976 se
rect 1256 973 1262 976
rect 454 930 506 958
rect 558 967 1262 973
rect 1314 967 1326 976
rect 1378 973 1384 976
tri 1384 973 1387 976 sw
rect 1378 967 1552 973
rect 558 933 570 967
rect 604 933 642 967
rect 676 933 714 967
rect 748 933 786 967
rect 820 933 858 967
rect 892 933 930 967
rect 964 933 1002 967
rect 1036 933 1074 967
rect 1108 933 1146 967
rect 1180 933 1218 967
rect 1252 933 1262 967
rect 1324 933 1326 967
rect 1396 933 1434 967
rect 1468 933 1506 967
rect 1540 933 1552 967
rect 1616 966 1835 999
tri 1762 964 1764 966 ne
rect 1764 964 1835 966
tri 1764 948 1780 964 ne
rect 1780 948 1835 964
tri 506 924 511 929 sw
rect 558 927 1262 933
tri 1253 924 1256 927 ne
rect 1256 924 1262 927
rect 1314 924 1326 933
rect 1378 927 1552 933
tri 1780 931 1797 948 ne
rect 1378 924 1384 927
tri 1384 924 1387 927 nw
rect 506 895 511 924
tri 511 895 540 924 sw
rect 506 889 1545 895
rect 506 878 1427 889
rect 454 857 1427 878
rect 454 850 466 857
rect 500 855 1427 857
rect 1461 855 1499 889
rect 1533 855 1545 889
rect 500 850 1545 855
rect 506 849 1545 850
rect 506 817 508 849
tri 508 817 540 849 nw
rect 506 816 507 817
tri 507 816 508 817 nw
tri 506 815 507 816 nw
rect 454 785 506 798
rect 454 770 466 785
rect 500 770 506 785
rect 558 811 1552 817
rect 558 777 570 811
rect 604 777 642 811
rect 676 777 714 811
rect 748 777 786 811
rect 820 777 858 811
rect 892 777 930 811
rect 964 777 1002 811
rect 1036 777 1074 811
rect 1108 777 1146 811
rect 1252 777 1290 811
rect 1324 777 1362 811
rect 1396 777 1434 811
rect 1468 777 1506 811
rect 1540 777 1552 811
tri 1780 779 1797 796 se
rect 1797 779 1835 948
rect 558 771 1174 777
tri 1140 742 1169 771 ne
rect 1169 759 1174 771
rect 1226 771 1552 777
tri 1777 776 1780 779 se
rect 1780 776 1835 779
tri 1772 771 1777 776 se
rect 1777 771 1835 776
rect 1226 759 1237 771
rect 1169 748 1237 759
tri 1237 748 1260 771 nw
tri 1749 748 1772 771 se
rect 1772 748 1835 771
rect 1169 747 1231 748
rect 1169 742 1174 747
tri 1169 737 1174 742 ne
rect 454 713 506 718
rect 454 690 466 713
rect 500 690 506 713
rect 699 699 751 705
tri 672 668 699 695 se
tri 665 661 672 668 se
rect 672 661 699 668
rect 454 610 466 638
rect 500 610 506 638
rect 558 655 699 661
rect 1226 742 1231 747
tri 1231 742 1237 748 nw
tri 1226 737 1231 742 nw
tri 751 689 757 695 sw
rect 1174 689 1226 695
rect 1616 736 1835 748
rect 1616 702 1622 736
rect 1656 702 1835 736
rect 751 668 757 689
tri 757 668 778 689 sw
rect 751 661 778 668
tri 778 661 785 668 sw
rect 751 655 1552 661
rect 558 621 570 655
rect 604 621 642 655
rect 676 647 699 655
rect 751 647 786 655
rect 676 629 714 647
rect 748 629 786 647
rect 676 621 699 629
rect 751 621 786 629
rect 820 621 858 655
rect 892 621 930 655
rect 964 621 1002 655
rect 1036 621 1074 655
rect 1108 621 1146 655
rect 1180 621 1218 655
rect 1252 621 1290 655
rect 1324 621 1362 655
rect 1396 621 1434 655
rect 1468 621 1506 655
rect 1540 621 1552 655
rect 558 615 699 621
tri 665 606 674 615 ne
rect 674 606 699 615
tri 674 594 686 606 ne
rect 686 594 699 606
tri 686 588 692 594 ne
rect 692 588 699 594
tri 692 581 699 588 ne
rect 751 615 1552 621
rect 1616 640 1835 702
rect 751 606 776 615
tri 776 606 785 615 nw
rect 1616 606 1622 640
rect 1656 606 1835 640
rect 751 594 764 606
tri 764 594 776 606 nw
rect 751 588 758 594
tri 758 588 764 594 nw
rect 751 587 757 588
tri 757 587 758 588 nw
tri 751 581 757 587 nw
rect 1174 581 1226 587
rect 699 571 751 577
rect 454 535 466 558
rect 500 535 506 558
rect 454 530 506 535
tri 1145 510 1174 539 se
rect 1616 544 1835 606
rect 1174 517 1226 529
tri 1140 505 1145 510 se
rect 1145 505 1174 510
rect 454 463 466 478
rect 500 463 506 478
rect 454 459 506 463
rect 558 499 1174 505
tri 1226 510 1255 539 sw
rect 1616 510 1622 544
rect 1656 510 1835 544
rect 1226 505 1255 510
tri 1255 505 1260 510 sw
rect 1226 499 1552 505
rect 558 465 570 499
rect 604 465 642 499
rect 676 465 714 499
rect 748 465 786 499
rect 820 465 858 499
rect 892 465 930 499
rect 964 465 1002 499
rect 1036 465 1074 499
rect 1108 465 1146 499
rect 1252 465 1290 499
rect 1324 465 1362 499
rect 1396 465 1434 499
rect 1468 465 1506 499
rect 1540 465 1552 499
rect 1616 498 1835 510
tri 1752 491 1759 498 ne
rect 1759 491 1835 498
tri 1759 484 1766 491 ne
rect 1766 484 1835 491
tri 1766 482 1768 484 ne
rect 1768 482 1835 484
tri 1768 480 1770 482 ne
rect 1770 480 1835 482
tri 1770 466 1784 480 ne
tri 506 459 508 461 sw
rect 558 459 1552 465
rect 454 450 508 459
rect 506 446 508 450
tri 508 446 521 459 sw
rect 506 444 521 446
tri 521 444 523 446 sw
rect 506 427 523 444
tri 523 427 540 444 sw
rect 506 421 1545 427
rect 506 398 1427 421
rect 454 391 466 398
rect 500 391 1427 398
rect 454 387 1427 391
rect 1461 387 1499 421
rect 1533 387 1545 421
rect 454 381 1545 387
rect 454 372 531 381
tri 531 372 540 381 nw
rect 454 370 511 372
rect 506 352 511 370
tri 511 352 531 372 nw
tri 506 347 511 352 nw
tri 698 349 701 352 se
rect 701 349 707 352
rect 454 290 506 318
rect 558 343 707 349
rect 558 309 570 343
rect 604 309 642 343
rect 676 309 707 343
rect 558 303 707 309
tri 698 300 701 303 ne
rect 701 300 707 303
rect 759 300 771 352
rect 823 349 829 352
tri 829 349 832 352 sw
rect 823 343 1552 349
rect 823 309 858 343
rect 892 309 930 343
rect 964 309 1002 343
rect 1036 309 1074 343
rect 1108 309 1146 343
rect 1180 309 1218 343
rect 1252 309 1290 343
rect 1324 309 1362 343
rect 1396 309 1434 343
rect 1468 309 1506 343
rect 1540 309 1552 343
rect 823 303 1552 309
tri 1761 303 1784 326 se
rect 1784 303 1835 480
rect 823 300 829 303
tri 829 300 832 303 nw
tri 1758 300 1761 303 se
rect 1761 300 1835 303
tri 1756 298 1758 300 se
rect 1758 298 1835 300
tri 1738 280 1756 298 se
rect 1756 280 1835 298
rect 454 210 506 238
rect 1616 268 1835 280
rect 617 230 669 236
tri 614 224 617 227 se
tri 593 203 614 224 se
rect 614 203 617 224
tri 583 193 593 203 se
rect 593 193 617 203
rect 454 137 506 158
rect 558 187 617 193
rect 1616 234 1622 268
rect 1656 234 1835 268
tri 669 224 672 227 sw
rect 669 203 672 224
tri 672 203 693 224 sw
rect 669 193 693 203
tri 693 193 703 203 sw
rect 669 187 1552 193
rect 558 153 570 187
rect 604 178 617 187
rect 604 160 642 178
rect 604 153 617 160
rect 676 153 714 187
rect 748 153 786 187
rect 820 153 858 187
rect 892 153 930 187
rect 964 153 1002 187
rect 1036 153 1074 187
rect 1108 153 1146 187
rect 1180 153 1218 187
rect 1252 153 1290 187
rect 1324 153 1362 187
rect 1396 153 1434 187
rect 1468 153 1506 187
rect 1540 153 1552 187
rect 558 147 617 153
tri 583 138 592 147 ne
rect 592 138 617 147
rect 454 130 466 137
rect 500 130 506 137
tri 592 131 599 138 ne
rect 599 131 617 138
tri 599 118 612 131 ne
rect 612 118 617 131
tri 612 113 617 118 ne
rect 669 147 1552 153
rect 1616 172 1835 234
rect 669 138 694 147
tri 694 138 703 147 nw
rect 1616 138 1622 172
rect 1656 138 1835 172
rect 669 131 687 138
tri 687 131 694 138 nw
rect 669 118 674 131
tri 674 118 687 131 nw
tri 669 113 674 118 nw
rect 617 102 669 108
rect 454 65 506 78
rect 454 50 466 65
rect 500 50 506 65
rect 1616 76 1835 138
rect 1616 42 1622 76
rect 1656 42 1835 76
tri 698 37 701 40 se
rect 701 37 707 40
rect 454 -7 506 -2
rect 558 31 707 37
rect 558 -3 570 31
rect 604 -3 642 31
rect 676 -3 707 31
rect 454 -30 466 -7
rect 500 -12 506 -7
tri 506 -12 511 -7 sw
rect 558 -9 707 -3
tri 698 -12 701 -9 ne
rect 701 -12 707 -9
rect 759 -12 771 40
rect 823 37 829 40
tri 829 37 832 40 sw
rect 823 31 1552 37
rect 823 -3 858 31
rect 892 -3 930 31
rect 964 -3 1002 31
rect 1036 -3 1074 31
rect 1108 -3 1146 31
rect 1180 -3 1218 31
rect 1252 -3 1290 31
rect 1324 -3 1362 31
rect 1396 -3 1434 31
rect 1468 -3 1506 31
rect 1540 -3 1552 31
rect 1616 30 1835 42
tri 1748 2 1776 30 ne
rect 1776 2 1835 30
rect 823 -9 1552 -3
tri 1776 -6 1784 2 ne
rect 823 -12 829 -9
tri 829 -12 832 -9 nw
rect 500 -13 511 -12
tri 511 -13 512 -12 sw
rect 500 -30 512 -13
rect 506 -38 512 -30
tri 512 -38 537 -13 sw
rect 506 -41 537 -38
tri 537 -41 540 -38 sw
rect 506 -47 1545 -41
rect 506 -81 1427 -47
rect 1461 -81 1499 -47
rect 1533 -81 1545 -47
rect 506 -82 1545 -81
rect 454 -110 466 -82
rect 500 -87 1545 -82
rect 500 -92 535 -87
tri 535 -92 540 -87 nw
rect 500 -103 524 -92
tri 524 -103 535 -92 nw
rect 500 -107 520 -103
tri 520 -107 524 -103 nw
rect 500 -110 515 -107
rect 506 -112 515 -110
tri 515 -112 520 -107 nw
rect 506 -119 508 -112
tri 508 -119 515 -112 nw
tri 506 -121 508 -119 nw
rect 454 -185 466 -162
rect 500 -185 506 -162
rect 558 -125 1552 -119
rect 558 -159 570 -125
rect 604 -159 642 -125
rect 676 -159 693 -125
rect 748 -159 786 -125
rect 820 -159 858 -125
rect 892 -159 930 -125
rect 964 -159 1002 -125
rect 1036 -159 1074 -125
rect 1108 -159 1146 -125
rect 1180 -159 1218 -125
rect 1252 -159 1290 -125
rect 1324 -159 1362 -125
rect 1396 -159 1434 -125
rect 1468 -159 1506 -125
rect 1540 -159 1552 -125
rect 558 -165 693 -159
tri 658 -176 669 -165 ne
rect 669 -176 693 -165
tri 669 -179 672 -176 ne
rect 672 -177 693 -176
rect 745 -165 1552 -159
tri 1772 -165 1784 -153 se
rect 1784 -165 1835 2
rect 745 -176 768 -165
tri 768 -176 779 -165 nw
tri 1761 -176 1772 -165 se
rect 1772 -176 1835 -165
rect 745 -177 765 -176
rect 672 -179 765 -177
tri 765 -179 768 -176 nw
tri 1758 -179 1761 -176 se
rect 1761 -179 1835 -176
rect 454 -190 506 -185
tri 672 -186 679 -179 ne
rect 679 -186 758 -179
tri 758 -186 765 -179 nw
tri 1751 -186 1758 -179 se
rect 1758 -186 1835 -179
tri 679 -200 693 -186 ne
rect 693 -188 756 -186
tri 756 -188 758 -186 nw
tri 1749 -188 1751 -186 se
rect 1751 -188 1835 -186
rect 693 -189 745 -188
rect 454 -257 466 -242
rect 500 -257 506 -242
rect 454 -270 506 -257
rect 454 -329 466 -322
rect 500 -329 506 -322
rect 454 -350 506 -329
rect 535 -237 587 -231
tri 745 -199 756 -188 nw
tri 587 -247 593 -241 sw
rect 693 -247 745 -241
rect 1616 -200 1835 -188
rect 1616 -234 1622 -200
rect 1656 -234 1835 -200
rect 587 -249 593 -247
tri 593 -249 595 -247 sw
rect 587 -251 595 -249
tri 595 -251 597 -249 sw
rect 587 -260 597 -251
tri 597 -260 606 -251 sw
rect 587 -275 606 -260
tri 606 -275 621 -260 sw
rect 587 -281 1552 -275
rect 535 -307 570 -289
rect 604 -315 642 -281
rect 676 -315 714 -281
rect 748 -315 786 -281
rect 820 -315 858 -281
rect 892 -315 930 -281
rect 964 -315 1002 -281
rect 1036 -315 1074 -281
rect 1108 -315 1146 -281
rect 1180 -315 1218 -281
rect 1252 -315 1290 -281
rect 1324 -315 1362 -281
rect 1396 -315 1434 -281
rect 1468 -315 1506 -281
rect 1540 -315 1552 -281
rect 587 -321 1552 -315
rect 1616 -285 1835 -234
rect 1616 -319 1622 -285
rect 1656 -319 1835 -285
rect 587 -322 620 -321
tri 620 -322 621 -321 nw
rect 587 -323 619 -322
tri 619 -323 620 -322 nw
rect 587 -332 610 -323
tri 610 -332 619 -323 nw
rect 587 -352 590 -332
tri 590 -352 610 -332 nw
tri 587 -355 590 -352 nw
rect 535 -365 587 -359
rect 687 -358 751 -352
rect 454 -430 506 -402
tri 682 -405 687 -400 se
rect 687 -405 693 -358
tri 674 -413 682 -405 se
rect 682 -410 693 -405
rect 745 -405 751 -358
rect 1616 -371 1835 -319
tri 751 -405 759 -397 sw
rect 1616 -405 1622 -371
rect 1656 -405 1835 -371
tri 1866 1230 1875 1239 se
rect 1875 1230 1930 1239
tri 1930 1230 1939 1239 nw
rect 1866 1220 1920 1230
tri 1920 1220 1930 1230 nw
tri 1982 1220 1983 1221 se
rect 1983 1220 2035 2582
tri 2035 2579 2038 2582 nw
tri 2105 2579 2108 2582 se
rect 2108 2579 6269 2582
tri 2083 2557 2105 2579 se
rect 2105 2557 6269 2579
rect 1866 212 1918 1220
tri 1918 1218 1920 1220 nw
tri 1980 1218 1982 1220 se
rect 1982 1218 2035 1220
rect 1866 144 1918 160
rect 1866 76 1918 92
tri 1950 1188 1980 1218 se
rect 1980 1199 2035 1218
rect 1980 1188 2024 1199
tri 2024 1188 2035 1199 nw
tri 2065 2539 2083 2557 se
rect 2083 2539 6269 2557
rect 2065 2533 6269 2539
rect 6321 2533 6349 2585
rect 6401 2533 6407 2585
rect 6449 2533 6455 2585
rect 6507 2533 6519 2585
rect 6571 2533 7303 2585
rect 7355 2533 7367 2585
rect 7419 2533 7427 2585
rect 7658 2533 7664 2585
rect 7716 2533 7728 2585
rect 7780 2538 8400 2585
rect 7780 2533 8074 2538
tri 8074 2533 8079 2538 nw
tri 8244 2533 8249 2538 ne
rect 8249 2533 8400 2538
rect 8476 2840 8522 2880
rect 8476 2806 8482 2840
rect 8516 2806 8522 2840
rect 8476 2766 8522 2806
rect 8476 2732 8482 2766
rect 8516 2732 8522 2766
rect 8476 2691 8522 2732
rect 8476 2657 8482 2691
rect 8516 2657 8522 2691
rect 8476 2616 8522 2657
rect 8476 2582 8482 2616
rect 8516 2582 8522 2616
rect 2065 2531 2141 2533
tri 2141 2531 2143 2533 nw
rect 2065 2523 2133 2531
tri 2133 2523 2141 2531 nw
tri 8468 2523 8476 2531 se
rect 8476 2523 8522 2582
rect 2065 2508 2118 2523
tri 2118 2508 2133 2523 nw
tri 8453 2508 8468 2523 se
rect 8468 2508 8522 2523
rect 1950 1186 2022 1188
tri 2022 1186 2024 1188 nw
rect 1950 76 2002 1186
tri 2002 1166 2022 1186 nw
rect 2065 221 2117 2508
tri 2117 2507 2118 2508 nw
tri 8089 2507 8090 2508 se
rect 8090 2507 8096 2508
tri 8087 2505 8089 2507 se
rect 8089 2505 8096 2507
tri 2174 2499 2180 2505 se
rect 2180 2499 8096 2505
rect 2065 157 2117 169
rect 2065 99 2117 105
tri 2145 2470 2174 2499 se
rect 2174 2470 2245 2499
rect 2145 2465 2245 2470
rect 2279 2465 2323 2499
rect 2357 2465 2400 2499
rect 2434 2465 2510 2499
rect 2544 2465 2583 2499
rect 2617 2465 2656 2499
rect 2690 2465 2729 2499
rect 2763 2465 2802 2499
rect 2836 2465 2875 2499
rect 2909 2465 2948 2499
rect 2982 2465 3021 2499
rect 3055 2465 3094 2499
rect 3128 2465 3167 2499
rect 3201 2465 3240 2499
rect 3274 2465 3313 2499
rect 3347 2465 3386 2499
rect 3420 2465 3459 2499
rect 3493 2465 3532 2499
rect 3566 2465 3605 2499
rect 3639 2465 3678 2499
rect 3712 2465 3751 2499
rect 3785 2465 3824 2499
rect 3858 2465 3897 2499
rect 3931 2465 3970 2499
rect 4004 2465 4043 2499
rect 4077 2465 4116 2499
rect 4150 2465 4189 2499
rect 4223 2465 4262 2499
rect 4296 2465 4335 2499
rect 4369 2465 4408 2499
rect 4442 2465 4481 2499
rect 4515 2465 4554 2499
rect 4588 2465 4627 2499
rect 4661 2465 4700 2499
rect 4734 2465 4773 2499
rect 4807 2465 4846 2499
rect 4880 2465 4919 2499
rect 4953 2465 4992 2499
rect 5026 2465 5065 2499
rect 5099 2465 5138 2499
rect 5172 2465 5211 2499
rect 5245 2465 5284 2499
rect 5318 2465 5357 2499
rect 5391 2465 5430 2499
rect 5464 2465 5503 2499
rect 5537 2465 5576 2499
rect 5610 2465 5649 2499
rect 5683 2465 5722 2499
rect 5756 2465 5795 2499
rect 5829 2465 5868 2499
rect 5902 2465 5941 2499
rect 5975 2465 6014 2499
rect 6048 2465 6087 2499
rect 6121 2465 6160 2499
rect 6194 2465 6233 2499
rect 6267 2465 6306 2499
rect 6340 2465 6379 2499
rect 6413 2465 6452 2499
rect 6486 2465 6525 2499
rect 6559 2465 6598 2499
rect 6632 2465 6671 2499
rect 6705 2465 6744 2499
rect 6778 2465 6816 2499
rect 6850 2465 6888 2499
rect 6922 2465 6960 2499
rect 6994 2465 7032 2499
rect 7066 2465 7104 2499
rect 7138 2465 7176 2499
rect 7210 2465 7248 2499
rect 7282 2465 7320 2499
rect 7354 2465 7392 2499
rect 7426 2465 7464 2499
rect 7498 2465 7536 2499
rect 7570 2465 7608 2499
rect 7642 2465 7680 2499
rect 7714 2465 7752 2499
rect 7786 2465 7824 2499
rect 7858 2465 7896 2499
rect 7930 2465 7968 2499
rect 8002 2465 8040 2499
rect 8074 2465 8096 2499
rect 2145 2459 8096 2465
rect 2145 2456 2221 2459
tri 2221 2456 2224 2459 nw
tri 8087 2456 8090 2459 ne
rect 8090 2456 8096 2459
rect 8148 2456 8160 2508
rect 8212 2507 8218 2508
tri 8218 2507 8219 2508 sw
tri 8452 2507 8453 2508 se
rect 8453 2507 8522 2508
rect 8212 2505 8219 2507
tri 8219 2505 8221 2507 sw
tri 8450 2505 8452 2507 se
rect 8452 2505 8522 2507
rect 8212 2499 8522 2505
rect 8218 2465 8256 2499
rect 8290 2465 8328 2499
rect 8362 2465 8400 2499
rect 8434 2496 8522 2499
rect 8434 2484 8510 2496
tri 8510 2484 8522 2496 nw
tri 8551 3292 8562 3303 se
rect 8562 3292 8601 3303
tri 8601 3292 8612 3303 nw
tri 8646 3292 8657 3303 se
rect 8657 3293 8697 3303
tri 8697 3293 8707 3303 nw
tri 8746 3293 8756 3303 se
rect 8756 3293 8812 3303
tri 8812 3293 8822 3303 nw
rect 8657 3292 8691 3293
rect 8551 3281 8590 3292
tri 8590 3281 8601 3292 nw
tri 8641 3287 8646 3292 se
rect 8646 3287 8691 3292
tri 8691 3287 8697 3293 nw
tri 8740 3287 8746 3293 se
rect 8746 3287 8800 3293
tri 8635 3281 8641 3287 se
rect 8641 3281 8685 3287
tri 8685 3281 8691 3287 nw
tri 8734 3281 8740 3287 se
rect 8740 3281 8800 3287
tri 8800 3281 8812 3293 nw
rect 8434 2465 8485 2484
rect 8212 2459 8485 2465
tri 8485 2459 8510 2484 nw
rect 8212 2456 8218 2459
tri 8218 2456 8221 2459 nw
rect 2145 2453 2218 2456
tri 2218 2453 2221 2456 nw
rect 2145 2450 2215 2453
tri 2215 2450 2218 2453 nw
tri 8548 2450 8551 2453 se
rect 8551 2450 8587 3281
tri 8587 3278 8590 3281 nw
tri 8632 3278 8635 3281 se
rect 8635 3278 8679 3281
tri 8629 3275 8632 3278 se
rect 8632 3275 8679 3278
tri 8679 3275 8685 3281 nw
tri 8728 3275 8734 3281 se
rect 8734 3275 8794 3281
tri 8794 3275 8800 3281 nw
tri 8619 3265 8629 3275 se
rect 8629 3265 8669 3275
tri 8669 3265 8679 3275 nw
tri 8718 3265 8728 3275 se
rect 8728 3265 8784 3275
tri 8784 3265 8794 3275 nw
rect 2145 2440 2205 2450
tri 2205 2440 2215 2450 nw
tri 8538 2440 8548 2450 se
rect 8548 2440 8587 2450
rect 2145 2435 2200 2440
tri 2200 2435 2205 2440 nw
tri 8533 2435 8538 2440 se
rect 8538 2435 8587 2440
rect 2145 2428 2193 2435
tri 2193 2428 2200 2435 nw
tri 8526 2428 8533 2435 se
rect 8533 2431 8587 2435
rect 8533 2428 8584 2431
tri 8584 2428 8587 2431 nw
tri 8618 3264 8619 3265 se
rect 8619 3264 8668 3265
tri 8668 3264 8669 3265 nw
tri 8717 3264 8718 3265 se
rect 8718 3264 8781 3265
rect 8618 3254 8658 3264
tri 8658 3254 8668 3264 nw
tri 8715 3262 8717 3264 se
rect 8717 3262 8781 3264
tri 8781 3262 8784 3265 nw
rect 8715 3254 8773 3262
tri 8773 3254 8781 3262 nw
rect 9935 3254 9981 3321
rect 2145 2402 2191 2428
tri 2191 2426 2193 2428 nw
tri 2256 2426 2258 2428 se
rect 2258 2426 8567 2428
tri 2252 2422 2256 2426 se
rect 2256 2422 8567 2426
tri 2241 2411 2252 2422 se
rect 2252 2411 8567 2422
tri 8567 2411 8584 2428 nw
rect 2145 2368 2151 2402
rect 2185 2368 2191 2402
rect 2145 2329 2191 2368
rect 2145 2295 2151 2329
rect 2185 2295 2191 2329
rect 2145 2256 2191 2295
rect 2145 2222 2151 2256
rect 2185 2222 2191 2256
rect 2145 2182 2191 2222
rect 2145 2148 2151 2182
rect 2185 2148 2191 2182
rect 2145 2108 2191 2148
rect 2145 2074 2151 2108
rect 2185 2074 2191 2108
rect 2145 2034 2191 2074
rect 2145 2000 2151 2034
rect 2185 2000 2191 2034
rect 2145 1960 2191 2000
rect 2145 1926 2151 1960
rect 2185 1926 2191 1960
rect 2145 1886 2191 1926
rect 2145 1852 2151 1886
rect 2185 1852 2191 1886
rect 2145 1812 2191 1852
rect 2145 1778 2151 1812
rect 2185 1778 2191 1812
rect 2145 1738 2191 1778
rect 2145 1704 2151 1738
rect 2185 1704 2191 1738
rect 2145 1664 2191 1704
rect 2145 1630 2151 1664
rect 2185 1630 2191 1664
rect 2145 1590 2191 1630
rect 2145 1556 2151 1590
rect 2185 1556 2191 1590
rect 2145 1516 2191 1556
rect 2145 1482 2151 1516
rect 2185 1482 2191 1516
rect 2145 1442 2191 1482
rect 2145 1408 2151 1442
rect 2185 1408 2191 1442
rect 2145 1368 2191 1408
rect 2145 1334 2151 1368
rect 2185 1334 2191 1368
rect 2145 1294 2191 1334
rect 2145 1260 2151 1294
rect 2185 1260 2191 1294
rect 2145 1220 2191 1260
rect 2145 1186 2151 1220
rect 2185 1186 2191 1220
rect 2145 1146 2191 1186
rect 2145 1112 2151 1146
rect 2185 1112 2191 1146
rect 2145 1072 2191 1112
rect 2145 1038 2151 1072
rect 2185 1038 2191 1072
rect 2145 998 2191 1038
rect 2145 964 2151 998
rect 2185 964 2191 998
rect 2145 924 2191 964
rect 2145 890 2151 924
rect 2185 890 2191 924
rect 2145 850 2191 890
rect 2145 816 2151 850
rect 2185 816 2191 850
rect 2145 776 2191 816
rect 2145 742 2151 776
rect 2185 742 2191 776
rect 2145 702 2191 742
rect 2145 668 2151 702
rect 2185 668 2191 702
rect 2145 628 2191 668
rect 2145 594 2151 628
rect 2185 594 2191 628
rect 2145 554 2191 594
rect 2145 520 2151 554
rect 2185 520 2191 554
rect 2145 480 2191 520
rect 2145 446 2151 480
rect 2185 446 2191 480
rect 2145 406 2191 446
rect 2145 372 2151 406
rect 2185 372 2191 406
rect 2145 332 2191 372
rect 2145 298 2151 332
rect 2185 298 2191 332
rect 2145 258 2191 298
rect 2145 224 2151 258
rect 2185 224 2191 258
rect 2145 184 2191 224
rect 2145 150 2151 184
rect 2185 150 2191 184
rect 2145 110 2191 150
tri 2002 76 2024 98 sw
rect 2145 76 2151 110
rect 2185 76 2191 110
rect 1950 69 2024 76
tri 2024 69 2031 76 sw
rect 1950 59 2031 69
tri 2031 59 2041 69 sw
rect 1950 54 2041 59
tri 2041 54 2046 59 sw
tri 1950 46 1958 54 ne
rect 1958 46 2046 54
tri 2046 46 2054 54 sw
tri 1958 36 1968 46 ne
rect 1968 36 2054 46
tri 2054 36 2064 46 sw
rect 2145 36 2191 76
rect 1866 8 1918 24
tri 1968 2 2002 36 ne
rect 2002 17 2064 36
tri 2064 17 2083 36 sw
rect 2002 2 2083 17
tri 2002 -13 2017 2 ne
rect 2017 -13 2083 2
tri 2017 -27 2031 -13 ne
rect 1866 -60 1918 -44
rect 1866 -128 1918 -112
rect 1866 -196 1918 -180
rect 1866 -265 1918 -248
rect 1866 -334 1918 -317
rect 1866 -392 1918 -386
rect 1948 -53 2000 -47
rect 1948 -117 2000 -105
rect 745 -410 759 -405
rect 682 -413 759 -410
tri 759 -413 767 -405 sw
tri 656 -431 674 -413 se
rect 674 -417 767 -413
tri 767 -417 771 -413 sw
rect 1616 -417 1835 -405
rect 674 -422 771 -417
rect 674 -431 693 -422
rect 558 -437 693 -431
rect 745 -431 771 -422
tri 771 -431 785 -417 sw
tri 1740 -431 1754 -417 ne
rect 1754 -431 1835 -417
rect 745 -437 1552 -431
tri 1754 -433 1756 -431 ne
rect 1756 -433 1835 -431
tri 1835 -433 1842 -426 sw
tri 1756 -434 1757 -433 ne
rect 1757 -434 1842 -433
tri 1842 -434 1843 -433 sw
rect 558 -471 570 -437
rect 604 -471 642 -437
rect 676 -471 693 -437
rect 748 -471 786 -437
rect 820 -471 858 -437
rect 892 -471 930 -437
rect 964 -471 1002 -437
rect 1036 -471 1074 -437
rect 1108 -471 1146 -437
rect 1180 -471 1218 -437
rect 1252 -471 1290 -437
rect 1324 -471 1362 -437
rect 1396 -471 1434 -437
rect 1468 -471 1506 -437
rect 1540 -471 1552 -437
tri 1757 -464 1787 -434 ne
rect 1787 -447 1843 -434
tri 1843 -447 1856 -434 sw
rect 558 -474 693 -471
rect 745 -474 1552 -471
rect 454 -488 506 -482
tri 506 -488 519 -475 sw
rect 558 -477 1552 -474
tri 690 -480 693 -477 ne
rect 693 -480 745 -477
tri 745 -480 748 -477 nw
rect 454 -505 519 -488
tri 519 -505 536 -488 sw
rect 454 -507 536 -505
tri 536 -507 538 -505 sw
rect 454 -509 538 -507
tri 538 -509 540 -507 sw
rect 454 -510 1545 -509
rect 506 -515 1545 -510
rect 506 -549 1427 -515
rect 1461 -549 1499 -515
rect 1533 -549 1545 -515
rect 506 -555 1545 -549
rect 1787 -531 1856 -447
rect 506 -562 530 -555
rect 454 -565 530 -562
tri 530 -565 540 -555 nw
rect 1787 -565 1802 -531
rect 1836 -565 1856 -531
rect 454 -577 518 -565
tri 518 -577 530 -565 nw
rect 454 -580 515 -577
tri 515 -580 518 -577 nw
rect 454 -587 506 -580
rect 454 -590 466 -587
rect 500 -590 506 -587
tri 506 -589 515 -580 nw
rect 558 -593 1552 -587
rect 558 -627 570 -593
rect 604 -627 642 -593
rect 676 -627 714 -593
rect 748 -627 786 -593
rect 820 -627 858 -593
rect 892 -627 930 -593
rect 964 -627 1002 -593
rect 1036 -627 1074 -593
rect 1180 -627 1218 -593
rect 1252 -627 1290 -593
rect 1324 -627 1362 -593
rect 1396 -627 1434 -593
rect 1468 -627 1506 -593
rect 1540 -627 1552 -593
rect 558 -633 1098 -627
tri 1064 -637 1068 -633 ne
rect 1068 -637 1098 -633
tri 1068 -638 1069 -637 ne
rect 1069 -638 1098 -637
rect 454 -660 506 -642
tri 1069 -649 1080 -638 ne
rect 1080 -645 1098 -638
rect 1150 -633 1552 -627
rect 1787 -603 1856 -565
rect 1150 -637 1180 -633
tri 1180 -637 1184 -633 nw
rect 1787 -637 1802 -603
rect 1836 -637 1856 -603
rect 1150 -638 1179 -637
tri 1179 -638 1180 -637 nw
rect 1150 -645 1168 -638
rect 1080 -649 1168 -645
tri 1168 -649 1179 -638 nw
tri 1080 -653 1084 -649 ne
rect 1084 -653 1164 -649
tri 1164 -653 1168 -649 nw
rect 1787 -651 1856 -637
rect 454 -670 466 -660
rect 500 -670 506 -660
tri 1084 -661 1092 -653 ne
rect 1092 -657 1150 -653
rect 1092 -661 1098 -657
rect 937 -667 989 -661
tri 1092 -667 1098 -661 ne
tri 933 -713 937 -709 se
tri 925 -721 933 -713 se
rect 933 -719 937 -713
tri 1150 -667 1164 -653 nw
tri 1934 -687 1948 -673 se
rect 1948 -687 2000 -169
tri 1912 -709 1934 -687 se
rect 1934 -709 2000 -687
tri 989 -713 993 -709 sw
rect 989 -715 993 -713
tri 993 -715 995 -713 sw
rect 1098 -715 1150 -709
tri 1727 -713 1731 -709 se
rect 1731 -713 2000 -709
tri 1725 -715 1727 -713 se
rect 1727 -715 2000 -713
rect 989 -719 995 -715
rect 933 -721 995 -719
tri 995 -721 1001 -715 sw
tri 1719 -721 1725 -715 se
rect 1725 -720 2000 -715
rect 1725 -721 1999 -720
tri 1999 -721 2000 -720 nw
rect 454 -733 506 -722
rect 454 -750 466 -733
rect 500 -750 506 -733
rect 454 -806 506 -802
rect 454 -830 466 -806
rect 500 -830 506 -806
rect 617 -727 669 -721
tri 919 -727 925 -721 se
rect 925 -727 1001 -721
tri 1001 -727 1007 -721 sw
tri 1713 -727 1719 -721 se
rect 1719 -727 1993 -721
tri 1993 -727 1999 -721 nw
tri 903 -743 919 -727 se
rect 919 -731 1007 -727
rect 919 -743 937 -731
rect 617 -791 669 -779
rect 824 -749 937 -743
rect 989 -743 1007 -731
tri 1007 -743 1023 -727 sw
tri 1712 -728 1713 -727 se
rect 1713 -728 1992 -727
tri 1992 -728 1993 -727 nw
rect 1712 -743 1977 -728
tri 1977 -743 1992 -728 nw
rect 989 -749 1552 -743
rect 824 -783 836 -749
rect 870 -783 911 -749
rect 1020 -783 1061 -749
rect 1095 -783 1136 -749
rect 1170 -783 1210 -749
rect 1244 -783 1284 -749
rect 1318 -783 1358 -749
rect 1392 -783 1432 -749
rect 1466 -783 1506 -749
rect 1540 -783 1552 -749
rect 1712 -752 1968 -743
tri 1968 -752 1977 -743 nw
rect 1712 -760 1756 -752
tri 1756 -760 1764 -752 nw
rect 1610 -766 1662 -760
rect 824 -789 1552 -783
tri 1604 -788 1610 -782 se
tri 1603 -789 1604 -788 se
rect 1604 -789 1610 -788
tri 1599 -793 1603 -789 se
rect 1603 -793 1610 -789
tri 1597 -795 1599 -793 se
rect 1599 -795 1610 -793
tri 1591 -801 1597 -795 se
rect 1597 -801 1610 -795
tri 1574 -818 1591 -801 se
rect 1591 -818 1610 -801
rect 669 -830 1662 -818
rect 669 -843 1610 -830
tri 506 -863 524 -845 sw
rect 617 -849 1610 -843
tri 1571 -863 1585 -849 ne
rect 1585 -863 1610 -849
rect 506 -877 524 -863
tri 524 -877 538 -863 sw
tri 1585 -877 1599 -863 ne
rect 1599 -877 1610 -863
rect 506 -880 669 -877
tri 669 -880 672 -877 sw
tri 1599 -880 1602 -877 ne
rect 1602 -880 1610 -877
rect 506 -882 1548 -880
rect 454 -910 466 -882
rect 500 -886 1548 -882
rect 500 -910 666 -886
rect 506 -920 666 -910
rect 700 -920 742 -886
rect 776 -920 818 -886
rect 852 -920 894 -886
rect 928 -920 970 -886
rect 1004 -920 1046 -886
rect 1080 -920 1122 -886
rect 1156 -920 1198 -886
rect 1232 -920 1274 -886
rect 1308 -920 1350 -886
rect 1384 -920 1426 -886
rect 1460 -920 1502 -886
rect 1536 -920 1548 -886
tri 1602 -888 1610 -880 ne
rect 1610 -888 1662 -882
rect 1712 -761 1755 -760
tri 1755 -761 1756 -760 nw
rect 506 -923 1548 -920
rect 506 -926 525 -923
tri 525 -926 528 -923 nw
tri 644 -926 647 -923 ne
rect 647 -926 1548 -923
rect 506 -935 516 -926
tri 516 -935 525 -926 nw
tri 506 -945 516 -935 nw
tri 1622 -945 1628 -939 se
rect 1628 -941 1680 -935
tri 1610 -957 1622 -945 se
rect 1622 -957 1628 -945
rect 454 -986 466 -962
rect 500 -986 506 -962
rect 454 -990 506 -986
rect 535 -1009 541 -957
rect 593 -1009 605 -957
rect 657 -993 1628 -957
rect 657 -995 1680 -993
rect 657 -998 1325 -995
tri 1325 -998 1328 -995 nw
tri 1589 -998 1592 -995 ne
rect 1592 -998 1680 -995
rect 657 -1009 663 -998
tri 1592 -1009 1603 -998 ne
rect 1603 -1005 1680 -998
rect 1603 -1009 1628 -1005
tri 1603 -1018 1612 -1009 ne
rect 1612 -1018 1628 -1009
tri 1612 -1024 1618 -1018 ne
rect 1618 -1024 1628 -1018
tri 1333 -1028 1337 -1024 se
rect 1337 -1028 1343 -1024
rect 454 -1059 466 -1042
rect 500 -1059 506 -1042
rect 454 -1070 506 -1059
rect 1091 -1034 1343 -1028
rect 1091 -1068 1103 -1034
rect 1137 -1068 1183 -1034
rect 1217 -1068 1263 -1034
rect 1297 -1068 1343 -1034
rect 1091 -1074 1343 -1068
tri 1333 -1076 1335 -1074 ne
rect 1335 -1076 1343 -1074
rect 1395 -1076 1415 -1024
rect 1467 -1076 1487 -1024
rect 1539 -1028 1545 -1024
tri 1545 -1028 1549 -1024 sw
rect 1539 -1074 1549 -1028
tri 1618 -1034 1628 -1024 ne
rect 1628 -1063 1680 -1057
rect 1539 -1076 1546 -1074
tri 1546 -1076 1548 -1074 nw
tri 1609 -1104 1616 -1097 se
rect 1616 -1104 1662 -1097
rect 454 -1132 466 -1122
rect 500 -1132 506 -1122
rect 454 -1150 506 -1132
rect 941 -1156 947 -1104
rect 999 -1156 1011 -1104
rect 1063 -1109 1662 -1104
rect 1063 -1143 1622 -1109
rect 1656 -1143 1662 -1109
rect 1063 -1156 1662 -1143
tri 1582 -1164 1590 -1156 ne
rect 1590 -1164 1662 -1156
tri 1590 -1184 1610 -1164 ne
rect 1610 -1184 1662 -1164
rect 454 -1205 466 -1202
rect 500 -1205 506 -1202
rect 454 -1230 506 -1205
rect 558 -1190 1552 -1184
tri 1610 -1190 1616 -1184 ne
rect 558 -1224 570 -1190
rect 604 -1224 642 -1190
rect 676 -1224 714 -1190
rect 748 -1224 786 -1190
rect 820 -1224 858 -1190
rect 892 -1224 930 -1190
rect 964 -1224 1002 -1190
rect 1036 -1224 1074 -1190
rect 1108 -1224 1146 -1190
rect 1180 -1224 1218 -1190
rect 1252 -1224 1256 -1190
rect 1324 -1224 1362 -1190
rect 1396 -1224 1434 -1190
rect 1468 -1224 1506 -1190
rect 1540 -1224 1552 -1190
rect 558 -1230 1256 -1224
tri 1222 -1231 1223 -1230 ne
rect 1223 -1231 1256 -1230
tri 1223 -1264 1256 -1231 ne
rect 1308 -1230 1552 -1224
rect 1308 -1231 1341 -1230
tri 1341 -1231 1342 -1230 nw
rect 1616 -1231 1662 -1184
rect 1256 -1254 1308 -1242
rect 454 -1310 506 -1282
tri 1308 -1264 1341 -1231 nw
rect 1616 -1265 1622 -1231
rect 1656 -1265 1662 -1231
rect 1616 -1277 1662 -1265
rect 1256 -1312 1308 -1306
rect 1609 -1319 1661 -1313
tri 1334 -1340 1337 -1337 se
rect 1337 -1340 1343 -1337
rect 454 -1390 506 -1362
rect 558 -1346 1343 -1340
rect 1395 -1346 1415 -1337
rect 1467 -1346 1487 -1337
rect 1539 -1340 1545 -1337
tri 1545 -1340 1548 -1337 sw
rect 1539 -1346 1552 -1340
rect 558 -1380 570 -1346
rect 604 -1380 642 -1346
rect 676 -1380 714 -1346
rect 748 -1380 786 -1346
rect 820 -1380 858 -1346
rect 892 -1380 930 -1346
rect 964 -1380 1002 -1346
rect 1036 -1380 1074 -1346
rect 1108 -1380 1146 -1346
rect 1180 -1380 1218 -1346
rect 1252 -1380 1290 -1346
rect 1324 -1380 1343 -1346
rect 1396 -1380 1415 -1346
rect 1468 -1380 1487 -1346
rect 1540 -1380 1552 -1346
rect 558 -1386 1343 -1380
tri 1334 -1389 1337 -1386 ne
rect 1337 -1389 1343 -1386
rect 1395 -1389 1415 -1380
rect 1467 -1389 1487 -1380
rect 1539 -1386 1552 -1380
rect 1539 -1389 1545 -1386
tri 1545 -1389 1548 -1386 nw
rect 1609 -1398 1661 -1371
rect 454 -1463 506 -1442
rect 454 -1470 466 -1463
rect 500 -1470 506 -1463
rect 950 -1468 956 -1416
rect 1008 -1468 1035 -1416
rect 1087 -1419 1326 -1416
tri 1326 -1419 1329 -1416 sw
rect 1087 -1450 1609 -1419
rect 1087 -1458 1661 -1450
rect 1087 -1468 1093 -1458
tri 1286 -1466 1294 -1458 ne
rect 1294 -1466 1661 -1458
tri 1129 -1496 1135 -1490 se
rect 1135 -1496 1141 -1490
rect 454 -1536 506 -1522
rect 454 -1550 466 -1536
rect 500 -1550 506 -1536
rect 558 -1502 1141 -1496
rect 558 -1536 570 -1502
rect 604 -1536 642 -1502
rect 676 -1536 714 -1502
rect 748 -1536 786 -1502
rect 820 -1536 858 -1502
rect 892 -1536 930 -1502
rect 964 -1536 1002 -1502
rect 1036 -1536 1074 -1502
rect 1108 -1536 1141 -1502
rect 558 -1542 1141 -1536
rect 1193 -1542 1205 -1490
rect 1257 -1496 1266 -1490
tri 1266 -1496 1272 -1490 sw
rect 1257 -1502 1552 -1496
rect 1257 -1536 1290 -1502
rect 1324 -1536 1362 -1502
rect 1396 -1536 1434 -1502
rect 1468 -1536 1506 -1502
rect 1540 -1536 1552 -1502
rect 1257 -1542 1552 -1536
rect 1613 -1501 1665 -1495
rect 454 -1609 506 -1602
rect 454 -1630 466 -1609
rect 500 -1630 506 -1609
rect 1613 -1580 1665 -1553
rect 1613 -1638 1665 -1632
tri 1331 -1652 1337 -1646 se
rect 1337 -1652 1343 -1646
rect 454 -1710 466 -1682
rect 500 -1710 506 -1682
rect 558 -1658 1343 -1652
rect 1395 -1658 1415 -1646
rect 1467 -1658 1487 -1646
rect 1539 -1652 1545 -1646
tri 1545 -1652 1551 -1646 sw
rect 1539 -1658 1552 -1652
rect 558 -1692 570 -1658
rect 604 -1692 642 -1658
rect 676 -1692 714 -1658
rect 748 -1692 786 -1658
rect 820 -1692 858 -1658
rect 892 -1692 930 -1658
rect 964 -1692 1002 -1658
rect 1036 -1692 1074 -1658
rect 1108 -1692 1146 -1658
rect 1180 -1692 1218 -1658
rect 1252 -1692 1290 -1658
rect 1324 -1692 1343 -1658
rect 1396 -1692 1415 -1658
rect 1468 -1692 1487 -1658
rect 1540 -1692 1552 -1658
rect 558 -1698 1343 -1692
rect 1395 -1698 1415 -1692
rect 1467 -1698 1487 -1692
rect 1539 -1698 1552 -1692
tri 1685 -1698 1712 -1671 se
rect 1712 -1698 1747 -761
tri 1747 -769 1755 -761 nw
tri 1662 -1721 1685 -1698 se
rect 1685 -1721 1747 -1698
rect 454 -1789 466 -1762
rect 500 -1789 506 -1762
rect 1616 -1733 1747 -1721
tri 773 -1767 777 -1763 se
rect 777 -1767 829 -1763
tri 829 -1767 833 -1763 sw
rect 1616 -1767 1622 -1733
rect 1656 -1767 1747 -1733
rect 454 -1790 506 -1789
tri 732 -1808 773 -1767 se
rect 773 -1769 833 -1767
rect 773 -1808 777 -1769
rect 454 -1862 466 -1842
rect 500 -1862 506 -1842
rect 558 -1814 777 -1808
rect 829 -1808 833 -1769
tri 833 -1808 874 -1767 sw
rect 829 -1814 1553 -1808
rect 558 -1848 570 -1814
rect 604 -1848 642 -1814
rect 676 -1848 714 -1814
rect 748 -1821 777 -1814
rect 829 -1821 858 -1814
rect 748 -1833 786 -1821
rect 820 -1833 858 -1821
rect 748 -1848 777 -1833
rect 829 -1848 858 -1833
rect 892 -1848 930 -1814
rect 964 -1848 1002 -1814
rect 1036 -1848 1074 -1814
rect 1108 -1848 1146 -1814
rect 1180 -1848 1218 -1814
rect 1252 -1848 1290 -1814
rect 1324 -1848 1362 -1814
rect 1396 -1848 1434 -1814
rect 1468 -1848 1501 -1814
rect 558 -1854 777 -1848
rect 454 -1870 506 -1862
tri 740 -1891 777 -1854 ne
rect 829 -1854 1501 -1848
rect 777 -1891 829 -1885
tri 829 -1891 866 -1854 nw
tri 1456 -1891 1493 -1854 ne
rect 1493 -1866 1501 -1854
rect 1493 -1878 1553 -1866
rect 1493 -1891 1501 -1878
tri 1493 -1899 1501 -1891 ne
rect 454 -1935 466 -1922
rect 500 -1935 506 -1922
rect 454 -1950 506 -1935
rect 1501 -1936 1553 -1930
rect 1616 -1818 1747 -1767
rect 1616 -1852 1622 -1818
rect 1656 -1852 1747 -1818
rect 1616 -1904 1747 -1852
rect 1616 -1938 1622 -1904
rect 1656 -1938 1747 -1904
rect 1616 -1950 1747 -1938
rect 1779 -801 1831 -795
rect 1779 -865 1831 -853
tri 1105 -1964 1111 -1958 se
rect 1111 -1964 1117 -1958
rect 454 -2008 466 -2002
rect 500 -2008 506 -2002
rect 454 -2031 506 -2008
rect 558 -1970 1117 -1964
rect 1169 -1970 1189 -1958
rect 1241 -1970 1261 -1958
rect 1313 -1964 1319 -1958
tri 1319 -1964 1325 -1958 sw
rect 1313 -1970 1552 -1964
rect 558 -2004 570 -1970
rect 604 -2004 642 -1970
rect 676 -2004 714 -1970
rect 748 -2004 786 -1970
rect 820 -2004 858 -1970
rect 892 -2004 930 -1970
rect 964 -2004 1002 -1970
rect 1036 -2004 1074 -1970
rect 1108 -2004 1117 -1970
rect 1180 -2004 1189 -1970
rect 1252 -2004 1261 -1970
rect 1324 -2004 1362 -1970
rect 1396 -2004 1434 -1970
rect 1468 -2004 1506 -1970
rect 1540 -2004 1552 -1970
rect 558 -2010 1117 -2004
rect 1169 -2010 1189 -2004
rect 1241 -2010 1261 -2004
rect 1313 -2010 1552 -2004
tri 1609 -2040 1616 -2033 se
rect 1616 -2040 1662 -2033
rect 454 -2112 506 -2083
tri 652 -2120 692 -2080 se
rect 692 -2085 745 -2079
rect 692 -2120 693 -2085
rect 454 -2391 506 -2164
rect 558 -2126 693 -2120
tri 745 -2092 758 -2079 sw
rect 859 -2092 865 -2040
rect 917 -2092 929 -2040
rect 981 -2045 1662 -2040
rect 981 -2079 1622 -2045
rect 1656 -2079 1662 -2045
rect 981 -2092 1662 -2079
rect 745 -2120 758 -2092
tri 758 -2120 786 -2092 sw
tri 1582 -2120 1610 -2092 ne
rect 1610 -2120 1662 -2092
rect 745 -2126 1057 -2120
tri 1610 -2126 1616 -2120 ne
rect 558 -2160 570 -2126
rect 604 -2160 644 -2126
rect 678 -2137 693 -2126
rect 678 -2149 718 -2137
rect 678 -2160 693 -2149
rect 752 -2160 792 -2126
rect 826 -2160 865 -2126
rect 899 -2160 938 -2126
rect 972 -2160 1011 -2126
rect 1045 -2160 1057 -2126
rect 1616 -2130 1662 -2120
tri 1104 -2150 1105 -2149 se
rect 1105 -2150 1319 -2149
tri 1319 -2150 1320 -2149 sw
rect 558 -2166 693 -2160
tri 652 -2170 656 -2166 ne
rect 656 -2170 693 -2166
tri 656 -2207 693 -2170 ne
rect 745 -2166 1057 -2160
tri 1100 -2154 1104 -2150 se
rect 1104 -2154 1110 -2150
rect 745 -2170 782 -2166
tri 782 -2170 786 -2166 nw
rect 745 -2201 750 -2170
rect 693 -2202 750 -2201
tri 750 -2202 782 -2170 nw
rect 1100 -2202 1110 -2154
rect 1162 -2202 1185 -2150
rect 1237 -2202 1260 -2150
rect 1312 -2153 1320 -2150
tri 1320 -2153 1323 -2150 sw
rect 1312 -2202 1323 -2153
rect 693 -2207 745 -2202
tri 745 -2207 750 -2202 nw
tri 1096 -2243 1100 -2239 se
rect 1100 -2243 1323 -2202
rect 1616 -2164 1622 -2130
rect 1656 -2164 1662 -2130
rect 1616 -2216 1662 -2164
tri 1089 -2250 1096 -2243 se
rect 1096 -2250 1323 -2243
tri 1323 -2250 1330 -2243 sw
rect 1616 -2250 1622 -2216
rect 1656 -2250 1662 -2216
tri 1063 -2276 1089 -2250 se
rect 1089 -2262 1330 -2250
tri 1330 -2262 1342 -2250 sw
rect 1616 -2262 1662 -2250
rect 1089 -2276 1342 -2262
tri 1342 -2276 1356 -2262 sw
rect 558 -2282 1552 -2276
rect 558 -2316 570 -2282
rect 604 -2316 642 -2282
rect 676 -2316 714 -2282
rect 748 -2316 786 -2282
rect 820 -2316 858 -2282
rect 892 -2316 930 -2282
rect 964 -2316 1002 -2282
rect 1036 -2316 1074 -2282
rect 1108 -2316 1146 -2282
rect 1180 -2316 1218 -2282
rect 1252 -2316 1290 -2282
rect 1324 -2316 1362 -2282
rect 1396 -2316 1434 -2282
rect 1468 -2316 1506 -2282
rect 1540 -2316 1552 -2282
rect 558 -2322 1552 -2316
tri 506 -2391 536 -2361 sw
rect 454 -2397 1574 -2391
rect 454 -2431 597 -2397
rect 631 -2431 675 -2397
rect 709 -2431 753 -2397
rect 787 -2431 831 -2397
rect 865 -2431 909 -2397
rect 943 -2431 987 -2397
rect 1021 -2431 1065 -2397
rect 1099 -2431 1143 -2397
rect 1177 -2431 1220 -2397
rect 1254 -2431 1297 -2397
rect 1331 -2431 1374 -2397
rect 1408 -2431 1451 -2397
rect 1485 -2431 1528 -2397
rect 1562 -2431 1574 -2397
rect 454 -2437 1574 -2431
tri 1753 -2469 1779 -2443 se
rect 1779 -2469 1831 -917
rect 478 -2474 1831 -2469
rect 478 -2499 1806 -2474
tri 1806 -2499 1831 -2474 nw
rect 1860 -896 1912 -890
rect 1860 -960 1912 -948
rect 401 -3243 447 -3231
rect 401 -3277 407 -3243
rect 441 -3277 447 -3243
rect 401 -3316 447 -3277
rect 401 -3350 407 -3316
rect 441 -3350 447 -3316
rect 401 -3389 447 -3350
tri 398 -3423 401 -3420 se
rect 401 -3423 407 -3389
rect 441 -3423 447 -3389
tri 395 -3426 398 -3423 se
rect 398 -3426 447 -3423
rect 395 -3432 447 -3426
rect 395 -3496 407 -3484
rect 441 -3496 447 -3484
rect 395 -3554 407 -3548
tri 395 -3560 401 -3554 ne
rect 401 -3569 407 -3554
rect 441 -3569 447 -3548
rect 401 -3608 447 -3569
rect 401 -3642 407 -3608
rect 441 -3642 447 -3608
rect 401 -3681 447 -3642
rect 401 -3715 407 -3681
rect 441 -3715 447 -3681
rect 401 -3754 447 -3715
rect 401 -3788 407 -3754
rect 441 -3788 447 -3754
rect 401 -3827 447 -3788
rect 401 -3861 407 -3827
rect 441 -3861 447 -3827
rect 401 -3900 447 -3861
rect 401 -3934 407 -3900
rect 441 -3934 447 -3900
rect 401 -3973 447 -3934
rect 401 -4007 407 -3973
rect 441 -4007 447 -3973
rect 401 -4046 447 -4007
rect 401 -4080 407 -4046
rect 441 -4080 447 -4046
rect 401 -4119 447 -4080
rect 401 -4153 407 -4119
rect 441 -4153 447 -4119
rect 401 -4192 447 -4153
tri 399 -4226 401 -4224 se
rect 401 -4226 407 -4192
rect 441 -4226 447 -4192
tri 398 -4227 399 -4226 se
rect 399 -4227 447 -4226
tri 447 -4227 450 -4224 sw
rect 398 -4233 450 -4227
rect 398 -4299 407 -4285
rect 441 -4299 450 -4285
rect 398 -4365 407 -4351
rect 441 -4365 450 -4351
rect 398 -4423 407 -4417
tri 398 -4426 401 -4423 ne
rect 401 -4445 407 -4423
rect 441 -4423 450 -4417
rect 441 -4445 447 -4423
tri 447 -4426 450 -4423 nw
rect 401 -4484 447 -4445
rect 401 -4518 407 -4484
rect 441 -4518 447 -4484
rect 401 -4557 447 -4518
rect 401 -4591 407 -4557
rect 441 -4591 447 -4557
rect 401 -4630 447 -4591
rect 401 -4664 407 -4630
rect 441 -4664 447 -4630
rect 401 -4703 447 -4664
rect 401 -4737 407 -4703
rect 441 -4737 447 -4703
rect 401 -4775 447 -4737
rect 401 -4809 407 -4775
rect 441 -4809 447 -4775
rect 401 -4847 447 -4809
rect 401 -4881 407 -4847
rect 441 -4881 447 -4847
rect 401 -4919 447 -4881
rect 401 -4953 407 -4919
rect 441 -4953 447 -4919
rect 401 -4991 447 -4953
rect 401 -5025 407 -4991
rect 441 -5025 447 -4991
rect 401 -5063 447 -5025
rect 401 -5097 407 -5063
rect 441 -5097 447 -5063
rect 401 -5135 447 -5097
rect 401 -5169 407 -5135
rect 441 -5169 447 -5135
rect 401 -5207 447 -5169
rect 401 -5241 407 -5207
rect 441 -5241 447 -5207
rect 401 -5279 447 -5241
rect 401 -5313 407 -5279
rect 441 -5313 447 -5279
rect 401 -5351 447 -5313
rect 401 -5385 407 -5351
rect 441 -5385 447 -5351
rect 401 -5423 447 -5385
rect 401 -5457 407 -5423
rect 441 -5457 447 -5423
rect 401 -5495 447 -5457
rect 401 -5529 407 -5495
rect 441 -5529 447 -5495
rect 401 -5567 447 -5529
rect 401 -5601 407 -5567
rect 441 -5601 447 -5567
rect 401 -5639 447 -5601
rect 401 -5673 407 -5639
rect 441 -5673 447 -5639
rect 401 -5711 447 -5673
rect 401 -5745 407 -5711
rect 441 -5745 447 -5711
rect 401 -5783 447 -5745
rect 401 -5817 407 -5783
rect 441 -5817 447 -5783
rect 401 -5855 447 -5817
rect 401 -5889 407 -5855
rect 441 -5889 447 -5855
rect 401 -5927 447 -5889
rect 401 -5961 407 -5927
rect 441 -5961 447 -5927
rect 401 -5999 447 -5961
rect 401 -6033 407 -5999
rect 441 -6033 447 -5999
rect 401 -6071 447 -6033
rect 401 -6105 407 -6071
rect 441 -6105 447 -6071
rect 401 -6143 447 -6105
rect 401 -6177 407 -6143
rect 441 -6177 447 -6143
rect 401 -6215 447 -6177
rect 401 -6249 407 -6215
rect 441 -6249 447 -6215
rect 401 -6287 447 -6249
rect 401 -6321 407 -6287
rect 441 -6321 447 -6287
rect 401 -6359 447 -6321
rect 401 -6393 407 -6359
rect 441 -6393 447 -6359
rect 401 -6431 447 -6393
rect 401 -6465 407 -6431
rect 441 -6465 447 -6431
rect 401 -6503 447 -6465
rect 401 -6537 407 -6503
rect 441 -6537 447 -6503
rect 401 -6575 447 -6537
rect 401 -6609 407 -6575
rect 441 -6609 447 -6575
rect 401 -6647 447 -6609
rect 401 -6681 407 -6647
rect 441 -6681 447 -6647
rect 401 -6719 447 -6681
rect 401 -6753 407 -6719
rect 441 -6753 447 -6719
rect 401 -6791 447 -6753
rect 401 -6825 407 -6791
rect 441 -6825 447 -6791
rect 401 -6863 447 -6825
rect 401 -6897 407 -6863
rect 441 -6897 447 -6863
rect 401 -6935 447 -6897
rect 401 -6969 407 -6935
rect 441 -6969 447 -6935
rect 401 -7007 447 -6969
rect 401 -7041 407 -7007
rect 441 -7041 447 -7007
rect 401 -7079 447 -7041
rect 401 -7113 407 -7079
rect 441 -7113 447 -7079
rect 401 -7151 447 -7113
rect 401 -7185 407 -7151
rect 441 -7185 447 -7151
rect 401 -7223 447 -7185
rect 401 -7257 407 -7223
rect 441 -7257 447 -7223
rect 401 -7295 447 -7257
rect 401 -7329 407 -7295
rect 441 -7329 447 -7295
rect 401 -7367 447 -7329
rect 401 -7401 407 -7367
rect 441 -7401 447 -7367
rect 401 -7439 447 -7401
rect 401 -7473 407 -7439
rect 441 -7473 447 -7439
rect 401 -7511 447 -7473
rect 401 -7545 407 -7511
rect 441 -7545 447 -7511
rect 401 -7583 447 -7545
rect 401 -7617 407 -7583
rect 441 -7617 447 -7583
rect 401 -7655 447 -7617
rect 401 -7689 407 -7655
rect 441 -7689 447 -7655
rect 401 -7727 447 -7689
rect 401 -7761 407 -7727
rect 441 -7761 447 -7727
rect 401 -7799 447 -7761
rect 401 -7833 407 -7799
rect 441 -7833 447 -7799
rect 401 -7871 447 -7833
rect 401 -7905 407 -7871
rect 441 -7905 447 -7871
rect 401 -7943 447 -7905
rect 401 -7977 407 -7943
rect 441 -7977 447 -7943
rect 401 -8015 447 -7977
rect 401 -8049 407 -8015
rect 441 -8049 447 -8015
rect 401 -8087 447 -8049
rect 401 -8121 407 -8087
rect 441 -8121 447 -8087
rect 401 -8159 447 -8121
rect 401 -8193 407 -8159
rect 441 -8193 447 -8159
rect 401 -8231 447 -8193
rect 401 -8265 407 -8231
rect 441 -8265 447 -8231
rect 401 -8303 447 -8265
rect 401 -8337 407 -8303
rect 441 -8337 447 -8303
rect 401 -8375 447 -8337
rect 401 -8409 407 -8375
rect 441 -8409 447 -8375
rect 401 -8447 447 -8409
rect 401 -8481 407 -8447
rect 441 -8481 447 -8447
rect 401 -8519 447 -8481
rect 401 -8553 407 -8519
rect 441 -8553 447 -8519
rect 401 -8591 447 -8553
rect 401 -8625 407 -8591
rect 441 -8625 447 -8591
rect 401 -8663 447 -8625
rect 401 -8697 407 -8663
rect 441 -8697 447 -8663
rect 401 -8735 447 -8697
rect 401 -8769 407 -8735
rect 441 -8769 447 -8735
rect 401 -8807 447 -8769
rect 401 -8841 407 -8807
rect 441 -8841 447 -8807
rect 401 -8879 447 -8841
rect 401 -8913 407 -8879
rect 441 -8913 447 -8879
rect 401 -8951 447 -8913
rect 401 -8985 407 -8951
rect 441 -8985 447 -8951
rect 401 -9023 447 -8985
rect 401 -9057 407 -9023
rect 441 -9057 447 -9023
rect 401 -9095 447 -9057
rect 401 -9129 407 -9095
rect 441 -9129 447 -9095
rect 401 -9167 447 -9129
rect 401 -9201 407 -9167
rect 441 -9201 447 -9167
rect 401 -9239 447 -9201
rect 401 -9273 407 -9239
rect 441 -9273 447 -9239
rect 401 -9311 447 -9273
rect 401 -9345 407 -9311
rect 441 -9345 447 -9311
rect 401 -9383 447 -9345
rect 401 -9417 407 -9383
rect 441 -9417 447 -9383
rect 401 -9455 447 -9417
rect 401 -9489 407 -9455
rect 441 -9489 447 -9455
rect 401 -9527 447 -9489
rect 401 -9561 407 -9527
rect 441 -9561 447 -9527
rect 401 -9599 447 -9561
rect 401 -9633 407 -9599
rect 441 -9633 447 -9599
rect 401 -9671 447 -9633
rect 401 -9705 407 -9671
rect 441 -9705 447 -9671
rect 401 -9743 447 -9705
rect 401 -9777 407 -9743
rect 441 -9777 447 -9743
rect 401 -9815 447 -9777
rect 401 -9849 407 -9815
rect 441 -9849 447 -9815
rect 401 -9887 447 -9849
rect 401 -9921 407 -9887
rect 441 -9921 447 -9887
rect 401 -9959 447 -9921
rect 401 -9993 407 -9959
rect 441 -9993 447 -9959
rect 401 -10031 447 -9993
rect 401 -10065 407 -10031
rect 441 -10065 447 -10031
rect 401 -10103 447 -10065
rect 401 -10137 407 -10103
rect 441 -10137 447 -10103
rect 401 -10175 447 -10137
rect 401 -10209 407 -10175
rect 441 -10209 447 -10175
rect 401 -10247 447 -10209
rect 401 -10281 407 -10247
rect 441 -10281 447 -10247
rect 401 -10319 447 -10281
rect 401 -10353 407 -10319
rect 441 -10353 447 -10319
rect 401 -10391 447 -10353
rect 401 -10425 407 -10391
rect 441 -10425 447 -10391
rect 401 -10463 447 -10425
rect 401 -10497 407 -10463
rect 441 -10497 447 -10463
rect 401 -10535 447 -10497
rect 401 -10569 407 -10535
rect 441 -10569 447 -10535
rect 401 -10607 447 -10569
rect 401 -10641 407 -10607
rect 441 -10641 447 -10607
rect 401 -10679 447 -10641
rect 401 -10713 407 -10679
rect 441 -10713 447 -10679
rect 401 -10751 447 -10713
rect 401 -10785 407 -10751
rect 441 -10785 447 -10751
rect 401 -10823 447 -10785
rect 401 -10857 407 -10823
rect 441 -10857 447 -10823
rect 401 -10895 447 -10857
rect 401 -10929 407 -10895
rect 441 -10929 447 -10895
rect 401 -10967 447 -10929
rect 401 -11001 407 -10967
rect 441 -11001 447 -10967
rect 401 -11039 447 -11001
rect 478 -10994 506 -2499
tri 506 -2526 533 -2499 nw
tri 1843 -2526 1860 -2509 se
rect 1860 -2526 1912 -1012
tri 1835 -2534 1843 -2526 se
rect 1843 -2534 1912 -2526
rect 542 -2580 1912 -2534
rect 1949 -987 2001 -981
rect 1949 -1051 2001 -1039
rect 542 -2584 610 -2580
tri 610 -2584 614 -2580 nw
rect 542 -10846 588 -2584
tri 588 -2606 610 -2584 nw
tri 1927 -2606 1949 -2584 se
rect 1949 -2606 2001 -1103
tri 1923 -2610 1927 -2606 se
rect 1927 -2610 2001 -2606
rect 542 -10880 548 -10846
rect 582 -10880 588 -10846
rect 542 -10918 588 -10880
rect 542 -10952 548 -10918
rect 582 -10952 588 -10918
rect 542 -10964 588 -10952
rect 624 -2612 2001 -2610
rect 624 -2638 1975 -2612
tri 1975 -2638 2001 -2612 nw
rect 624 -2644 672 -2638
tri 672 -2644 678 -2638 nw
tri 506 -10994 532 -10968 sw
tri 598 -10994 624 -10968 se
rect 624 -10994 652 -2644
tri 652 -2664 672 -2644 nw
tri 2011 -2664 2031 -2644 se
rect 2031 -2664 2083 -13
rect 2145 2 2151 36
rect 2185 2 2191 36
rect 2145 -38 2191 2
rect 2145 -72 2151 -38
rect 2185 -72 2191 -38
rect 2145 -112 2191 -72
rect 2145 -146 2151 -112
rect 2185 -146 2191 -112
rect 2145 -186 2191 -146
tri 2221 2391 2241 2411 se
rect 2241 2398 8554 2411
tri 8554 2398 8567 2411 nw
rect 2241 2391 2284 2398
tri 2284 2391 2291 2398 nw
tri 8613 2391 8618 2396 se
rect 8618 2391 8648 3254
tri 8648 3244 8658 3254 nw
rect 8715 3244 8763 3254
tri 8763 3244 8773 3254 nw
rect 2221 2377 2270 2391
tri 2270 2377 2284 2391 nw
tri 8599 2377 8613 2391 se
rect 8613 2377 8648 2391
rect 2221 -40 2257 2377
tri 2257 2364 2270 2377 nw
tri 8592 2370 8599 2377 se
rect 8599 2370 8648 2377
tri 2331 2364 2337 2370 se
rect 2337 2364 8648 2370
tri 2330 2363 2331 2364 se
rect 2331 2363 8648 2364
tri 2305 2338 2330 2363 se
rect 2330 2362 8648 2363
rect 2330 2340 8626 2362
tri 8626 2340 8648 2362 nw
rect 2330 2338 2364 2340
tri 2364 2338 2366 2340 nw
tri 2302 2335 2305 2338 se
rect 2305 2335 2361 2338
tri 2361 2335 2364 2338 nw
rect 2302 2308 2334 2335
tri 2334 2308 2361 2335 nw
tri 2257 -40 2266 -31 sw
rect 2221 -47 2266 -40
tri 2266 -47 2273 -40 sw
rect 2221 -53 2273 -47
rect 2221 -117 2273 -105
rect 2221 -175 2273 -169
rect 2145 -220 2151 -186
rect 2185 -220 2191 -186
tri 2280 -215 2302 -193 se
rect 2302 -215 2332 2308
tri 2332 2306 2334 2308 nw
rect 7459 2256 7465 2308
rect 7517 2256 7529 2308
rect 7581 2256 7587 2308
tri 8601 2278 8604 2281 se
rect 8604 2278 8650 2281
tri 8650 2278 8653 2281 sw
rect 8601 2272 8653 2278
tri 7657 2245 7658 2246 se
rect 7658 2245 7664 2246
tri 7655 2243 7657 2245 se
rect 7657 2243 7664 2245
tri 4382 2237 4386 2241 se
rect 4386 2237 4392 2241
rect 2431 2231 2758 2237
rect 2431 2197 2443 2231
rect 2477 2197 2535 2231
rect 2569 2197 2627 2231
rect 2661 2225 2758 2231
rect 3060 2231 4392 2237
rect 4444 2231 4476 2241
rect 4528 2231 4560 2241
rect 4612 2231 4644 2241
rect 4696 2240 4702 2241
tri 4702 2240 4703 2241 sw
rect 4696 2237 4703 2240
tri 4703 2237 4706 2240 sw
tri 7138 2237 7141 2240 se
rect 7141 2237 7147 2240
rect 4696 2231 7147 2237
rect 3060 2225 3138 2231
rect 2661 2219 3138 2225
rect 2661 2197 2790 2219
rect 2431 2191 2790 2197
rect 2712 2185 2790 2191
rect 2824 2185 2882 2219
rect 2916 2185 2974 2219
rect 3008 2197 3138 2219
rect 3172 2197 3211 2231
rect 3245 2197 3284 2231
rect 3318 2197 3357 2231
rect 3391 2197 3430 2231
rect 3464 2197 3503 2231
rect 3537 2197 3576 2231
rect 3610 2197 3649 2231
rect 3683 2197 3722 2231
rect 3756 2197 3795 2231
rect 3829 2197 3868 2231
rect 3902 2197 3941 2231
rect 3975 2197 4014 2231
rect 4048 2197 4087 2231
rect 4121 2197 4160 2231
rect 4194 2197 4233 2231
rect 4267 2197 4306 2231
rect 4340 2197 4379 2231
rect 4444 2197 4452 2231
rect 4559 2197 4560 2231
rect 4632 2197 4644 2231
rect 4705 2197 4744 2231
rect 4778 2197 4817 2231
rect 4851 2197 4890 2231
rect 4924 2197 4963 2231
rect 4997 2197 5036 2231
rect 5070 2197 5109 2231
rect 5143 2197 5182 2231
rect 5216 2197 5255 2231
rect 5289 2197 5328 2231
rect 5362 2197 5401 2231
rect 5435 2197 5474 2231
rect 5508 2197 5547 2231
rect 5581 2197 5620 2231
rect 5654 2197 5693 2231
rect 5727 2197 5766 2231
rect 5800 2197 5839 2231
rect 5873 2197 5912 2231
rect 5946 2197 5985 2231
rect 6019 2197 6058 2231
rect 6092 2197 6131 2231
rect 6165 2197 6204 2231
rect 6238 2197 6277 2231
rect 6311 2197 6350 2231
rect 6384 2197 6423 2231
rect 6457 2197 6496 2231
rect 6530 2197 6569 2231
rect 6603 2197 6641 2231
rect 6675 2197 6713 2231
rect 6747 2197 6785 2231
rect 6819 2197 6857 2231
rect 6891 2197 6929 2231
rect 6963 2197 7147 2231
rect 3008 2191 4392 2197
rect 3008 2185 3106 2191
tri 4382 2189 4384 2191 ne
rect 4384 2189 4392 2191
rect 4444 2189 4476 2197
rect 4528 2189 4560 2197
rect 4612 2189 4644 2197
rect 4696 2191 7147 2197
rect 4696 2189 4702 2191
tri 4702 2189 4704 2191 nw
tri 7138 2189 7140 2191 ne
rect 7140 2189 7147 2191
tri 7140 2188 7141 2189 ne
rect 7141 2188 7147 2189
rect 7199 2188 7211 2240
rect 7263 2237 7269 2240
tri 7269 2237 7272 2240 sw
rect 7263 2191 7272 2237
rect 7655 2197 7664 2243
tri 7655 2194 7658 2197 ne
rect 7658 2194 7664 2197
rect 7716 2194 7728 2246
rect 7780 2245 7786 2246
tri 7786 2245 7787 2246 sw
rect 7780 2243 7787 2245
tri 7787 2243 7789 2245 sw
rect 7780 2237 8544 2243
rect 7780 2203 7821 2237
rect 7855 2203 7898 2237
rect 7932 2203 7975 2237
rect 8009 2203 8052 2237
rect 8086 2203 8129 2237
rect 8163 2203 8206 2237
rect 8240 2203 8283 2237
rect 8317 2203 8359 2237
rect 8393 2203 8435 2237
rect 8469 2203 8544 2237
rect 7780 2197 8544 2203
rect 7780 2194 7786 2197
tri 7786 2194 7789 2197 nw
tri 8473 2194 8476 2197 ne
rect 8476 2194 8544 2197
rect 7263 2188 7269 2191
tri 7269 2188 7272 2191 nw
tri 8476 2188 8482 2194 ne
rect 8482 2188 8544 2194
rect 2712 2179 3106 2185
tri 8482 2179 8491 2188 ne
rect 8491 2179 8544 2188
tri 8491 2173 8497 2179 ne
rect 8497 2173 8544 2179
tri 8497 2172 8498 2173 ne
tri 6047 2145 6048 2146 se
rect 6048 2145 6054 2146
tri 3036 2143 3038 2145 se
rect 3038 2143 3044 2145
rect 2408 2137 3044 2143
rect 3096 2137 3115 2145
rect 3167 2137 3186 2145
rect 3238 2137 3256 2145
rect 3308 2143 3314 2145
tri 3314 2143 3316 2145 sw
tri 6045 2143 6047 2145 se
rect 6047 2143 6054 2145
rect 3308 2137 4410 2143
rect 2408 2103 2420 2137
rect 2454 2103 2492 2137
rect 2526 2103 2564 2137
rect 2598 2103 2636 2137
rect 2670 2103 2708 2137
rect 2742 2103 2780 2137
rect 2814 2103 2852 2137
rect 2886 2103 2924 2137
rect 2958 2103 2996 2137
rect 3030 2103 3044 2137
rect 3102 2103 3115 2137
rect 3174 2103 3186 2137
rect 3246 2103 3256 2137
rect 3318 2103 3356 2137
rect 3390 2103 3428 2137
rect 3462 2103 3500 2137
rect 3534 2103 3572 2137
rect 3606 2103 3644 2137
rect 3678 2103 3716 2137
rect 3750 2103 3788 2137
rect 3822 2103 3860 2137
rect 3894 2103 3932 2137
rect 3966 2103 4004 2137
rect 4038 2103 4076 2137
rect 4110 2103 4148 2137
rect 4182 2103 4220 2137
rect 4254 2103 4292 2137
rect 4326 2103 4364 2137
rect 4398 2103 4410 2137
rect 2408 2097 3044 2103
tri 3033 2093 3037 2097 ne
rect 3037 2093 3044 2097
rect 3096 2093 3115 2103
rect 3167 2093 3186 2103
rect 3238 2093 3256 2103
rect 3308 2097 4410 2103
rect 4676 2137 6054 2143
rect 4676 2103 4688 2137
rect 4722 2103 4760 2137
rect 4794 2103 4832 2137
rect 4866 2103 4904 2137
rect 4938 2103 4976 2137
rect 5010 2103 5048 2137
rect 5082 2103 5120 2137
rect 5154 2103 5192 2137
rect 5226 2103 5264 2137
rect 5298 2103 5336 2137
rect 5370 2103 5408 2137
rect 5442 2103 5480 2137
rect 5514 2103 5552 2137
rect 5586 2103 5624 2137
rect 5658 2103 5696 2137
rect 5730 2103 5768 2137
rect 5802 2103 5840 2137
rect 5874 2103 5912 2137
rect 5946 2103 5984 2137
rect 6018 2103 6054 2137
rect 4676 2097 6054 2103
rect 3308 2094 3315 2097
tri 3315 2094 3318 2097 nw
tri 6045 2094 6048 2097 ne
rect 6048 2094 6054 2097
rect 6106 2094 6118 2146
rect 6170 2143 6176 2146
tri 6176 2143 6179 2146 sw
rect 6170 2137 7094 2143
rect 6170 2103 6200 2137
rect 6234 2103 6272 2137
rect 6306 2103 6344 2137
rect 6378 2103 6416 2137
rect 6450 2103 6488 2137
rect 6522 2103 6560 2137
rect 6594 2103 6632 2137
rect 6666 2103 7094 2137
rect 6170 2097 7094 2103
rect 6170 2094 6176 2097
tri 6176 2094 6179 2097 nw
tri 7014 2094 7017 2097 ne
rect 7017 2094 7094 2097
rect 3308 2093 3314 2094
tri 3314 2093 3315 2094 nw
rect 4463 2088 4515 2094
rect 4463 2022 4515 2036
rect 4463 1955 4515 1970
rect 2408 1901 2422 1910
rect 2474 1901 2493 1910
rect 2408 1867 2420 1901
rect 2474 1867 2492 1901
rect 2408 1858 2422 1867
rect 2474 1858 2493 1867
rect 2545 1858 2564 1910
rect 2616 1858 2634 1910
rect 2686 1907 2692 1910
tri 2692 1907 2695 1910 sw
tri 3860 1907 3863 1910 se
rect 3863 1907 3869 1910
rect 2686 1901 3869 1907
rect 3921 1901 3940 1910
rect 3992 1901 4011 1910
rect 4063 1901 4081 1910
rect 4133 1907 4139 1910
tri 4139 1907 4142 1910 sw
rect 4133 1901 4410 1907
rect 2686 1867 2708 1901
rect 2742 1867 2780 1901
rect 2814 1867 2852 1901
rect 2886 1867 2924 1901
rect 2958 1867 2996 1901
rect 3030 1867 3068 1901
rect 3102 1867 3140 1901
rect 3174 1867 3212 1901
rect 3246 1867 3284 1901
rect 3318 1867 3356 1901
rect 3390 1867 3428 1901
rect 3462 1867 3500 1901
rect 3534 1867 3572 1901
rect 3606 1867 3644 1901
rect 3678 1867 3716 1901
rect 3750 1867 3788 1901
rect 3822 1867 3860 1901
rect 3921 1867 3932 1901
rect 3992 1867 4004 1901
rect 4063 1867 4076 1901
rect 4133 1867 4148 1901
rect 4182 1867 4220 1901
rect 4254 1867 4292 1901
rect 4326 1867 4364 1901
rect 4398 1867 4410 1901
rect 2686 1861 3869 1867
rect 2686 1858 2693 1861
tri 2693 1858 2696 1861 nw
tri 3860 1858 3863 1861 ne
rect 3863 1858 3869 1861
rect 3921 1858 3940 1867
rect 3992 1858 4011 1867
rect 4063 1858 4081 1867
rect 4133 1861 4410 1867
rect 4463 1894 4472 1903
rect 4506 1894 4515 1903
rect 4463 1888 4515 1894
rect 4133 1858 4139 1861
tri 4139 1858 4142 1861 nw
rect 4463 1821 4472 1836
rect 4506 1821 4515 1836
rect 4463 1754 4472 1769
rect 4506 1754 4515 1769
rect 4463 1697 4515 1702
rect 4463 1687 4472 1697
rect 4506 1687 4515 1697
tri 3035 1671 3038 1674 se
rect 3038 1671 3044 1674
rect 2408 1665 3044 1671
rect 3096 1665 3115 1674
rect 3167 1665 3186 1674
rect 3238 1665 3256 1674
rect 3308 1671 3314 1674
tri 3314 1671 3317 1674 sw
rect 3308 1665 4410 1671
rect 2408 1631 2420 1665
rect 2454 1631 2492 1665
rect 2526 1631 2564 1665
rect 2598 1631 2636 1665
rect 2670 1631 2708 1665
rect 2742 1631 2780 1665
rect 2814 1631 2852 1665
rect 2886 1631 2924 1665
rect 2958 1631 2996 1665
rect 3030 1631 3044 1665
rect 3102 1631 3115 1665
rect 3174 1631 3186 1665
rect 3246 1631 3256 1665
rect 3318 1631 3356 1665
rect 3390 1631 3428 1665
rect 3462 1631 3500 1665
rect 3534 1631 3572 1665
rect 3606 1631 3644 1665
rect 3678 1631 3716 1665
rect 3750 1631 3788 1665
rect 3822 1631 3860 1665
rect 3894 1631 3932 1665
rect 3966 1631 4004 1665
rect 4038 1631 4076 1665
rect 4110 1631 4148 1665
rect 4182 1631 4220 1665
rect 4254 1631 4292 1665
rect 4326 1631 4364 1665
rect 4398 1631 4410 1665
rect 2408 1625 3044 1631
tri 3035 1622 3038 1625 ne
rect 3038 1622 3044 1625
rect 3096 1622 3115 1631
rect 3167 1622 3186 1631
rect 3238 1622 3256 1631
rect 3308 1625 4410 1631
rect 4568 2088 4620 2094
tri 7017 2087 7024 2094 ne
rect 7024 2087 7094 2094
rect 8498 2119 8544 2173
rect 8601 2211 8613 2220
rect 8647 2211 8653 2220
rect 8601 2208 8653 2211
rect 8601 2149 8613 2156
tri 8601 2143 8607 2149 ne
rect 8607 2139 8613 2149
rect 8647 2139 8653 2156
tri 8544 2119 8558 2133 sw
rect 8607 2127 8653 2139
rect 8498 2113 8558 2119
tri 8558 2113 8564 2119 sw
tri 8498 2087 8524 2113 ne
rect 8524 2087 8564 2113
tri 7024 2085 7026 2087 ne
rect 7026 2085 7094 2087
tri 7026 2081 7030 2085 ne
rect 7030 2081 7094 2085
tri 7030 2063 7048 2081 ne
rect 4568 2018 4620 2036
rect 4568 1955 4580 1966
rect 4614 1955 4620 1966
rect 4568 1947 4620 1955
rect 6823 1958 6869 1970
rect 6823 1924 6829 1958
rect 6863 1924 6869 1958
tri 6648 1908 6650 1910 se
rect 6650 1908 6659 1910
tri 6647 1907 6648 1908 se
rect 6648 1907 6659 1908
rect 4568 1876 4580 1895
rect 4614 1876 4620 1895
rect 4676 1901 6659 1907
rect 4676 1867 4688 1901
rect 4722 1867 4760 1901
rect 4794 1867 4832 1901
rect 4866 1867 4904 1901
rect 4938 1867 4976 1901
rect 5010 1867 5048 1901
rect 5082 1867 5120 1901
rect 5154 1867 5192 1901
rect 5226 1867 5264 1901
rect 5298 1867 5336 1901
rect 5370 1867 5408 1901
rect 5442 1867 5480 1901
rect 5514 1867 5552 1901
rect 5586 1867 5624 1901
rect 5658 1867 5696 1901
rect 5730 1867 5768 1901
rect 5802 1867 5840 1901
rect 5874 1867 5912 1901
rect 5946 1867 5984 1901
rect 6018 1867 6056 1901
rect 6090 1867 6128 1901
rect 6162 1867 6200 1901
rect 6234 1867 6272 1901
rect 6306 1867 6344 1901
rect 6378 1867 6416 1901
rect 6450 1867 6488 1901
rect 6522 1867 6560 1901
rect 6594 1867 6632 1901
rect 4676 1861 6659 1867
tri 6647 1858 6650 1861 ne
rect 6650 1858 6659 1861
rect 6711 1858 6723 1910
rect 6775 1858 6781 1910
tri 6699 1852 6705 1858 ne
rect 6705 1852 6781 1858
tri 6705 1846 6711 1852 ne
rect 6711 1846 6781 1852
tri 6711 1836 6721 1846 ne
rect 6721 1836 6781 1846
tri 6721 1829 6728 1836 ne
rect 6728 1829 6781 1836
rect 4568 1811 4620 1824
tri 6728 1823 6734 1829 ne
rect 6734 1823 6781 1829
tri 6734 1822 6735 1823 ne
rect 4568 1805 4580 1811
rect 4614 1805 4620 1811
rect 4568 1734 4620 1753
rect 4568 1676 4620 1682
tri 6045 1671 6048 1674 se
rect 6048 1671 6054 1674
rect 3308 1622 3314 1625
tri 3314 1622 3317 1625 nw
rect 4463 1620 4515 1635
rect 4676 1665 6054 1671
rect 4676 1631 4688 1665
rect 4722 1631 4760 1665
rect 4794 1631 4832 1665
rect 4866 1631 4904 1665
rect 4938 1631 4976 1665
rect 5010 1631 5048 1665
rect 5082 1631 5120 1665
rect 5154 1631 5192 1665
rect 5226 1631 5264 1665
rect 5298 1631 5336 1665
rect 5370 1631 5408 1665
rect 5442 1631 5480 1665
rect 5514 1631 5552 1665
rect 5586 1631 5624 1665
rect 5658 1631 5696 1665
rect 5730 1631 5768 1665
rect 5802 1631 5840 1665
rect 5874 1631 5912 1665
rect 5946 1631 5984 1665
rect 6018 1631 6054 1665
rect 4676 1625 6054 1631
tri 6045 1622 6048 1625 ne
rect 6048 1622 6054 1625
rect 6106 1622 6118 1674
rect 6170 1671 6176 1674
tri 6176 1671 6179 1674 sw
rect 6170 1665 6678 1671
rect 6170 1631 6200 1665
rect 6234 1631 6272 1665
rect 6306 1631 6344 1665
rect 6378 1631 6416 1665
rect 6450 1631 6488 1665
rect 6522 1631 6560 1665
rect 6594 1631 6632 1665
rect 6666 1631 6678 1665
rect 6170 1625 6678 1631
rect 6735 1640 6781 1823
rect 6823 1886 6869 1924
rect 6823 1852 6829 1886
rect 6863 1852 6869 1886
tri 7037 1852 7048 1863 se
rect 7048 1852 7094 2081
rect 7487 2085 8481 2087
tri 8524 2086 8525 2087 ne
rect 8525 2086 8564 2087
tri 8481 2085 8482 2086 sw
tri 8525 2085 8526 2086 ne
rect 8526 2085 8564 2086
tri 8564 2085 8592 2113 sw
rect 7487 2081 8482 2085
rect 7487 2047 7499 2081
rect 7533 2047 7571 2081
rect 7605 2047 7643 2081
rect 7677 2047 7715 2081
rect 7749 2047 7787 2081
rect 7821 2047 7859 2081
rect 7893 2047 7931 2081
rect 7965 2047 8003 2081
rect 8037 2047 8075 2081
rect 8109 2047 8147 2081
rect 8181 2047 8219 2081
rect 8253 2047 8291 2081
rect 8325 2047 8363 2081
rect 8397 2047 8435 2081
rect 8469 2066 8482 2081
tri 8482 2066 8501 2085 sw
tri 8526 2066 8545 2085 ne
rect 8545 2079 8592 2085
tri 8592 2079 8598 2085 sw
rect 8545 2066 8598 2079
tri 8598 2066 8611 2079 sw
rect 8469 2062 8501 2066
tri 8501 2062 8505 2066 sw
tri 8545 2062 8549 2066 ne
rect 8549 2062 8611 2066
tri 8611 2062 8615 2066 sw
rect 8469 2047 8505 2062
tri 8505 2047 8520 2062 sw
tri 8549 2047 8564 2062 ne
rect 8564 2047 8615 2062
tri 8615 2047 8630 2062 sw
rect 7487 2042 8520 2047
tri 8520 2042 8525 2047 sw
rect 7487 2041 8525 2042
tri 8342 2013 8370 2041 ne
rect 8370 2013 8525 2041
tri 8564 2013 8598 2047 ne
rect 8598 2027 8630 2047
tri 8630 2027 8650 2047 sw
tri 8370 2012 8371 2013 ne
rect 8371 2012 8525 2013
tri 8371 1987 8396 2012 ne
rect 8396 1987 8525 2012
tri 8396 1979 8404 1987 ne
rect 7297 1919 7303 1971
rect 7355 1919 7367 1971
rect 7419 1919 8143 1971
rect 8195 1919 8207 1971
rect 8259 1919 8266 1971
rect 8404 1958 8525 1987
rect 8404 1924 8485 1958
rect 8519 1924 8525 1958
rect 8404 1915 8525 1924
tri 8404 1912 8407 1915 ne
rect 8407 1912 8525 1915
tri 8407 1908 8411 1912 ne
rect 8411 1908 8525 1912
tri 8411 1886 8433 1908 ne
rect 8433 1886 8525 1908
tri 8433 1863 8456 1886 ne
rect 8456 1863 8485 1886
tri 7094 1852 7105 1863 sw
tri 8456 1852 8467 1863 ne
rect 8467 1852 8485 1863
rect 8519 1852 8525 1886
rect 6823 1758 6869 1852
tri 7031 1846 7037 1852 se
rect 7037 1846 7105 1852
tri 7105 1846 7111 1852 sw
tri 8467 1846 8473 1852 ne
rect 8473 1846 8525 1852
tri 7021 1836 7031 1846 se
rect 7031 1840 7111 1846
tri 7111 1840 7117 1846 sw
tri 8473 1840 8479 1846 ne
rect 8479 1840 8525 1846
rect 7031 1836 7117 1840
tri 7117 1836 7121 1840 sw
tri 7014 1829 7021 1836 se
rect 7021 1835 7121 1836
tri 7121 1835 7122 1836 sw
rect 7021 1829 7122 1835
tri 7122 1829 7128 1835 sw
tri 7884 1829 7890 1835 se
rect 7890 1829 7896 1835
rect 6955 1823 7896 1829
rect 7948 1823 7977 1835
rect 8029 1829 8035 1835
tri 8035 1829 8041 1835 sw
rect 8029 1823 8447 1829
rect 6955 1789 6967 1823
rect 7001 1789 7043 1823
rect 7077 1789 7119 1823
rect 7153 1789 7195 1823
rect 7229 1789 7271 1823
rect 7305 1789 7347 1823
rect 7381 1789 7423 1823
rect 7457 1789 7499 1823
rect 7533 1789 7575 1823
rect 7609 1789 7651 1823
rect 7685 1789 7726 1823
rect 7760 1789 7801 1823
rect 7835 1789 7876 1823
rect 7948 1789 7951 1823
rect 8060 1789 8101 1823
rect 8135 1789 8176 1823
rect 8210 1789 8251 1823
rect 8285 1789 8326 1823
rect 8360 1789 8401 1823
rect 8435 1789 8447 1823
rect 6955 1783 7896 1789
rect 7948 1783 7977 1789
rect 8029 1783 8447 1789
rect 8598 1774 8650 2027
tri 8477 1768 8479 1770 se
rect 8479 1768 8525 1770
tri 8467 1758 8477 1768 se
rect 8477 1758 8525 1768
rect 6823 1724 6829 1758
rect 6863 1724 6869 1758
tri 8456 1747 8467 1758 se
rect 8467 1747 8485 1758
tri 7362 1740 7369 1747 se
rect 7369 1740 8485 1747
rect 6823 1686 6869 1724
rect 6823 1652 6829 1686
rect 6863 1652 6869 1686
tri 6781 1640 6783 1642 sw
rect 6823 1640 6869 1652
rect 6966 1724 8485 1740
rect 8519 1724 8525 1758
rect 6966 1715 8525 1724
rect 6966 1663 7007 1715
rect 7059 1663 7105 1715
rect 7157 1663 7202 1715
rect 7254 1686 8525 1715
rect 7254 1663 8485 1686
rect 6966 1652 8485 1663
rect 8519 1652 8525 1686
rect 8598 1710 8650 1722
rect 8598 1652 8650 1658
rect 6966 1646 8525 1652
rect 6966 1640 7471 1646
tri 7471 1640 7477 1646 nw
tri 8324 1640 8330 1646 ne
rect 8330 1640 8525 1646
rect 6735 1639 6783 1640
tri 6783 1639 6784 1640 sw
rect 6966 1639 7470 1640
tri 7470 1639 7471 1640 nw
tri 8330 1639 8331 1640 ne
rect 8331 1639 8525 1640
rect 6735 1637 6784 1639
tri 6784 1637 6786 1639 sw
rect 6735 1635 6786 1637
tri 6786 1635 6788 1637 sw
rect 6170 1622 6176 1625
tri 6176 1622 6179 1625 nw
rect 6735 1622 6788 1635
tri 6788 1622 6801 1635 sw
tri 8702 1622 8715 1635 se
rect 8715 1622 8761 3244
tri 8761 3242 8763 3244 nw
rect 9935 3220 9941 3254
rect 9975 3220 9981 3254
tri 9559 3203 9565 3209 se
rect 9565 3203 9572 3209
rect 8877 3197 9572 3203
rect 9624 3197 9640 3209
rect 9692 3208 9698 3209
tri 9698 3208 9699 3209 sw
rect 9935 3208 9981 3220
rect 10064 3337 10110 3349
rect 10064 3303 10070 3337
rect 10104 3303 10110 3337
rect 10174 3336 10186 3370
rect 10220 3336 10258 3370
rect 10292 3336 10330 3370
rect 10364 3336 10402 3370
rect 10436 3336 10474 3370
rect 10508 3336 10546 3370
rect 10580 3336 10618 3370
rect 10652 3336 10690 3370
rect 10724 3336 10762 3370
rect 10796 3336 10834 3370
rect 10868 3336 10906 3370
rect 10940 3336 10978 3370
rect 11012 3336 11050 3370
rect 11084 3336 11122 3370
rect 11156 3359 11298 3370
rect 11332 3359 11379 3393
rect 11156 3336 11379 3359
rect 10174 3330 11379 3336
tri 10174 3324 10180 3330 ne
rect 10180 3324 11379 3330
tri 11262 3315 11271 3324 ne
rect 11271 3315 11379 3324
rect 10064 3265 10110 3303
tri 11271 3296 11290 3315 ne
rect 10064 3231 10070 3265
rect 10104 3231 10110 3265
rect 10064 3219 10110 3231
rect 11290 3281 11298 3315
rect 11332 3281 11379 3315
rect 11290 3237 11379 3281
rect 10064 3214 10105 3219
tri 10105 3214 10110 3219 nw
rect 10174 3214 10797 3220
rect 10849 3214 10869 3220
rect 10921 3214 10941 3220
rect 10993 3214 11012 3220
rect 11064 3214 11083 3220
rect 11135 3214 11168 3220
rect 9692 3203 9699 3208
tri 9699 3203 9704 3208 sw
rect 9692 3197 9871 3203
rect 8877 3163 8889 3197
rect 8923 3163 8961 3197
rect 8995 3163 9033 3197
rect 9067 3163 9105 3197
rect 9139 3163 9177 3197
rect 9211 3163 9249 3197
rect 9283 3163 9321 3197
rect 9355 3163 9393 3197
rect 9427 3163 9465 3197
rect 9499 3163 9537 3197
rect 9571 3163 9572 3197
rect 9715 3163 9753 3197
rect 9787 3163 9825 3197
rect 9859 3163 9871 3197
rect 8877 3157 9572 3163
rect 9624 3157 9640 3163
rect 9692 3157 9871 3163
rect 8875 3075 8881 3127
rect 8933 3075 8945 3127
rect 8997 3079 9893 3127
rect 8997 3075 9003 3079
tri 9003 3075 9007 3079 nw
tri 9883 3075 9887 3079 ne
rect 9887 3075 9893 3079
rect 9945 3075 9957 3127
rect 10009 3075 10015 3127
rect 10064 3125 10100 3214
tri 10100 3209 10105 3214 nw
rect 10174 3180 10186 3214
rect 10220 3180 10258 3214
rect 10292 3180 10330 3214
rect 10364 3180 10402 3214
rect 10436 3180 10474 3214
rect 10508 3180 10546 3214
rect 10580 3180 10618 3214
rect 10652 3180 10690 3214
rect 10724 3180 10762 3214
rect 10796 3180 10797 3214
rect 10868 3180 10869 3214
rect 10940 3180 10941 3214
rect 11156 3180 11168 3214
rect 10174 3174 10797 3180
tri 10785 3168 10791 3174 ne
rect 10791 3168 10797 3174
rect 10849 3168 10869 3180
rect 10921 3168 10941 3180
rect 10993 3168 11012 3180
rect 11064 3168 11083 3180
rect 11135 3174 11168 3180
rect 11290 3203 11298 3237
rect 11332 3203 11379 3237
rect 11135 3168 11141 3174
tri 11141 3168 11147 3174 nw
rect 11290 3159 11379 3203
tri 10100 3125 10110 3135 sw
rect 11290 3125 11298 3159
rect 11332 3125 11379 3159
rect 10064 3107 10110 3125
tri 10110 3107 10128 3125 sw
tri 11273 3107 11290 3124 se
rect 11290 3107 11379 3125
rect 10064 3055 10070 3107
rect 10122 3055 10134 3107
rect 10186 3055 10192 3107
tri 11262 3096 11273 3107 se
rect 11273 3096 11379 3107
tri 11259 3093 11262 3096 se
rect 11262 3093 11379 3096
rect 10284 3087 11379 3093
rect 10284 3053 10362 3087
rect 10396 3053 10434 3087
rect 10468 3053 10506 3087
rect 10540 3053 10578 3087
rect 10612 3053 10650 3087
rect 10684 3053 10722 3087
rect 10756 3053 10794 3087
rect 10828 3053 10866 3087
rect 10900 3053 10938 3087
rect 10972 3053 11010 3087
rect 11044 3053 11082 3087
rect 11116 3053 11154 3087
rect 11188 3053 11226 3087
rect 11260 3053 11379 3087
tri 11438 3758 11444 3764 se
rect 11444 3758 11490 4491
tri 11490 4480 11501 4491 nw
rect 11552 4439 11591 4491
rect 11643 4439 11656 4491
rect 11708 4486 14402 4491
tri 14402 4486 14407 4491 sw
tri 14591 4486 14596 4491 se
rect 14596 4486 17684 4491
rect 11708 4457 17684 4486
rect 17718 4457 17728 4491
tri 18388 4458 18392 4462 se
rect 18392 4458 18427 4587
tri 18427 4576 18438 4587 nw
rect 11708 4445 17728 4457
tri 18376 4446 18388 4458 se
rect 18388 4446 18427 4458
rect 19359 4564 19667 4576
rect 19359 4530 19365 4564
rect 19399 4530 19627 4564
rect 19661 4530 19667 4564
rect 19359 4492 19667 4530
rect 19359 4458 19365 4492
rect 19399 4458 19627 4492
rect 19661 4458 19667 4492
rect 19359 4446 19667 4458
rect 19964 4556 20016 4569
rect 19964 4491 20016 4504
tri 18375 4445 18376 4446 se
rect 18376 4445 18427 4446
rect 11708 4441 11716 4445
tri 11716 4441 11720 4445 nw
tri 18371 4441 18375 4445 se
rect 18375 4441 18427 4445
rect 11708 4439 11714 4441
tri 11714 4439 11716 4441 nw
tri 18369 4439 18371 4441 se
rect 18371 4439 18427 4441
rect 11552 4323 11587 4439
tri 18349 4419 18369 4439 se
rect 18369 4419 18427 4439
rect 19964 4426 20016 4439
tri 18347 4417 18349 4419 se
rect 18349 4417 18427 4419
tri 11757 4411 11763 4417 se
rect 11763 4411 13817 4417
rect 11630 4359 11636 4411
rect 11688 4359 11700 4411
rect 11752 4371 13817 4411
rect 14713 4411 18164 4417
rect 14713 4377 14725 4411
rect 14759 4377 14797 4411
rect 14831 4377 18164 4411
rect 14713 4371 18164 4377
rect 18172 4371 18427 4417
rect 18457 4417 18587 4419
tri 18587 4417 18589 4419 sw
rect 18457 4411 19490 4417
rect 18457 4377 18469 4411
rect 18503 4377 18541 4411
rect 18575 4405 19490 4411
rect 18575 4377 19450 4405
rect 18457 4371 19450 4377
rect 19484 4371 19490 4405
rect 11752 4368 11767 4371
tri 11767 4368 11770 4371 nw
tri 13737 4368 13740 4371 ne
rect 13740 4368 13817 4371
tri 19410 4368 19413 4371 ne
rect 19413 4368 19490 4371
rect 11752 4359 11758 4368
tri 11758 4359 11767 4368 nw
tri 13740 4359 13749 4368 ne
rect 13749 4359 13817 4368
tri 19413 4359 19422 4368 ne
rect 19422 4359 19490 4368
tri 13749 4343 13765 4359 ne
rect 13765 4343 13817 4359
tri 19422 4343 19438 4359 ne
rect 19438 4343 19490 4359
tri 13765 4337 13771 4343 ne
tri 11587 4323 11601 4337 sw
rect 11552 4317 11841 4323
tri 11552 4311 11558 4317 ne
rect 11558 4311 11841 4317
tri 11558 4286 11583 4311 ne
rect 11583 4286 11801 4311
rect 11795 4277 11801 4286
rect 11835 4277 11841 4311
rect 11795 4239 11841 4277
rect 13771 4299 13817 4343
rect 13921 4337 19161 4343
tri 19438 4337 19444 4343 ne
rect 13921 4303 13933 4337
rect 13967 4303 14005 4337
rect 14039 4303 19043 4337
rect 19077 4303 19115 4337
rect 19149 4303 19161 4337
tri 13817 4299 13821 4303 sw
rect 13921 4299 19161 4303
rect 13771 4297 13821 4299
tri 13821 4297 13823 4299 sw
rect 13921 4297 14051 4299
tri 14051 4297 14053 4299 nw
tri 19028 4297 19030 4299 ne
rect 19030 4297 19161 4299
rect 13771 4296 13823 4297
tri 13823 4296 13824 4297 sw
tri 19030 4296 19031 4297 ne
rect 19031 4296 19161 4297
rect 19444 4333 19490 4343
rect 19444 4299 19450 4333
rect 19484 4299 19490 4333
rect 13771 4295 13824 4296
tri 13824 4295 13825 4296 sw
rect 13771 4287 13825 4295
tri 13825 4287 13833 4295 sw
rect 19444 4287 19490 4299
rect 19964 4368 19973 4374
rect 20007 4368 20016 4374
rect 19964 4361 20016 4368
rect 19964 4296 19973 4309
rect 20007 4296 20016 4309
rect 13771 4271 13833 4287
tri 13833 4271 13849 4287 sw
rect 13771 4269 13849 4271
tri 13849 4269 13851 4271 sw
rect 13771 4263 15228 4269
rect 11795 4205 11801 4239
rect 11835 4205 11841 4239
rect 13238 4211 13247 4263
rect 13299 4211 13311 4263
rect 13363 4211 13369 4263
rect 13771 4229 15110 4263
rect 15144 4229 15182 4263
rect 15216 4229 15228 4263
rect 13771 4223 15228 4229
rect 16456 4265 17790 4271
rect 16456 4231 16468 4265
rect 16502 4231 16540 4265
rect 16574 4231 17672 4265
rect 17706 4231 17744 4265
rect 17778 4231 17790 4265
rect 16456 4225 17790 4231
rect 19964 4231 19973 4244
rect 20007 4231 20016 4244
rect 11795 4193 11841 4205
rect 15517 4189 19769 4195
rect 10284 3051 11379 3053
rect 10284 3049 11377 3051
tri 11377 3049 11379 3051 nw
tri 11434 3049 11438 3053 se
rect 11438 3049 11490 3758
rect 11560 4160 11620 4172
rect 11560 4126 11580 4160
rect 11614 4126 11620 4160
rect 11560 4088 11620 4126
rect 12388 4157 12518 4163
rect 12388 4151 12400 4157
rect 12434 4151 12472 4157
rect 12506 4151 12518 4157
rect 12388 4099 12394 4151
rect 12446 4099 12460 4151
rect 12512 4099 12518 4151
rect 15517 4155 15529 4189
rect 15563 4155 15601 4189
rect 15635 4183 19769 4189
rect 15635 4157 19729 4183
rect 15635 4155 15647 4157
rect 15517 4149 15647 4155
tri 15647 4149 15655 4157 nw
tri 19689 4149 19697 4157 ne
rect 19697 4149 19729 4157
rect 19763 4149 19769 4183
tri 19697 4129 19717 4149 ne
rect 19717 4129 19769 4149
rect 11560 4054 11580 4088
rect 11614 4054 11620 4088
rect 13077 4068 13083 4120
rect 13135 4068 13147 4120
rect 13199 4114 15984 4120
rect 13199 4080 14089 4114
rect 14123 4080 14161 4114
rect 14195 4080 14890 4114
rect 14924 4080 14962 4114
rect 14996 4080 15721 4114
rect 15755 4080 15794 4114
rect 15828 4080 15866 4114
rect 15900 4080 15938 4114
rect 15972 4080 15984 4114
rect 13199 4074 15984 4080
rect 16305 4080 16316 4127
tri 16305 4075 16310 4080 ne
rect 16310 4075 16316 4080
rect 16368 4075 16380 4127
rect 16432 4075 16438 4127
rect 16837 4121 16889 4127
rect 16990 4125 16996 4129
rect 13199 4073 13210 4074
tri 13210 4073 13211 4074 nw
rect 13199 4068 13205 4073
tri 13205 4068 13210 4073 nw
rect 16931 4119 16996 4125
rect 17048 4119 17062 4129
rect 16931 4085 16943 4119
rect 16977 4085 16996 4119
rect 17049 4085 17062 4119
rect 16931 4079 16996 4085
rect 16990 4077 16996 4079
rect 17048 4077 17062 4085
rect 17114 4077 17120 4129
tri 19717 4127 19719 4129 ne
rect 19719 4127 19769 4129
tri 19719 4123 19723 4127 ne
rect 19723 4111 19769 4127
rect 18593 4099 19311 4105
rect 11560 4042 11620 4054
rect 11560 3498 11602 4042
tri 11602 4024 11620 4042 nw
rect 12436 4015 12442 4067
rect 12494 4015 12506 4067
rect 12558 4015 12566 4067
rect 12733 4056 12779 4068
rect 12733 4022 12739 4056
rect 12773 4022 12779 4056
rect 16837 4055 16889 4069
tri 12729 4015 12733 4019 se
rect 12733 4015 12779 4022
tri 12779 4015 12786 4022 sw
tri 12723 4009 12729 4015 se
rect 12729 4009 12786 4015
tri 12786 4009 12792 4015 sw
rect 17675 4062 17727 4068
tri 17673 4024 17675 4026 se
tri 16953 4018 16959 4024 se
rect 16959 4018 17438 4024
tri 17438 4018 17444 4024 sw
tri 17667 4018 17673 4024 se
rect 17673 4018 17675 4024
tri 12721 4007 12723 4009 se
rect 12723 4007 12792 4009
tri 12792 4007 12794 4009 sw
tri 12717 4003 12721 4007 se
rect 12721 4003 12794 4007
tri 12794 4003 12798 4007 sw
tri 16938 4003 16953 4018 se
rect 16953 4013 17444 4018
tri 17444 4013 17449 4018 sw
tri 17662 4013 17667 4018 se
rect 17667 4013 17675 4018
rect 16953 4003 17449 4013
tri 17449 4003 17459 4013 sw
tri 17652 4003 17662 4013 se
rect 17662 4010 17675 4013
rect 17759 4030 17765 4082
rect 17817 4030 17839 4082
rect 17891 4030 17912 4082
rect 17964 4079 17970 4082
rect 17964 4073 17977 4079
rect 17965 4039 17977 4073
rect 18593 4065 18605 4099
rect 18639 4065 18677 4099
rect 18711 4098 19311 4099
rect 18711 4065 19259 4098
tri 18075 4056 18084 4065 ne
rect 18084 4056 18168 4065
tri 18168 4056 18177 4065 nw
rect 18593 4059 19259 4065
tri 19234 4056 19237 4059 ne
rect 19237 4056 19259 4059
rect 19723 4077 19729 4111
rect 19763 4077 19769 4111
rect 19723 4065 19769 4077
rect 19964 4166 19973 4179
rect 20007 4166 20016 4179
rect 19964 4110 20016 4114
rect 19964 4100 19973 4110
rect 20007 4100 20016 4110
rect 17964 4033 17977 4039
tri 18084 4037 18103 4056 ne
rect 18103 4037 18149 4056
tri 18149 4037 18168 4056 nw
tri 19237 4037 19256 4056 ne
rect 19256 4046 19259 4056
rect 19256 4037 19311 4046
tri 18103 4033 18107 4037 ne
rect 18107 4033 18143 4037
rect 17964 4030 17970 4033
tri 18107 4031 18109 4033 ne
rect 18109 4031 18143 4033
tri 18143 4031 18149 4037 nw
tri 19256 4034 19259 4037 ne
rect 19259 4034 19311 4037
rect 17662 4003 17727 4010
tri 12712 3998 12717 4003 se
rect 12717 3998 12798 4003
rect 11632 3994 11760 3998
rect 11632 3942 11638 3994
rect 11690 3942 11702 3994
rect 11754 3985 11760 3994
tri 11760 3985 11773 3998 sw
tri 12699 3985 12712 3998 se
rect 12712 3997 12798 3998
tri 12798 3997 12804 4003 sw
rect 16837 3997 16889 4003
tri 16932 3997 16938 4003 se
rect 16938 3997 17459 4003
tri 17459 3997 17465 4003 sw
tri 17646 3997 17652 4003 se
rect 17652 3998 17727 4003
rect 17652 3997 17675 3998
rect 12712 3985 12804 3997
rect 11754 3984 12804 3985
tri 12804 3984 12817 3997 sw
tri 16919 3984 16932 3997 se
rect 16932 3984 17465 3997
tri 17465 3984 17478 3997 sw
tri 17633 3984 17646 3997 se
rect 17646 3984 17675 3997
rect 11754 3950 12739 3984
rect 12773 3969 16512 3984
tri 16512 3969 16527 3984 sw
tri 16904 3969 16919 3984 se
rect 16919 3980 17675 3984
rect 16919 3969 17015 3980
tri 17015 3969 17026 3980 nw
tri 17208 3969 17219 3980 ne
rect 17219 3969 17675 3980
rect 12773 3965 16527 3969
tri 16527 3965 16531 3969 sw
tri 16900 3965 16904 3969 se
rect 16904 3965 17011 3969
tri 17011 3965 17015 3969 nw
tri 17219 3965 17223 3969 ne
rect 17223 3965 17675 3969
rect 12773 3964 17010 3965
tri 17010 3964 17011 3965 nw
tri 17223 3964 17224 3965 ne
rect 17224 3964 17675 3965
rect 12773 3961 17007 3964
tri 17007 3961 17010 3964 nw
tri 17224 3961 17227 3964 ne
rect 17227 3961 17675 3964
rect 12773 3955 17001 3961
tri 17001 3955 17007 3961 nw
tri 17227 3955 17233 3961 ne
rect 17233 3955 17675 3961
rect 12773 3950 16986 3955
rect 11754 3942 16986 3950
rect 11632 3940 16986 3942
tri 16986 3940 17001 3955 nw
tri 17233 3940 17248 3955 ne
rect 17248 3946 17675 3955
rect 18417 4003 18588 4013
rect 18417 3969 18429 4003
rect 18463 3969 18501 4003
rect 18535 3969 18588 4003
rect 18417 3961 18588 3969
rect 18640 3961 18652 4013
rect 18704 3961 18710 4013
rect 17248 3940 17727 3946
tri 19254 3940 19259 3945 se
rect 19259 3940 19311 3982
rect 11632 3939 12782 3940
tri 12782 3939 12783 3940 nw
tri 16475 3939 16476 3940 ne
rect 16476 3939 16984 3940
rect 11632 3938 11761 3939
tri 11761 3938 11762 3939 nw
tri 12727 3938 12728 3939 ne
rect 12728 3938 12781 3939
tri 12781 3938 12782 3939 nw
tri 16476 3938 16477 3939 ne
rect 16477 3938 16984 3939
tri 16984 3938 16986 3940 nw
tri 19252 3938 19254 3940 se
rect 19254 3938 19311 3940
tri 16477 3930 16485 3938 ne
rect 16485 3930 16976 3938
tri 16976 3930 16984 3938 nw
rect 17107 3932 17159 3938
tri 16485 3926 16489 3930 ne
rect 16489 3926 16972 3930
tri 16972 3926 16976 3930 nw
tri 19244 3930 19252 3938 se
rect 19252 3930 19311 3938
tri 16489 3921 16494 3926 ne
rect 16494 3921 16967 3926
tri 16967 3921 16972 3926 nw
rect 11777 3852 11783 3904
rect 11835 3852 11847 3904
rect 11899 3898 14416 3904
rect 11899 3864 14298 3898
rect 14332 3864 14370 3898
rect 14404 3864 14416 3898
rect 11899 3858 14416 3864
tri 19237 3923 19244 3930 se
rect 19244 3923 19311 3930
tri 19224 3910 19237 3923 se
rect 19237 3910 19298 3923
tri 19298 3910 19311 3923 nw
rect 19964 4037 20016 4048
rect 19964 4034 19973 4037
rect 20007 4034 20016 4037
rect 19964 3968 20016 3982
tri 19205 3891 19224 3910 se
rect 19224 3891 19279 3910
tri 19279 3891 19298 3910 nw
rect 19964 3902 20016 3916
tri 19202 3888 19205 3891 se
rect 19205 3888 19276 3891
tri 19276 3888 19279 3891 nw
rect 17107 3866 17159 3880
rect 11899 3857 11910 3858
tri 11910 3857 11911 3858 nw
rect 11899 3854 11907 3857
tri 11907 3854 11910 3857 nw
rect 11899 3852 11905 3854
tri 11905 3852 11907 3854 nw
rect 18760 3836 18766 3888
rect 18818 3836 18833 3888
rect 18885 3836 19009 3888
rect 19036 3857 19245 3888
tri 19245 3857 19276 3888 nw
rect 19036 3836 19224 3857
tri 19224 3836 19245 3857 nw
rect 19964 3836 20016 3850
rect 17107 3808 17159 3814
rect 19023 3771 19109 3773
rect 19023 3745 19088 3771
rect 18630 3719 19088 3745
rect 19140 3719 19165 3771
rect 19217 3719 19242 3771
rect 19294 3719 19300 3771
rect 18630 3701 19300 3719
rect 18630 3649 19088 3701
rect 19140 3649 19165 3701
rect 19217 3649 19242 3701
rect 19294 3649 19300 3701
rect 18630 3631 19300 3649
rect 18630 3590 19088 3631
rect 19023 3579 19088 3590
rect 19140 3579 19165 3631
rect 19217 3579 19242 3631
rect 19294 3579 19300 3631
rect 19964 3770 20016 3784
rect 19964 3711 19973 3718
rect 20007 3711 20016 3718
rect 19964 3704 20016 3711
rect 19964 3638 19973 3652
rect 20007 3638 20016 3652
rect 19023 3571 19109 3579
rect 19964 3572 19973 3586
rect 20007 3572 20016 3586
rect 11574 3412 11580 3464
rect 11632 3412 11644 3464
rect 11696 3412 13083 3464
rect 13135 3412 13147 3464
rect 13199 3412 13205 3464
rect 13241 3412 13247 3464
rect 13299 3412 13311 3464
rect 13363 3412 18767 3464
rect 18819 3412 18833 3464
rect 18885 3412 18891 3464
rect 19460 3431 19539 3510
rect 19964 3506 19973 3520
rect 20007 3506 20016 3520
rect 19964 3440 19973 3454
rect 20007 3440 20016 3454
tri 19939 3383 19964 3408 se
rect 19964 3383 20016 3388
rect 11553 3382 20016 3383
rect 11553 3377 17298 3382
rect 11553 3343 11565 3377
rect 11599 3343 11638 3377
rect 11672 3343 11711 3377
rect 11745 3343 11784 3377
rect 11818 3343 11857 3377
rect 11891 3343 11930 3377
rect 11964 3343 12003 3377
rect 12037 3343 12076 3377
rect 12110 3343 12149 3377
rect 12183 3343 12222 3377
rect 12256 3343 12295 3377
rect 12329 3343 12368 3377
rect 12402 3343 12441 3377
rect 12475 3343 12514 3377
rect 12548 3343 12587 3377
rect 12621 3343 12660 3377
rect 12694 3343 12733 3377
rect 12767 3343 12806 3377
rect 12840 3343 12879 3377
rect 12913 3343 12952 3377
rect 12986 3343 13025 3377
rect 13059 3343 13098 3377
rect 13132 3343 13171 3377
rect 13205 3343 13244 3377
rect 13278 3343 13317 3377
rect 13351 3343 13390 3377
rect 13424 3343 13463 3377
rect 13497 3343 13536 3377
rect 13570 3343 13609 3377
rect 13643 3343 13682 3377
rect 13716 3343 13755 3377
rect 13789 3343 13828 3377
rect 13862 3343 13901 3377
rect 13935 3343 13974 3377
rect 14008 3343 14047 3377
rect 14081 3343 14120 3377
rect 14154 3343 14193 3377
rect 14227 3343 14266 3377
rect 14300 3343 14339 3377
rect 14373 3343 14412 3377
rect 14446 3343 14485 3377
rect 14519 3343 14558 3377
rect 14592 3343 14631 3377
rect 14665 3343 14704 3377
rect 14738 3343 14777 3377
rect 14811 3343 14849 3377
rect 14883 3343 14921 3377
rect 14955 3343 14993 3377
rect 15027 3343 15065 3377
rect 15099 3343 15137 3377
rect 15171 3343 15209 3377
rect 15243 3343 15281 3377
rect 15315 3343 15353 3377
rect 15387 3343 15425 3377
rect 15459 3343 15497 3377
rect 15531 3343 15569 3377
rect 15603 3343 15641 3377
rect 15675 3343 15713 3377
rect 15747 3343 15785 3377
rect 15819 3343 15857 3377
rect 15891 3343 15929 3377
rect 15963 3343 16001 3377
rect 16035 3343 16073 3377
rect 16107 3343 16145 3377
rect 16179 3343 16217 3377
rect 16251 3343 16289 3377
rect 16323 3343 16361 3377
rect 16395 3343 16433 3377
rect 16467 3343 16505 3377
rect 16539 3343 16577 3377
rect 16611 3343 16649 3377
rect 16683 3343 16721 3377
rect 16755 3343 16793 3377
rect 16827 3343 16865 3377
rect 16899 3343 16937 3377
rect 16971 3343 17009 3377
rect 17043 3343 17081 3377
rect 17115 3343 17153 3377
rect 17187 3343 17225 3377
rect 17259 3343 17297 3377
rect 11553 3337 17298 3343
rect 17286 3336 17298 3337
tri 17286 3330 17292 3336 ne
rect 17292 3330 17298 3336
rect 17350 3330 17362 3382
rect 17414 3377 20016 3382
rect 17414 3343 17441 3377
rect 17475 3343 17513 3377
rect 17547 3343 17585 3377
rect 17619 3343 17657 3377
rect 17691 3343 17729 3377
rect 17763 3343 17801 3377
rect 17835 3343 17873 3377
rect 17907 3343 17945 3377
rect 17979 3343 18017 3377
rect 18051 3343 18089 3377
rect 18123 3343 18161 3377
rect 18195 3343 18233 3377
rect 18267 3343 18305 3377
rect 18339 3343 18377 3377
rect 18411 3343 18449 3377
rect 18483 3343 18521 3377
rect 18555 3343 18593 3377
rect 18627 3343 18665 3377
rect 18699 3343 18737 3377
rect 18771 3343 18809 3377
rect 18843 3343 18881 3377
rect 18915 3343 18953 3377
rect 18987 3343 19025 3377
rect 19059 3343 19097 3377
rect 19131 3343 19169 3377
rect 19203 3343 19241 3377
rect 19275 3343 19313 3377
rect 19347 3343 19385 3377
rect 19419 3343 19457 3377
rect 19491 3343 19529 3377
rect 19563 3343 19601 3377
rect 19635 3343 19673 3377
rect 19707 3343 19745 3377
rect 19779 3343 19817 3377
rect 19851 3343 19889 3377
rect 19923 3343 20016 3377
rect 17414 3337 20016 3343
rect 17414 3336 17427 3337
rect 17414 3330 17421 3336
tri 17421 3330 17427 3336 nw
rect 17920 3336 18972 3337
tri 17920 3330 17926 3336 ne
rect 17926 3330 18000 3336
tri 17926 3308 17948 3330 ne
rect 17948 3308 18000 3330
tri 18000 3308 18028 3336 nw
tri 18369 3308 18397 3336 ne
rect 18397 3308 18511 3336
tri 18511 3308 18539 3336 nw
tri 18864 3308 18892 3336 ne
rect 18892 3308 18944 3336
tri 18944 3308 18972 3336 nw
tri 19940 3310 19967 3337 ne
rect 17948 3305 17997 3308
tri 17997 3305 18000 3308 nw
tri 18397 3305 18400 3308 ne
rect 18400 3306 18509 3308
tri 18509 3306 18511 3308 nw
tri 18892 3306 18894 3308 ne
rect 18400 3305 18508 3306
tri 18508 3305 18509 3306 nw
rect 18894 3305 18940 3308
tri 11581 3275 11606 3300 se
rect 11606 3275 17765 3300
rect 10284 3047 11375 3049
tri 11375 3047 11377 3049 nw
tri 11432 3047 11434 3049 se
rect 11434 3047 11490 3049
tri 10259 3014 10284 3039 se
rect 10284 3014 10343 3047
rect 8845 2962 8851 3014
rect 8903 2962 8915 3014
rect 8967 3013 8973 3014
tri 8973 3013 8974 3014 sw
tri 10258 3013 10259 3014 se
rect 10259 3013 10343 3014
tri 10343 3013 10377 3047 nw
tri 11398 3013 11432 3047 se
rect 11432 3013 11490 3047
rect 8967 3008 8974 3013
tri 8974 3008 8979 3013 sw
tri 10253 3008 10258 3013 se
rect 10258 3008 10338 3013
tri 10338 3008 10343 3013 nw
tri 11393 3008 11398 3013 se
rect 11398 3008 11490 3013
rect 8967 3002 10337 3008
tri 10337 3007 10338 3008 nw
tri 11392 3007 11393 3008 se
rect 11393 3007 11490 3008
rect 8976 2968 9017 3002
rect 9051 2968 9092 3002
rect 9126 2968 9167 3002
rect 9201 2968 9242 3002
rect 9276 2968 9317 3002
rect 9351 2968 9392 3002
rect 9426 2968 9467 3002
rect 9501 2968 9542 3002
rect 9576 2968 9617 3002
rect 9651 2968 9692 3002
rect 9726 2968 9767 3002
rect 9801 2968 9842 3002
rect 9876 2968 9917 3002
rect 9951 2968 9992 3002
rect 10026 2968 10067 3002
rect 10101 2968 10142 3002
rect 10176 2968 10217 3002
rect 10251 2968 10291 3002
rect 10325 2968 10337 3002
tri 11383 2998 11392 3007 se
rect 11392 3006 11490 3007
rect 11392 2998 11482 3006
tri 11482 2998 11490 3006 nw
tri 11558 3252 11581 3275 se
rect 11581 3254 17765 3275
rect 11581 3252 16999 3254
tri 16999 3252 17001 3254 nw
tri 17603 3252 17605 3254 ne
rect 17605 3252 17765 3254
rect 11558 3248 16995 3252
tri 16995 3248 16999 3252 nw
tri 17605 3248 17609 3252 ne
rect 17609 3248 17765 3252
rect 17817 3248 17839 3300
rect 17891 3248 17897 3300
rect 17948 3275 17994 3305
tri 17994 3302 17997 3305 nw
tri 18400 3302 18403 3305 ne
rect 18403 3304 18507 3305
tri 18507 3304 18508 3305 nw
rect 18403 3302 18503 3304
tri 18403 3300 18405 3302 ne
rect 18405 3300 18503 3302
tri 18503 3300 18507 3304 nw
tri 18405 3275 18430 3300 ne
rect 18430 3275 18478 3300
tri 18478 3275 18503 3300 nw
rect 11558 3241 11637 3248
tri 11637 3241 11644 3248 nw
rect 17948 3241 17954 3275
rect 17988 3241 17994 3275
tri 18430 3273 18432 3275 ne
rect 11558 3233 11629 3241
tri 11629 3233 11637 3241 nw
rect 11558 3218 11614 3233
tri 11614 3218 11629 3233 nw
rect 11558 3216 11612 3218
tri 11612 3216 11614 3218 nw
tri 11678 3216 11680 3218 se
rect 11680 3216 16930 3218
tri 11380 2995 11383 2998 se
rect 11383 2995 11479 2998
tri 11479 2995 11482 2998 nw
tri 10410 2976 10429 2995 se
rect 10429 2976 11460 2995
tri 11460 2976 11479 2995 nw
rect 8967 2962 10337 2968
tri 10396 2962 10410 2976 se
rect 10410 2962 11433 2976
tri 10376 2942 10396 2962 se
rect 10396 2949 11433 2962
tri 11433 2949 11460 2976 nw
rect 10396 2942 10461 2949
tri 10461 2942 10468 2949 nw
tri 10360 2926 10376 2942 se
rect 10376 2926 10445 2942
tri 10445 2926 10461 2942 nw
tri 10352 2918 10360 2926 se
rect 10360 2918 10437 2926
tri 10437 2918 10445 2926 nw
rect 9189 2866 9195 2918
rect 9247 2866 9259 2918
rect 9311 2892 10411 2918
tri 10411 2892 10437 2918 nw
rect 9311 2883 10402 2892
tri 10402 2883 10411 2892 nw
rect 9311 2868 10387 2883
tri 10387 2868 10402 2883 nw
rect 9311 2866 10385 2868
tri 10385 2866 10387 2868 nw
tri 10767 2866 10769 2868 se
rect 10769 2866 10775 2868
tri 10763 2862 10767 2866 se
rect 10767 2862 10775 2866
rect 10476 2856 10775 2862
rect 10827 2856 10839 2868
rect 10891 2862 10897 2868
tri 10897 2862 10903 2868 sw
rect 10891 2856 11325 2862
rect 10476 2822 10488 2856
rect 10522 2822 10568 2856
rect 10602 2822 10647 2856
rect 10681 2822 10726 2856
rect 10760 2822 10775 2856
rect 10918 2822 10963 2856
rect 10997 2822 11042 2856
rect 11076 2822 11121 2856
rect 11155 2822 11200 2856
rect 11234 2822 11279 2856
rect 11313 2822 11325 2856
rect 10476 2816 10775 2822
rect 10827 2816 10839 2822
rect 10891 2816 11325 2822
rect 11477 2780 11529 2786
tri 11463 2710 11477 2724 se
rect 11477 2716 11529 2728
rect 8862 2658 8868 2710
rect 8920 2658 8932 2710
rect 8984 2703 8990 2710
tri 8990 2703 8997 2710 sw
tri 11456 2703 11463 2710 se
rect 11463 2703 11477 2710
rect 8984 2690 8997 2703
tri 8997 2690 9010 2703 sw
tri 11443 2690 11456 2703 se
rect 11456 2690 11477 2703
rect 8984 2664 11477 2690
rect 8984 2658 11529 2664
rect 8856 2578 8865 2630
rect 8917 2578 8929 2630
rect 8981 2578 10098 2630
rect 10150 2578 10206 2630
rect 10258 2578 10314 2630
rect 10366 2578 10372 2630
rect 10596 2578 10602 2630
rect 10654 2578 10673 2630
rect 10725 2578 10731 2630
tri 11553 2579 11558 2584 se
rect 11558 2579 11610 3216
tri 11610 3214 11612 3216 nw
tri 11676 3214 11678 3216 se
rect 11678 3214 16930 3216
tri 11644 3182 11676 3214 se
rect 11676 3182 16930 3214
tri 11552 2578 11553 2579 se
rect 11553 2578 11610 2579
tri 11531 2557 11552 2578 se
rect 11552 2557 11610 2578
tri 11524 2550 11531 2557 se
rect 11531 2550 11610 2557
tri 8802 2524 8828 2550 se
rect 8828 2536 11610 2550
rect 8828 2524 11597 2536
tri 8801 2523 8802 2524 se
rect 8802 2523 11597 2524
tri 11597 2523 11610 2536 nw
tri 11639 3177 11644 3182 se
rect 11644 3177 16930 3182
rect 11639 3166 16930 3177
rect 16982 3166 16994 3218
rect 17046 3166 17052 3218
rect 17092 3216 17298 3222
rect 17350 3216 17362 3222
rect 17414 3216 17571 3222
rect 17092 3182 17104 3216
rect 17138 3182 17189 3216
rect 17223 3182 17273 3216
rect 17350 3182 17357 3216
rect 17414 3182 17441 3216
rect 17475 3182 17525 3216
rect 17559 3182 17571 3216
rect 17092 3170 17298 3182
rect 17350 3170 17362 3182
rect 17414 3170 17571 3182
rect 17613 3202 17659 3214
rect 17613 3168 17619 3202
rect 17653 3168 17659 3202
rect 17948 3203 17994 3241
tri 17739 3187 17742 3190 se
rect 17742 3187 17838 3190
tri 17730 3178 17739 3187 se
rect 17739 3178 17838 3187
rect 11639 3144 11703 3166
tri 11703 3144 11725 3166 nw
rect 11639 3136 11695 3144
tri 11695 3136 11703 3144 nw
rect 4463 1553 4515 1568
rect 6735 1616 6801 1622
tri 6801 1616 6807 1622 sw
tri 8696 1616 8702 1622 se
rect 8702 1616 8761 1622
rect 6735 1610 6807 1616
tri 6807 1610 6813 1616 sw
tri 7507 1610 7513 1616 se
rect 7513 1610 8301 1616
tri 8301 1610 8307 1616 sw
tri 8690 1610 8696 1616 se
rect 8696 1610 8761 1616
rect 6735 1609 6813 1610
tri 6813 1609 6814 1610 sw
tri 7506 1609 7507 1610 se
rect 7507 1609 8307 1610
tri 8307 1609 8308 1610 sw
tri 8689 1609 8690 1610 se
rect 8690 1609 8761 1610
rect 6735 1590 8761 1609
rect 6735 1570 8741 1590
tri 8741 1570 8761 1590 nw
tri 8790 2512 8801 2523 se
rect 8801 2512 11586 2523
tri 11586 2512 11597 2523 nw
rect 8790 2507 11581 2512
tri 11581 2507 11586 2512 nw
rect 8790 2498 11572 2507
tri 11572 2498 11581 2507 nw
tri 11635 2498 11639 2502 se
rect 11639 2498 11691 3136
tri 11691 3132 11695 3136 nw
tri 11758 3132 11762 3136 se
rect 11762 3132 15831 3136
tri 11756 3130 11758 3132 se
rect 11758 3130 15831 3132
tri 11722 3096 11756 3130 se
rect 11756 3096 15831 3130
rect 8790 2484 8862 2498
tri 8862 2484 8876 2498 nw
tri 11621 2484 11635 2498 se
rect 11635 2484 11691 2498
rect 8790 2468 8846 2484
tri 8846 2468 8862 2484 nw
tri 11605 2468 11621 2484 se
rect 11621 2468 11691 2484
rect 6735 1563 7559 1570
tri 7559 1563 7566 1570 nw
tri 8248 1563 8255 1570 ne
rect 8255 1563 8734 1570
tri 8734 1563 8741 1570 nw
tri 8787 1558 8790 1561 se
rect 8790 1558 8842 2468
tri 8842 2464 8846 2468 nw
tri 8899 2464 8903 2468 se
rect 8903 2464 11691 2468
tri 8885 2450 8899 2464 se
rect 8899 2456 11691 2464
rect 8899 2450 11685 2456
tri 11685 2450 11691 2456 nw
tri 11720 3094 11722 3096 se
rect 11722 3094 15831 3096
rect 11720 3084 15831 3094
rect 15883 3084 15895 3136
rect 15947 3084 16316 3136
rect 16368 3084 16380 3136
rect 16432 3084 16438 3136
rect 17613 3134 17659 3168
tri 17712 3160 17730 3178 se
rect 17730 3160 17798 3178
tri 17711 3159 17712 3160 se
rect 17712 3159 17798 3160
rect 17711 3144 17798 3159
rect 17832 3144 17838 3178
rect 17948 3169 17954 3203
rect 17988 3169 17994 3203
rect 17948 3157 17994 3169
rect 18432 3208 18478 3275
rect 18432 3174 18438 3208
rect 18472 3174 18478 3208
rect 18894 3271 18900 3305
rect 18934 3271 18940 3305
tri 18940 3304 18944 3308 nw
rect 18894 3233 18940 3271
rect 19967 3294 20016 3337
tri 20016 3294 20042 3320 sw
rect 18894 3199 18900 3233
rect 18934 3199 18940 3233
tri 19941 3222 19967 3248 se
rect 19967 3222 20042 3294
tri 19935 3216 19941 3222 se
rect 19941 3216 20042 3222
tri 19933 3214 19935 3216 se
rect 19935 3214 20002 3216
tri 19920 3201 19933 3214 se
rect 19933 3201 20002 3214
rect 18894 3187 18940 3199
rect 17613 3130 17665 3134
rect 17451 3123 17503 3129
rect 11720 3072 11794 3084
tri 11794 3072 11806 3084 nw
rect 11720 3054 11776 3072
tri 11776 3054 11794 3072 nw
rect 17451 3059 17503 3071
tri 8785 1556 8787 1558 se
rect 8787 1556 8842 1558
tri 8771 1542 8785 1556 se
rect 8785 1542 8842 1556
tri 7898 1535 7905 1542 se
rect 7905 1535 8227 1542
tri 8227 1535 8234 1542 sw
tri 8764 1535 8771 1542 se
rect 8771 1535 8842 1542
rect 4463 1495 4515 1501
rect 6740 1532 8842 1535
rect 6740 1514 8824 1532
tri 8824 1514 8842 1532 nw
tri 8871 2436 8885 2450 se
rect 8885 2436 11671 2450
tri 11671 2436 11685 2450 nw
rect 8871 2435 11670 2436
tri 11670 2435 11671 2436 nw
rect 8871 2420 11655 2435
tri 11655 2420 11670 2435 nw
rect 8871 2416 11651 2420
tri 11651 2416 11655 2420 nw
tri 11716 2416 11720 2420 se
rect 11720 2416 11772 3054
tri 11772 3050 11776 3054 nw
tri 11837 3050 11841 3054 se
rect 11841 3050 17037 3054
tri 11834 3047 11837 3050 se
rect 11837 3047 17037 3050
rect 8871 2411 8952 2416
tri 8952 2411 8957 2416 nw
tri 11711 2411 11716 2416 se
rect 11716 2411 11772 2416
rect 8871 2386 8927 2411
tri 8927 2386 8952 2411 nw
tri 11686 2386 11711 2411 se
rect 11711 2386 11772 2411
rect 6740 1513 7939 1514
tri 7939 1513 7940 1514 nw
tri 8192 1513 8193 1514 ne
rect 8193 1513 8823 1514
tri 8823 1513 8824 1514 nw
rect 6740 1507 7933 1513
tri 7933 1507 7939 1513 nw
tri 8193 1507 8199 1513 ne
rect 8199 1507 8817 1513
tri 8817 1507 8823 1513 nw
rect 6740 1479 6790 1507
tri 6790 1479 6818 1507 nw
tri 8855 1479 8871 1495 se
rect 8871 1479 8923 2386
tri 8923 2382 8927 2386 nw
tri 8981 2382 8985 2386 se
rect 8985 2382 11772 2386
tri 8976 2377 8981 2382 se
rect 8981 2377 11772 2382
tri 8962 2363 8976 2377 se
rect 8976 2374 11772 2377
rect 8976 2363 11761 2374
tri 11761 2363 11772 2374 nw
tri 11802 3015 11834 3047 se
rect 11834 3015 17037 3047
rect 11802 3002 17037 3015
rect 17089 3002 17101 3054
rect 17153 3002 17159 3054
rect 17195 3047 17451 3053
rect 17195 3013 17207 3047
rect 17241 3013 17291 3047
rect 17325 3013 17374 3047
rect 17408 3013 17451 3047
rect 17195 3007 17451 3013
rect 11802 2998 11884 3002
tri 11884 2998 11888 3002 nw
rect 17195 3001 17503 3007
rect 17613 3128 17619 3130
rect 17653 3128 17665 3130
rect 17613 3064 17665 3076
rect 17613 3006 17665 3012
rect 17711 3106 17838 3144
rect 17711 3072 17798 3106
rect 17832 3072 17838 3106
rect 17711 3060 17838 3072
rect 18104 3154 18156 3160
rect 18104 3088 18156 3102
rect 17711 3054 17776 3060
tri 17776 3054 17782 3060 nw
rect 17711 3042 17764 3054
tri 17764 3042 17776 3054 nw
rect 11802 2976 11862 2998
tri 11862 2976 11884 2998 nw
tri 17703 2982 17711 2990 se
rect 17711 2982 17757 3042
tri 17757 3035 17764 3042 nw
rect 18104 3030 18156 3036
rect 18273 3154 18325 3160
rect 18273 3088 18325 3102
rect 18273 3030 18325 3036
rect 18432 3136 18478 3174
rect 19996 3182 20002 3201
rect 20036 3182 20042 3216
tri 20042 3201 20087 3246 sw
rect 18432 3102 18438 3136
rect 18472 3102 18478 3136
rect 18432 3064 18478 3102
rect 18432 3030 18438 3064
rect 18472 3030 18478 3064
rect 18583 3154 18635 3160
rect 18583 3088 18635 3102
rect 18583 3030 18635 3036
rect 18733 3154 18785 3160
rect 19050 3159 19096 3160
rect 18733 3088 18785 3102
rect 18733 3030 18785 3036
rect 18821 3153 19096 3159
rect 18873 3148 19096 3153
rect 18873 3114 19056 3148
rect 19090 3114 19096 3148
rect 18873 3101 19096 3114
rect 18821 3091 19096 3101
rect 18821 3087 18897 3091
rect 18873 3076 18897 3087
tri 18897 3076 18912 3091 nw
tri 19022 3076 19037 3091 ne
rect 19037 3076 19096 3091
tri 18873 3052 18897 3076 nw
tri 19037 3063 19050 3076 ne
rect 18432 3018 18478 3030
rect 18821 3029 18873 3035
rect 19050 3042 19056 3076
rect 19090 3042 19096 3076
rect 19050 3030 19096 3042
rect 19996 3143 20042 3182
rect 19996 3109 20002 3143
rect 20036 3109 20042 3143
rect 19996 3070 20042 3109
rect 19996 3036 20002 3070
rect 20036 3036 20042 3070
rect 19996 2998 20042 3036
tri 19947 2982 19963 2998 ne
rect 19963 2982 20002 2998
tri 17697 2976 17703 2982 se
rect 17703 2976 17757 2982
rect 2408 1429 2422 1439
rect 2474 1429 2493 1439
rect 2408 1395 2420 1429
rect 2474 1395 2492 1429
rect 2408 1387 2422 1395
rect 2474 1387 2493 1395
rect 2545 1387 2564 1439
rect 2616 1387 2634 1439
rect 2686 1435 2692 1439
tri 2692 1435 2696 1439 sw
tri 3859 1435 3863 1439 se
rect 3863 1435 3869 1439
rect 2686 1429 3869 1435
rect 3921 1429 3940 1439
rect 3992 1429 4011 1439
rect 4063 1429 4081 1439
rect 4133 1435 4139 1439
tri 4139 1435 4143 1439 sw
rect 4133 1429 6678 1435
rect 2686 1395 2708 1429
rect 2742 1395 2780 1429
rect 2814 1395 2852 1429
rect 2886 1395 2924 1429
rect 2958 1395 2996 1429
rect 3030 1395 3068 1429
rect 3102 1395 3140 1429
rect 3174 1395 3212 1429
rect 3246 1395 3284 1429
rect 3318 1395 3356 1429
rect 3390 1395 3428 1429
rect 3462 1395 3500 1429
rect 3534 1395 3572 1429
rect 3606 1395 3644 1429
rect 3678 1395 3716 1429
rect 3750 1395 3788 1429
rect 3822 1395 3860 1429
rect 3921 1395 3932 1429
rect 3992 1395 4004 1429
rect 4063 1395 4076 1429
rect 4133 1395 4148 1429
rect 4182 1395 4220 1429
rect 4254 1395 4292 1429
rect 4326 1395 4364 1429
rect 4398 1395 4688 1429
rect 4722 1395 4760 1429
rect 4794 1395 4832 1429
rect 4866 1395 4904 1429
rect 4938 1395 4976 1429
rect 5010 1395 5048 1429
rect 5082 1395 5120 1429
rect 5154 1395 5192 1429
rect 5226 1395 5264 1429
rect 5298 1395 5336 1429
rect 5370 1395 5408 1429
rect 5442 1395 5480 1429
rect 5514 1395 5552 1429
rect 5586 1395 5624 1429
rect 5658 1395 5696 1429
rect 5730 1395 5768 1429
rect 5802 1395 5840 1429
rect 5874 1395 5912 1429
rect 5946 1395 5984 1429
rect 6018 1395 6056 1429
rect 6090 1395 6128 1429
rect 6162 1395 6200 1429
rect 6234 1395 6272 1429
rect 6306 1395 6344 1429
rect 6378 1395 6416 1429
rect 6450 1395 6488 1429
rect 6522 1395 6560 1429
rect 6594 1395 6632 1429
rect 6666 1395 6678 1429
rect 2686 1389 3869 1395
rect 2686 1387 2694 1389
tri 2694 1387 2696 1389 nw
tri 3860 1387 3862 1389 ne
rect 3862 1387 3869 1389
rect 3921 1387 3940 1395
rect 3992 1387 4011 1395
rect 4063 1387 4081 1395
rect 4133 1389 6678 1395
rect 4133 1387 4140 1389
tri 4140 1387 4142 1389 nw
rect 4467 1355 4604 1361
tri 6734 1355 6740 1361 se
rect 6740 1355 6785 1479
tri 6785 1474 6790 1479 nw
rect 7325 1473 7827 1479
rect 7325 1439 7511 1473
rect 7545 1439 7601 1473
rect 7635 1439 7691 1473
rect 7725 1439 7781 1473
rect 7815 1439 7827 1473
tri 8845 1469 8855 1479 se
rect 8855 1469 8923 1479
tri 7961 1456 7974 1469 se
rect 7974 1456 8923 1469
rect 4520 1321 4558 1355
rect 4592 1321 4604 1355
rect 4519 1303 4604 1321
rect 4467 1291 4604 1303
rect 4519 1273 4604 1291
rect 4520 1239 4558 1273
rect 4592 1239 4604 1273
rect 4467 1233 4604 1239
rect 6204 1349 6256 1355
tri 6256 1328 6283 1355 sw
tri 6707 1328 6734 1355 se
rect 6734 1328 6785 1355
rect 7141 1433 7260 1439
rect 7141 1381 7142 1433
rect 7194 1381 7208 1433
rect 7141 1364 7260 1381
rect 6256 1297 6785 1328
rect 6204 1285 6785 1297
rect 6256 1246 6785 1285
rect 6996 1323 7048 1329
rect 6996 1259 7048 1271
rect 6256 1245 6274 1246
tri 6274 1245 6275 1246 nw
rect 6204 1227 6256 1233
tri 6256 1227 6274 1245 nw
tri 6799 1202 6802 1205 se
rect 6802 1202 6808 1205
tri 3034 1199 3037 1202 se
rect 3037 1199 3044 1202
rect 2408 1193 3044 1199
rect 3096 1193 3115 1202
rect 3167 1193 3186 1202
rect 3238 1193 3256 1202
rect 3308 1199 3322 1202
tri 3322 1199 3325 1202 sw
tri 6796 1199 6799 1202 se
rect 6799 1199 6808 1202
rect 3308 1193 6808 1199
rect 2408 1159 2420 1193
rect 2454 1159 2492 1193
rect 2526 1159 2564 1193
rect 2598 1159 2636 1193
rect 2670 1159 2708 1193
rect 2742 1159 2780 1193
rect 2814 1159 2852 1193
rect 2886 1159 2924 1193
rect 2958 1159 2996 1193
rect 3030 1159 3044 1193
rect 3102 1159 3115 1193
rect 3174 1159 3186 1193
rect 3246 1159 3256 1193
rect 3318 1159 3356 1193
rect 3390 1159 3428 1193
rect 3462 1159 3500 1193
rect 3534 1159 3572 1193
rect 3606 1159 3644 1193
rect 3678 1159 3716 1193
rect 3750 1159 3788 1193
rect 3822 1159 3860 1193
rect 3894 1159 3932 1193
rect 3966 1159 4004 1193
rect 4038 1159 4076 1193
rect 4110 1159 4148 1193
rect 4182 1159 4220 1193
rect 4254 1159 4292 1193
rect 4326 1159 4364 1193
rect 4398 1159 4688 1193
rect 4722 1159 4760 1193
rect 4794 1159 4832 1193
rect 4866 1159 4904 1193
rect 4938 1159 4976 1193
rect 5010 1159 5048 1193
rect 5082 1159 5120 1193
rect 5154 1159 5192 1193
rect 5226 1159 5264 1193
rect 5298 1159 5336 1193
rect 5370 1159 5408 1193
rect 5442 1159 5480 1193
rect 5514 1159 5552 1193
rect 5586 1159 5624 1193
rect 5658 1159 5696 1193
rect 5730 1159 5768 1193
rect 5802 1159 5840 1193
rect 5874 1159 5912 1193
rect 5946 1159 5984 1193
rect 6018 1159 6056 1193
rect 6090 1159 6128 1193
rect 6162 1159 6200 1193
rect 6234 1159 6272 1193
rect 6306 1159 6344 1193
rect 6378 1159 6416 1193
rect 6450 1159 6488 1193
rect 6522 1159 6560 1193
rect 6594 1159 6632 1193
rect 6666 1159 6808 1193
rect 2408 1153 3044 1159
tri 3033 1150 3036 1153 ne
rect 3036 1150 3044 1153
rect 3096 1150 3115 1159
rect 3167 1150 3186 1159
rect 3238 1150 3256 1159
rect 3308 1153 6808 1159
rect 6860 1153 6872 1205
rect 6924 1153 6930 1205
rect 6996 1200 7048 1207
tri 6996 1194 7002 1200 ne
rect 3308 1150 3322 1153
tri 3322 1150 3325 1153 nw
tri 5726 1118 5733 1125 se
rect 5733 1118 5739 1125
tri 3858 1114 3861 1117 se
rect 3861 1114 3867 1117
tri 3848 1104 3858 1114 se
rect 3858 1104 3867 1114
rect 2454 1098 3007 1104
rect 2454 1064 2466 1098
rect 2500 1064 2549 1098
rect 2583 1064 2632 1098
rect 2666 1064 2715 1098
rect 2749 1064 2797 1098
rect 2831 1064 2879 1098
rect 2913 1064 2961 1098
rect 2995 1064 3007 1098
rect 2454 1058 3007 1064
rect 3082 1098 3633 1104
rect 3082 1064 3094 1098
rect 3128 1064 3177 1098
rect 3211 1064 3259 1098
rect 3293 1064 3341 1098
rect 3375 1064 3423 1098
rect 3457 1064 3505 1098
rect 3539 1064 3587 1098
rect 3621 1064 3633 1098
rect 3082 1058 3633 1064
rect 3830 1098 3867 1104
rect 3830 1064 3842 1098
rect 3919 1065 3931 1117
rect 3983 1114 3989 1117
tri 3989 1114 3992 1117 sw
rect 3983 1104 3992 1114
tri 3992 1104 4002 1114 sw
rect 3983 1098 4069 1104
rect 3983 1065 4023 1098
rect 3876 1064 3933 1065
rect 3967 1064 4023 1065
rect 4057 1064 4069 1098
rect 3830 1058 4069 1064
tri 2596 1056 2598 1058 ne
rect 2598 1056 2713 1058
tri 2713 1056 2715 1058 nw
tri 3223 1056 3225 1058 ne
rect 3225 1056 3337 1058
tri 3337 1056 3339 1058 nw
tri 3830 1056 3832 1058 ne
rect 3832 1056 3920 1058
tri 3920 1056 3922 1058 nw
tri 3980 1056 3982 1058 ne
rect 3982 1057 4068 1058
tri 4068 1057 4069 1058 nw
rect 4135 1097 5479 1103
rect 4135 1063 4147 1097
rect 4181 1063 4252 1097
rect 4286 1063 4357 1097
rect 4391 1063 4603 1097
rect 4637 1063 4677 1097
rect 4711 1063 4751 1097
rect 4785 1063 4825 1097
rect 4859 1063 5071 1097
rect 5105 1063 5144 1097
rect 5178 1063 5217 1097
rect 5251 1063 5289 1097
rect 5323 1063 5361 1097
rect 5395 1063 5433 1097
rect 5467 1063 5479 1097
rect 5512 1066 5518 1118
rect 5570 1066 5582 1118
rect 5634 1066 5640 1118
tri 5722 1114 5726 1118 se
rect 5726 1114 5739 1118
tri 5531 1064 5533 1066 ne
rect 5533 1064 5640 1066
rect 4135 1057 5479 1063
tri 5533 1062 5535 1064 ne
rect 5535 1062 5640 1064
tri 5535 1058 5539 1062 ne
rect 5539 1058 5640 1062
tri 5718 1110 5722 1114 se
rect 5722 1110 5739 1114
rect 5718 1098 5739 1110
rect 5718 1064 5730 1098
rect 5791 1073 5803 1125
rect 5855 1123 5866 1125
tri 5866 1123 5868 1125 sw
rect 5855 1114 5868 1123
tri 5868 1114 5877 1123 sw
rect 5855 1104 5877 1114
tri 5877 1104 5887 1114 sw
rect 5855 1098 5930 1104
rect 5855 1073 5884 1098
rect 5764 1064 5807 1073
rect 5841 1064 5884 1073
rect 5918 1064 5930 1098
rect 6048 1071 6054 1123
rect 6106 1071 6118 1123
rect 6170 1071 6176 1123
tri 6100 1064 6107 1071 ne
rect 6107 1064 6176 1071
rect 5718 1058 5930 1064
tri 6107 1062 6109 1064 ne
rect 6109 1062 6176 1064
tri 6109 1058 6113 1062 ne
rect 6113 1058 6176 1062
tri 5539 1057 5540 1058 ne
rect 5540 1057 5640 1058
rect 3982 1056 4067 1057
tri 4067 1056 4068 1057 nw
tri 4212 1056 4213 1057 ne
rect 4213 1056 4313 1057
tri 4313 1056 4314 1057 nw
tri 5148 1056 5149 1057 ne
rect 5149 1056 5249 1057
tri 5249 1056 5250 1057 nw
tri 5540 1056 5541 1057 ne
rect 5541 1056 5640 1057
tri 6113 1056 6115 1058 ne
rect 6115 1056 6176 1058
tri 2598 1042 2612 1056 ne
rect 2612 1042 2699 1056
tri 2699 1042 2713 1056 nw
tri 3225 1042 3239 1056 ne
rect 3239 1042 3323 1056
tri 3323 1042 3337 1056 nw
tri 3832 1042 3846 1056 ne
rect 3846 1042 3906 1056
tri 3906 1042 3920 1056 nw
tri 3982 1042 3996 1056 ne
rect 3996 1042 4053 1056
tri 4053 1042 4067 1056 nw
tri 4213 1042 4227 1056 ne
rect 4227 1042 4299 1056
tri 4299 1042 4313 1056 nw
tri 5149 1042 5163 1056 ne
rect 5163 1042 5235 1056
tri 5235 1042 5249 1056 nw
tri 5541 1042 5555 1056 ne
rect 5555 1051 5640 1056
rect 5555 1042 5631 1051
tri 5631 1042 5640 1051 nw
tri 6115 1042 6129 1056 ne
rect 6129 1042 6176 1056
tri 2612 1033 2621 1042 ne
rect 2621 1033 2690 1042
tri 2690 1033 2699 1042 nw
tri 3239 1033 3248 1042 ne
rect 3248 1033 3314 1042
tri 3314 1033 3323 1042 nw
tri 3846 1039 3849 1042 ne
tri 2621 1029 2625 1033 ne
rect 2625 1029 2686 1033
tri 2686 1029 2690 1033 nw
tri 3248 1029 3252 1033 ne
rect 3252 1029 3310 1033
tri 3310 1029 3314 1033 nw
tri 2625 1024 2630 1029 ne
rect 2400 982 2446 994
rect 2400 948 2406 982
rect 2440 948 2446 982
rect 2400 910 2446 948
rect 2400 876 2406 910
rect 2440 876 2446 910
rect 2400 838 2446 876
rect 2400 804 2406 838
rect 2440 804 2446 838
rect 2400 766 2446 804
rect 2400 732 2406 766
rect 2440 732 2446 766
rect 2400 694 2446 732
rect 2400 660 2406 694
rect 2440 660 2446 694
rect 2400 622 2446 660
rect 2400 588 2406 622
rect 2440 588 2446 622
rect 2400 550 2446 588
tri 2372 516 2400 544 se
rect 2400 516 2406 550
rect 2440 544 2446 550
rect 2556 982 2602 994
rect 2556 948 2562 982
rect 2596 948 2602 982
rect 2556 910 2602 948
rect 2556 876 2562 910
rect 2596 876 2602 910
rect 2556 838 2602 876
rect 2556 804 2562 838
rect 2596 804 2602 838
rect 2556 766 2602 804
rect 2556 732 2562 766
rect 2596 732 2602 766
rect 2556 694 2602 732
rect 2556 660 2562 694
rect 2596 660 2602 694
rect 2556 622 2602 660
rect 2556 588 2562 622
rect 2596 588 2602 622
rect 2556 550 2602 588
tri 2446 544 2451 549 sw
rect 2440 516 2451 544
tri 2451 516 2479 544 sw
rect 2556 516 2562 550
rect 2596 516 2602 550
tri 2371 515 2372 516 se
rect 2372 515 2479 516
tri 2479 515 2480 516 sw
rect 2371 463 2377 515
rect 2429 478 2441 515
rect 2440 463 2441 478
rect 2493 463 2499 515
rect 2556 478 2602 516
tri 2371 444 2390 463 ne
rect 2390 444 2406 463
rect 2440 444 2461 463
tri 2461 444 2480 463 nw
rect 2556 444 2562 478
rect 2596 444 2602 478
tri 2390 434 2400 444 ne
rect 2400 434 2451 444
tri 2451 434 2461 444 nw
rect 2400 406 2446 434
tri 2446 429 2451 434 nw
rect 2400 372 2406 406
rect 2440 372 2446 406
rect 2400 334 2446 372
rect 2400 300 2406 334
rect 2440 300 2446 334
rect 2400 262 2446 300
rect 2400 228 2406 262
rect 2440 228 2446 262
rect 2400 190 2446 228
rect 2400 156 2406 190
rect 2440 156 2446 190
rect 2556 406 2602 444
rect 2556 372 2562 406
rect 2596 372 2602 406
rect 2556 334 2602 372
rect 2556 300 2562 334
rect 2596 300 2602 334
rect 2556 262 2602 300
rect 2556 228 2562 262
rect 2596 228 2602 262
rect 2556 190 2602 228
rect 2630 318 2681 1029
tri 2681 1024 2686 1029 nw
tri 3252 1024 3257 1029 ne
rect 2712 982 2758 994
rect 2712 948 2718 982
rect 2752 948 2758 982
rect 2712 910 2758 948
rect 2712 876 2718 910
rect 2752 876 2758 910
rect 2712 838 2758 876
rect 2712 804 2718 838
rect 2752 804 2758 838
rect 2712 766 2758 804
rect 2712 732 2718 766
rect 2752 732 2758 766
rect 2712 694 2758 732
rect 2712 660 2718 694
rect 2752 660 2758 694
rect 2712 622 2758 660
rect 2712 588 2718 622
rect 2752 588 2758 622
rect 2712 550 2758 588
rect 2712 516 2718 550
rect 2752 516 2758 550
rect 2868 982 2914 994
rect 2868 948 2874 982
rect 2908 948 2914 982
rect 2868 910 2914 948
rect 2868 876 2874 910
rect 2908 876 2914 910
rect 2868 838 2914 876
rect 2868 804 2874 838
rect 2908 804 2914 838
rect 2868 766 2914 804
rect 2868 732 2874 766
rect 2908 732 2914 766
rect 2868 694 2914 732
rect 2868 660 2874 694
rect 2908 660 2914 694
rect 2868 622 2914 660
rect 2868 588 2874 622
rect 2908 588 2914 622
rect 2868 550 2914 588
tri 2758 516 2791 549 sw
rect 2868 516 2874 550
rect 2908 516 2914 550
rect 3024 982 3070 994
rect 3024 948 3030 982
rect 3064 948 3070 982
rect 3024 910 3070 948
rect 3024 876 3030 910
rect 3064 876 3070 910
rect 3024 838 3070 876
rect 3024 804 3030 838
rect 3064 804 3070 838
rect 3024 766 3070 804
rect 3024 732 3030 766
rect 3064 732 3070 766
rect 3024 694 3070 732
rect 3024 660 3030 694
rect 3064 660 3070 694
rect 3180 982 3226 994
rect 3180 948 3186 982
rect 3220 948 3226 982
rect 3180 910 3226 948
rect 3180 876 3186 910
rect 3220 876 3226 910
rect 3180 838 3226 876
rect 3180 804 3186 838
rect 3220 804 3226 838
rect 3180 766 3226 804
rect 3180 732 3186 766
rect 3220 732 3226 766
rect 3180 694 3226 732
rect 3024 622 3070 660
rect 3024 588 3030 622
rect 3064 588 3070 622
rect 3024 550 3070 588
tri 2991 516 3024 549 se
rect 3024 516 3030 550
rect 3064 543 3070 550
tri 3177 674 3180 677 se
rect 3180 674 3186 694
rect 3177 668 3186 674
rect 3220 674 3226 694
tri 3226 674 3229 677 sw
rect 3220 668 3229 674
rect 3177 604 3186 616
rect 3220 604 3229 616
rect 3177 550 3229 552
tri 3070 543 3076 549 sw
rect 3177 546 3186 550
tri 3177 543 3180 546 ne
rect 3064 516 3076 543
tri 3076 516 3103 543 sw
rect 3180 516 3186 546
rect 3220 546 3229 550
rect 3220 516 3226 546
tri 3226 543 3229 546 nw
rect 2712 515 2791 516
tri 2791 515 2792 516 sw
rect 2712 444 2718 515
rect 2770 463 2782 515
rect 2834 463 2840 515
rect 2868 478 2914 516
tri 2990 515 2991 516 se
rect 2991 515 3103 516
tri 3103 515 3104 516 sw
rect 2752 444 2773 463
tri 2773 444 2792 463 nw
rect 2868 444 2874 478
rect 2908 444 2914 478
rect 2988 463 2994 515
rect 3046 478 3058 515
rect 3110 463 3116 515
rect 3180 478 3226 516
tri 2990 444 3009 463 ne
rect 3009 444 3030 463
rect 3064 444 3085 463
tri 3085 444 3104 463 nw
rect 3180 444 3186 478
rect 3220 444 3226 478
rect 2712 406 2758 444
tri 2758 429 2773 444 nw
rect 2712 372 2718 406
rect 2752 372 2758 406
rect 2712 334 2758 372
tri 2681 318 2682 319 sw
rect 2630 312 2682 318
rect 2630 248 2682 260
rect 2630 190 2682 196
rect 2712 300 2718 334
rect 2752 300 2758 334
rect 2712 262 2758 300
rect 2712 228 2718 262
rect 2752 228 2758 262
rect 2712 190 2758 228
rect 2400 118 2446 156
rect 2400 84 2406 118
rect 2440 84 2446 118
rect 2400 46 2446 84
rect 2400 12 2406 46
rect 2440 12 2446 46
rect 2400 0 2446 12
tri 2553 160 2556 163 se
rect 2556 160 2562 190
rect 2553 156 2562 160
rect 2596 160 2602 190
tri 2602 160 2605 163 sw
rect 2596 156 2605 160
rect 2553 154 2605 156
rect 2553 89 2562 102
rect 2596 89 2605 102
rect 2553 24 2562 37
rect 2596 24 2605 37
tri 2531 -40 2553 -18 se
rect 2712 156 2718 190
rect 2752 156 2758 190
rect 2868 406 2914 444
tri 3009 429 3024 444 ne
rect 2868 372 2874 406
rect 2908 372 2914 406
rect 2868 334 2914 372
rect 2868 300 2874 334
rect 2908 300 2914 334
rect 2868 262 2914 300
rect 2868 228 2874 262
rect 2908 228 2914 262
rect 2868 190 2914 228
rect 2712 118 2758 156
rect 2712 84 2718 118
rect 2752 84 2758 118
rect 2712 46 2758 84
rect 2712 12 2718 46
rect 2752 12 2758 46
rect 2712 0 2758 12
tri 2865 160 2868 163 se
rect 2868 160 2874 190
rect 2865 156 2874 160
rect 2908 160 2914 190
rect 3024 406 3070 444
tri 3070 429 3085 444 nw
rect 3024 372 3030 406
rect 3064 372 3070 406
rect 3024 334 3070 372
rect 3024 300 3030 334
rect 3064 300 3070 334
rect 3024 262 3070 300
rect 3024 228 3030 262
rect 3064 228 3070 262
rect 3024 190 3070 228
tri 2914 160 2917 163 sw
rect 2908 156 2917 160
rect 2865 154 2917 156
rect 2865 89 2874 102
rect 2908 89 2917 102
rect 2865 24 2874 37
rect 2908 24 2917 37
tri 2864 -13 2865 -12 se
tri 2859 -18 2864 -13 se
rect 2864 -18 2865 -13
rect 2553 -40 2605 -28
tri 2605 -40 2627 -18 sw
tri 2837 -40 2859 -18 se
rect 2859 -28 2865 -18
rect 3024 156 3030 190
rect 3064 156 3070 190
rect 3024 118 3070 156
rect 3024 84 3030 118
rect 3064 84 3070 118
rect 3024 46 3070 84
rect 3024 12 3030 46
rect 3064 12 3070 46
rect 3024 0 3070 12
rect 3180 406 3226 444
rect 3180 372 3186 406
rect 3220 372 3226 406
rect 3180 334 3226 372
rect 3180 300 3186 334
rect 3220 300 3226 334
rect 3180 262 3226 300
tri 3254 400 3257 403 se
rect 3257 400 3305 1029
tri 3305 1024 3310 1029 nw
rect 3336 982 3382 994
rect 3336 948 3342 982
rect 3376 948 3382 982
rect 3336 910 3382 948
rect 3336 876 3342 910
rect 3376 876 3382 910
rect 3336 838 3382 876
rect 3336 804 3342 838
rect 3376 804 3382 838
rect 3336 766 3382 804
rect 3336 732 3342 766
rect 3376 732 3382 766
rect 3336 694 3382 732
rect 3336 660 3342 694
rect 3376 660 3382 694
rect 3492 982 3538 994
rect 3492 948 3498 982
rect 3532 948 3538 982
rect 3492 910 3538 948
rect 3492 876 3498 910
rect 3532 876 3538 910
rect 3492 838 3538 876
rect 3492 804 3498 838
rect 3532 804 3538 838
rect 3492 766 3538 804
rect 3492 732 3498 766
rect 3532 732 3538 766
rect 3492 694 3538 732
rect 3336 622 3382 660
rect 3336 588 3342 622
rect 3376 588 3382 622
rect 3336 550 3382 588
rect 3336 516 3342 550
rect 3376 543 3382 550
tri 3489 674 3492 677 se
rect 3492 674 3498 694
rect 3489 668 3498 674
rect 3532 674 3538 694
rect 3648 982 3694 994
rect 3648 948 3654 982
rect 3688 948 3694 982
rect 3648 910 3694 948
rect 3648 876 3654 910
rect 3688 876 3694 910
rect 3648 838 3694 876
rect 3648 804 3654 838
rect 3688 804 3694 838
rect 3648 766 3694 804
rect 3648 732 3654 766
rect 3688 732 3694 766
rect 3648 694 3694 732
tri 3538 674 3541 677 sw
rect 3532 668 3541 674
rect 3489 604 3498 616
rect 3532 604 3541 616
rect 3489 550 3541 552
tri 3382 543 3388 549 sw
rect 3489 546 3498 550
tri 3489 543 3492 546 ne
rect 3376 516 3388 543
tri 3388 516 3415 543 sw
rect 3492 516 3498 546
rect 3532 546 3541 550
rect 3648 660 3654 694
rect 3688 660 3694 694
rect 3648 622 3694 660
rect 3648 588 3654 622
rect 3688 588 3694 622
rect 3648 550 3694 588
rect 3532 516 3538 546
tri 3538 543 3541 546 nw
tri 3642 543 3648 549 se
rect 3648 543 3654 550
tri 3615 516 3642 543 se
rect 3642 516 3654 543
rect 3688 543 3694 550
rect 3772 982 3818 994
rect 3772 948 3778 982
rect 3812 948 3818 982
rect 3772 910 3818 948
rect 3772 876 3778 910
rect 3812 876 3818 910
rect 3772 838 3818 876
rect 3772 804 3778 838
rect 3812 804 3818 838
rect 3772 766 3818 804
rect 3772 732 3778 766
rect 3812 732 3818 766
rect 3772 694 3818 732
rect 3772 660 3778 694
rect 3812 660 3818 694
rect 3772 622 3818 660
rect 3772 588 3778 622
rect 3812 588 3818 622
rect 3772 550 3818 588
tri 3694 543 3700 549 sw
rect 3688 516 3700 543
tri 3700 516 3727 543 sw
rect 3772 516 3778 550
rect 3812 516 3818 550
rect 3336 515 3415 516
tri 3415 515 3416 516 sw
rect 3336 444 3342 515
rect 3394 463 3406 515
rect 3458 463 3464 515
rect 3492 478 3538 516
tri 3614 515 3615 516 se
rect 3615 515 3727 516
tri 3727 515 3728 516 sw
rect 3376 444 3397 463
tri 3397 444 3416 463 nw
rect 3492 444 3498 478
rect 3532 444 3538 478
rect 3612 463 3618 515
rect 3670 478 3682 515
rect 3734 463 3740 515
rect 3772 478 3818 516
tri 3848 484 3849 485 se
rect 3849 484 3897 1042
tri 3897 1033 3906 1042 nw
tri 3996 1033 4005 1042 ne
rect 3928 982 3974 994
rect 3928 948 3934 982
rect 3968 948 3974 982
rect 3928 910 3974 948
rect 3928 876 3934 910
rect 3968 876 3974 910
rect 3928 838 3974 876
rect 3928 804 3934 838
rect 3968 804 3974 838
rect 3928 766 3974 804
rect 3928 732 3934 766
rect 3968 732 3974 766
rect 3928 694 3974 732
tri 3925 674 3928 677 se
rect 3928 674 3934 694
rect 3925 668 3934 674
rect 3968 674 3974 694
tri 3974 674 3977 677 sw
rect 3968 668 3977 674
rect 3925 604 3934 616
rect 3968 604 3977 616
rect 3925 550 3977 552
rect 3925 546 3934 550
tri 3925 543 3928 546 ne
tri 3614 444 3633 463 ne
rect 3633 444 3654 463
rect 3688 444 3709 463
tri 3709 444 3728 463 nw
rect 3772 444 3778 478
rect 3812 444 3818 478
rect 3336 406 3382 444
tri 3382 429 3397 444 nw
tri 3305 400 3306 401 sw
rect 3254 394 3306 400
rect 3254 330 3306 342
rect 3254 272 3306 278
tri 3254 269 3257 272 ne
rect 3257 269 3303 272
tri 3303 269 3306 272 nw
rect 3336 372 3342 406
rect 3376 372 3382 406
rect 3336 334 3382 372
rect 3336 300 3342 334
rect 3376 300 3382 334
rect 3180 228 3186 262
rect 3220 228 3226 262
rect 3180 190 3226 228
rect 3180 156 3186 190
rect 3220 156 3226 190
rect 3180 118 3226 156
rect 3180 84 3186 118
rect 3220 84 3226 118
rect 3180 46 3226 84
rect 3180 12 3186 46
rect 3220 12 3226 46
rect 3180 0 3226 12
rect 3336 262 3382 300
rect 3336 228 3342 262
rect 3376 228 3382 262
rect 3336 190 3382 228
rect 3336 156 3342 190
rect 3376 156 3382 190
rect 3336 118 3382 156
rect 3336 84 3342 118
rect 3376 84 3382 118
rect 3336 46 3382 84
rect 3336 12 3342 46
rect 3376 12 3382 46
rect 3336 0 3382 12
rect 3492 406 3538 444
tri 3633 429 3648 444 ne
rect 3492 372 3498 406
rect 3532 372 3538 406
rect 3492 334 3538 372
rect 3492 300 3498 334
rect 3532 300 3538 334
rect 3492 262 3538 300
rect 3492 228 3498 262
rect 3532 228 3538 262
rect 3492 190 3538 228
rect 3492 156 3498 190
rect 3532 156 3538 190
rect 3492 118 3538 156
rect 3492 84 3498 118
rect 3532 84 3538 118
rect 3492 46 3538 84
rect 3492 12 3498 46
rect 3532 12 3538 46
rect 3492 0 3538 12
rect 3648 406 3694 444
tri 3694 429 3709 444 nw
rect 3648 372 3654 406
rect 3688 372 3694 406
rect 3648 334 3694 372
rect 3648 300 3654 334
rect 3688 300 3694 334
rect 3648 262 3694 300
rect 3648 228 3654 262
rect 3688 228 3694 262
rect 3648 190 3694 228
rect 3648 156 3654 190
rect 3688 156 3694 190
rect 3772 406 3818 444
rect 3772 372 3778 406
rect 3812 372 3818 406
rect 3772 334 3818 372
tri 3846 482 3848 484 se
rect 3848 482 3897 484
rect 3928 516 3934 546
rect 3968 546 3977 550
rect 3968 516 3974 546
tri 3974 543 3977 546 nw
tri 3897 482 3898 483 sw
rect 3846 476 3898 482
rect 3846 412 3898 424
rect 3846 354 3898 360
tri 3846 351 3849 354 ne
rect 3849 351 3895 354
tri 3895 351 3898 354 nw
rect 3928 478 3974 516
rect 4005 484 4053 1042
tri 4227 1033 4236 1042 ne
rect 4236 1033 4290 1042
tri 4290 1033 4299 1042 nw
tri 5163 1033 5172 1042 ne
rect 5172 1033 5226 1042
tri 5226 1033 5235 1042 nw
tri 5555 1033 5564 1042 ne
rect 5564 1033 5622 1042
tri 5622 1033 5631 1042 nw
tri 6129 1041 6130 1042 ne
tri 4236 1032 4237 1033 ne
rect 4084 982 4130 994
rect 4084 948 4090 982
rect 4124 948 4130 982
rect 4084 910 4130 948
rect 4084 876 4090 910
rect 4124 876 4130 910
rect 4084 838 4130 876
rect 4084 804 4090 838
rect 4124 804 4130 838
rect 4084 766 4130 804
rect 4084 732 4090 766
rect 4124 732 4130 766
rect 4084 694 4130 732
rect 4084 660 4090 694
rect 4124 660 4130 694
rect 4084 622 4130 660
rect 4084 588 4090 622
rect 4124 588 4130 622
rect 4084 550 4130 588
rect 4084 516 4090 550
rect 4124 516 4130 550
tri 4053 484 4054 485 sw
rect 3928 444 3934 478
rect 3968 444 3974 478
rect 3928 406 3974 444
rect 3928 372 3934 406
rect 3968 372 3974 406
rect 3772 300 3778 334
rect 3812 300 3818 334
rect 3772 262 3818 300
rect 3772 228 3778 262
rect 3812 228 3818 262
rect 3772 190 3818 228
rect 3648 118 3694 156
rect 3648 84 3654 118
rect 3688 84 3694 118
rect 3648 46 3694 84
rect 3648 12 3654 46
rect 3688 12 3694 46
rect 3648 0 3694 12
tri 3769 160 3772 163 se
rect 3772 160 3778 190
rect 3769 156 3778 160
rect 3812 160 3818 190
rect 3928 334 3974 372
tri 4004 482 4005 483 se
rect 4005 482 4054 484
tri 4054 482 4056 484 sw
rect 4004 476 4056 482
rect 4004 412 4056 424
rect 4004 354 4056 360
tri 4004 351 4007 354 ne
rect 4007 351 4053 354
tri 4053 351 4056 354 nw
rect 4084 478 4130 516
rect 4084 444 4090 478
rect 4124 444 4130 478
rect 4084 406 4130 444
rect 4084 372 4090 406
rect 4124 372 4130 406
rect 3928 300 3934 334
rect 3968 300 3974 334
rect 3928 262 3974 300
rect 3928 228 3934 262
rect 3968 228 3974 262
rect 3928 190 3974 228
tri 3818 160 3821 163 sw
rect 3812 156 3821 160
rect 3769 154 3821 156
rect 3769 89 3778 102
rect 3812 89 3821 102
rect 3769 24 3778 37
rect 3812 24 3821 37
tri 2917 -13 2918 -12 sw
tri 3768 -13 3769 -12 se
rect 2917 -28 2918 -13
rect 2859 -40 2918 -28
tri 2918 -40 2945 -13 sw
tri 3741 -40 3768 -13 se
rect 3768 -28 3769 -13
rect 3928 156 3934 190
rect 3968 156 3974 190
rect 4084 334 4130 372
rect 4084 300 4090 334
rect 4124 300 4130 334
rect 4084 262 4130 300
rect 4084 228 4090 262
rect 4124 228 4130 262
rect 4084 190 4130 228
rect 3928 118 3974 156
rect 3928 84 3934 118
rect 3968 84 3974 118
rect 3928 46 3974 84
rect 3928 12 3934 46
rect 3968 12 3974 46
rect 3928 0 3974 12
tri 4081 160 4084 163 se
rect 4084 160 4090 190
rect 4081 156 4090 160
rect 4124 160 4130 190
rect 4237 982 4289 1033
tri 4289 1032 4290 1033 nw
tri 5172 1032 5173 1033 ne
rect 4237 971 4246 982
rect 4280 971 4289 982
rect 4237 910 4289 919
rect 4237 907 4246 910
rect 4280 907 4289 910
rect 4237 838 4289 855
rect 4237 804 4246 838
rect 4280 804 4289 838
rect 4237 766 4289 804
rect 4237 732 4246 766
rect 4280 732 4289 766
rect 4237 694 4289 732
rect 4237 660 4246 694
rect 4280 660 4289 694
rect 4237 622 4289 660
rect 4237 588 4246 622
rect 4280 588 4289 622
rect 4237 550 4289 588
rect 4237 516 4246 550
rect 4280 516 4289 550
rect 4237 478 4289 516
rect 4237 444 4246 478
rect 4280 444 4289 478
rect 4237 406 4289 444
rect 4237 372 4246 406
rect 4280 372 4289 406
rect 4237 334 4289 372
rect 4237 300 4246 334
rect 4280 300 4289 334
rect 4237 262 4289 300
rect 4237 228 4246 262
rect 4280 228 4289 262
rect 4237 190 4289 228
tri 4130 160 4133 163 sw
rect 4124 156 4133 160
rect 4081 154 4133 156
rect 4081 89 4090 102
rect 4124 89 4133 102
rect 4081 24 4090 37
rect 4124 24 4133 37
tri 3821 -13 3822 -12 sw
tri 4080 -13 4081 -12 se
rect 3821 -28 3822 -13
rect 3768 -40 3822 -28
tri 3822 -40 3849 -13 sw
tri 4053 -40 4080 -13 se
rect 4080 -28 4081 -13
rect 4237 156 4246 190
rect 4280 156 4289 190
rect 4396 982 4442 994
rect 4396 948 4402 982
rect 4436 948 4442 982
rect 4396 910 4442 948
rect 4396 876 4402 910
rect 4436 876 4442 910
rect 4396 838 4442 876
rect 4396 804 4402 838
rect 4436 804 4442 838
rect 4396 766 4442 804
rect 4396 732 4402 766
rect 4436 732 4442 766
rect 4396 694 4442 732
rect 4396 660 4402 694
rect 4436 660 4442 694
rect 4396 622 4442 660
rect 4396 588 4402 622
rect 4436 588 4442 622
rect 4396 550 4442 588
rect 4396 516 4402 550
rect 4436 516 4442 550
rect 4396 478 4442 516
rect 4396 444 4402 478
rect 4436 444 4442 478
rect 4396 406 4442 444
rect 4396 372 4402 406
rect 4436 372 4442 406
rect 4396 334 4442 372
rect 4396 300 4402 334
rect 4436 300 4442 334
rect 4396 262 4442 300
rect 4396 228 4402 262
rect 4436 228 4442 262
rect 4396 190 4442 228
rect 4237 118 4289 156
rect 4237 84 4246 118
rect 4280 84 4289 118
rect 4237 46 4289 84
rect 4237 12 4246 46
rect 4280 12 4289 46
rect 4237 0 4289 12
tri 4393 160 4396 163 se
rect 4396 160 4402 190
rect 4393 156 4402 160
rect 4436 160 4442 190
rect 4552 982 4598 994
rect 4552 948 4558 982
rect 4592 948 4598 982
rect 4552 910 4598 948
rect 4552 876 4558 910
rect 4592 876 4598 910
rect 4552 838 4598 876
rect 4552 804 4558 838
rect 4592 804 4598 838
rect 4552 766 4598 804
rect 4552 732 4558 766
rect 4592 732 4598 766
rect 4552 694 4598 732
rect 4552 660 4558 694
rect 4592 660 4598 694
rect 4552 622 4598 660
rect 4552 588 4558 622
rect 4592 588 4598 622
rect 4552 550 4598 588
rect 4552 516 4558 550
rect 4592 516 4598 550
rect 4552 478 4598 516
rect 4552 444 4558 478
rect 4592 444 4598 478
rect 4552 406 4598 444
rect 4552 372 4558 406
rect 4592 372 4598 406
rect 4552 334 4598 372
rect 4552 300 4558 334
rect 4592 300 4598 334
rect 4552 262 4598 300
rect 4552 228 4558 262
rect 4592 228 4598 262
rect 4552 190 4598 228
tri 4442 160 4445 163 sw
rect 4436 156 4445 160
rect 4393 154 4445 156
rect 4393 89 4402 102
rect 4436 89 4445 102
rect 4393 24 4402 37
rect 4436 24 4445 37
tri 4133 -13 4134 -12 sw
tri 4392 -13 4393 -12 se
rect 4133 -28 4134 -13
rect 4080 -34 4134 -28
tri 4134 -34 4155 -13 sw
tri 4371 -34 4392 -13 se
rect 4392 -28 4393 -13
tri 4549 160 4552 163 se
rect 4552 160 4558 190
rect 4549 156 4558 160
rect 4592 160 4598 190
rect 4703 982 4759 994
rect 4703 948 4714 982
rect 4748 948 4759 982
rect 4703 910 4759 948
rect 4703 876 4714 910
rect 4748 876 4759 910
rect 4703 838 4759 876
rect 4703 804 4714 838
rect 4748 804 4759 838
rect 4703 766 4759 804
rect 4703 732 4714 766
rect 4748 732 4759 766
rect 4703 694 4759 732
rect 4703 660 4714 694
rect 4748 660 4759 694
rect 4703 622 4759 660
rect 4703 588 4714 622
rect 4748 588 4759 622
rect 4703 550 4759 588
rect 4703 516 4714 550
rect 4748 516 4759 550
rect 4864 982 4910 994
rect 4864 948 4870 982
rect 4904 948 4910 982
rect 4864 910 4910 948
rect 4864 876 4870 910
rect 4904 876 4910 910
rect 4864 838 4910 876
rect 4864 804 4870 838
rect 4904 804 4910 838
rect 4864 766 4910 804
rect 4864 732 4870 766
rect 4904 732 4910 766
rect 4864 694 4910 732
rect 4864 660 4870 694
rect 4904 660 4910 694
rect 4864 622 4910 660
rect 4864 588 4870 622
rect 4904 588 4910 622
rect 4864 550 4910 588
tri 4759 516 4784 541 sw
rect 4864 516 4870 550
rect 4904 516 4910 550
rect 4703 507 4784 516
tri 4784 507 4793 516 sw
rect 4703 455 4709 507
rect 4761 455 4773 507
rect 4825 455 4831 507
rect 4864 478 4910 516
rect 4703 444 4714 455
rect 4748 444 4782 455
tri 4782 444 4793 455 nw
rect 4864 444 4870 478
rect 4904 444 4910 478
rect 4703 433 4771 444
tri 4771 433 4782 444 nw
rect 4703 406 4759 433
tri 4759 421 4771 433 nw
rect 4703 372 4714 406
rect 4748 372 4759 406
rect 4703 334 4759 372
rect 4703 300 4714 334
rect 4748 300 4759 334
rect 4703 262 4759 300
rect 4703 228 4714 262
rect 4748 228 4759 262
rect 4703 190 4759 228
tri 4598 160 4601 163 sw
rect 4592 156 4601 160
rect 4549 154 4601 156
rect 4549 89 4558 102
rect 4592 89 4601 102
rect 4549 24 4558 37
rect 4592 24 4601 37
tri 4445 -13 4446 -12 sw
tri 4548 -13 4549 -12 se
rect 4445 -28 4446 -13
rect 4392 -34 4446 -28
tri 4446 -34 4467 -13 sw
tri 4527 -34 4548 -13 se
rect 4548 -28 4549 -13
rect 4703 156 4714 190
rect 4748 156 4759 190
rect 4864 406 4910 444
rect 4864 372 4870 406
rect 4904 372 4910 406
rect 4864 334 4910 372
rect 4864 300 4870 334
rect 4904 300 4910 334
rect 4864 262 4910 300
rect 4864 228 4870 262
rect 4904 228 4910 262
rect 4864 190 4910 228
rect 4703 118 4759 156
rect 4703 84 4714 118
rect 4748 84 4759 118
rect 4703 46 4759 84
rect 4703 12 4714 46
rect 4748 12 4759 46
rect 4703 0 4759 12
tri 4861 160 4864 163 se
rect 4864 160 4870 190
rect 4861 156 4870 160
rect 4904 160 4910 190
rect 5020 982 5066 994
rect 5020 948 5026 982
rect 5060 948 5066 982
rect 5020 910 5066 948
rect 5020 876 5026 910
rect 5060 876 5066 910
rect 5020 838 5066 876
rect 5173 982 5225 1033
tri 5225 1032 5226 1033 nw
tri 5564 1032 5565 1033 ne
rect 5565 1032 5619 1033
tri 5565 1030 5567 1032 ne
rect 5567 1030 5619 1032
tri 5619 1030 5622 1033 nw
rect 5567 1029 5618 1030
tri 5618 1029 5619 1030 nw
rect 5173 971 5182 982
rect 5216 971 5225 982
rect 5173 910 5225 919
rect 5173 907 5182 910
rect 5216 907 5225 910
rect 5173 849 5225 855
tri 5173 846 5176 849 ne
rect 5020 804 5026 838
rect 5060 804 5066 838
rect 5020 766 5066 804
rect 5020 732 5026 766
rect 5060 732 5066 766
rect 5020 694 5066 732
rect 5020 660 5026 694
rect 5060 660 5066 694
rect 5020 622 5066 660
rect 5020 588 5026 622
rect 5060 588 5066 622
rect 5020 550 5066 588
rect 5020 516 5026 550
rect 5060 516 5066 550
rect 5020 478 5066 516
rect 5020 444 5026 478
rect 5060 444 5066 478
rect 5020 406 5066 444
rect 5020 372 5026 406
rect 5060 372 5066 406
rect 5020 334 5066 372
rect 5020 300 5026 334
rect 5060 300 5066 334
rect 5020 262 5066 300
rect 5020 228 5026 262
rect 5060 228 5066 262
rect 5020 190 5066 228
tri 4910 160 4913 163 sw
rect 4904 156 4913 160
rect 4861 154 4913 156
rect 4861 89 4870 102
rect 4904 89 4913 102
rect 4861 24 4870 37
rect 4904 24 4913 37
tri 4601 -13 4602 -12 sw
tri 4860 -13 4861 -12 se
rect 4601 -28 4602 -13
rect 4548 -34 4602 -28
tri 4602 -34 4623 -13 sw
tri 4839 -34 4860 -13 se
rect 4860 -28 4861 -13
tri 5017 160 5020 163 se
rect 5020 160 5026 190
rect 5017 156 5026 160
rect 5060 160 5066 190
rect 5176 838 5222 849
tri 5222 846 5225 849 nw
rect 5332 982 5378 994
rect 5488 982 5534 994
rect 5332 948 5338 982
rect 5372 948 5378 982
rect 5332 910 5378 948
rect 5332 876 5338 910
rect 5372 876 5378 910
rect 5176 804 5182 838
rect 5216 804 5222 838
rect 5176 766 5222 804
rect 5176 732 5182 766
rect 5216 732 5222 766
rect 5176 694 5222 732
rect 5176 660 5182 694
rect 5216 660 5222 694
rect 5176 622 5222 660
rect 5176 588 5182 622
rect 5216 588 5222 622
rect 5176 550 5222 588
rect 5176 516 5182 550
rect 5216 516 5222 550
rect 5176 478 5222 516
rect 5176 444 5182 478
rect 5216 444 5222 478
rect 5176 406 5222 444
rect 5176 372 5182 406
rect 5216 372 5222 406
rect 5176 334 5222 372
rect 5176 300 5182 334
rect 5216 300 5222 334
rect 5176 262 5222 300
rect 5176 228 5182 262
rect 5216 228 5222 262
rect 5176 190 5222 228
tri 5066 160 5069 163 sw
rect 5060 156 5069 160
rect 5017 154 5069 156
rect 5017 89 5026 102
rect 5060 89 5069 102
rect 5017 24 5026 37
rect 5060 24 5069 37
tri 4913 -13 4914 -12 sw
tri 5016 -13 5017 -12 se
rect 4913 -28 4914 -13
rect 4860 -34 4914 -28
tri 4914 -34 4935 -13 sw
tri 4995 -34 5016 -13 se
rect 5016 -28 5017 -13
rect 5176 156 5182 190
rect 5216 156 5222 190
rect 5332 838 5378 876
tri 5483 977 5488 982 se
rect 5488 977 5494 982
rect 5483 971 5494 977
rect 5528 977 5534 982
tri 5534 977 5535 978 sw
rect 5528 971 5535 977
rect 5483 910 5535 919
rect 5483 907 5494 910
rect 5528 907 5535 910
rect 5483 849 5535 855
tri 5483 846 5486 849 ne
rect 5486 846 5534 849
tri 5534 848 5535 849 nw
tri 5486 844 5488 846 ne
rect 5332 804 5338 838
rect 5372 804 5378 838
rect 5332 766 5378 804
rect 5332 732 5338 766
rect 5372 732 5378 766
rect 5332 694 5378 732
rect 5332 660 5338 694
rect 5372 660 5378 694
rect 5332 622 5378 660
rect 5332 588 5338 622
rect 5372 588 5378 622
rect 5332 550 5378 588
rect 5332 516 5338 550
rect 5372 516 5378 550
rect 5332 478 5378 516
rect 5332 444 5338 478
rect 5372 444 5378 478
rect 5332 406 5378 444
rect 5332 372 5338 406
rect 5372 372 5378 406
rect 5332 334 5378 372
rect 5332 300 5338 334
rect 5372 300 5378 334
rect 5332 262 5378 300
rect 5332 228 5338 262
rect 5372 228 5378 262
rect 5332 190 5378 228
rect 5176 118 5222 156
rect 5176 84 5182 118
rect 5216 84 5222 118
rect 5176 46 5222 84
rect 5176 12 5182 46
rect 5216 12 5222 46
rect 5176 0 5222 12
tri 5329 160 5332 163 se
rect 5332 160 5338 190
rect 5329 156 5338 160
rect 5372 160 5378 190
rect 5488 838 5534 846
rect 5488 804 5494 838
rect 5528 804 5534 838
rect 5488 766 5534 804
rect 5488 732 5494 766
rect 5528 732 5534 766
rect 5488 694 5534 732
rect 5488 660 5494 694
rect 5528 660 5534 694
rect 5488 622 5534 660
rect 5488 588 5494 622
rect 5528 588 5534 622
rect 5488 550 5534 588
rect 5488 516 5494 550
rect 5528 516 5534 550
rect 5488 478 5534 516
rect 5488 444 5494 478
rect 5528 444 5534 478
rect 5488 406 5534 444
rect 5567 564 5617 1029
tri 5617 1028 5618 1029 nw
rect 5662 982 5708 994
rect 5662 948 5668 982
rect 5702 948 5708 982
rect 5662 910 5708 948
rect 5662 876 5668 910
rect 5702 876 5708 910
rect 5662 838 5708 876
rect 5662 804 5668 838
rect 5702 804 5708 838
rect 5662 779 5708 804
rect 5818 982 5864 994
rect 5818 948 5824 982
rect 5858 948 5864 982
rect 5818 910 5864 948
rect 5818 876 5824 910
rect 5858 876 5864 910
rect 5818 838 5864 876
rect 5818 804 5824 838
rect 5858 804 5864 838
tri 5708 779 5717 788 sw
rect 5662 770 5717 779
tri 5717 770 5726 779 sw
rect 5662 766 5726 770
tri 5726 766 5730 770 sw
rect 5818 766 5864 804
tri 5656 754 5662 760 se
rect 5662 754 5668 766
rect 5702 760 5730 766
tri 5730 760 5736 766 sw
rect 5702 754 5736 760
tri 5736 754 5742 760 sw
rect 5656 702 5662 754
rect 5714 702 5729 754
rect 5781 702 5787 754
rect 5818 732 5824 766
rect 5858 732 5864 766
tri 5656 698 5660 702 ne
rect 5660 698 5738 702
tri 5738 698 5742 702 nw
tri 5660 696 5662 698 ne
rect 5662 696 5736 698
tri 5736 696 5738 698 nw
rect 5662 694 5734 696
tri 5734 694 5736 696 nw
rect 5818 694 5864 732
rect 5662 660 5668 694
rect 5702 689 5729 694
tri 5729 689 5734 694 nw
rect 5702 660 5708 689
tri 5708 668 5729 689 nw
rect 5662 622 5708 660
rect 5662 588 5668 622
rect 5702 588 5708 622
tri 5617 564 5619 566 sw
rect 5567 558 5619 564
rect 5567 494 5619 506
rect 5567 436 5619 442
tri 5567 433 5570 436 ne
rect 5570 433 5616 436
tri 5616 433 5619 436 nw
rect 5662 550 5708 588
rect 5662 516 5668 550
rect 5702 516 5708 550
rect 5662 478 5708 516
rect 5662 444 5668 478
rect 5702 444 5708 478
rect 5488 372 5494 406
rect 5528 372 5534 406
rect 5488 334 5534 372
rect 5488 300 5494 334
rect 5528 300 5534 334
rect 5488 262 5534 300
rect 5488 228 5494 262
rect 5528 228 5534 262
rect 5488 190 5534 228
tri 5378 160 5381 163 sw
rect 5372 156 5381 160
rect 5329 154 5381 156
rect 5329 89 5338 102
rect 5372 89 5381 102
rect 5329 24 5338 37
rect 5372 24 5381 37
tri 5069 -13 5070 -12 sw
tri 5328 -13 5329 -12 se
rect 5069 -28 5070 -13
rect 5016 -34 5070 -28
rect 4080 -40 4155 -34
tri 4155 -40 4161 -34 sw
tri 4365 -40 4371 -34 se
rect 4371 -40 4467 -34
tri 4467 -40 4473 -34 sw
tri 4521 -40 4527 -34 se
rect 4527 -40 4623 -34
tri 4623 -40 4629 -34 sw
tri 4833 -40 4839 -34 se
rect 4839 -40 4935 -34
tri 4935 -40 4941 -34 sw
tri 4989 -40 4995 -34 se
rect 4995 -40 5070 -34
tri 5070 -40 5097 -13 sw
tri 5301 -40 5328 -13 se
rect 5328 -28 5329 -13
rect 5488 156 5494 190
rect 5528 156 5534 190
rect 5488 118 5534 156
rect 5488 84 5494 118
rect 5528 84 5534 118
rect 5488 46 5534 84
rect 5488 12 5494 46
rect 5528 12 5534 46
rect 5488 0 5534 12
rect 5662 406 5708 444
rect 5662 372 5668 406
rect 5702 372 5708 406
rect 5662 334 5708 372
rect 5662 300 5668 334
rect 5702 300 5708 334
rect 5662 262 5708 300
rect 5662 228 5668 262
rect 5702 228 5708 262
rect 5662 190 5708 228
rect 5662 156 5668 190
rect 5702 156 5708 190
rect 5818 660 5824 694
rect 5858 660 5864 694
rect 5974 982 6020 994
rect 5974 948 5980 982
rect 6014 948 6020 982
rect 5974 910 6020 948
rect 5974 876 5980 910
rect 6014 876 6020 910
rect 5974 838 6020 876
rect 5974 804 5980 838
rect 6014 804 6020 838
rect 5974 766 6020 804
rect 5974 732 5980 766
rect 6014 732 6020 766
rect 5974 694 6020 732
tri 5947 662 5974 689 se
rect 5974 662 5980 694
tri 5945 660 5947 662 se
rect 5947 660 5980 662
rect 6014 660 6020 694
rect 6130 982 6176 1042
rect 6204 1114 6256 1116
tri 6256 1114 6258 1116 sw
rect 6204 1110 6258 1114
rect 6256 1108 6258 1110
tri 6258 1108 6264 1114 sw
rect 6256 1104 6264 1108
tri 6264 1104 6268 1108 sw
rect 6256 1098 6344 1104
rect 6260 1064 6298 1098
rect 6332 1064 6344 1098
rect 6256 1058 6344 1064
rect 6430 1096 6455 1108
rect 6507 1096 6519 1108
rect 6571 1102 6579 1108
tri 6579 1102 6585 1108 sw
rect 6571 1096 6782 1102
rect 6430 1062 6442 1096
rect 6507 1062 6516 1096
rect 6571 1062 6590 1096
rect 6624 1062 6663 1096
rect 6697 1062 6736 1096
rect 6770 1062 6782 1096
rect 6919 1090 6965 1102
rect 6204 1056 6279 1058
tri 6279 1056 6281 1058 nw
rect 6430 1056 6455 1062
rect 6507 1056 6519 1062
rect 6571 1056 6782 1062
tri 6908 1056 6919 1067 se
rect 6919 1056 6925 1090
rect 6959 1056 6965 1090
rect 6204 1046 6265 1056
rect 6256 1042 6265 1046
tri 6265 1042 6279 1056 nw
tri 6894 1042 6908 1056 se
rect 6908 1042 6965 1056
tri 6256 1033 6265 1042 nw
tri 6885 1033 6894 1042 se
rect 6894 1033 6965 1042
tri 6881 1029 6885 1033 se
rect 6885 1029 6965 1033
tri 6878 1026 6881 1029 se
rect 6881 1026 6965 1029
tri 6689 1025 6690 1026 se
rect 6690 1025 6736 1026
rect 6204 988 6256 994
tri 6285 1022 6288 1025 se
rect 6288 1022 6334 1025
tri 6334 1022 6337 1025 sw
rect 6285 1016 6337 1022
rect 6130 948 6136 982
rect 6170 948 6176 982
rect 6130 910 6176 948
rect 6130 876 6136 910
rect 6170 876 6176 910
tri 6687 1023 6689 1025 se
rect 6689 1023 6736 1025
tri 6736 1023 6739 1026 sw
tri 6875 1023 6878 1026 se
rect 6878 1023 6965 1026
rect 6687 1017 6739 1023
rect 6285 952 6292 964
rect 6326 952 6337 964
rect 6285 894 6292 900
tri 6285 893 6286 894 ne
rect 6130 838 6176 876
rect 6130 804 6136 838
rect 6170 804 6176 838
rect 6130 766 6176 804
rect 6130 732 6136 766
rect 6170 732 6176 766
rect 6130 694 6176 732
tri 6020 660 6022 662 sw
rect 6130 660 6136 694
rect 6170 660 6176 694
rect 5818 622 5864 660
tri 5940 655 5945 660 se
rect 5945 656 6022 660
tri 6022 656 6026 660 sw
rect 5945 655 6026 656
tri 6026 655 6027 656 sw
rect 5818 588 5824 622
rect 5858 588 5864 622
rect 5896 603 5902 655
rect 5954 603 5969 655
rect 6021 603 6027 655
tri 5940 596 5947 603 ne
rect 5947 596 5980 603
tri 5947 588 5955 596 ne
rect 5955 588 5980 596
rect 6014 588 6020 603
tri 6020 596 6027 603 nw
rect 6130 622 6176 660
rect 5818 550 5864 588
tri 5955 569 5974 588 ne
rect 5818 516 5824 550
rect 5858 516 5864 550
rect 5818 478 5864 516
rect 5818 444 5824 478
rect 5858 444 5864 478
rect 5818 406 5864 444
rect 5818 372 5824 406
rect 5858 372 5864 406
rect 5818 334 5864 372
rect 5818 300 5824 334
rect 5858 300 5864 334
rect 5818 262 5864 300
rect 5818 228 5824 262
rect 5858 228 5864 262
rect 5818 190 5864 228
tri 5817 163 5818 164 se
rect 5818 163 5824 190
rect 5662 118 5708 156
rect 5662 84 5668 118
rect 5702 84 5708 118
rect 5662 46 5708 84
rect 5662 12 5668 46
rect 5702 12 5708 46
rect 5662 0 5708 12
tri 5814 160 5817 163 se
rect 5817 160 5824 163
rect 5814 156 5824 160
rect 5858 160 5864 190
rect 5974 550 6020 588
rect 5974 516 5980 550
rect 6014 516 6020 550
rect 6130 588 6136 622
rect 6170 588 6176 622
rect 6130 550 6176 588
tri 6128 522 6130 524 se
rect 6130 522 6136 550
tri 6125 519 6128 522 se
rect 6128 519 6136 522
tri 6122 516 6125 519 se
rect 6125 516 6136 519
rect 6170 516 6176 550
rect 6286 876 6292 894
rect 6326 894 6337 900
rect 6326 892 6335 894
tri 6335 892 6337 894 nw
rect 6410 982 6456 994
rect 6410 948 6416 982
rect 6450 948 6456 982
rect 6410 910 6456 948
rect 6326 876 6332 892
tri 6332 889 6335 892 nw
rect 6286 838 6332 876
rect 6286 804 6292 838
rect 6326 804 6332 838
rect 6286 766 6332 804
rect 6286 732 6292 766
rect 6326 732 6332 766
rect 6286 694 6332 732
rect 6286 660 6292 694
rect 6326 660 6332 694
rect 6286 622 6332 660
rect 6286 588 6292 622
rect 6326 588 6332 622
rect 6286 550 6332 588
tri 6176 516 6179 519 sw
rect 6286 516 6292 550
rect 6326 516 6332 550
rect 5974 478 6020 516
tri 6097 491 6122 516 se
rect 6122 491 6179 516
tri 6179 491 6204 516 sw
tri 6096 490 6097 491 se
rect 6097 490 6204 491
tri 6204 490 6205 491 sw
rect 5974 444 5980 478
rect 6014 444 6020 478
rect 5974 406 6020 444
rect 6079 438 6085 490
rect 6137 478 6149 490
rect 6137 438 6149 444
rect 6201 438 6207 490
rect 6286 478 6332 516
rect 6286 444 6292 478
rect 6326 444 6332 478
tri 6096 433 6101 438 ne
rect 6101 433 6200 438
tri 6200 433 6205 438 nw
tri 6101 421 6113 433 ne
rect 6113 421 6188 433
tri 6188 421 6200 433 nw
tri 6113 419 6115 421 ne
rect 6115 419 6186 421
tri 6186 419 6188 421 nw
tri 6115 410 6124 419 ne
rect 6124 410 6177 419
tri 6177 410 6186 419 nw
tri 6124 409 6125 410 ne
rect 6125 409 6176 410
tri 6176 409 6177 410 nw
tri 6125 406 6128 409 ne
rect 6128 406 6176 409
rect 5974 372 5980 406
rect 6014 372 6020 406
tri 6128 404 6130 406 ne
rect 5974 334 6020 372
rect 5974 300 5980 334
rect 6014 300 6020 334
rect 5974 262 6020 300
rect 5974 228 5980 262
rect 6014 228 6020 262
rect 5974 190 6020 228
tri 5864 160 5866 162 sw
rect 5858 156 5866 160
rect 5814 154 5866 156
rect 5814 89 5824 102
rect 5858 89 5866 102
rect 5814 24 5824 37
rect 5858 24 5866 37
tri 5381 -13 5382 -12 sw
tri 5813 -13 5814 -12 se
rect 5381 -28 5382 -13
rect 5328 -40 5382 -28
tri 5382 -40 5409 -13 sw
tri 5786 -40 5813 -13 se
rect 5813 -28 5814 -13
rect 5974 156 5980 190
rect 6014 156 6020 190
rect 5974 118 6020 156
rect 5974 84 5980 118
rect 6014 84 6020 118
rect 5974 46 6020 84
rect 5974 12 5980 46
rect 6014 12 6020 46
rect 5974 0 6020 12
rect 6130 372 6136 406
rect 6170 372 6176 406
rect 6130 334 6176 372
rect 6130 300 6136 334
rect 6170 300 6176 334
rect 6130 262 6176 300
rect 6130 228 6136 262
rect 6170 228 6176 262
rect 6130 190 6176 228
rect 6130 156 6136 190
rect 6170 156 6176 190
rect 6130 118 6176 156
rect 6130 84 6136 118
rect 6170 84 6176 118
rect 6130 46 6176 84
rect 6130 12 6136 46
rect 6170 12 6176 46
rect 6130 0 6176 12
rect 6286 406 6332 444
rect 6286 372 6292 406
rect 6326 372 6332 406
rect 6286 334 6332 372
rect 6286 300 6292 334
rect 6326 300 6332 334
rect 6286 262 6332 300
rect 6286 228 6292 262
rect 6326 228 6332 262
rect 6286 190 6332 228
rect 6286 156 6292 190
rect 6326 156 6332 190
rect 6410 876 6416 910
rect 6450 876 6456 910
rect 6410 838 6456 876
rect 6410 804 6416 838
rect 6450 804 6456 838
rect 6410 766 6456 804
rect 6410 732 6416 766
rect 6450 732 6456 766
rect 6410 694 6456 732
rect 6410 660 6416 694
rect 6450 660 6456 694
rect 6410 622 6456 660
rect 6566 982 6612 994
rect 6566 948 6572 982
rect 6606 948 6612 982
rect 6566 910 6612 948
rect 6566 876 6572 910
rect 6606 876 6612 910
tri 6866 1014 6875 1023 se
rect 6875 1014 6965 1023
rect 6687 953 6696 965
rect 6730 953 6739 965
rect 6687 895 6696 901
tri 6687 894 6688 895 ne
rect 6688 894 6696 895
tri 6688 892 6690 894 ne
rect 6566 838 6612 876
rect 6566 804 6572 838
rect 6606 804 6612 838
rect 6566 766 6612 804
rect 6566 732 6572 766
rect 6606 732 6612 766
rect 6566 694 6612 732
rect 6566 660 6572 694
rect 6606 660 6612 694
tri 6565 655 6566 656 se
rect 6566 655 6612 660
rect 6690 876 6696 894
rect 6730 895 6739 901
rect 6730 876 6736 895
tri 6736 892 6739 895 nw
tri 6846 994 6866 1014 se
rect 6866 994 6925 1014
rect 6846 982 6925 994
rect 6846 948 6852 982
rect 6886 980 6925 982
rect 6959 980 6965 1014
rect 6886 968 6965 980
rect 7002 982 7048 1200
rect 6886 948 6924 968
tri 6924 948 6944 968 nw
rect 7002 948 7008 982
rect 7042 948 7048 982
rect 6846 923 6899 948
tri 6899 923 6924 948 nw
rect 6846 910 6892 923
tri 6892 916 6899 923 nw
rect 6690 838 6736 876
rect 6690 804 6696 838
rect 6730 804 6736 838
rect 6690 766 6736 804
rect 6690 732 6696 766
rect 6730 732 6736 766
rect 6690 694 6736 732
rect 6690 660 6696 694
rect 6730 660 6736 694
tri 6612 655 6613 656 sw
rect 6410 588 6416 622
rect 6450 588 6456 622
rect 6410 550 6456 588
rect 6410 516 6416 550
rect 6450 516 6456 550
tri 6563 653 6565 655 se
rect 6565 653 6613 655
tri 6613 653 6615 655 sw
rect 6563 647 6615 653
rect 6563 588 6572 595
rect 6606 588 6615 595
rect 6563 583 6615 588
rect 6563 525 6572 531
tri 6563 522 6566 525 ne
rect 6410 478 6456 516
rect 6410 444 6416 478
rect 6450 444 6456 478
rect 6410 406 6456 444
rect 6410 372 6416 406
rect 6450 372 6456 406
rect 6410 334 6456 372
rect 6410 300 6416 334
rect 6450 300 6456 334
rect 6410 262 6456 300
rect 6410 228 6416 262
rect 6450 228 6456 262
rect 6410 190 6456 228
rect 6286 118 6332 156
rect 6286 84 6292 118
rect 6326 84 6332 118
rect 6286 46 6332 84
rect 6286 12 6292 46
rect 6326 12 6332 46
rect 6286 0 6332 12
tri 6407 160 6410 163 se
rect 6410 160 6416 190
rect 6407 156 6416 160
rect 6450 160 6456 190
rect 6566 516 6572 525
rect 6606 525 6615 531
rect 6606 516 6612 525
tri 6612 522 6615 525 nw
rect 6690 622 6736 660
rect 6690 588 6696 622
rect 6730 588 6736 622
rect 6690 550 6736 588
rect 6566 478 6612 516
rect 6566 444 6572 478
rect 6606 444 6612 478
rect 6566 406 6612 444
rect 6566 372 6572 406
rect 6606 372 6612 406
rect 6566 334 6612 372
rect 6566 300 6572 334
rect 6606 300 6612 334
rect 6566 262 6612 300
rect 6566 228 6572 262
rect 6606 228 6612 262
rect 6566 190 6612 228
tri 6456 160 6459 163 sw
rect 6450 156 6459 160
rect 6407 154 6459 156
rect 6407 89 6416 102
rect 6450 89 6459 102
rect 6407 24 6416 37
rect 6450 24 6459 37
tri 5866 -13 5867 -12 sw
tri 6406 -13 6407 -12 se
rect 5866 -28 5867 -13
rect 5813 -40 5867 -28
tri 5867 -40 5894 -13 sw
tri 6379 -40 6406 -13 se
rect 6406 -28 6407 -13
rect 6566 156 6572 190
rect 6606 156 6612 190
rect 6566 118 6612 156
rect 6566 84 6572 118
rect 6606 84 6612 118
rect 6566 46 6612 84
rect 6566 12 6572 46
rect 6606 12 6612 46
rect 6566 0 6612 12
rect 6690 516 6696 550
rect 6730 516 6736 550
rect 6690 478 6736 516
rect 6690 444 6696 478
rect 6730 444 6736 478
rect 6690 406 6736 444
rect 6690 372 6696 406
rect 6730 372 6736 406
rect 6690 334 6736 372
rect 6690 300 6696 334
rect 6730 300 6736 334
rect 6690 262 6736 300
rect 6690 228 6696 262
rect 6730 228 6736 262
rect 6690 190 6736 228
rect 6690 156 6696 190
rect 6730 156 6736 190
rect 6846 876 6852 910
rect 6886 876 6892 910
rect 6846 838 6892 876
rect 6846 804 6852 838
rect 6886 804 6892 838
rect 6846 766 6892 804
rect 6846 732 6852 766
rect 6886 732 6892 766
rect 6846 694 6892 732
rect 6846 660 6852 694
rect 6886 660 6892 694
rect 6846 622 6892 660
rect 6846 588 6852 622
rect 6886 588 6892 622
rect 6846 550 6892 588
rect 6846 516 6852 550
rect 6886 516 6892 550
rect 6846 478 6892 516
rect 6846 444 6852 478
rect 6886 444 6892 478
rect 6846 406 6892 444
rect 6846 372 6852 406
rect 6886 372 6892 406
rect 6846 334 6892 372
rect 6846 300 6852 334
rect 6886 300 6892 334
rect 6846 262 6892 300
rect 6846 228 6852 262
rect 6886 228 6892 262
rect 6846 190 6892 228
rect 6690 118 6736 156
rect 6690 84 6696 118
rect 6730 84 6736 118
rect 6690 46 6736 84
rect 6690 12 6696 46
rect 6730 12 6736 46
rect 6690 0 6736 12
tri 6843 160 6846 163 se
rect 6846 160 6852 190
rect 6843 156 6852 160
rect 6886 160 6892 190
rect 7002 910 7048 948
rect 7002 876 7008 910
rect 7042 876 7048 910
rect 7002 838 7048 876
rect 7002 804 7008 838
rect 7042 804 7048 838
rect 7002 766 7048 804
rect 7002 732 7008 766
rect 7042 732 7048 766
rect 7002 694 7048 732
rect 7002 660 7008 694
rect 7042 660 7048 694
rect 7002 622 7048 660
rect 7002 588 7008 622
rect 7042 588 7048 622
rect 7002 550 7048 588
rect 7002 516 7008 550
rect 7042 516 7048 550
rect 7002 478 7048 516
rect 7002 444 7008 478
rect 7042 444 7048 478
rect 7002 406 7048 444
rect 7002 372 7008 406
rect 7042 372 7048 406
rect 7002 334 7048 372
rect 7002 300 7008 334
rect 7042 300 7048 334
rect 7002 262 7048 300
rect 7002 228 7008 262
rect 7042 228 7048 262
rect 7002 190 7048 228
tri 6892 160 6895 163 sw
rect 6886 156 6895 160
rect 6843 154 6895 156
rect 6843 89 6852 102
rect 6886 89 6895 102
rect 6843 24 6852 37
rect 6886 24 6895 37
tri 6459 -13 6460 -12 sw
tri 6842 -13 6843 -12 se
rect 6459 -28 6460 -13
rect 6406 -40 6460 -28
tri 6460 -40 6487 -13 sw
tri 6815 -40 6842 -13 se
rect 6842 -28 6843 -13
rect 7002 156 7008 190
rect 7042 156 7048 190
rect 7002 118 7048 156
rect 7002 84 7008 118
rect 7042 84 7048 118
rect 7002 46 7048 84
rect 7002 12 7008 46
rect 7042 12 7048 46
rect 7002 0 7048 12
rect 7141 1312 7142 1364
rect 7194 1312 7208 1364
rect 7141 1294 7260 1312
rect 7141 1242 7142 1294
rect 7194 1242 7208 1294
rect 7141 1224 7260 1242
rect 7141 1172 7142 1224
rect 7194 1172 7208 1224
rect 7141 154 7260 1172
rect 7325 1433 7827 1439
tri 7939 1434 7961 1456 se
rect 7961 1446 8923 1456
rect 7961 1434 8911 1446
tri 8911 1434 8923 1446 nw
tri 8952 2353 8962 2363 se
rect 8962 2353 11751 2363
tri 11751 2353 11761 2363 nw
rect 8952 2338 11736 2353
tri 11736 2338 11751 2353 nw
rect 8952 2334 11732 2338
tri 11732 2334 11736 2338 nw
tri 11798 2334 11802 2338 se
rect 11802 2334 11854 2976
tri 11854 2968 11862 2976 nw
tri 17693 2972 17697 2976 se
rect 17697 2972 17757 2976
tri 12855 2961 12856 2962 se
rect 12856 2961 12862 2962
tri 11908 2942 11927 2961 se
rect 11927 2942 12862 2961
tri 11892 2926 11908 2942 se
rect 11908 2926 12862 2942
rect 8952 2304 9008 2334
tri 9008 2304 9038 2334 nw
tri 11768 2304 11798 2334 se
rect 11798 2304 11854 2334
tri 7938 1433 7939 1434 se
rect 7939 1433 8901 1434
rect 7325 1413 7384 1433
tri 7384 1413 7404 1433 nw
tri 7929 1424 7938 1433 se
rect 7938 1424 8901 1433
tri 8901 1424 8911 1434 nw
rect 7929 1417 8894 1424
tri 8894 1417 8901 1424 nw
rect 7929 1413 8003 1417
tri 8003 1413 8007 1417 nw
rect 7325 647 7377 1413
tri 7377 1406 7384 1413 nw
rect 7929 1406 7996 1413
tri 7996 1406 8003 1413 nw
tri 8945 1406 8952 1413 se
rect 8952 1406 9004 2304
tri 9004 2300 9008 2304 nw
tri 9059 2300 9063 2304 se
rect 9063 2300 11854 2304
tri 9037 2278 9059 2300 se
rect 9059 2289 11854 2300
rect 9059 2278 11843 2289
tri 11843 2278 11854 2289 nw
tri 11886 2920 11892 2926 se
rect 11892 2920 12862 2926
rect 11886 2910 12862 2920
rect 12914 2910 12926 2962
rect 12978 2961 12984 2962
tri 12984 2961 12985 2962 sw
rect 12978 2910 16301 2961
rect 11886 2909 16301 2910
rect 16353 2909 16365 2961
rect 16417 2909 16423 2961
rect 16766 2920 16772 2972
rect 16824 2920 16836 2972
rect 16888 2920 17757 2972
rect 17789 2930 17795 2982
rect 17847 2976 17859 2982
rect 17911 2976 19045 2982
rect 17847 2942 17855 2976
rect 17911 2942 17954 2976
rect 17988 2942 18053 2976
rect 18087 2942 18339 2976
rect 18373 2942 18438 2976
rect 18472 2942 18537 2976
rect 18571 2942 18801 2976
rect 18835 2942 18900 2976
rect 18934 2942 18999 2976
rect 19033 2942 19045 2976
tri 19963 2968 19977 2982 ne
rect 19977 2968 20002 2982
tri 19977 2964 19981 2968 ne
rect 19981 2964 20002 2968
rect 20036 2964 20042 2998
tri 19981 2962 19983 2964 ne
rect 19983 2962 20042 2964
tri 19983 2961 19984 2962 ne
rect 19984 2961 20042 2962
tri 19984 2949 19996 2961 ne
rect 17847 2930 17859 2942
rect 17911 2936 19045 2942
rect 17911 2930 17917 2936
tri 17917 2930 17923 2936 nw
rect 11886 2895 11958 2909
tri 11958 2895 11972 2909 nw
rect 11886 2892 11955 2895
tri 11955 2892 11958 2895 nw
rect 11886 2883 11946 2892
tri 11946 2883 11955 2892 nw
rect 18405 2883 18953 2895
rect 19005 2883 19044 2895
tri 9035 2276 9037 2278 se
rect 9037 2276 11841 2278
tri 11841 2276 11843 2278 nw
rect 7418 1389 7464 1401
rect 7418 1355 7424 1389
rect 7458 1355 7464 1389
rect 7418 1317 7464 1355
rect 7418 1283 7424 1317
rect 7458 1283 7464 1317
rect 7504 1389 7550 1401
rect 7504 1355 7510 1389
rect 7544 1355 7550 1389
rect 7504 1317 7550 1355
rect 7418 1245 7464 1283
rect 7418 1211 7424 1245
rect 7458 1211 7464 1245
rect 7418 1173 7464 1211
rect 7418 1139 7424 1173
rect 7458 1139 7464 1173
tri 7501 1299 7504 1302 se
rect 7504 1299 7510 1317
rect 7501 1293 7510 1299
rect 7544 1299 7550 1317
rect 7590 1389 7636 1401
rect 7590 1355 7596 1389
rect 7630 1355 7636 1389
rect 7590 1317 7636 1355
tri 7550 1299 7553 1302 sw
rect 7544 1293 7553 1299
rect 7501 1229 7510 1241
rect 7544 1229 7553 1241
rect 7501 1173 7553 1177
rect 7501 1171 7510 1173
tri 7501 1168 7504 1171 ne
rect 7418 1101 7464 1139
rect 7418 1067 7424 1101
rect 7458 1067 7464 1101
rect 7418 1029 7464 1067
rect 7418 995 7424 1029
rect 7458 995 7464 1029
rect 7418 957 7464 995
rect 7418 923 7424 957
rect 7458 923 7464 957
rect 7418 885 7464 923
rect 7418 851 7424 885
rect 7458 851 7464 885
rect 7418 813 7464 851
rect 7418 779 7424 813
rect 7458 779 7464 813
rect 7418 741 7464 779
rect 7418 707 7424 741
rect 7458 707 7464 741
rect 7418 669 7464 707
rect 7418 635 7424 669
rect 7458 635 7464 669
rect 7325 583 7377 595
rect 7325 525 7377 531
tri 7414 610 7418 614 se
rect 7418 610 7464 635
rect 7504 1139 7510 1171
rect 7544 1171 7553 1173
rect 7544 1139 7550 1171
tri 7550 1168 7553 1171 nw
rect 7590 1283 7596 1317
rect 7630 1283 7636 1317
rect 7676 1389 7722 1401
rect 7676 1355 7682 1389
rect 7716 1355 7722 1389
rect 7676 1317 7722 1355
rect 7590 1245 7636 1283
rect 7590 1211 7596 1245
rect 7630 1211 7636 1245
rect 7590 1173 7636 1211
rect 7504 1101 7550 1139
rect 7504 1067 7510 1101
rect 7544 1067 7550 1101
rect 7504 1029 7550 1067
rect 7504 995 7510 1029
rect 7544 995 7550 1029
rect 7504 957 7550 995
rect 7504 923 7510 957
rect 7544 923 7550 957
rect 7504 885 7550 923
rect 7504 851 7510 885
rect 7544 851 7550 885
rect 7504 813 7550 851
rect 7504 779 7510 813
rect 7544 779 7550 813
rect 7504 741 7550 779
rect 7504 707 7510 741
rect 7544 707 7550 741
rect 7504 669 7550 707
rect 7504 635 7510 669
rect 7544 635 7550 669
tri 7464 610 7466 612 sw
rect 7414 604 7466 610
rect 7414 540 7466 552
rect 7414 482 7466 488
tri 7414 480 7416 482 ne
rect 7416 480 7466 482
tri 7416 478 7418 480 ne
rect 7141 102 7142 154
rect 7194 102 7208 154
rect 7141 84 7260 102
rect 7141 32 7142 84
rect 7194 32 7208 84
rect 7141 13 7260 32
rect 6842 -40 6895 -28
tri 6895 -40 6902 -33 sw
rect 7141 -39 7142 13
rect 7194 -39 7208 13
tri 2519 -52 2531 -40 se
rect 2531 -46 2627 -40
tri 2627 -46 2633 -40 sw
tri 2831 -46 2837 -40 se
rect 2837 -46 2945 -40
tri 2945 -46 2951 -40 sw
tri 3735 -46 3741 -40 se
rect 3741 -46 3849 -40
tri 3849 -46 3855 -40 sw
tri 4047 -46 4053 -40 se
rect 4053 -46 4161 -40
tri 4161 -46 4167 -40 sw
tri 4359 -46 4365 -40 se
rect 4365 -46 4473 -40
tri 4473 -46 4479 -40 sw
tri 4515 -46 4521 -40 se
rect 4521 -46 4629 -40
tri 4629 -46 4635 -40 sw
tri 4827 -46 4833 -40 se
rect 4833 -46 4941 -40
tri 4941 -46 4947 -40 sw
tri 4983 -46 4989 -40 se
rect 4989 -46 5097 -40
tri 5097 -46 5103 -40 sw
tri 5295 -46 5301 -40 se
rect 5301 -46 5409 -40
tri 5409 -46 5415 -40 sw
tri 5780 -46 5786 -40 se
rect 5786 -46 5894 -40
tri 5894 -46 5900 -40 sw
tri 6373 -46 6379 -40 se
rect 6379 -46 6487 -40
tri 6487 -46 6493 -40 sw
tri 6809 -46 6815 -40 se
rect 6815 -46 6902 -40
tri 6902 -46 6908 -40 sw
rect 2531 -52 2633 -46
tri 2633 -52 2639 -46 sw
tri 2736 -52 2742 -46 se
rect 2742 -52 2748 -46
rect 2398 -58 2748 -52
rect 2800 -58 2813 -46
rect 2865 -58 2878 -46
rect 2930 -58 2943 -46
rect 2995 -58 3008 -46
rect 3060 -58 3073 -46
rect 2398 -92 2410 -58
rect 2444 -92 2483 -58
rect 2517 -92 2556 -58
rect 2590 -92 2629 -58
rect 2663 -92 2702 -58
rect 2736 -92 2748 -58
rect 2809 -92 2813 -58
rect 3060 -92 3067 -58
rect 2398 -98 2748 -92
rect 2800 -98 2813 -92
rect 2865 -98 2878 -92
rect 2930 -98 2943 -92
rect 2995 -98 3008 -92
rect 3060 -98 3073 -92
rect 3125 -98 3138 -46
rect 3190 -98 3203 -46
rect 3255 -98 3268 -46
rect 3320 -98 3333 -46
rect 3385 -58 3398 -46
rect 3450 -58 3463 -46
rect 3515 -58 3528 -46
rect 3580 -58 3593 -46
rect 3645 -58 3658 -46
rect 3393 -92 3398 -58
rect 3645 -92 3651 -58
rect 3385 -98 3398 -92
rect 3450 -98 3463 -92
rect 3515 -98 3528 -92
rect 3580 -98 3593 -92
rect 3645 -98 3658 -92
rect 3710 -98 3723 -46
rect 3775 -98 3788 -46
rect 3840 -98 3853 -46
rect 3905 -98 3918 -46
rect 3970 -58 3983 -46
rect 4035 -58 4048 -46
rect 4100 -58 4113 -46
rect 4165 -58 4178 -46
rect 4230 -58 4243 -46
rect 4295 -58 4308 -46
rect 3977 -92 3983 -58
rect 4230 -92 4233 -58
rect 4295 -92 4305 -58
rect 3970 -98 3983 -92
rect 4035 -98 4048 -92
rect 4100 -98 4113 -92
rect 4165 -98 4178 -92
rect 4230 -98 4243 -92
rect 4295 -98 4308 -92
rect 4360 -98 4373 -46
rect 4425 -98 4438 -46
rect 4490 -98 4503 -46
rect 4555 -98 4568 -46
rect 4620 -58 4632 -46
rect 4684 -58 4696 -46
rect 4748 -58 4760 -46
rect 4812 -58 4824 -46
rect 4876 -58 4888 -46
rect 4627 -92 4632 -58
rect 4876 -92 4881 -58
rect 4620 -98 4632 -92
rect 4684 -98 4696 -92
rect 4748 -98 4760 -92
rect 4812 -98 4824 -92
rect 4876 -98 4888 -92
rect 4940 -98 4952 -46
rect 5004 -98 5016 -46
rect 5068 -98 5080 -46
rect 5132 -98 5144 -46
rect 5196 -58 5208 -46
rect 5260 -58 5272 -46
rect 5324 -58 5336 -46
rect 5388 -58 5400 -46
rect 5452 -58 5464 -46
rect 5203 -92 5208 -58
rect 5452 -92 5457 -58
rect 5196 -98 5208 -92
rect 5260 -98 5272 -92
rect 5324 -98 5336 -92
rect 5388 -98 5400 -92
rect 5452 -98 5464 -92
rect 5516 -98 5528 -46
rect 5580 -98 5592 -46
rect 5644 -98 5680 -46
rect 5732 -98 5745 -46
rect 5797 -98 5810 -46
rect 5862 -58 5875 -46
rect 5927 -58 5940 -46
rect 5992 -58 6005 -46
rect 6057 -58 6070 -46
rect 6122 -58 6135 -46
rect 5868 -92 5875 -58
rect 6122 -92 6129 -58
rect 5862 -98 5875 -92
rect 5927 -98 5940 -92
rect 5992 -98 6005 -92
rect 6057 -98 6070 -92
rect 6122 -98 6135 -92
rect 6187 -98 6200 -46
rect 6252 -98 6265 -46
rect 6317 -98 6330 -46
rect 6382 -98 6395 -46
rect 6447 -58 6460 -46
rect 6512 -58 6525 -46
rect 6577 -58 6590 -46
rect 6642 -58 6655 -46
rect 6707 -58 6720 -46
rect 6455 -92 6460 -58
rect 6707 -92 6713 -58
rect 6447 -98 6460 -92
rect 6512 -98 6525 -92
rect 6577 -98 6590 -92
rect 6642 -98 6655 -92
rect 6707 -98 6720 -92
rect 6772 -98 6785 -46
rect 6837 -98 6850 -46
rect 6902 -98 6908 -46
rect 7141 -58 7260 -39
rect 7141 -110 7142 -58
rect 7194 -110 7208 -58
rect 7141 -116 7260 -110
rect 7418 453 7464 480
tri 7464 478 7466 480 nw
rect 7504 597 7550 635
rect 7590 1139 7596 1173
rect 7630 1139 7636 1173
tri 7673 1299 7676 1302 se
rect 7676 1299 7682 1317
rect 7673 1293 7682 1299
rect 7716 1299 7722 1317
rect 7762 1389 7808 1401
rect 7762 1355 7768 1389
rect 7802 1355 7808 1389
rect 7762 1317 7808 1355
tri 7722 1299 7725 1302 sw
rect 7716 1293 7725 1299
rect 7673 1229 7682 1241
rect 7716 1229 7725 1241
rect 7673 1173 7725 1177
rect 7673 1171 7682 1173
tri 7673 1168 7676 1171 ne
rect 7590 1101 7636 1139
rect 7590 1067 7596 1101
rect 7630 1067 7636 1101
rect 7590 1029 7636 1067
rect 7590 995 7596 1029
rect 7630 995 7636 1029
rect 7590 957 7636 995
rect 7590 923 7596 957
rect 7630 923 7636 957
rect 7590 885 7636 923
rect 7590 851 7596 885
rect 7630 851 7636 885
rect 7590 813 7636 851
rect 7590 779 7596 813
rect 7630 779 7636 813
rect 7590 741 7636 779
rect 7590 707 7596 741
rect 7630 707 7636 741
rect 7590 669 7636 707
rect 7590 635 7596 669
rect 7630 635 7636 669
rect 7504 563 7510 597
rect 7544 563 7550 597
rect 7504 525 7550 563
rect 7504 491 7510 525
rect 7544 491 7550 525
rect 7418 419 7424 453
rect 7458 419 7464 453
rect 7418 381 7464 419
rect 7418 347 7424 381
rect 7458 347 7464 381
rect 7418 309 7464 347
rect 7418 275 7424 309
rect 7458 275 7464 309
rect 7418 237 7464 275
rect 7418 203 7424 237
rect 7458 203 7464 237
rect 7418 165 7464 203
rect 7418 131 7424 165
rect 7458 131 7464 165
rect 7418 93 7464 131
rect 7418 59 7424 93
rect 7458 59 7464 93
rect 7418 21 7464 59
rect 7418 -13 7424 21
rect 7458 -13 7464 21
rect 7418 -167 7464 -13
rect 7504 453 7550 491
tri 7586 610 7590 614 se
rect 7590 610 7636 635
rect 7676 1139 7682 1171
rect 7716 1171 7725 1173
rect 7716 1139 7722 1171
tri 7722 1168 7725 1171 nw
rect 7762 1283 7768 1317
rect 7802 1283 7808 1317
rect 7848 1389 7894 1401
rect 7848 1355 7854 1389
rect 7888 1355 7894 1389
rect 7848 1317 7894 1355
rect 7762 1245 7808 1283
rect 7762 1211 7768 1245
rect 7802 1211 7808 1245
rect 7762 1173 7808 1211
rect 7676 1101 7722 1139
rect 7676 1067 7682 1101
rect 7716 1067 7722 1101
rect 7676 1029 7722 1067
rect 7676 995 7682 1029
rect 7716 995 7722 1029
rect 7676 957 7722 995
rect 7676 923 7682 957
rect 7716 923 7722 957
rect 7676 885 7722 923
rect 7676 851 7682 885
rect 7716 851 7722 885
rect 7676 813 7722 851
rect 7676 779 7682 813
rect 7716 779 7722 813
rect 7676 741 7722 779
rect 7676 707 7682 741
rect 7716 707 7722 741
rect 7762 1139 7768 1173
rect 7802 1139 7808 1173
tri 7845 1299 7848 1302 se
rect 7848 1299 7854 1317
rect 7845 1293 7854 1299
rect 7888 1300 7894 1317
rect 7929 1400 7990 1406
tri 7990 1400 7996 1406 nw
tri 8939 1400 8945 1406 se
rect 8945 1400 9004 1406
rect 7929 1399 7989 1400
tri 7989 1399 7990 1400 nw
tri 8938 1399 8939 1400 se
rect 8939 1399 9004 1400
tri 7894 1300 7896 1302 sw
rect 7888 1299 7896 1300
tri 7896 1299 7897 1300 sw
rect 7888 1293 7897 1299
rect 7845 1229 7854 1241
rect 7888 1229 7897 1241
rect 7845 1173 7897 1177
rect 7845 1171 7854 1173
tri 7845 1168 7848 1171 ne
rect 7762 1101 7808 1139
rect 7762 1067 7768 1101
rect 7802 1067 7808 1101
rect 7762 1029 7808 1067
rect 7762 995 7768 1029
rect 7802 995 7808 1029
rect 7762 957 7808 995
rect 7762 923 7768 957
rect 7802 923 7808 957
rect 7762 885 7808 923
rect 7762 851 7768 885
rect 7802 851 7808 885
rect 7762 813 7808 851
rect 7762 779 7768 813
rect 7802 779 7808 813
rect 7762 741 7808 779
rect 7676 669 7722 707
rect 7676 635 7682 669
rect 7716 635 7722 669
tri 7636 610 7638 612 sw
rect 7586 604 7638 610
rect 7586 540 7638 552
rect 7586 482 7638 488
tri 7586 480 7588 482 ne
rect 7588 480 7638 482
tri 7588 478 7590 480 ne
rect 7504 419 7510 453
rect 7544 419 7550 453
rect 7504 381 7550 419
rect 7504 347 7510 381
rect 7544 347 7550 381
rect 7504 309 7550 347
rect 7504 275 7510 309
rect 7544 275 7550 309
rect 7504 237 7550 275
rect 7504 203 7510 237
rect 7544 203 7550 237
rect 7504 165 7550 203
rect 7504 131 7510 165
rect 7544 131 7550 165
rect 7504 93 7550 131
rect 7504 59 7510 93
rect 7544 59 7550 93
rect 7504 21 7550 59
rect 7504 -13 7510 21
rect 7544 -13 7550 21
rect 7504 -25 7550 -13
rect 7590 453 7636 480
tri 7636 478 7638 480 nw
rect 7676 597 7722 635
rect 7676 563 7682 597
rect 7716 563 7722 597
tri 7758 720 7762 724 se
rect 7762 720 7768 741
rect 7758 714 7768 720
rect 7802 720 7808 741
rect 7848 1139 7854 1171
rect 7888 1171 7897 1173
rect 7888 1139 7894 1171
tri 7894 1168 7897 1171 nw
rect 7848 1101 7894 1139
rect 7848 1067 7854 1101
rect 7888 1067 7894 1101
rect 7848 1029 7894 1067
rect 7848 995 7854 1029
rect 7888 995 7894 1029
rect 7848 957 7894 995
rect 7848 923 7854 957
rect 7888 923 7894 957
rect 7848 885 7894 923
rect 7848 851 7854 885
rect 7888 851 7894 885
rect 7848 813 7894 851
rect 7848 779 7854 813
rect 7888 779 7894 813
rect 7848 741 7894 779
tri 7808 720 7810 722 sw
rect 7802 714 7810 720
rect 7758 650 7768 662
rect 7802 650 7810 662
rect 7758 597 7810 598
rect 7758 592 7768 597
tri 7758 590 7760 592 ne
rect 7760 590 7768 592
tri 7760 588 7762 590 ne
rect 7676 525 7722 563
rect 7676 491 7682 525
rect 7716 491 7722 525
rect 7590 419 7596 453
rect 7630 419 7636 453
rect 7590 381 7636 419
rect 7590 347 7596 381
rect 7630 347 7636 381
rect 7590 309 7636 347
rect 7590 275 7596 309
rect 7630 275 7636 309
rect 7590 237 7636 275
rect 7590 203 7596 237
rect 7630 203 7636 237
rect 7590 165 7636 203
rect 7590 131 7596 165
rect 7630 131 7636 165
rect 7590 93 7636 131
rect 7590 59 7596 93
rect 7630 59 7636 93
rect 7590 21 7636 59
rect 7590 -13 7596 21
rect 7630 -13 7636 21
tri 7464 -167 7489 -142 sw
tri 7565 -167 7590 -142 se
rect 7590 -167 7636 -13
rect 7676 453 7722 491
rect 7676 419 7682 453
rect 7716 419 7722 453
rect 7676 381 7722 419
rect 7676 347 7682 381
rect 7716 347 7722 381
rect 7676 309 7722 347
rect 7676 275 7682 309
rect 7716 275 7722 309
rect 7676 237 7722 275
rect 7676 203 7682 237
rect 7716 203 7722 237
rect 7676 165 7722 203
rect 7676 131 7682 165
rect 7716 131 7722 165
rect 7676 93 7722 131
rect 7676 59 7682 93
rect 7716 59 7722 93
rect 7676 21 7722 59
rect 7676 -13 7682 21
rect 7716 -13 7722 21
rect 7676 -25 7722 -13
rect 7762 563 7768 590
rect 7802 590 7810 597
rect 7802 563 7808 590
tri 7808 588 7810 590 nw
rect 7848 707 7854 741
rect 7888 707 7894 741
rect 7848 669 7894 707
rect 7848 635 7854 669
rect 7888 635 7894 669
rect 7848 597 7894 635
rect 7762 525 7808 563
rect 7762 491 7768 525
rect 7802 491 7808 525
rect 7762 453 7808 491
rect 7762 419 7768 453
rect 7802 419 7808 453
rect 7762 381 7808 419
rect 7762 347 7768 381
rect 7802 347 7808 381
rect 7762 309 7808 347
rect 7762 275 7768 309
rect 7802 275 7808 309
rect 7762 237 7808 275
rect 7762 203 7768 237
rect 7802 203 7808 237
rect 7762 165 7808 203
rect 7762 131 7768 165
rect 7802 131 7808 165
rect 7762 93 7808 131
rect 7762 59 7768 93
rect 7802 59 7808 93
rect 7762 21 7808 59
rect 7762 -13 7768 21
rect 7802 -13 7808 21
tri 7636 -167 7661 -142 sw
tri 7737 -167 7762 -142 se
rect 7762 -167 7808 -13
rect 7848 563 7854 597
rect 7888 563 7894 597
rect 7848 525 7894 563
rect 7848 491 7854 525
rect 7888 491 7894 525
rect 7848 453 7894 491
rect 7848 419 7854 453
rect 7888 419 7894 453
rect 7848 381 7894 419
rect 7929 530 7981 1399
tri 7981 1391 7989 1399 nw
tri 8930 1391 8938 1399 se
rect 8938 1391 9004 1399
tri 8926 1387 8930 1391 se
rect 8930 1387 9004 1391
tri 8041 1378 8050 1387 se
rect 8050 1378 9004 1387
tri 8018 1355 8041 1378 se
rect 8041 1362 9004 1378
rect 8041 1355 8997 1362
tri 8997 1355 9004 1362 nw
tri 9034 2275 9035 2276 se
rect 9035 2275 11840 2276
tri 11840 2275 11841 2276 nw
rect 9034 2265 11830 2275
tri 11830 2265 11840 2275 nw
rect 9034 2252 11817 2265
tri 11817 2252 11830 2265 nw
rect 9034 2236 9104 2252
tri 9104 2236 9120 2252 nw
rect 9034 2231 9099 2236
tri 9099 2231 9104 2236 nw
rect 9034 2222 9090 2231
tri 9090 2222 9099 2231 nw
rect 7929 466 7981 478
rect 7929 408 7981 414
tri 8010 1347 8018 1355 se
rect 8018 1347 8989 1355
tri 8989 1347 8997 1355 nw
rect 8010 1335 8977 1347
tri 8977 1335 8989 1347 nw
rect 8010 1321 8074 1335
tri 8074 1321 8088 1335 nw
tri 9026 1321 9034 1329 se
rect 9034 1321 9086 2222
tri 9086 2218 9090 2222 nw
tri 9148 2218 9152 2222 se
rect 9152 2218 10607 2222
tri 9143 2213 9148 2218 se
rect 9148 2213 10607 2218
rect 8010 1315 8068 1321
tri 8068 1315 8074 1321 nw
tri 9020 1315 9026 1321 se
rect 9026 1315 9086 1321
rect 8010 446 8062 1315
tri 8062 1309 8068 1315 nw
tri 9014 1309 9020 1315 se
rect 9020 1309 9086 1315
tri 9008 1303 9014 1309 se
rect 9014 1303 9086 1309
tri 8126 1300 8129 1303 se
rect 8129 1300 9086 1303
tri 8092 1266 8126 1300 se
rect 8126 1291 9086 1300
rect 8126 1266 9061 1291
tri 9061 1266 9086 1291 nw
tri 9118 2188 9143 2213 se
rect 9143 2188 10607 2213
rect 9118 2170 10607 2188
rect 10659 2170 10671 2222
rect 10723 2170 10731 2222
tri 11884 2170 11886 2172 se
rect 11886 2170 11938 2883
tri 11938 2875 11946 2883 nw
rect 12241 2849 16569 2855
rect 12241 2815 12253 2849
rect 12287 2815 12325 2849
rect 12359 2815 12397 2849
rect 12431 2815 12469 2849
rect 12503 2815 12542 2849
rect 12576 2815 12615 2849
rect 12649 2815 12688 2849
rect 12722 2815 12761 2849
rect 12795 2815 12834 2849
rect 12868 2815 12907 2849
rect 12941 2815 12980 2849
rect 13014 2815 13053 2849
rect 13087 2815 13126 2849
rect 13160 2815 13199 2849
rect 13233 2815 13272 2849
rect 13306 2815 13345 2849
rect 13379 2815 13418 2849
rect 13452 2815 13491 2849
rect 13525 2815 13564 2849
rect 13598 2815 13637 2849
rect 13671 2815 13710 2849
rect 13744 2815 13783 2849
rect 13817 2815 13856 2849
rect 13890 2815 13929 2849
rect 13963 2815 14002 2849
rect 14036 2815 14075 2849
rect 14109 2815 14148 2849
rect 14182 2815 14221 2849
rect 14255 2815 14294 2849
rect 14328 2815 14367 2849
rect 14401 2815 14440 2849
rect 14474 2815 14513 2849
rect 14547 2815 14586 2849
rect 14620 2815 14659 2849
rect 14693 2815 14732 2849
rect 14766 2815 14805 2849
rect 14839 2815 14878 2849
rect 14912 2815 14951 2849
rect 14985 2815 15024 2849
rect 15058 2815 15097 2849
rect 15131 2815 15170 2849
rect 15204 2815 15243 2849
rect 15277 2815 15316 2849
rect 15350 2815 15389 2849
rect 15423 2815 15462 2849
rect 15496 2815 15535 2849
rect 15569 2815 15608 2849
rect 15642 2815 15681 2849
rect 15715 2815 15754 2849
rect 15788 2815 15827 2849
rect 15861 2815 15900 2849
rect 15934 2815 15973 2849
rect 16007 2815 16046 2849
rect 16080 2815 16119 2849
rect 16153 2815 16192 2849
rect 16226 2815 16265 2849
rect 16299 2815 16338 2849
rect 16372 2815 16569 2849
rect 16758 2831 16764 2883
rect 16816 2831 16828 2883
rect 16880 2831 18066 2883
rect 18118 2831 18132 2883
rect 18184 2831 18190 2883
rect 18405 2849 18417 2883
rect 18451 2849 18497 2883
rect 18531 2849 18577 2883
rect 18611 2849 18657 2883
rect 18691 2849 18737 2883
rect 18771 2849 18817 2883
rect 18851 2849 18897 2883
rect 18931 2849 18953 2883
rect 19011 2849 19044 2883
rect 18405 2843 18953 2849
rect 19005 2843 19044 2849
rect 19096 2843 19102 2895
rect 12241 2809 16569 2815
tri 16370 2782 16397 2809 ne
rect 16397 2782 16569 2809
tri 16397 2778 16401 2782 ne
rect 16401 2778 16569 2782
tri 16401 2776 16403 2778 ne
rect 16403 2776 16569 2778
tri 16403 2775 16404 2776 ne
rect 16404 2742 16410 2776
rect 16444 2742 16569 2776
rect 16404 2703 16569 2742
rect 17126 2737 17132 2789
rect 17184 2737 17196 2789
rect 17248 2778 18053 2789
rect 17248 2744 17935 2778
rect 17969 2744 18007 2778
rect 18041 2744 18053 2778
rect 17248 2738 18053 2744
rect 17248 2737 18052 2738
tri 18052 2737 18053 2738 nw
rect 16404 2669 16410 2703
rect 16444 2669 16569 2703
rect 16404 2638 16569 2669
rect 16767 2640 16773 2692
rect 16825 2640 16837 2692
rect 16889 2640 18218 2692
rect 18270 2640 18282 2692
rect 18334 2640 18340 2692
rect 18395 2687 18401 2739
rect 18453 2727 18492 2739
rect 18544 2727 19102 2739
rect 18464 2693 18492 2727
rect 18544 2693 18588 2727
rect 18622 2693 18666 2727
rect 18700 2693 18744 2727
rect 18778 2693 18822 2727
rect 18856 2693 18900 2727
rect 18934 2693 18978 2727
rect 19012 2693 19056 2727
rect 19090 2693 19102 2727
rect 18453 2687 18492 2693
rect 18544 2687 19102 2693
tri 16569 2638 16571 2640 sw
rect 16404 2630 16571 2638
rect 16404 2596 16410 2630
rect 16444 2612 16571 2630
tri 16571 2612 16597 2638 sw
rect 16444 2606 16597 2612
tri 16597 2606 16603 2612 sw
rect 16444 2596 16603 2606
rect 16404 2585 16603 2596
tri 16603 2585 16624 2606 sw
rect 16404 2579 17258 2585
rect 16404 2557 16601 2579
rect 16404 2523 16410 2557
rect 16444 2545 16601 2557
rect 16635 2545 16675 2579
rect 16709 2545 16749 2579
rect 16783 2545 16823 2579
rect 16857 2545 16897 2579
rect 16931 2545 16971 2579
rect 17005 2545 17045 2579
rect 17079 2545 17119 2579
rect 17153 2545 17192 2579
rect 17226 2545 17258 2579
rect 17286 2566 17298 2612
tri 17286 2560 17292 2566 ne
rect 17292 2560 17298 2566
rect 17350 2560 17362 2612
rect 17414 2606 19086 2612
rect 17414 2572 17805 2606
rect 17839 2572 17878 2606
rect 17912 2572 17951 2606
rect 17985 2572 18024 2606
rect 18058 2572 18097 2606
rect 18131 2572 18170 2606
rect 18204 2572 18243 2606
rect 18277 2572 18316 2606
rect 18350 2572 18389 2606
rect 18423 2572 18462 2606
rect 18496 2572 18535 2606
rect 18569 2572 18608 2606
rect 18642 2572 18680 2606
rect 18714 2572 18752 2606
rect 18786 2572 18824 2606
rect 18858 2572 18896 2606
rect 18930 2572 18968 2606
rect 19002 2572 19040 2606
rect 19074 2572 19086 2606
rect 17414 2566 19086 2572
rect 17414 2560 17421 2566
tri 17421 2560 17427 2566 nw
rect 16444 2523 17258 2545
rect 16404 2507 17258 2523
rect 16404 2484 16601 2507
rect 16404 2450 16410 2484
rect 16444 2473 16601 2484
rect 16635 2473 16675 2507
rect 16709 2473 16749 2507
rect 16783 2473 16823 2507
rect 16857 2473 16897 2507
rect 16931 2473 16971 2507
rect 17005 2473 17045 2507
rect 17079 2473 17119 2507
rect 17153 2473 17192 2507
rect 17226 2473 17258 2507
rect 16444 2450 17258 2473
rect 16404 2435 17258 2450
rect 16404 2411 16601 2435
rect 16404 2377 16410 2411
rect 16444 2401 16601 2411
rect 16635 2401 16675 2435
rect 16709 2401 16749 2435
rect 16783 2401 16823 2435
rect 16857 2401 16897 2435
rect 16931 2401 16971 2435
rect 17005 2401 17045 2435
rect 17079 2401 17119 2435
rect 17153 2401 17192 2435
rect 17226 2401 17258 2435
rect 16444 2395 17258 2401
rect 16444 2388 16963 2395
tri 16963 2388 16970 2395 nw
rect 16444 2377 16925 2388
rect 16404 2363 16925 2377
rect 16404 2338 16590 2363
rect 16404 2304 16410 2338
rect 16444 2329 16590 2338
rect 16624 2329 16662 2363
rect 16696 2329 16734 2363
rect 16768 2329 16806 2363
rect 16840 2350 16925 2363
tri 16925 2350 16963 2388 nw
rect 16840 2329 16891 2350
rect 16444 2316 16891 2329
tri 16891 2316 16925 2350 nw
rect 16444 2304 16874 2316
rect 16404 2276 16874 2304
tri 16874 2299 16891 2316 nw
rect 16404 2265 16590 2276
tri 16399 2231 16404 2236 se
rect 16404 2231 16410 2265
rect 16444 2242 16590 2265
rect 16624 2242 16662 2276
rect 16696 2242 16734 2276
rect 16768 2242 16806 2276
rect 16840 2242 16874 2276
rect 16444 2231 16874 2242
tri 16374 2206 16399 2231 se
rect 16399 2206 16874 2231
tri 16360 2192 16374 2206 se
rect 16374 2192 16874 2206
rect 9118 2158 9192 2170
tri 9192 2158 9204 2170 nw
tri 11872 2158 11884 2170 se
rect 11884 2158 11938 2170
tri 16326 2158 16360 2192 se
rect 16360 2158 16410 2192
rect 16444 2188 16874 2192
rect 16444 2158 16590 2188
rect 9118 2154 9188 2158
tri 9188 2154 9192 2158 nw
tri 11868 2154 11872 2158 se
rect 11872 2154 11938 2158
tri 16322 2154 16326 2158 se
rect 16326 2154 16590 2158
rect 16624 2154 16662 2188
rect 16696 2154 16734 2188
rect 16768 2154 16806 2188
rect 16840 2154 16874 2188
rect 9118 2138 9172 2154
tri 9172 2138 9188 2154 nw
tri 11852 2138 11868 2154 se
rect 11868 2138 11938 2154
rect 7848 347 7854 381
rect 7888 347 7894 381
rect 7848 309 7894 347
rect 8010 382 8062 394
rect 8010 324 8062 330
tri 8090 1264 8092 1266 se
rect 8092 1264 9059 1266
tri 9059 1264 9061 1266 nw
rect 8090 1251 9046 1264
tri 9046 1251 9059 1264 nw
rect 8090 1250 8167 1251
tri 8167 1250 8168 1251 nw
rect 7848 275 7854 309
rect 7888 275 7894 309
rect 7848 237 7894 275
rect 7848 203 7854 237
rect 7888 203 7894 237
rect 7848 165 7894 203
rect 8090 312 8142 1250
tri 8142 1225 8167 1250 nw
rect 9118 1216 9170 2138
tri 9170 2136 9172 2138 nw
tri 9233 2136 9235 2138 se
rect 9235 2136 9929 2138
tri 9231 2134 9233 2136 se
rect 9233 2134 9929 2136
tri 9216 2119 9231 2134 se
rect 9231 2119 9929 2134
tri 9201 2104 9216 2119 se
rect 9216 2104 9929 2119
rect 9201 2086 9929 2104
rect 9981 2086 9993 2138
rect 10045 2115 11938 2138
tri 16302 2134 16322 2154 se
rect 16322 2134 16874 2154
tri 16287 2119 16302 2134 se
rect 16302 2119 16874 2134
rect 10045 2086 11909 2115
tri 11909 2086 11938 2115 nw
tri 16254 2086 16287 2119 se
rect 16287 2086 16410 2119
rect 9201 2085 9286 2086
tri 9286 2085 9287 2086 nw
tri 16253 2085 16254 2086 se
rect 16254 2085 16410 2086
rect 16444 2100 16874 2119
tri 19871 2100 19902 2131 se
rect 19902 2100 19954 2937
rect 16444 2085 16590 2100
rect 9201 2066 9267 2085
tri 9267 2066 9286 2085 nw
tri 16234 2066 16253 2085 se
rect 16253 2066 16590 2085
rect 16624 2066 16662 2100
rect 16696 2066 16734 2100
rect 16768 2066 16806 2100
rect 16840 2066 16874 2100
tri 19859 2088 19871 2100 se
rect 19871 2088 19954 2100
rect 9201 2062 9263 2066
tri 9263 2062 9267 2066 nw
tri 16230 2062 16234 2066 se
rect 16234 2062 16874 2066
tri 16874 2062 16900 2088 sw
tri 19833 2062 19859 2088 se
rect 19859 2062 19954 2088
rect 9201 2053 9254 2062
tri 9254 2053 9263 2062 nw
tri 16221 2053 16230 2062 se
rect 16230 2053 16900 2062
rect 9201 1984 9253 2053
tri 9253 2052 9254 2053 nw
rect 10488 2052 16900 2053
rect 10488 2047 10775 2052
rect 9201 1920 9253 1932
rect 9201 1862 9253 1868
rect 9401 2013 9454 2019
rect 9453 1961 9454 2013
rect 10488 2013 10500 2047
rect 10534 2013 10573 2047
rect 10607 2013 10646 2047
rect 10680 2013 10719 2047
rect 10753 2013 10775 2047
rect 10488 2000 10775 2013
rect 10827 2000 10839 2052
rect 10891 2047 10927 2052
rect 10899 2013 10927 2047
rect 10891 2000 10927 2013
rect 10979 2000 10992 2052
rect 11044 2000 11057 2052
rect 11109 2047 11122 2052
rect 11174 2047 11187 2052
rect 11239 2047 11252 2052
rect 11304 2047 11317 2052
rect 11369 2047 11382 2052
rect 11434 2047 11447 2052
rect 11116 2013 11122 2047
rect 11369 2013 11370 2047
rect 11434 2013 11442 2047
rect 11109 2000 11122 2013
rect 11174 2000 11187 2013
rect 11239 2000 11252 2013
rect 11304 2000 11317 2013
rect 11369 2000 11382 2013
rect 11434 2000 11447 2013
rect 11499 2000 11512 2052
rect 11564 2000 11577 2052
rect 11629 2000 11642 2052
rect 11694 2000 11707 2052
rect 11759 2047 11772 2052
rect 11824 2047 11837 2052
rect 11889 2047 11901 2052
rect 11953 2047 11965 2052
rect 12017 2047 12029 2052
rect 12081 2047 12093 2052
rect 11764 2013 11772 2047
rect 11836 2013 11837 2047
rect 12017 2013 12018 2047
rect 12081 2013 12090 2047
rect 11759 2000 11772 2013
rect 11824 2000 11837 2013
rect 11889 2000 11901 2013
rect 11953 2000 11965 2013
rect 12017 2000 12029 2013
rect 12081 2000 12093 2013
rect 12145 2000 12157 2052
rect 12209 2000 12221 2052
rect 12273 2000 12285 2052
rect 12337 2047 12349 2052
rect 12401 2047 12413 2052
rect 12465 2047 12477 2052
rect 12529 2047 12541 2052
rect 12593 2047 12605 2052
rect 12657 2047 12669 2052
rect 12340 2013 12349 2047
rect 12412 2013 12413 2047
rect 12593 2013 12594 2047
rect 12657 2013 12666 2047
rect 12337 2000 12349 2013
rect 12401 2000 12413 2013
rect 12465 2000 12477 2013
rect 12529 2000 12541 2013
rect 12593 2000 12605 2013
rect 12657 2000 12669 2013
rect 12721 2000 12733 2052
rect 12785 2000 12797 2052
rect 12849 2000 12861 2052
rect 12913 2047 12925 2052
rect 12977 2047 12989 2052
rect 13041 2047 13053 2052
rect 13105 2047 13117 2052
rect 13169 2047 13181 2052
rect 13233 2047 13245 2052
rect 12916 2013 12925 2047
rect 12988 2013 12989 2047
rect 13169 2013 13170 2047
rect 13233 2013 13242 2047
rect 12913 2000 12925 2013
rect 12977 2000 12989 2013
rect 13041 2000 13053 2013
rect 13105 2000 13117 2013
rect 13169 2000 13181 2013
rect 13233 2000 13245 2013
rect 13297 2000 13309 2052
rect 13361 2000 13373 2052
rect 13425 2000 13437 2052
rect 13489 2051 16900 2052
tri 16900 2051 16911 2062 sw
tri 19822 2051 19833 2062 se
rect 19833 2051 19954 2062
rect 19996 2926 20042 2961
rect 19996 2892 20002 2926
rect 20036 2892 20042 2926
tri 20042 2913 20127 2998 nw
rect 19996 2854 20042 2892
rect 19996 2820 20002 2854
rect 20036 2820 20042 2854
rect 19996 2782 20042 2820
rect 19996 2748 20002 2782
rect 20036 2748 20042 2782
rect 19996 2710 20042 2748
rect 19996 2676 20002 2710
rect 20036 2676 20042 2710
rect 19996 2638 20042 2676
rect 19996 2604 20002 2638
rect 20036 2604 20042 2638
rect 19996 2566 20042 2604
rect 19996 2532 20002 2566
rect 20036 2532 20042 2566
rect 19996 2494 20042 2532
rect 19996 2460 20002 2494
rect 20036 2460 20042 2494
rect 19996 2422 20042 2460
rect 19996 2388 20002 2422
rect 20036 2388 20042 2422
rect 19996 2350 20042 2388
rect 19996 2316 20002 2350
rect 20036 2316 20042 2350
rect 19996 2278 20042 2316
rect 19996 2244 20002 2278
rect 20036 2244 20042 2278
rect 19996 2206 20042 2244
rect 19996 2172 20002 2206
rect 20036 2172 20042 2206
rect 19996 2134 20042 2172
rect 19996 2100 20002 2134
rect 20036 2100 20042 2134
rect 19996 2062 20042 2100
rect 13489 2047 16911 2051
rect 13492 2013 13530 2047
rect 13564 2013 13602 2047
rect 13636 2013 13674 2047
rect 13708 2013 13746 2047
rect 13780 2013 13818 2047
rect 13852 2013 13890 2047
rect 13924 2013 13962 2047
rect 13996 2013 14034 2047
rect 14068 2013 14106 2047
rect 14140 2013 14178 2047
rect 14212 2013 14250 2047
rect 14284 2013 14322 2047
rect 14356 2013 14394 2047
rect 14428 2013 14466 2047
rect 14500 2013 14538 2047
rect 14572 2013 14610 2047
rect 14644 2013 14682 2047
rect 14716 2013 14754 2047
rect 14788 2013 14826 2047
rect 14860 2013 14898 2047
rect 14932 2013 14970 2047
rect 15004 2013 15042 2047
rect 15076 2013 15114 2047
rect 15148 2013 15186 2047
rect 15220 2013 15258 2047
rect 15292 2013 15330 2047
rect 15364 2013 15402 2047
rect 15436 2013 15474 2047
rect 15508 2013 15546 2047
rect 15580 2013 15618 2047
rect 15652 2013 15690 2047
rect 15724 2013 15762 2047
rect 15796 2013 15834 2047
rect 15868 2013 15906 2047
rect 15940 2013 15978 2047
rect 16012 2013 16050 2047
rect 16084 2013 16122 2047
rect 16156 2013 16194 2047
rect 16228 2013 16266 2047
rect 16300 2013 16338 2047
rect 16372 2028 16911 2047
tri 16911 2028 16934 2051 sw
rect 19996 2028 20002 2062
rect 20036 2028 20042 2062
tri 25297 2047 25325 2075 se
rect 25325 2047 25334 2075
rect 16372 2025 16934 2028
tri 16934 2025 16937 2028 sw
rect 16372 2013 16937 2025
rect 13489 2012 16937 2013
rect 13489 2000 16590 2012
tri 12587 1978 12609 2000 ne
rect 12609 1978 16590 2000
rect 16624 1978 16662 2012
rect 16696 1978 16734 2012
rect 16768 1978 16806 2012
rect 16840 2007 16937 2012
tri 16937 2007 16955 2025 sw
rect 16840 2000 16955 2007
tri 16955 2000 16962 2007 sw
rect 16840 1991 16962 2000
tri 16962 1991 16971 2000 sw
rect 16840 1990 16971 1991
tri 16971 1990 16972 1991 sw
rect 19996 1990 20042 2028
rect 16840 1978 16972 1990
rect 9401 1953 9411 1961
rect 9445 1953 9454 1961
tri 12609 1956 12631 1978 ne
rect 12631 1956 16972 1978
tri 16972 1956 17006 1990 sw
rect 19996 1956 20002 1990
rect 20036 1956 20042 1990
rect 24033 2025 24695 2031
rect 24033 1991 24045 2025
rect 24079 1991 24121 2025
rect 24155 1991 24197 2025
rect 24231 1991 24273 2025
rect 24307 1991 24349 2025
rect 24383 1991 24424 2025
rect 24458 1991 24499 2025
rect 24533 1991 24574 2025
rect 24608 1991 24649 2025
rect 24683 1991 24695 2025
rect 24033 1985 24695 1991
rect 25297 2023 25334 2047
rect 25386 2023 25398 2075
rect 25450 2023 25456 2075
rect 9401 1932 9454 1953
rect 9453 1880 9454 1932
tri 12631 1927 12660 1956 ne
rect 12660 1927 17006 1956
rect 9401 1874 9411 1880
rect 9445 1874 9454 1880
rect 9401 1850 9454 1874
rect 9453 1798 9454 1850
rect 9401 1795 9411 1798
rect 9445 1795 9454 1798
rect 9401 1792 9454 1795
tri 9401 1788 9405 1792 ne
rect 9405 1791 9454 1792
rect 9203 1774 9255 1780
rect 9203 1710 9255 1722
rect 9203 1300 9255 1658
rect 9405 1750 9451 1791
tri 9451 1788 9454 1791 nw
rect 9722 1918 12417 1927
rect 9722 1884 9734 1918
rect 9768 1884 9808 1918
rect 9842 1884 9882 1918
rect 9916 1884 9956 1918
rect 9990 1884 10030 1918
rect 10064 1884 10104 1918
rect 10138 1884 10178 1918
rect 10212 1884 10252 1918
rect 10286 1884 10326 1918
rect 10360 1884 10400 1918
rect 10434 1884 10473 1918
rect 10507 1884 10546 1918
rect 10580 1884 10619 1918
rect 10653 1884 10692 1918
rect 10726 1885 10765 1918
rect 10799 1885 10838 1918
rect 10872 1885 10911 1918
rect 10945 1885 10984 1918
rect 11018 1885 11057 1918
rect 11091 1885 11130 1918
rect 11164 1885 11203 1918
rect 11237 1885 11276 1918
rect 11310 1885 11349 1918
rect 11383 1885 11422 1918
rect 11456 1885 11495 1918
rect 11529 1885 11568 1918
rect 11602 1885 11641 1918
rect 11675 1885 11714 1918
rect 11748 1885 11787 1918
rect 11821 1885 11860 1918
rect 11894 1885 11933 1918
rect 11967 1885 12006 1918
rect 12040 1885 12079 1918
rect 12113 1885 12152 1918
rect 12186 1885 12225 1918
rect 12259 1885 12298 1918
rect 12332 1885 12371 1918
rect 12405 1885 12417 1918
tri 12660 1911 12676 1927 ne
rect 12676 1924 17006 1927
tri 17006 1924 17038 1956 sw
tri 19967 1924 19996 1953 se
rect 19996 1924 20042 1956
rect 24462 1927 24664 1938
rect 12676 1911 17038 1924
rect 10726 1884 10762 1885
rect 9722 1836 10762 1884
rect 9722 1802 9734 1836
rect 9768 1802 9808 1836
rect 9842 1802 9882 1836
rect 9916 1802 9956 1836
rect 9990 1802 10030 1836
rect 10064 1802 10104 1836
rect 10138 1802 10178 1836
rect 10212 1802 10252 1836
rect 10286 1802 10326 1836
rect 10360 1802 10400 1836
rect 10434 1802 10473 1836
rect 10507 1802 10546 1836
rect 10580 1802 10619 1836
rect 10653 1802 10692 1836
rect 10726 1833 10762 1836
rect 10814 1833 10829 1885
rect 10881 1833 10896 1885
rect 10948 1833 10963 1885
rect 11018 1884 11030 1885
rect 11091 1884 11097 1885
rect 11417 1884 11422 1885
rect 11484 1884 11495 1885
rect 11015 1836 11030 1884
rect 11082 1836 11097 1884
rect 11149 1836 11164 1884
rect 11216 1836 11231 1884
rect 11283 1836 11298 1884
rect 11350 1836 11365 1884
rect 11417 1836 11432 1884
rect 11484 1836 11499 1884
rect 11018 1833 11030 1836
rect 11091 1833 11097 1836
rect 11417 1833 11422 1836
rect 11484 1833 11495 1836
rect 11551 1833 11566 1885
rect 11618 1833 11633 1885
rect 11685 1833 11699 1885
rect 11751 1833 11765 1885
rect 11821 1884 11831 1885
rect 11894 1884 11897 1885
rect 12147 1884 12152 1885
rect 12213 1884 12225 1885
rect 11817 1836 11831 1884
rect 11883 1836 11897 1884
rect 11949 1836 11963 1884
rect 12015 1836 12029 1884
rect 12081 1836 12095 1884
rect 12147 1836 12161 1884
rect 12213 1836 12227 1884
rect 11821 1833 11831 1836
rect 11894 1833 11897 1836
rect 12147 1833 12152 1836
rect 12213 1833 12225 1836
rect 12279 1833 12293 1885
rect 12345 1833 12359 1885
rect 12411 1833 12417 1885
tri 12676 1877 12710 1911 ne
rect 12710 1877 12756 1911
rect 12790 1877 12830 1911
rect 12864 1877 12904 1911
rect 12938 1877 12978 1911
rect 13012 1877 13052 1911
rect 13086 1877 13126 1911
rect 13160 1877 13200 1911
rect 13234 1877 13274 1911
rect 13308 1877 13348 1911
rect 13382 1877 13422 1911
rect 13456 1877 13496 1911
rect 13530 1877 13569 1911
rect 13603 1877 13642 1911
rect 13676 1877 13715 1911
rect 13749 1877 13788 1911
rect 13822 1877 13861 1911
rect 13895 1877 13934 1911
rect 13968 1877 14007 1911
rect 14041 1877 14080 1911
rect 14114 1877 14153 1911
rect 14187 1877 14226 1911
rect 14260 1877 14299 1911
rect 14333 1877 14372 1911
rect 14406 1877 14445 1911
rect 14479 1877 14518 1911
rect 14552 1877 14591 1911
rect 14625 1877 14664 1911
rect 14698 1877 14737 1911
rect 14771 1877 14810 1911
rect 14844 1877 14883 1911
rect 14917 1877 14956 1911
rect 14990 1877 15029 1911
rect 15063 1877 15102 1911
rect 15136 1877 15175 1911
rect 15209 1877 15248 1911
rect 15282 1877 15321 1911
rect 15355 1877 15394 1911
rect 15428 1877 15467 1911
rect 15501 1877 15540 1911
rect 15574 1877 15613 1911
rect 15647 1877 15686 1911
rect 15720 1877 15759 1911
rect 15793 1877 15832 1911
rect 15866 1877 15905 1911
rect 15939 1877 15978 1911
rect 16012 1877 16051 1911
rect 16085 1877 16124 1911
rect 16158 1877 16197 1911
rect 16231 1877 16270 1911
rect 16304 1877 16343 1911
rect 16377 1877 16416 1911
rect 16450 1877 16489 1911
rect 16523 1877 16562 1911
rect 16596 1877 16635 1911
rect 16669 1877 16708 1911
rect 16742 1909 17038 1911
tri 17038 1909 17053 1924 sw
rect 16742 1902 19197 1909
rect 16742 1877 16847 1902
tri 12710 1868 12719 1877 ne
rect 12719 1868 16847 1877
rect 16881 1868 16919 1902
rect 16953 1868 16991 1902
rect 17025 1868 17063 1902
rect 17097 1868 17135 1902
rect 17169 1868 17207 1902
rect 17241 1868 17279 1902
rect 17313 1868 17351 1902
rect 17385 1868 17423 1902
rect 17457 1868 17495 1902
rect 17529 1868 17567 1902
rect 17601 1868 17639 1902
rect 17673 1868 17711 1902
rect 17745 1868 17783 1902
rect 17817 1868 17855 1902
rect 17889 1868 17927 1902
rect 17961 1868 17999 1902
rect 18033 1868 18071 1902
rect 18105 1868 18143 1902
rect 18177 1868 18215 1902
rect 18249 1868 18287 1902
rect 18321 1868 18359 1902
rect 18393 1868 18431 1902
rect 18465 1868 18503 1902
rect 18537 1868 18575 1902
rect 18609 1868 18647 1902
rect 18681 1868 18719 1902
rect 18753 1868 18791 1902
rect 18825 1868 18863 1902
rect 18897 1868 18935 1902
rect 18969 1868 19007 1902
rect 19041 1868 19079 1902
rect 19113 1868 19151 1902
rect 19185 1868 19197 1902
tri 12719 1846 12741 1868 ne
rect 12741 1846 19197 1868
tri 12741 1843 12744 1846 ne
rect 12744 1844 19197 1846
rect 12744 1843 16450 1844
tri 16450 1843 16451 1844 nw
tri 16770 1843 16771 1844 ne
rect 16771 1843 19197 1844
rect 10726 1805 10765 1833
rect 10799 1805 10838 1833
rect 10872 1805 10911 1833
rect 10945 1805 10984 1833
rect 11018 1805 11057 1833
rect 11091 1805 11130 1833
rect 11164 1805 11203 1833
rect 11237 1805 11276 1833
rect 11310 1805 11349 1833
rect 11383 1805 11422 1833
rect 11456 1805 11495 1833
rect 11529 1805 11568 1833
rect 11602 1805 11641 1833
rect 11675 1805 11714 1833
rect 11748 1805 11787 1833
rect 11821 1805 11860 1833
rect 11894 1805 11933 1833
rect 11967 1805 12006 1833
rect 12040 1805 12079 1833
rect 12113 1805 12152 1833
rect 12186 1805 12225 1833
rect 12259 1805 12298 1833
rect 12332 1805 12371 1833
rect 12405 1805 12417 1833
tri 16771 1816 16798 1843 ne
rect 16798 1816 19197 1843
rect 10726 1802 10762 1805
rect 9405 1716 9411 1750
rect 9445 1716 9451 1750
rect 9405 1671 9451 1716
rect 9405 1637 9411 1671
rect 9445 1637 9451 1671
rect 9405 1592 9451 1637
rect 9405 1558 9411 1592
rect 9445 1558 9451 1592
rect 9405 1513 9451 1558
rect 9722 1754 10762 1802
rect 9722 1720 9734 1754
rect 9768 1720 9808 1754
rect 9842 1720 9882 1754
rect 9916 1720 9956 1754
rect 9990 1720 10030 1754
rect 10064 1720 10104 1754
rect 10138 1720 10178 1754
rect 10212 1720 10252 1754
rect 10286 1720 10326 1754
rect 10360 1720 10400 1754
rect 10434 1720 10473 1754
rect 10507 1720 10546 1754
rect 10580 1720 10619 1754
rect 10653 1720 10692 1754
rect 10726 1753 10762 1754
rect 10814 1753 10829 1805
rect 10881 1753 10896 1805
rect 10948 1753 10963 1805
rect 11018 1802 11030 1805
rect 11091 1802 11097 1805
rect 11417 1802 11422 1805
rect 11484 1802 11495 1805
rect 11015 1754 11030 1802
rect 11082 1754 11097 1802
rect 11149 1754 11164 1802
rect 11216 1754 11231 1802
rect 11283 1754 11298 1802
rect 11350 1754 11365 1802
rect 11417 1754 11432 1802
rect 11484 1754 11499 1802
rect 11018 1753 11030 1754
rect 11091 1753 11097 1754
rect 11417 1753 11422 1754
rect 11484 1753 11495 1754
rect 11551 1753 11566 1805
rect 11618 1753 11633 1805
rect 11685 1753 11699 1805
rect 11751 1753 11765 1805
rect 11821 1802 11831 1805
rect 11894 1802 11897 1805
rect 12147 1802 12152 1805
rect 12213 1802 12225 1805
rect 11817 1754 11831 1802
rect 11883 1754 11897 1802
rect 11949 1754 11963 1802
rect 12015 1754 12029 1802
rect 12081 1754 12095 1802
rect 12147 1754 12161 1802
rect 12213 1754 12227 1802
rect 11821 1753 11831 1754
rect 11894 1753 11897 1754
rect 12147 1753 12152 1754
rect 12213 1753 12225 1754
rect 12279 1753 12293 1805
rect 12345 1753 12359 1805
rect 12411 1753 12417 1805
tri 16798 1782 16832 1816 ne
rect 16832 1782 16847 1816
rect 16881 1782 16919 1816
rect 16953 1782 16991 1816
rect 17025 1782 17063 1816
rect 17097 1782 17135 1816
rect 17169 1782 17207 1816
rect 17241 1782 17279 1816
rect 17313 1782 17351 1816
rect 17385 1782 17423 1816
rect 17457 1782 17495 1816
rect 17529 1782 17567 1816
rect 17601 1782 17639 1816
rect 17673 1782 17711 1816
rect 17745 1782 17783 1816
rect 17817 1782 17855 1816
rect 17889 1782 17927 1816
rect 17961 1782 17999 1816
rect 18033 1782 18071 1816
rect 18105 1782 18143 1816
rect 18177 1782 18215 1816
rect 18249 1782 18287 1816
rect 18321 1782 18359 1816
rect 18393 1782 18431 1816
rect 18465 1782 18503 1816
rect 18537 1782 18575 1816
rect 18609 1782 18647 1816
rect 18681 1782 18719 1816
rect 18753 1782 18791 1816
rect 18825 1782 18863 1816
rect 18897 1782 18935 1816
rect 18969 1782 19007 1816
rect 19041 1782 19079 1816
rect 19113 1782 19151 1816
rect 19185 1782 19197 1816
tri 16832 1779 16835 1782 ne
rect 10726 1725 10765 1753
rect 10799 1725 10838 1753
rect 10872 1725 10911 1753
rect 10945 1725 10984 1753
rect 11018 1725 11057 1753
rect 11091 1725 11130 1753
rect 11164 1725 11203 1753
rect 11237 1725 11276 1753
rect 11310 1725 11349 1753
rect 11383 1725 11422 1753
rect 11456 1725 11495 1753
rect 11529 1725 11568 1753
rect 11602 1725 11641 1753
rect 11675 1725 11714 1753
rect 11748 1725 11787 1753
rect 11821 1725 11860 1753
rect 11894 1725 11933 1753
rect 11967 1725 12006 1753
rect 12040 1725 12079 1753
rect 12113 1725 12152 1753
rect 12186 1725 12225 1753
rect 12259 1725 12298 1753
rect 12332 1725 12371 1753
rect 12405 1725 12417 1753
tri 12710 1734 12742 1766 se
rect 12742 1760 16773 1766
rect 12742 1734 16535 1760
tri 12706 1730 12710 1734 se
rect 12710 1730 16535 1734
rect 10726 1720 10762 1725
rect 9722 1673 10762 1720
rect 10814 1673 10829 1725
rect 10881 1673 10896 1725
rect 10948 1673 10963 1725
rect 11018 1720 11030 1725
rect 11091 1720 11097 1725
rect 11417 1720 11422 1725
rect 11484 1720 11495 1725
rect 11015 1673 11030 1720
rect 11082 1673 11097 1720
rect 11149 1673 11164 1720
rect 11216 1673 11231 1720
rect 11283 1673 11298 1720
rect 11350 1673 11365 1720
rect 11417 1673 11432 1720
rect 11484 1673 11499 1720
rect 11551 1673 11566 1725
rect 11618 1673 11633 1725
rect 11685 1673 11699 1725
rect 11751 1673 11765 1725
rect 11821 1720 11831 1725
rect 11894 1720 11897 1725
rect 12147 1720 12152 1725
rect 12213 1720 12225 1725
rect 11817 1673 11831 1720
rect 11883 1673 11897 1720
rect 11949 1673 11963 1720
rect 12015 1673 12029 1720
rect 12081 1673 12095 1720
rect 12147 1673 12161 1720
rect 12213 1673 12227 1720
rect 12279 1673 12293 1725
rect 12345 1673 12359 1725
rect 12411 1673 12417 1725
tri 12672 1696 12706 1730 se
rect 12706 1708 16535 1730
rect 16587 1708 16611 1760
rect 16663 1708 16687 1760
rect 16739 1708 16773 1760
rect 12706 1696 16773 1708
tri 12666 1690 12672 1696 se
rect 12672 1690 16773 1696
rect 9722 1672 12417 1673
rect 9722 1638 9734 1672
rect 9768 1638 9808 1672
rect 9842 1638 9882 1672
rect 9916 1638 9956 1672
rect 9990 1638 10030 1672
rect 10064 1638 10104 1672
rect 10138 1638 10178 1672
rect 10212 1638 10252 1672
rect 10286 1638 10326 1672
rect 10360 1638 10400 1672
rect 10434 1638 10473 1672
rect 10507 1638 10546 1672
rect 10580 1638 10619 1672
rect 10653 1638 10692 1672
rect 10726 1645 10765 1672
rect 10799 1645 10838 1672
rect 10872 1645 10911 1672
rect 10945 1645 10984 1672
rect 11018 1645 11057 1672
rect 11091 1645 11130 1672
rect 11164 1645 11203 1672
rect 11237 1645 11276 1672
rect 11310 1645 11349 1672
rect 11383 1645 11422 1672
rect 11456 1645 11495 1672
rect 11529 1645 11568 1672
rect 11602 1645 11641 1672
rect 11675 1645 11714 1672
rect 11748 1645 11787 1672
rect 11821 1645 11860 1672
rect 11894 1645 11933 1672
rect 11967 1645 12006 1672
rect 12040 1645 12079 1672
rect 12113 1645 12152 1672
rect 12186 1645 12225 1672
rect 12259 1645 12298 1672
rect 12332 1645 12371 1672
rect 12405 1645 12417 1672
tri 12632 1656 12666 1690 se
rect 12666 1681 16773 1690
rect 12666 1656 16535 1681
rect 10726 1638 10762 1645
rect 9722 1593 10762 1638
rect 10814 1593 10829 1645
rect 10881 1593 10896 1645
rect 10948 1593 10963 1645
rect 11018 1638 11030 1645
rect 11091 1638 11097 1645
rect 11417 1638 11422 1645
rect 11484 1638 11495 1645
rect 11015 1593 11030 1638
rect 11082 1593 11097 1638
rect 11149 1593 11164 1638
rect 11216 1593 11231 1638
rect 11283 1593 11298 1638
rect 11350 1593 11365 1638
rect 11417 1593 11432 1638
rect 11484 1593 11499 1638
rect 11551 1593 11566 1645
rect 11618 1593 11633 1645
rect 11685 1593 11699 1645
rect 11751 1593 11765 1645
rect 11821 1638 11831 1645
rect 11894 1638 11897 1645
rect 12147 1638 12152 1645
rect 12213 1638 12225 1645
rect 11817 1593 11831 1638
rect 11883 1593 11897 1638
rect 11949 1593 11963 1638
rect 12015 1593 12029 1638
rect 12081 1593 12095 1638
rect 12147 1593 12161 1638
rect 12213 1593 12227 1638
rect 12279 1593 12293 1645
rect 12345 1593 12359 1645
rect 12411 1593 12417 1645
tri 12620 1644 12632 1656 se
rect 12632 1644 16535 1656
tri 12586 1610 12620 1644 se
rect 12620 1629 16535 1644
rect 16587 1629 16611 1681
rect 16663 1629 16687 1681
rect 16739 1629 16773 1681
rect 12620 1610 16773 1629
rect 9722 1590 12417 1593
rect 9722 1556 9734 1590
rect 9768 1556 9808 1590
rect 9842 1556 9882 1590
rect 9916 1556 9956 1590
rect 9990 1556 10030 1590
rect 10064 1556 10104 1590
rect 10138 1556 10178 1590
rect 10212 1556 10252 1590
rect 10286 1556 10326 1590
rect 10360 1556 10400 1590
rect 10434 1556 10473 1590
rect 10507 1556 10546 1590
rect 10580 1556 10619 1590
rect 10653 1556 10692 1590
rect 10726 1556 10765 1590
rect 10799 1556 10838 1590
rect 10872 1556 10911 1590
rect 10945 1556 10984 1590
rect 11018 1556 11057 1590
rect 11091 1556 11130 1590
rect 11164 1556 11203 1590
rect 11237 1556 11276 1590
rect 11310 1556 11349 1590
rect 11383 1556 11422 1590
rect 11456 1556 11495 1590
rect 11529 1556 11568 1590
rect 11602 1556 11641 1590
rect 11675 1556 11714 1590
rect 11748 1556 11787 1590
rect 11821 1556 11860 1590
rect 11894 1556 11933 1590
rect 11967 1556 12006 1590
rect 12040 1556 12079 1590
rect 12113 1556 12152 1590
rect 12186 1556 12225 1590
rect 12259 1556 12298 1590
rect 12332 1556 12371 1590
rect 12405 1556 12417 1590
tri 12554 1578 12586 1610 se
rect 12586 1602 16773 1610
rect 16835 1755 19197 1782
rect 16835 1730 18875 1755
rect 18927 1730 18941 1755
rect 16835 1696 16847 1730
rect 16881 1696 16919 1730
rect 16953 1696 16991 1730
rect 17025 1696 17063 1730
rect 17097 1696 17135 1730
rect 17169 1696 17207 1730
rect 17241 1696 17279 1730
rect 17313 1696 17351 1730
rect 17385 1696 17423 1730
rect 17457 1696 17495 1730
rect 17529 1696 17567 1730
rect 17601 1696 17639 1730
rect 17673 1696 17711 1730
rect 17745 1696 17783 1730
rect 17817 1696 17855 1730
rect 17889 1696 17927 1730
rect 17961 1696 17999 1730
rect 18033 1696 18071 1730
rect 18105 1696 18143 1730
rect 18177 1696 18215 1730
rect 18249 1696 18287 1730
rect 18321 1696 18359 1730
rect 18393 1696 18431 1730
rect 18465 1696 18503 1730
rect 18537 1696 18575 1730
rect 18609 1696 18647 1730
rect 18681 1696 18719 1730
rect 18753 1696 18791 1730
rect 18825 1696 18863 1730
rect 18927 1703 18935 1730
rect 18993 1703 19007 1755
rect 19059 1703 19073 1755
rect 19125 1703 19139 1755
rect 19191 1703 19197 1755
rect 18897 1696 18935 1703
rect 18969 1696 19007 1703
rect 19041 1696 19079 1703
rect 19113 1696 19151 1703
rect 19185 1696 19197 1703
rect 16835 1655 19197 1696
rect 16835 1644 18875 1655
rect 18927 1644 18941 1655
rect 16835 1610 16847 1644
rect 16881 1610 16919 1644
rect 16953 1610 16991 1644
rect 17025 1610 17063 1644
rect 17097 1610 17135 1644
rect 17169 1610 17207 1644
rect 17241 1610 17279 1644
rect 17313 1610 17351 1644
rect 17385 1610 17423 1644
rect 17457 1610 17495 1644
rect 17529 1610 17567 1644
rect 17601 1610 17639 1644
rect 17673 1610 17711 1644
rect 17745 1610 17783 1644
rect 17817 1610 17855 1644
rect 17889 1610 17927 1644
rect 17961 1610 17999 1644
rect 18033 1610 18071 1644
rect 18105 1610 18143 1644
rect 18177 1610 18215 1644
rect 18249 1610 18287 1644
rect 18321 1610 18359 1644
rect 18393 1610 18431 1644
rect 18465 1610 18503 1644
rect 18537 1610 18575 1644
rect 18609 1610 18647 1644
rect 18681 1610 18719 1644
rect 18753 1610 18791 1644
rect 18825 1610 18863 1644
rect 18927 1610 18935 1644
rect 16835 1603 18875 1610
rect 18927 1603 18941 1610
rect 18993 1603 19007 1655
rect 19059 1603 19073 1655
rect 19125 1603 19139 1655
rect 19191 1603 19197 1655
rect 19967 1878 20042 1924
rect 24437 1888 24695 1927
rect 19967 1846 20013 1878
tri 20013 1849 20042 1878 nw
rect 19967 1812 19973 1846
rect 20007 1812 20013 1846
rect 19967 1768 20013 1812
rect 19967 1734 19973 1768
rect 20007 1734 20013 1768
rect 19967 1690 20013 1734
rect 19967 1656 19973 1690
rect 20007 1656 20013 1690
rect 19967 1612 20013 1656
rect 12586 1578 16535 1602
rect 9722 1547 12417 1556
tri 12523 1547 12554 1578 se
rect 12554 1550 16535 1578
rect 16587 1550 16611 1602
rect 16663 1550 16687 1602
rect 16739 1550 16773 1602
rect 12554 1547 16773 1550
tri 12520 1544 12523 1547 se
rect 12523 1544 16773 1547
rect 19967 1578 19973 1612
rect 20007 1578 20013 1612
tri 12513 1537 12520 1544 se
rect 12520 1537 12883 1544
tri 12883 1537 12890 1544 nw
tri 12510 1534 12513 1537 se
rect 12513 1534 12880 1537
tri 12880 1534 12883 1537 nw
tri 17293 1534 17296 1537 se
rect 17296 1534 17619 1537
rect 9405 1479 9411 1513
rect 9445 1479 9451 1513
tri 12476 1500 12510 1534 se
rect 12510 1514 12860 1534
tri 12860 1514 12880 1534 nw
tri 17273 1514 17293 1534 se
rect 17293 1514 17619 1534
rect 12510 1500 12846 1514
tri 12846 1500 12860 1514 nw
tri 12901 1500 12915 1514 se
rect 12915 1500 14443 1514
tri 12472 1496 12476 1500 se
rect 12476 1496 12842 1500
tri 12842 1496 12846 1500 nw
tri 12897 1496 12901 1500 se
rect 12901 1496 14443 1500
tri 12461 1485 12472 1496 se
rect 12472 1485 12831 1496
tri 12831 1485 12842 1496 nw
tri 12886 1485 12897 1496 se
rect 12897 1485 14443 1496
rect 9405 1434 9451 1479
rect 9405 1400 9411 1434
rect 9445 1400 9451 1434
rect 9405 1378 9451 1400
tri 12437 1461 12461 1485 se
rect 12461 1461 12807 1485
tri 12807 1461 12831 1485 nw
tri 12863 1462 12886 1485 se
rect 12886 1475 14443 1485
rect 12886 1462 12926 1475
tri 12926 1462 12939 1475 nw
tri 14423 1462 14436 1475 ne
rect 14436 1462 14443 1475
rect 14495 1462 14507 1514
rect 14559 1485 17619 1514
rect 17671 1485 17683 1537
rect 17735 1485 17741 1537
rect 19967 1534 20013 1578
rect 19967 1500 19973 1534
rect 20007 1500 20013 1534
rect 14559 1475 17325 1485
tri 17325 1475 17335 1485 nw
rect 14559 1462 14566 1475
tri 14566 1462 14579 1475 nw
tri 12862 1461 12863 1462 se
rect 12863 1461 12925 1462
tri 12925 1461 12926 1462 nw
rect 12437 1456 12802 1461
tri 12802 1456 12807 1461 nw
rect 12862 1456 12920 1461
tri 12920 1456 12925 1461 nw
rect 19967 1456 20013 1500
rect 12437 1422 12768 1456
tri 12768 1422 12802 1456 nw
rect 12437 1399 12745 1422
tri 12745 1399 12768 1422 nw
rect 12437 1397 12743 1399
tri 12743 1397 12745 1399 nw
tri 9451 1378 9470 1397 sw
rect 12437 1378 12724 1397
tri 12724 1378 12743 1397 nw
rect 9405 1361 9470 1378
tri 9470 1361 9487 1378 sw
tri 12252 1361 12258 1367 se
rect 12258 1361 12264 1367
rect 9405 1355 12264 1361
rect 12316 1355 12328 1367
rect 9405 1321 9483 1355
rect 9517 1321 9556 1355
rect 9590 1321 9629 1355
rect 9663 1321 9702 1355
rect 9736 1321 9775 1355
rect 9809 1321 9848 1355
rect 9882 1321 9921 1355
rect 9955 1321 9994 1355
rect 10028 1321 10067 1355
rect 10101 1321 10140 1355
rect 10174 1321 10213 1355
rect 10247 1321 10286 1355
rect 10320 1321 10359 1355
rect 10393 1321 10432 1355
rect 10466 1321 10505 1355
rect 10539 1321 10578 1355
rect 10612 1321 10651 1355
rect 10685 1321 10724 1355
rect 10758 1321 10797 1355
rect 10831 1321 10870 1355
rect 10904 1321 10943 1355
rect 10977 1321 11016 1355
rect 11050 1321 11089 1355
rect 11123 1321 11162 1355
rect 11196 1321 11235 1355
rect 11269 1321 11308 1355
rect 11342 1321 11381 1355
rect 11415 1321 11454 1355
rect 11488 1321 11527 1355
rect 11561 1321 11600 1355
rect 11634 1321 11672 1355
rect 11706 1321 11744 1355
rect 11778 1321 11816 1355
rect 11850 1321 11888 1355
rect 11922 1321 11960 1355
rect 11994 1321 12032 1355
rect 12066 1321 12104 1355
rect 12138 1321 12176 1355
rect 12210 1321 12248 1355
rect 12316 1321 12320 1355
rect 9405 1315 12264 1321
rect 12316 1315 12328 1321
rect 12380 1315 12386 1367
tri 9255 1300 9263 1308 sw
rect 9203 1282 9263 1300
tri 9263 1282 9281 1300 sw
rect 9203 1261 12291 1282
tri 9203 1250 9214 1261 ne
rect 9214 1250 12291 1261
tri 9214 1230 9234 1250 ne
rect 9234 1230 12291 1250
tri 10687 1225 10692 1230 ne
rect 10692 1225 12291 1230
tri 9170 1216 9179 1225 sw
tri 10692 1216 10701 1225 ne
rect 10701 1216 12291 1225
rect 8341 1164 8431 1216
rect 8483 1164 8509 1216
rect 8561 1164 8587 1216
rect 8639 1164 8665 1216
rect 8717 1164 8743 1216
rect 8795 1164 8871 1216
tri 8340 1039 8341 1040 se
rect 8341 1039 8871 1164
rect 9118 1199 9179 1216
tri 9179 1199 9196 1216 sw
tri 10701 1199 10718 1216 ne
rect 10718 1199 12291 1216
rect 9118 1183 9785 1199
tri 10718 1188 10729 1199 ne
rect 10729 1188 12291 1199
tri 9118 1147 9154 1183 ne
rect 9154 1147 9785 1183
tri 9707 1144 9710 1147 ne
rect 9710 1144 9785 1147
tri 10729 1144 10773 1188 ne
rect 10773 1144 12291 1188
tri 9710 1135 9719 1144 ne
rect 9719 1135 9785 1144
tri 10773 1135 10782 1144 ne
rect 10782 1135 12291 1144
tri 9719 1121 9733 1135 ne
rect 8340 1033 8871 1039
rect 9733 1042 9785 1135
tri 10782 1124 10793 1135 ne
tri 9785 1042 9805 1062 sw
rect 9733 1036 9805 1042
tri 9805 1036 9811 1042 sw
rect 8340 999 8352 1033
rect 8386 999 8431 1033
rect 8465 999 8510 1033
rect 8544 999 8589 1033
rect 8623 999 8668 1033
rect 8702 999 8747 1033
rect 8781 999 8825 1033
rect 8859 999 8871 1033
rect 8340 993 8871 999
rect 8955 1030 9677 1036
rect 8955 996 8967 1030
rect 9001 996 9041 1030
rect 9075 996 9115 1030
rect 9149 996 9189 1030
rect 9223 996 9263 1030
rect 9297 996 9337 1030
rect 9371 996 9411 1030
rect 9445 996 9485 1030
rect 9519 996 9558 1030
rect 9592 996 9631 1030
rect 9665 996 9677 1030
rect 8955 990 9677 996
rect 9733 1030 10520 1036
rect 9733 996 9745 1030
rect 9779 996 9819 1030
rect 9853 996 9893 1030
rect 9927 996 9967 1030
rect 10001 996 10041 1030
rect 10075 996 10116 1030
rect 10150 996 10191 1030
rect 10225 996 10266 1030
rect 10300 996 10341 1030
rect 10375 996 10416 1030
rect 10450 996 10520 1030
rect 10793 1030 12291 1135
rect 9733 990 10520 996
tri 9032 977 9045 990 ne
rect 9045 977 9117 990
tri 9117 977 9130 990 nw
tri 9344 977 9357 990 ne
rect 9357 977 9429 990
tri 9429 977 9442 990 nw
tri 9812 977 9825 990 ne
rect 9825 977 9897 990
tri 9897 977 9910 990 nw
tri 10124 977 10137 990 ne
rect 10137 977 10209 990
tri 10209 977 10222 990 nw
tri 10436 977 10449 990 ne
rect 10449 977 10520 990
tri 9045 964 9058 977 ne
rect 8090 248 8142 260
rect 8090 190 8142 196
rect 8171 914 8327 926
rect 8171 880 8177 914
rect 8211 880 8284 914
rect 8318 880 8327 914
rect 8171 842 8327 880
rect 8171 838 8284 842
rect 8171 804 8177 838
rect 8211 808 8284 838
rect 8318 808 8327 842
rect 8434 914 8480 926
rect 8434 880 8440 914
rect 8474 880 8480 914
rect 8434 842 8480 880
rect 8211 804 8327 808
rect 8171 770 8327 804
rect 8171 762 8284 770
rect 8171 728 8177 762
rect 8211 736 8284 762
rect 8318 736 8327 770
rect 8211 728 8327 736
rect 8171 698 8327 728
rect 8171 686 8284 698
rect 8171 652 8177 686
rect 8211 664 8284 686
rect 8318 664 8327 698
tri 8431 814 8434 817 se
rect 8434 814 8440 842
rect 8431 808 8440 814
rect 8474 814 8480 842
rect 8590 914 8636 926
rect 8590 880 8596 914
rect 8630 880 8636 914
rect 8590 842 8636 880
tri 8480 814 8483 817 sw
rect 8474 808 8483 814
rect 8431 744 8440 756
rect 8474 744 8483 756
rect 8431 686 8440 692
tri 8431 683 8434 686 ne
rect 8211 652 8327 664
rect 8171 626 8327 652
rect 8171 610 8284 626
rect 8171 576 8177 610
rect 8211 592 8284 610
rect 8318 592 8327 626
rect 8211 576 8327 592
rect 8171 554 8327 576
rect 8171 533 8284 554
rect 8171 499 8177 533
rect 8211 520 8284 533
rect 8318 520 8327 554
rect 8211 499 8327 520
rect 8171 482 8327 499
rect 8171 456 8284 482
rect 8171 422 8177 456
rect 8211 448 8284 456
rect 8318 448 8327 482
rect 8211 422 8327 448
rect 8171 410 8327 422
rect 8171 379 8284 410
rect 8171 345 8177 379
rect 8211 376 8284 379
rect 8318 376 8327 410
rect 8211 345 8327 376
rect 8171 338 8327 345
rect 8171 304 8284 338
rect 8318 304 8327 338
rect 8171 302 8327 304
rect 8171 268 8177 302
rect 8211 268 8327 302
rect 8171 266 8327 268
rect 8171 232 8284 266
rect 8318 232 8327 266
rect 8171 225 8327 232
rect 8171 191 8177 225
rect 8211 194 8327 225
rect 8211 191 8284 194
rect 7848 131 7854 165
rect 7888 131 7894 165
rect 7848 93 7894 131
rect 7848 59 7854 93
rect 7888 59 7894 93
rect 7848 21 7894 59
rect 7848 -13 7854 21
rect 7888 -13 7894 21
rect 7848 -25 7894 -13
rect 8171 160 8284 191
rect 8318 160 8327 194
rect 8171 154 8327 160
rect 8223 102 8275 154
rect 8171 88 8284 102
rect 8318 88 8327 102
rect 8171 72 8327 88
rect 8223 20 8275 72
rect 8171 16 8284 20
rect 8318 16 8327 20
rect 8171 -6 8327 16
rect 8171 -11 8177 -6
rect 8211 -11 8327 -6
rect 8223 -63 8275 -11
rect 8171 -69 8327 -63
rect 8434 664 8440 686
rect 8474 686 8483 692
rect 8474 664 8480 686
tri 8480 683 8483 686 nw
rect 8590 808 8596 842
rect 8630 808 8636 842
rect 8746 914 8792 926
rect 8746 880 8752 914
rect 8786 880 8792 914
rect 8746 842 8792 880
rect 8590 770 8636 808
rect 8590 736 8596 770
rect 8630 736 8636 770
rect 8590 698 8636 736
rect 8434 626 8480 664
rect 8434 592 8440 626
rect 8474 592 8480 626
rect 8434 554 8480 592
rect 8434 520 8440 554
rect 8474 520 8480 554
rect 8434 482 8480 520
rect 8434 448 8440 482
rect 8474 448 8480 482
rect 8434 410 8480 448
rect 8434 376 8440 410
rect 8474 376 8480 410
rect 8434 338 8480 376
rect 8434 304 8440 338
rect 8474 304 8480 338
rect 8434 266 8480 304
rect 8434 232 8440 266
rect 8474 232 8480 266
rect 8434 194 8480 232
rect 8434 160 8440 194
rect 8474 160 8480 194
rect 8590 664 8596 698
rect 8630 664 8636 698
tri 8743 814 8746 817 se
rect 8746 814 8752 842
rect 8743 808 8752 814
rect 8786 814 8792 842
rect 8902 914 8948 926
rect 8902 880 8908 914
rect 8942 880 8948 914
rect 8902 842 8948 880
tri 8792 814 8795 817 sw
rect 8786 808 8795 814
rect 8743 744 8752 756
rect 8786 744 8795 756
rect 8743 686 8752 692
tri 8743 683 8746 686 ne
rect 8590 626 8636 664
rect 8590 592 8596 626
rect 8630 592 8636 626
rect 8590 554 8636 592
rect 8590 520 8596 554
rect 8630 520 8636 554
rect 8590 482 8636 520
rect 8590 448 8596 482
rect 8630 448 8636 482
rect 8590 410 8636 448
rect 8590 376 8596 410
rect 8630 376 8636 410
rect 8590 338 8636 376
rect 8590 304 8596 338
rect 8630 304 8636 338
rect 8590 266 8636 304
rect 8590 232 8596 266
rect 8630 232 8636 266
rect 8590 194 8636 232
rect 8434 122 8480 160
rect 8434 88 8440 122
rect 8474 88 8480 122
rect 8434 50 8480 88
rect 8434 16 8440 50
rect 8474 16 8480 50
rect 8434 -22 8480 16
rect 8434 -56 8440 -22
rect 8474 -56 8480 -22
rect 8434 -68 8480 -56
tri 8587 160 8590 163 se
rect 8590 160 8596 194
rect 8630 160 8636 194
rect 8746 664 8752 686
rect 8786 686 8795 692
rect 8786 664 8792 686
tri 8792 683 8795 686 nw
rect 8902 808 8908 842
rect 8942 808 8948 842
rect 8902 770 8948 808
rect 8902 736 8908 770
rect 8942 736 8948 770
rect 8902 698 8948 736
rect 8746 626 8792 664
rect 8746 592 8752 626
rect 8786 592 8792 626
rect 8746 554 8792 592
rect 8746 520 8752 554
rect 8786 520 8792 554
rect 8746 482 8792 520
rect 8746 448 8752 482
rect 8786 448 8792 482
rect 8746 410 8792 448
rect 8746 376 8752 410
rect 8786 376 8792 410
rect 8746 338 8792 376
rect 8746 304 8752 338
rect 8786 304 8792 338
rect 8746 266 8792 304
rect 8746 232 8752 266
rect 8786 232 8792 266
rect 8746 194 8792 232
tri 8636 160 8639 163 sw
rect 8587 154 8639 160
rect 8587 88 8596 102
rect 8630 88 8639 102
rect 8587 72 8639 88
rect 8587 16 8596 20
rect 8630 16 8639 20
rect 8587 -11 8639 16
rect 8587 -69 8639 -63
rect 8746 160 8752 194
rect 8786 160 8792 194
rect 8902 664 8908 698
rect 8942 664 8948 698
rect 8902 626 8948 664
rect 9058 914 9104 977
tri 9104 964 9117 977 nw
tri 9357 964 9370 977 ne
rect 9058 880 9064 914
rect 9098 880 9104 914
rect 9058 842 9104 880
rect 9058 808 9064 842
rect 9098 808 9104 842
rect 9058 770 9104 808
rect 9058 736 9064 770
rect 9098 736 9104 770
rect 9058 698 9104 736
rect 9058 664 9064 698
rect 9098 664 9104 698
tri 9057 626 9058 627 se
rect 9058 626 9104 664
rect 9214 914 9260 926
rect 9214 880 9220 914
rect 9254 880 9260 914
rect 9214 842 9260 880
rect 9214 808 9220 842
rect 9254 808 9260 842
rect 9214 770 9260 808
rect 9214 736 9220 770
rect 9254 736 9260 770
rect 9214 698 9260 736
rect 9214 664 9220 698
rect 9254 664 9260 698
tri 9104 626 9105 627 sw
rect 9214 626 9260 664
rect 9370 914 9416 977
tri 9416 964 9429 977 nw
tri 9825 964 9838 977 ne
rect 9370 880 9376 914
rect 9410 880 9416 914
rect 9370 842 9416 880
rect 9370 808 9376 842
rect 9410 808 9416 842
rect 9370 770 9416 808
rect 9370 736 9376 770
rect 9410 736 9416 770
rect 9370 698 9416 736
rect 9370 664 9376 698
rect 9410 664 9416 698
tri 9369 626 9370 627 se
rect 9370 626 9416 664
rect 9526 914 9572 926
rect 9526 880 9532 914
rect 9566 880 9572 914
rect 9526 842 9572 880
rect 9526 808 9532 842
rect 9566 808 9572 842
rect 9526 770 9572 808
rect 9526 736 9532 770
rect 9566 736 9572 770
rect 9526 698 9572 736
rect 9526 664 9532 698
rect 9566 664 9572 698
tri 9416 626 9417 627 sw
rect 9526 626 9572 664
rect 9682 914 9728 926
rect 9682 880 9688 914
rect 9722 880 9728 914
rect 9682 842 9728 880
rect 9682 808 9688 842
rect 9722 808 9728 842
rect 9682 770 9728 808
rect 9682 736 9688 770
rect 9722 736 9728 770
rect 9682 698 9728 736
rect 9682 664 9688 698
rect 9722 664 9728 698
tri 9681 626 9682 627 se
rect 9682 626 9728 664
rect 9838 914 9884 977
tri 9884 964 9897 977 nw
tri 10137 964 10150 977 ne
rect 9838 880 9844 914
rect 9878 880 9884 914
rect 9838 842 9884 880
rect 9838 808 9844 842
rect 9878 808 9884 842
rect 9838 770 9884 808
rect 9838 736 9844 770
rect 9878 736 9884 770
rect 9838 698 9884 736
rect 9838 664 9844 698
rect 9878 664 9884 698
tri 9728 626 9729 627 sw
rect 9838 626 9884 664
rect 9994 914 10040 926
rect 9994 880 10000 914
rect 10034 880 10040 914
rect 9994 842 10040 880
rect 9994 808 10000 842
rect 10034 808 10040 842
rect 9994 770 10040 808
rect 9994 736 10000 770
rect 10034 736 10040 770
rect 9994 698 10040 736
rect 9994 664 10000 698
rect 10034 664 10040 698
tri 9993 626 9994 627 se
rect 9994 626 10040 664
rect 10150 914 10196 977
tri 10196 964 10209 977 nw
tri 10449 964 10462 977 ne
rect 10150 880 10156 914
rect 10190 880 10196 914
rect 10150 842 10196 880
rect 10150 808 10156 842
rect 10190 808 10196 842
rect 10150 770 10196 808
rect 10150 736 10156 770
rect 10190 736 10196 770
rect 10150 698 10196 736
rect 10150 664 10156 698
rect 10190 664 10196 698
tri 10040 626 10041 627 sw
rect 10150 626 10196 664
rect 10306 914 10352 926
rect 10306 880 10312 914
rect 10346 880 10352 914
rect 10306 842 10352 880
rect 10306 808 10312 842
rect 10346 808 10352 842
rect 10306 770 10352 808
rect 10306 736 10312 770
rect 10346 736 10352 770
rect 10306 698 10352 736
rect 10306 664 10312 698
rect 10346 664 10352 698
tri 10305 626 10306 627 se
rect 10306 626 10352 664
rect 10462 914 10520 977
rect 10462 880 10468 914
rect 10502 880 10520 914
rect 10462 842 10520 880
rect 10462 808 10468 842
rect 10502 808 10520 842
rect 10462 770 10520 808
rect 10462 736 10468 770
rect 10502 736 10520 770
rect 10462 698 10520 736
rect 10462 664 10468 698
rect 10502 664 10520 698
tri 10352 626 10353 627 sw
rect 10462 626 10520 664
rect 8902 592 8908 626
rect 8942 592 8948 626
rect 8902 554 8948 592
rect 8902 520 8908 554
rect 8942 520 8948 554
rect 8902 482 8948 520
tri 9055 624 9057 626 se
rect 9057 624 9064 626
rect 9055 618 9064 624
rect 9098 624 9105 626
tri 9105 624 9107 626 sw
rect 9098 618 9107 624
rect 9055 554 9107 566
rect 9055 496 9107 502
tri 9055 493 9058 496 ne
rect 8902 448 8908 482
rect 8942 448 8948 482
rect 8902 410 8948 448
rect 8902 376 8908 410
rect 8942 376 8948 410
rect 8902 338 8948 376
rect 8902 304 8908 338
rect 8942 304 8948 338
rect 8902 266 8948 304
rect 8902 232 8908 266
rect 8942 232 8948 266
rect 8902 194 8948 232
rect 8746 122 8792 160
rect 8746 88 8752 122
rect 8786 88 8792 122
rect 8746 50 8792 88
rect 8746 16 8752 50
rect 8786 16 8792 50
rect 8746 -22 8792 16
rect 8746 -56 8752 -22
rect 8786 -56 8792 -22
rect 8746 -68 8792 -56
tri 8899 160 8902 163 se
rect 8902 160 8908 194
rect 8942 160 8948 194
rect 9058 482 9104 496
tri 9104 493 9107 496 nw
rect 9214 592 9220 626
rect 9254 592 9260 626
rect 9214 554 9260 592
rect 9214 520 9220 554
rect 9254 520 9260 554
rect 9058 448 9064 482
rect 9098 448 9104 482
rect 9058 410 9104 448
rect 9058 376 9064 410
rect 9098 376 9104 410
rect 9058 338 9104 376
rect 9058 304 9064 338
rect 9098 304 9104 338
rect 9058 266 9104 304
rect 9058 232 9064 266
rect 9098 232 9104 266
rect 9058 194 9104 232
tri 8948 160 8951 163 sw
rect 8899 154 8951 160
rect 8899 88 8908 102
rect 8942 88 8951 102
rect 8899 72 8951 88
rect 8899 16 8908 20
rect 8942 16 8951 20
rect 8899 -11 8951 16
rect 8899 -69 8951 -63
rect 9058 160 9064 194
rect 9098 160 9104 194
rect 9214 482 9260 520
tri 9367 624 9369 626 se
rect 9369 624 9376 626
rect 9367 618 9376 624
rect 9410 624 9417 626
tri 9417 624 9419 626 sw
rect 9410 618 9419 624
rect 9367 554 9419 566
rect 9367 496 9419 502
tri 9367 493 9370 496 ne
rect 9214 448 9220 482
rect 9254 448 9260 482
rect 9214 410 9260 448
rect 9214 376 9220 410
rect 9254 376 9260 410
rect 9214 338 9260 376
rect 9214 304 9220 338
rect 9254 304 9260 338
rect 9214 266 9260 304
rect 9214 232 9220 266
rect 9254 232 9260 266
rect 9214 194 9260 232
rect 9058 122 9104 160
rect 9058 88 9064 122
rect 9098 88 9104 122
rect 9058 50 9104 88
rect 9058 16 9064 50
rect 9098 16 9104 50
rect 9058 -22 9104 16
rect 9058 -56 9064 -22
rect 9098 -56 9104 -22
rect 9058 -68 9104 -56
tri 9211 160 9214 163 se
rect 9214 160 9220 194
rect 9254 160 9260 194
rect 9370 482 9416 496
tri 9416 493 9419 496 nw
rect 9526 592 9532 626
rect 9566 592 9572 626
rect 9526 554 9572 592
rect 9526 520 9532 554
rect 9566 520 9572 554
rect 9370 448 9376 482
rect 9410 448 9416 482
rect 9370 410 9416 448
rect 9370 376 9376 410
rect 9410 376 9416 410
rect 9370 338 9416 376
rect 9370 304 9376 338
rect 9410 304 9416 338
rect 9370 266 9416 304
rect 9370 232 9376 266
rect 9410 232 9416 266
rect 9370 194 9416 232
tri 9260 160 9263 163 sw
rect 9211 154 9263 160
rect 9211 88 9220 102
rect 9254 88 9263 102
rect 9211 72 9263 88
rect 9211 16 9220 20
rect 9254 16 9263 20
rect 9211 -11 9263 16
rect 9211 -69 9263 -63
rect 9370 160 9376 194
rect 9410 160 9416 194
rect 9526 482 9572 520
tri 9679 624 9681 626 se
rect 9681 624 9688 626
rect 9679 618 9688 624
rect 9722 624 9729 626
tri 9729 624 9731 626 sw
rect 9722 618 9731 624
rect 9679 554 9731 566
rect 9679 496 9731 502
tri 9679 493 9682 496 ne
rect 9526 448 9532 482
rect 9566 448 9572 482
rect 9526 410 9572 448
rect 9526 376 9532 410
rect 9566 376 9572 410
rect 9526 338 9572 376
rect 9526 304 9532 338
rect 9566 304 9572 338
rect 9526 266 9572 304
rect 9526 232 9532 266
rect 9566 232 9572 266
rect 9526 194 9572 232
rect 9370 122 9416 160
rect 9370 88 9376 122
rect 9410 88 9416 122
rect 9370 50 9416 88
rect 9370 16 9376 50
rect 9410 16 9416 50
rect 9370 -22 9416 16
rect 9370 -56 9376 -22
rect 9410 -56 9416 -22
rect 9370 -68 9416 -56
tri 9523 160 9526 163 se
rect 9526 160 9532 194
rect 9566 160 9572 194
rect 9682 482 9728 496
tri 9728 493 9731 496 nw
rect 9838 592 9844 626
rect 9878 592 9884 626
rect 9838 554 9884 592
rect 9838 520 9844 554
rect 9878 520 9884 554
rect 9682 448 9688 482
rect 9722 448 9728 482
rect 9682 410 9728 448
rect 9838 482 9884 520
tri 9991 624 9993 626 se
rect 9993 624 10000 626
rect 9991 618 10000 624
rect 10034 624 10041 626
tri 10041 624 10043 626 sw
rect 10034 618 10043 624
rect 9991 554 10043 566
rect 9991 496 10043 502
tri 9991 493 9994 496 ne
rect 9838 448 9844 482
rect 9878 448 9884 482
tri 9835 428 9838 431 se
rect 9838 428 9884 448
rect 9994 482 10040 496
tri 10040 493 10043 496 nw
rect 10150 592 10156 626
rect 10190 592 10196 626
rect 10150 554 10196 592
rect 10150 520 10156 554
rect 10190 520 10196 554
rect 9994 448 10000 482
rect 10034 448 10040 482
rect 9682 376 9688 410
rect 9722 376 9728 410
rect 9682 338 9728 376
rect 9682 304 9688 338
rect 9722 304 9728 338
rect 9682 266 9728 304
tri 9834 427 9835 428 se
rect 9835 427 9884 428
rect 9834 426 9884 427
tri 9884 426 9886 428 sw
rect 9834 420 9886 426
rect 9834 350 9886 368
rect 9834 292 9886 298
tri 9834 288 9838 292 ne
rect 9682 232 9688 266
rect 9722 232 9728 266
rect 9682 194 9728 232
tri 9572 160 9575 163 sw
rect 9523 154 9575 160
rect 9523 88 9532 102
rect 9566 88 9575 102
rect 9523 72 9575 88
rect 9523 16 9532 20
rect 9566 16 9575 20
rect 9523 -11 9575 16
rect 9523 -69 9575 -63
rect 9682 160 9688 194
rect 9722 160 9728 194
rect 9682 122 9728 160
rect 9682 88 9688 122
rect 9722 88 9728 122
rect 9682 50 9728 88
rect 9682 16 9688 50
rect 9722 16 9728 50
rect 9682 -22 9728 16
rect 9682 -56 9688 -22
rect 9722 -56 9728 -22
rect 9682 -68 9728 -56
rect 9838 266 9884 292
tri 9884 290 9886 292 nw
rect 9994 410 10040 448
rect 10150 482 10196 520
tri 10303 624 10305 626 se
rect 10305 624 10312 626
rect 10303 618 10312 624
rect 10346 624 10353 626
tri 10353 624 10355 626 sw
rect 10346 618 10355 624
rect 10303 554 10355 566
rect 10303 496 10355 502
tri 10303 493 10306 496 ne
rect 10150 448 10156 482
rect 10190 448 10196 482
tri 10147 428 10150 431 se
rect 10150 428 10196 448
rect 10306 482 10352 496
tri 10352 493 10355 496 nw
rect 10462 592 10468 626
rect 10502 592 10520 626
rect 10462 554 10520 592
rect 10462 520 10468 554
rect 10502 520 10520 554
rect 10306 448 10312 482
rect 10346 448 10352 482
rect 9994 376 10000 410
rect 10034 376 10040 410
rect 9994 338 10040 376
rect 9994 304 10000 338
rect 10034 304 10040 338
rect 9838 232 9844 266
rect 9878 232 9884 266
rect 9838 194 9884 232
rect 9838 160 9844 194
rect 9878 160 9884 194
rect 9838 122 9884 160
rect 9838 88 9844 122
rect 9878 88 9884 122
rect 9838 50 9884 88
rect 9838 16 9844 50
rect 9878 16 9884 50
rect 9838 -22 9884 16
rect 9838 -56 9844 -22
rect 9878 -56 9884 -22
rect 9838 -68 9884 -56
rect 9994 266 10040 304
tri 10146 427 10147 428 se
rect 10147 427 10196 428
rect 10146 426 10196 427
tri 10196 426 10198 428 sw
rect 10146 420 10198 426
rect 10146 350 10198 368
rect 10146 292 10198 298
tri 10146 290 10148 292 ne
rect 10148 290 10196 292
tri 10196 290 10198 292 nw
rect 10306 410 10352 448
rect 10462 482 10520 520
rect 10462 448 10468 482
rect 10502 448 10520 482
tri 10460 428 10462 430 se
rect 10462 428 10520 448
rect 10306 376 10312 410
rect 10346 376 10352 410
rect 10306 338 10352 376
rect 10306 304 10312 338
rect 10346 304 10352 338
tri 10148 288 10150 290 ne
rect 9994 232 10000 266
rect 10034 232 10040 266
rect 9994 194 10040 232
rect 9994 160 10000 194
rect 10034 160 10040 194
rect 9994 122 10040 160
rect 9994 88 10000 122
rect 10034 88 10040 122
rect 9994 50 10040 88
rect 9994 16 10000 50
rect 10034 16 10040 50
rect 9994 -22 10040 16
rect 9994 -56 10000 -22
rect 10034 -56 10040 -22
rect 9994 -68 10040 -56
rect 10150 266 10196 290
rect 10150 232 10156 266
rect 10190 232 10196 266
rect 10150 194 10196 232
rect 10150 160 10156 194
rect 10190 160 10196 194
rect 10150 122 10196 160
rect 10150 88 10156 122
rect 10190 88 10196 122
rect 10150 50 10196 88
rect 10150 16 10156 50
rect 10190 16 10196 50
rect 10150 -22 10196 16
rect 10150 -56 10156 -22
rect 10190 -56 10196 -22
rect 10150 -68 10196 -56
rect 10306 266 10352 304
tri 10458 426 10460 428 se
rect 10460 426 10520 428
rect 10458 420 10520 426
rect 10510 368 10520 420
rect 10458 350 10520 368
rect 10510 298 10520 350
rect 10458 292 10520 298
tri 10458 290 10460 292 ne
rect 10460 290 10520 292
tri 10460 288 10462 290 ne
rect 10306 232 10312 266
rect 10346 232 10352 266
rect 10306 194 10352 232
rect 10306 160 10312 194
rect 10346 160 10352 194
rect 10306 122 10352 160
rect 10306 88 10312 122
rect 10346 88 10352 122
rect 10306 50 10352 88
rect 10306 16 10312 50
rect 10346 16 10352 50
rect 10306 -22 10352 16
rect 10306 -56 10312 -22
rect 10346 -56 10352 -22
rect 10306 -68 10352 -56
rect 10462 266 10520 290
rect 10462 232 10468 266
rect 10502 232 10520 266
rect 10462 194 10520 232
rect 10462 160 10468 194
rect 10502 160 10520 194
rect 10598 1011 10644 1023
rect 10598 977 10604 1011
rect 10638 977 10644 1011
rect 10793 996 10805 1030
rect 10839 996 10877 1030
rect 10911 996 10949 1030
rect 10983 996 11021 1030
rect 11055 996 11093 1030
rect 11127 996 11165 1030
rect 11199 996 11237 1030
rect 11271 996 11309 1030
rect 11343 996 11381 1030
rect 11415 996 11453 1030
rect 11487 996 11525 1030
rect 11559 996 11597 1030
rect 11631 996 11669 1030
rect 11703 996 11741 1030
rect 11775 996 11813 1030
rect 11847 996 11885 1030
rect 11919 996 11957 1030
rect 11991 996 12029 1030
rect 12063 996 12101 1030
rect 12135 996 12173 1030
rect 12207 996 12245 1030
rect 12279 996 12291 1030
rect 10793 990 12291 996
rect 10598 936 10644 977
rect 10598 902 10604 936
rect 10638 902 10644 936
rect 12437 979 12718 1378
tri 12718 1372 12724 1378 nw
rect 12862 1114 12908 1456
tri 12908 1444 12920 1456 nw
tri 13001 1432 13012 1443 se
rect 13012 1432 14361 1443
tri 14361 1432 14372 1443 sw
tri 14618 1432 14629 1443 se
rect 14629 1432 15831 1443
tri 12991 1422 13001 1432 se
rect 13001 1422 15831 1432
tri 12968 1399 12991 1422 se
rect 12991 1399 15831 1422
tri 12966 1397 12968 1399 se
rect 12968 1398 15831 1399
rect 12968 1397 13464 1398
tri 12955 1386 12966 1397 se
rect 12966 1391 13464 1397
tri 13464 1391 13471 1398 nw
tri 13654 1391 13661 1398 ne
rect 13661 1391 15831 1398
rect 15883 1391 15895 1443
rect 15947 1391 17381 1443
rect 17433 1391 17445 1443
rect 17497 1391 17503 1443
rect 19967 1422 19973 1456
rect 20007 1422 20013 1456
rect 12966 1386 13012 1391
tri 13012 1386 13017 1391 nw
rect 12862 1080 12868 1114
rect 12902 1080 12908 1114
rect 12862 1042 12908 1080
rect 12862 1008 12868 1042
rect 12902 1008 12908 1042
rect 12862 996 12908 1008
tri 12953 1384 12955 1386 se
rect 12955 1384 13010 1386
tri 13010 1384 13012 1386 nw
rect 12953 1378 13004 1384
tri 13004 1378 13010 1384 nw
rect 19967 1378 20013 1422
tri 12718 979 12719 980 sw
rect 12437 945 12719 979
tri 12719 945 12753 979 sw
rect 12437 940 12753 945
tri 12753 940 12758 945 sw
rect 12437 939 12758 940
rect 12437 927 12823 939
rect 10598 861 10644 902
rect 10598 827 10604 861
rect 10638 827 10644 861
rect 10598 786 10644 827
rect 10598 752 10604 786
rect 10638 752 10644 786
rect 10598 710 10644 752
rect 10598 676 10604 710
rect 10638 676 10644 710
rect 10598 634 10644 676
rect 10598 600 10604 634
rect 10638 600 10644 634
rect 10598 558 10644 600
rect 10598 524 10604 558
rect 10638 524 10644 558
rect 10598 482 10644 524
rect 10598 448 10604 482
rect 10638 448 10644 482
rect 10598 406 10644 448
rect 10598 372 10604 406
rect 10638 372 10644 406
rect 10598 330 10644 372
rect 10598 296 10604 330
rect 10638 296 10644 330
rect 10598 254 10644 296
rect 10598 220 10604 254
rect 10638 220 10644 254
rect 10598 178 10644 220
rect 10462 122 10520 160
rect 10462 88 10468 122
rect 10502 88 10520 122
rect 10462 50 10520 88
rect 10462 16 10468 50
rect 10502 16 10520 50
rect 10462 -22 10520 16
rect 10462 -56 10468 -22
rect 10502 -56 10520 -22
rect 10462 -68 10520 -56
tri 10595 160 10598 163 se
rect 10598 160 10604 178
rect 10595 151 10604 160
rect 10638 160 10644 178
rect 10731 914 10777 926
rect 10731 880 10737 914
rect 10771 880 10777 914
rect 10731 842 10777 880
rect 10731 808 10737 842
rect 10771 808 10777 842
rect 10731 770 10777 808
rect 10731 736 10737 770
rect 10771 736 10777 770
rect 10731 698 10777 736
rect 10731 664 10737 698
rect 10771 664 10777 698
rect 10731 626 10777 664
rect 10731 592 10737 626
rect 10771 592 10777 626
rect 10731 554 10777 592
rect 10731 520 10737 554
rect 10771 520 10777 554
rect 10731 482 10777 520
rect 10731 448 10737 482
rect 10771 448 10777 482
rect 10731 410 10777 448
rect 10731 376 10737 410
rect 10771 376 10777 410
rect 10731 338 10777 376
rect 10731 304 10737 338
rect 10771 304 10777 338
rect 10731 266 10777 304
rect 10731 232 10737 266
rect 10771 232 10777 266
rect 10731 194 10777 232
tri 10644 160 10647 163 sw
rect 10638 151 10647 160
rect 10595 68 10604 99
rect 10638 68 10647 99
rect 10595 57 10647 68
rect 10595 -8 10604 5
rect 10638 -8 10647 5
rect 10595 -38 10647 -8
rect 10595 -96 10647 -90
tri 10728 160 10731 163 se
rect 10731 160 10737 194
rect 10771 160 10777 194
rect 11187 914 11233 926
rect 11187 880 11193 914
rect 11227 880 11233 914
rect 11187 842 11233 880
rect 11187 808 11193 842
rect 11227 808 11233 842
rect 11187 770 11233 808
rect 11187 736 11193 770
rect 11227 736 11233 770
rect 11187 698 11233 736
rect 11187 664 11193 698
rect 11227 664 11233 698
rect 11187 626 11233 664
rect 11187 592 11193 626
rect 11227 592 11233 626
rect 11187 554 11233 592
rect 11187 520 11193 554
rect 11227 520 11233 554
rect 11187 482 11233 520
rect 11187 448 11193 482
rect 11227 448 11233 482
rect 11187 410 11233 448
rect 11187 376 11193 410
rect 11227 376 11233 410
rect 11187 338 11233 376
rect 11187 304 11193 338
rect 11227 304 11233 338
rect 11187 266 11233 304
rect 11187 232 11193 266
rect 11227 232 11233 266
rect 11187 194 11233 232
tri 10777 160 10780 163 sw
rect 10728 151 10780 160
rect 10728 88 10737 99
rect 10771 88 10780 99
rect 10728 57 10780 88
rect 10728 -22 10780 5
rect 10728 -38 10737 -22
rect 10771 -38 10780 -22
rect 10728 -96 10780 -90
tri 11184 160 11187 163 se
rect 11187 160 11193 194
rect 11227 160 11233 194
rect 11643 914 11689 926
rect 11643 880 11649 914
rect 11683 880 11689 914
rect 11643 842 11689 880
rect 11643 808 11649 842
rect 11683 808 11689 842
rect 11643 770 11689 808
rect 11643 736 11649 770
rect 11683 736 11689 770
rect 11643 698 11689 736
rect 11643 664 11649 698
rect 11683 664 11689 698
rect 11643 626 11689 664
rect 11643 592 11649 626
rect 11683 592 11689 626
rect 11643 554 11689 592
rect 11643 520 11649 554
rect 11683 520 11689 554
rect 11643 482 11689 520
rect 11643 448 11649 482
rect 11683 448 11689 482
rect 11643 410 11689 448
rect 11643 376 11649 410
rect 11683 376 11689 410
rect 11643 338 11689 376
rect 11643 304 11649 338
rect 11683 304 11689 338
rect 11643 266 11689 304
rect 11643 232 11649 266
rect 11683 232 11689 266
rect 11643 194 11689 232
tri 11233 160 11236 163 sw
rect 11184 151 11236 160
rect 11184 88 11193 99
rect 11227 88 11236 99
rect 11184 57 11236 88
rect 11184 -22 11236 5
rect 11184 -38 11193 -22
rect 11227 -38 11236 -22
rect 11184 -96 11236 -90
tri 11640 160 11643 163 se
rect 11643 160 11649 194
rect 11683 160 11689 194
rect 12099 914 12145 926
rect 12099 880 12105 914
rect 12139 880 12145 914
rect 12099 842 12145 880
rect 12099 808 12105 842
rect 12139 808 12145 842
rect 12099 770 12145 808
rect 12099 736 12105 770
rect 12139 736 12145 770
rect 12099 698 12145 736
rect 12099 664 12105 698
rect 12139 664 12145 698
rect 12099 626 12145 664
rect 12099 592 12105 626
rect 12139 592 12145 626
rect 12099 554 12145 592
rect 12099 520 12105 554
rect 12139 520 12145 554
rect 12099 482 12145 520
rect 12099 448 12105 482
rect 12139 448 12145 482
rect 12099 410 12145 448
rect 12099 376 12105 410
rect 12139 376 12145 410
rect 12099 338 12145 376
rect 12099 304 12105 338
rect 12139 304 12145 338
rect 12099 266 12145 304
rect 12099 232 12105 266
rect 12139 232 12145 266
rect 12099 194 12145 232
tri 11689 160 11692 163 sw
rect 11640 151 11692 160
rect 11640 88 11649 99
rect 11683 88 11692 99
rect 11640 57 11692 88
rect 11640 -22 11692 5
rect 11640 -38 11649 -22
rect 11683 -38 11692 -22
rect 11640 -96 11692 -90
tri 12097 160 12099 162 se
rect 12099 160 12105 194
rect 12139 160 12145 194
rect 12437 914 12783 927
rect 12437 880 12561 914
rect 12595 893 12783 914
rect 12817 893 12823 927
rect 12595 880 12823 893
rect 12437 842 12823 880
rect 12437 808 12561 842
rect 12595 808 12823 842
rect 12437 805 12823 808
rect 12437 771 12783 805
rect 12817 771 12823 805
rect 12437 770 12823 771
rect 12437 736 12561 770
rect 12595 759 12823 770
rect 12953 927 12999 1378
tri 12999 1373 13004 1378 nw
rect 13494 1315 13501 1367
rect 13553 1355 13565 1367
rect 13617 1361 13623 1367
tri 13623 1361 13629 1367 sw
rect 13617 1355 18903 1361
rect 13560 1321 13565 1355
rect 13633 1321 13672 1355
rect 13706 1321 13745 1355
rect 13779 1321 13818 1355
rect 13852 1321 13891 1355
rect 13925 1321 13964 1355
rect 13998 1321 14037 1355
rect 14071 1321 14110 1355
rect 14144 1321 14183 1355
rect 14217 1321 14255 1355
rect 14289 1321 14327 1355
rect 14361 1321 14399 1355
rect 14433 1321 14471 1355
rect 14505 1321 14543 1355
rect 14577 1321 14615 1355
rect 14649 1321 14687 1355
rect 14721 1321 14759 1355
rect 14793 1321 14831 1355
rect 14865 1321 14903 1355
rect 14937 1321 14975 1355
rect 15009 1321 15047 1355
rect 15081 1321 15119 1355
rect 15153 1321 15191 1355
rect 15225 1321 15263 1355
rect 15297 1321 15335 1355
rect 15369 1321 15407 1355
rect 15441 1321 15479 1355
rect 15513 1321 15551 1355
rect 15585 1321 15623 1355
rect 15657 1321 15695 1355
rect 15729 1321 15767 1355
rect 15801 1321 15839 1355
rect 15873 1321 15911 1355
rect 15945 1321 15983 1355
rect 16017 1321 16055 1355
rect 16089 1321 16127 1355
rect 16161 1321 16199 1355
rect 16233 1321 16271 1355
rect 16305 1321 16343 1355
rect 16377 1321 16415 1355
rect 16449 1321 16487 1355
rect 16521 1321 16559 1355
rect 16593 1321 16631 1355
rect 16665 1321 16703 1355
rect 16737 1321 16775 1355
rect 16809 1321 16847 1355
rect 16881 1321 16919 1355
rect 16953 1321 16991 1355
rect 17025 1321 17063 1355
rect 17097 1321 17135 1355
rect 17169 1321 17207 1355
rect 17241 1321 17279 1355
rect 17313 1321 17351 1355
rect 17385 1321 17423 1355
rect 17457 1321 17495 1355
rect 17529 1321 17567 1355
rect 17601 1321 17639 1355
rect 17673 1321 17711 1355
rect 17745 1321 17783 1355
rect 17817 1321 17855 1355
rect 17889 1321 17927 1355
rect 17961 1321 17999 1355
rect 18033 1321 18071 1355
rect 18105 1321 18143 1355
rect 18177 1321 18215 1355
rect 18249 1321 18287 1355
rect 18321 1321 18359 1355
rect 18393 1321 18431 1355
rect 18465 1321 18503 1355
rect 18537 1321 18575 1355
rect 18609 1321 18647 1355
rect 18681 1321 18719 1355
rect 18753 1321 18791 1355
rect 18825 1321 18903 1355
rect 13553 1315 13565 1321
rect 13617 1315 18903 1321
tri 18828 1300 18843 1315 ne
rect 18843 1300 18903 1315
tri 18843 1286 18857 1300 ne
tri 16974 1266 16983 1275 se
rect 16983 1266 17939 1275
tri 16958 1250 16974 1266 se
rect 16974 1250 17939 1266
tri 16949 1241 16958 1250 se
rect 16958 1241 17939 1250
rect 16949 1223 17939 1241
rect 17991 1223 18003 1275
rect 18055 1223 18061 1275
rect 18857 1250 18903 1300
rect 16949 1216 17018 1223
tri 17018 1216 17025 1223 nw
rect 18857 1216 18863 1250
rect 18897 1216 18903 1250
rect 15116 1135 15867 1141
rect 15116 1101 15219 1135
rect 15253 1101 15411 1135
rect 15445 1101 15506 1135
rect 15540 1101 15644 1135
rect 15678 1101 15736 1135
rect 15770 1101 15867 1135
rect 15116 1095 15867 1101
tri 13511 1075 13515 1079 se
rect 13515 1075 13805 1079
rect 13060 1069 13805 1075
rect 13857 1069 13873 1079
rect 13925 1069 13941 1079
rect 13060 1035 13072 1069
rect 13106 1035 13144 1069
rect 13178 1035 13216 1069
rect 13250 1035 13288 1069
rect 13322 1035 13360 1069
rect 13394 1035 13432 1069
rect 13466 1035 13504 1069
rect 13538 1035 13576 1069
rect 13610 1035 13648 1069
rect 13682 1035 13720 1069
rect 13754 1035 13792 1069
rect 13857 1035 13864 1069
rect 13925 1035 13936 1069
rect 13060 1029 13805 1035
tri 13511 1027 13513 1029 ne
rect 13513 1027 13805 1029
rect 13857 1027 13873 1035
rect 13925 1027 13941 1035
rect 13993 1027 14008 1079
rect 14060 1027 14075 1079
rect 14127 1027 14142 1079
rect 14194 1027 14209 1079
rect 14261 1027 14276 1079
rect 14328 1069 14343 1079
rect 14395 1069 14410 1079
rect 14462 1069 14477 1079
rect 14529 1069 14544 1079
rect 14596 1069 14611 1079
rect 14663 1069 14678 1079
rect 14730 1069 14745 1079
rect 14797 1069 14812 1079
rect 14864 1069 14879 1079
rect 14931 1069 14946 1079
rect 14998 1069 15062 1079
rect 14330 1035 14343 1069
rect 14402 1035 14410 1069
rect 14474 1035 14477 1069
rect 14797 1035 14800 1069
rect 14864 1035 14872 1069
rect 14931 1035 14944 1069
rect 14998 1035 15016 1069
rect 15050 1035 15062 1069
rect 14328 1027 14343 1035
rect 14395 1027 14410 1035
rect 14462 1027 14477 1035
rect 14529 1027 14544 1035
rect 14596 1027 14611 1035
rect 14663 1027 14678 1035
rect 14730 1027 14745 1035
rect 14797 1027 14812 1035
rect 14864 1027 14879 1035
rect 14931 1027 14946 1035
rect 14998 1027 15062 1035
rect 15116 1073 15169 1095
tri 15169 1073 15191 1095 nw
tri 15282 1073 15304 1095 ne
rect 15304 1073 15364 1095
tri 15364 1073 15386 1095 nw
tri 15537 1073 15559 1095 ne
rect 15559 1073 15619 1095
tri 15619 1073 15641 1095 nw
tri 15792 1073 15814 1095 ne
rect 15814 1073 15867 1095
rect 15116 1057 15162 1073
tri 15162 1066 15169 1073 nw
tri 15304 1066 15311 1073 ne
rect 15311 1067 15358 1073
tri 15358 1067 15364 1073 nw
tri 15559 1067 15565 1073 ne
rect 15565 1067 15612 1073
rect 12953 893 12959 927
rect 12993 893 12999 927
rect 12953 805 12999 893
rect 15116 1023 15122 1057
rect 15156 1023 15162 1057
rect 15311 1063 15357 1067
tri 15357 1066 15358 1067 nw
rect 15116 979 15162 1023
rect 15116 945 15122 979
rect 15156 945 15162 979
rect 15116 901 15162 945
rect 15116 867 15122 901
rect 15156 867 15162 901
rect 12953 771 12959 805
rect 12993 771 12999 805
rect 13060 833 13289 842
rect 13060 799 13072 833
rect 13106 799 13144 833
rect 13178 799 13216 833
rect 13250 799 13288 833
rect 13060 790 13289 799
rect 13341 790 13354 842
rect 13406 790 13419 842
rect 13471 790 13484 842
rect 13536 833 13549 842
rect 13601 833 13614 842
rect 13666 833 13678 842
rect 13730 839 13736 842
tri 13736 839 13739 842 sw
tri 14474 839 14477 842 se
rect 14477 839 14484 842
rect 13730 833 14484 839
rect 14536 833 14555 842
rect 14607 833 14626 842
rect 14678 833 14697 842
rect 14749 833 14768 842
rect 14820 833 14838 842
rect 14890 833 14908 842
rect 14960 839 14966 842
tri 14966 839 14969 842 sw
rect 14960 833 15062 839
rect 13538 799 13549 833
rect 13610 799 13614 833
rect 13754 799 13792 833
rect 13826 799 13864 833
rect 13898 799 13936 833
rect 13970 799 14008 833
rect 14042 799 14080 833
rect 14114 799 14152 833
rect 14186 799 14224 833
rect 14258 799 14296 833
rect 14330 799 14368 833
rect 14402 799 14440 833
rect 14474 799 14484 833
rect 14546 799 14555 833
rect 14618 799 14626 833
rect 14690 799 14697 833
rect 14762 799 14768 833
rect 14834 799 14838 833
rect 14906 799 14908 833
rect 14978 799 15016 833
rect 15050 799 15062 833
rect 13536 790 13549 799
rect 13601 790 13614 799
rect 13666 790 13678 799
rect 13730 793 14484 799
rect 13730 790 13736 793
tri 13736 790 13739 793 nw
tri 14474 790 14477 793 ne
rect 14477 790 14484 793
rect 14536 790 14555 799
rect 14607 790 14626 799
rect 14678 790 14697 799
rect 14749 790 14768 799
rect 14820 790 14838 799
rect 14890 790 14908 799
rect 14960 793 15062 799
rect 15116 823 15162 867
rect 14960 790 14966 793
tri 14966 790 14969 793 nw
rect 12953 759 12999 771
rect 15116 789 15122 823
rect 15156 789 15162 823
rect 12595 748 12747 759
tri 12747 748 12758 759 nw
rect 12595 745 12744 748
tri 12744 745 12747 748 nw
rect 15116 745 15162 789
rect 12595 736 12718 745
rect 12437 698 12718 736
tri 12718 719 12744 745 nw
rect 12437 664 12561 698
rect 12595 664 12718 698
rect 12437 636 12718 664
rect 12437 626 12678 636
rect 12437 592 12561 626
rect 12595 602 12678 626
rect 12712 602 12718 636
rect 15116 711 15122 745
rect 15156 711 15162 745
rect 15116 667 15162 711
rect 15116 633 15122 667
rect 15156 633 15162 667
tri 13796 603 13799 606 se
rect 13799 603 13805 606
rect 12595 592 12718 602
rect 12437 560 12718 592
rect 12437 554 12678 560
rect 12437 520 12561 554
rect 12595 526 12678 554
rect 12712 526 12718 560
rect 13060 597 13805 603
rect 13857 597 13876 606
rect 13928 597 13947 606
rect 13999 597 14018 606
rect 14070 597 14089 606
rect 14141 597 14159 606
rect 14211 597 14229 606
rect 14281 597 14299 606
rect 14351 603 14357 606
tri 14357 603 14360 606 sw
rect 14351 597 15062 603
rect 13060 563 13072 597
rect 13106 563 13144 597
rect 13178 563 13216 597
rect 13250 563 13288 597
rect 13322 563 13360 597
rect 13394 563 13432 597
rect 13466 563 13504 597
rect 13538 563 13576 597
rect 13610 563 13648 597
rect 13682 563 13720 597
rect 13754 563 13792 597
rect 13857 563 13864 597
rect 13928 563 13936 597
rect 13999 563 14008 597
rect 14070 563 14080 597
rect 14141 563 14152 597
rect 14211 563 14224 597
rect 14281 563 14296 597
rect 14351 563 14368 597
rect 14402 563 14440 597
rect 14474 563 14512 597
rect 14546 563 14584 597
rect 14618 563 14656 597
rect 14690 563 14728 597
rect 14762 563 14800 597
rect 14834 563 14872 597
rect 14906 563 14944 597
rect 14978 563 15016 597
rect 15050 563 15062 597
rect 13060 557 13805 563
tri 13796 555 13798 557 ne
rect 13798 555 13805 557
tri 13798 554 13799 555 ne
rect 13799 554 13805 555
rect 13857 554 13876 563
rect 13928 554 13947 563
rect 13999 554 14018 563
rect 14070 554 14089 563
rect 14141 554 14159 563
rect 14211 554 14229 563
rect 14281 554 14299 563
rect 14351 557 15062 563
rect 15116 589 15162 633
rect 14351 556 14359 557
tri 14359 556 14360 557 nw
rect 14351 555 14358 556
tri 14358 555 14359 556 nw
tri 15115 555 15116 556 se
rect 15116 555 15122 589
rect 15156 555 15162 589
rect 14351 554 14357 555
tri 14357 554 14358 555 nw
tri 15114 554 15115 555 se
rect 15115 554 15162 555
tri 15107 547 15114 554 se
rect 15114 547 15162 554
tri 15103 543 15107 547 se
rect 15107 543 15162 547
rect 12595 520 12718 526
tri 15082 522 15103 543 se
rect 15103 522 15162 543
rect 15214 1038 15266 1050
rect 15214 1004 15223 1038
rect 15257 1004 15266 1038
rect 15214 966 15266 1004
rect 15214 932 15223 966
rect 15257 932 15266 966
rect 15214 894 15266 932
rect 15214 860 15223 894
rect 15257 860 15266 894
rect 15214 671 15266 860
rect 15214 597 15266 619
rect 15214 523 15266 545
rect 12437 484 12718 520
rect 12437 482 12678 484
rect 12437 448 12561 482
rect 12595 450 12678 482
rect 12712 450 12718 484
rect 12595 448 12718 450
rect 12437 410 12718 448
rect 12437 376 12561 410
rect 12595 408 12718 410
rect 12595 376 12678 408
rect 12437 374 12678 376
rect 12712 374 12718 408
rect 12437 338 12718 374
rect 12437 304 12561 338
rect 12595 332 12718 338
rect 12595 304 12678 332
rect 12437 298 12678 304
rect 12712 298 12718 332
rect 12437 266 12718 298
rect 12758 516 15162 522
rect 12810 482 12816 516
rect 12850 482 12889 516
rect 12923 482 12962 516
rect 12810 464 12962 482
rect 12758 444 12962 464
rect 12758 433 12816 444
rect 12810 410 12816 433
rect 12850 410 12889 444
rect 12923 410 12962 444
rect 15084 514 15162 516
tri 15162 514 15170 522 sw
rect 15084 511 15170 514
rect 15084 477 15122 511
rect 15156 510 15170 511
tri 15170 510 15174 514 sw
rect 15156 477 15174 510
rect 15084 433 15174 477
rect 15084 410 15122 433
rect 12810 404 15122 410
rect 12810 399 12952 404
tri 12952 399 12957 404 nw
tri 15075 399 15080 404 ne
rect 15080 399 15122 404
rect 15156 399 15174 433
rect 12810 392 12945 399
tri 12945 392 12952 399 nw
tri 15080 392 15087 399 ne
rect 15087 392 15174 399
rect 12810 381 12923 392
rect 12758 370 12923 381
tri 12923 370 12945 392 nw
tri 15087 370 15109 392 ne
rect 12758 361 12914 370
tri 12914 361 12923 370 nw
tri 13281 367 13283 369 se
rect 13283 367 13289 369
rect 13060 361 13289 367
rect 12758 350 12880 361
rect 12810 327 12880 350
tri 12880 327 12914 361 nw
rect 13060 327 13072 361
rect 13106 327 13144 361
rect 13178 327 13216 361
rect 13250 327 13288 361
rect 12810 298 12875 327
tri 12875 322 12880 327 nw
rect 13060 321 13289 327
tri 13279 320 13280 321 ne
rect 13280 320 13289 321
tri 13280 317 13283 320 ne
rect 13283 317 13289 320
rect 13341 317 13354 369
rect 13406 317 13419 369
rect 13471 317 13484 369
rect 13536 361 13549 369
rect 13601 361 13614 369
rect 13666 361 13678 369
rect 13730 367 13830 369
tri 13830 367 13832 369 sw
tri 14475 367 14477 369 se
rect 14477 367 14484 369
rect 13730 361 14484 367
rect 14536 361 14555 369
rect 14607 361 14626 369
rect 14678 361 14697 369
rect 14749 361 14768 369
rect 14820 361 14838 369
rect 14890 361 14908 369
rect 14960 367 14966 369
tri 14966 367 14968 369 sw
rect 14960 361 15062 367
rect 13538 327 13549 361
rect 13610 327 13614 361
rect 13754 327 13792 361
rect 13826 327 13864 361
rect 13898 327 13936 361
rect 13970 327 14008 361
rect 14042 327 14080 361
rect 14114 327 14152 361
rect 14186 327 14224 361
rect 14258 327 14296 361
rect 14330 327 14368 361
rect 14402 327 14440 361
rect 14474 327 14484 361
rect 14546 327 14555 361
rect 14618 327 14626 361
rect 14690 327 14697 361
rect 14762 327 14768 361
rect 14834 327 14838 361
rect 14906 327 14908 361
rect 14978 327 15016 361
rect 15050 327 15062 361
rect 13536 317 13549 327
rect 13601 317 13614 327
rect 13666 317 13678 327
rect 13730 321 14484 327
rect 13730 320 13833 321
tri 13833 320 13834 321 nw
tri 14474 320 14475 321 ne
rect 14475 320 14484 321
rect 13730 317 13830 320
tri 13830 317 13833 320 nw
tri 14475 317 14478 320 ne
rect 14478 317 14484 320
rect 14536 317 14555 327
rect 14607 317 14626 327
rect 14678 317 14697 327
rect 14749 317 14768 327
rect 14820 317 14838 327
rect 14890 317 14908 327
rect 14960 321 15062 327
rect 15109 354 15174 392
rect 14960 320 14970 321
tri 14970 320 14971 321 nw
rect 15109 320 15122 354
rect 15156 320 15174 354
rect 14960 317 14967 320
tri 14967 317 14970 320 nw
rect 12758 292 12875 298
rect 12437 232 12561 266
rect 12595 256 12718 266
rect 12595 232 12678 256
rect 12437 222 12678 232
rect 12712 222 12718 256
rect 15109 275 15174 320
rect 15109 241 15122 275
rect 15156 241 15174 275
tri 13155 226 13157 228 se
rect 13157 226 13805 228
rect 12437 194 12718 222
tri 12145 160 12148 163 sw
rect 12437 160 12561 194
rect 12595 180 12718 194
tri 13121 192 13155 226 se
rect 13155 192 13805 226
tri 13119 190 13121 192 se
rect 13121 190 13805 192
rect 12595 160 12678 180
rect 12097 159 12148 160
tri 12148 159 12149 160 sw
rect 12097 151 12149 159
rect 12097 88 12105 99
rect 12139 88 12149 99
rect 12097 57 12149 88
rect 12097 -22 12149 5
rect 12097 -38 12105 -22
rect 12139 -38 12149 -22
rect 12097 -96 12149 -90
rect 12437 151 12678 160
rect 12712 168 12718 180
tri 13105 176 13119 190 se
rect 13119 176 13805 190
rect 13857 176 13876 228
rect 13928 176 13947 228
rect 13999 176 14018 228
rect 14070 176 14089 228
rect 14141 176 14159 228
rect 14211 176 14229 228
rect 14281 176 14299 228
rect 14351 176 15062 228
tri 12718 168 12726 176 sw
tri 13097 168 13105 176 se
rect 13105 168 15062 176
rect 12712 160 12726 168
tri 12726 160 12734 168 sw
tri 13089 160 13097 168 se
rect 13097 160 15062 168
rect 12712 157 12734 160
tri 12734 157 12737 160 sw
tri 13086 157 13089 160 se
rect 13089 157 15062 160
rect 12712 151 12737 157
tri 13083 154 13086 157 se
rect 13086 154 15062 157
rect 12437 99 12438 151
rect 12490 99 12520 151
rect 12572 122 12602 151
rect 12595 99 12602 122
rect 12654 146 12678 151
rect 12654 104 12684 146
rect 12654 99 12678 104
rect 12736 99 12737 151
rect 12437 88 12561 99
rect 12595 88 12678 99
rect 12437 70 12678 88
rect 12712 70 12737 99
tri 13060 131 13083 154 se
rect 13083 131 15062 154
rect 13060 125 15062 131
rect 13060 91 13072 125
rect 13106 91 13144 125
rect 13178 91 13216 125
rect 13250 91 13288 125
rect 13322 91 13360 125
rect 13394 91 13432 125
rect 13466 91 13504 125
rect 13538 91 13576 125
rect 13610 91 13648 125
rect 13682 91 13720 125
rect 13754 91 13792 125
rect 13826 91 13864 125
rect 13898 91 13936 125
rect 13970 91 14008 125
rect 14042 91 14080 125
rect 14114 91 14152 125
rect 14186 91 14224 125
rect 14258 91 14296 125
rect 14330 91 14368 125
rect 14402 91 14440 125
rect 14474 91 14512 125
rect 14546 91 14584 125
rect 14618 91 14656 125
rect 14690 91 14728 125
rect 14762 91 14800 125
rect 14834 91 14872 125
rect 14906 91 14944 125
rect 14978 91 15016 125
rect 15050 91 15062 125
rect 13060 85 15062 91
rect 12437 57 12737 70
rect 12437 5 12438 57
rect 12490 5 12520 57
rect 12572 50 12602 57
rect 12595 16 12602 50
rect 12572 5 12602 16
rect 12654 27 12684 57
rect 12654 5 12678 27
rect 12736 5 12737 57
rect 15109 77 15174 241
rect 15214 448 15266 471
rect 15214 373 15266 396
rect 15214 298 15266 321
rect 15214 264 15223 298
rect 15257 264 15266 298
rect 15214 226 15266 264
rect 15214 192 15223 226
rect 15257 192 15266 226
rect 15214 154 15266 192
rect 15214 120 15223 154
rect 15257 120 15266 154
rect 15214 108 15266 120
rect 15311 1029 15317 1063
rect 15351 1029 15357 1063
rect 15311 983 15357 1029
rect 15311 949 15317 983
rect 15351 949 15357 983
rect 15311 903 15357 949
rect 15311 869 15317 903
rect 15351 869 15357 903
rect 15311 823 15357 869
rect 15311 789 15317 823
rect 15351 789 15357 823
rect 15311 743 15357 789
rect 15311 709 15317 743
rect 15351 709 15357 743
rect 15311 663 15357 709
rect 15311 629 15317 663
rect 15351 629 15357 663
rect 15311 584 15357 629
rect 15311 550 15317 584
rect 15351 550 15357 584
rect 15311 505 15357 550
rect 15311 471 15317 505
rect 15351 471 15357 505
rect 15311 426 15357 471
rect 15311 392 15317 426
rect 15351 392 15357 426
tri 15309 105 15311 107 se
rect 15311 105 15357 392
rect 15452 1061 15504 1067
tri 15565 1066 15566 1067 ne
rect 15452 1004 15459 1009
rect 15493 1004 15504 1009
rect 15452 996 15504 1004
rect 15452 932 15459 944
rect 15493 932 15504 944
rect 15452 931 15504 932
rect 15452 866 15459 879
rect 15493 866 15504 879
rect 15452 800 15504 814
rect 15452 653 15504 748
rect 15452 619 15459 653
rect 15493 619 15504 653
rect 15452 581 15504 619
rect 15452 547 15459 581
rect 15493 547 15504 581
rect 15452 509 15504 547
rect 15452 475 15459 509
rect 15493 475 15504 509
rect 15452 298 15504 475
rect 15452 264 15459 298
rect 15493 264 15504 298
rect 15452 226 15504 264
rect 15452 192 15459 226
rect 15493 192 15504 226
rect 15452 154 15504 192
rect 15452 120 15459 154
rect 15493 120 15504 154
rect 15452 108 15504 120
rect 15566 1058 15612 1067
tri 15612 1066 15619 1073 nw
tri 15814 1066 15821 1073 ne
rect 15566 1024 15572 1058
rect 15606 1024 15612 1058
rect 15821 1063 15867 1073
rect 16346 1073 16392 1085
rect 15566 981 15612 1024
rect 15566 947 15572 981
rect 15606 947 15612 981
rect 15566 904 15612 947
rect 15566 870 15572 904
rect 15606 870 15612 904
rect 15566 826 15612 870
rect 15566 792 15572 826
rect 15606 792 15612 826
rect 15566 748 15612 792
rect 15566 714 15572 748
rect 15606 714 15612 748
rect 15566 670 15612 714
rect 15689 1038 15735 1050
rect 15689 1004 15695 1038
rect 15729 1004 15735 1038
rect 15689 966 15735 1004
rect 15689 932 15695 966
rect 15729 932 15735 966
rect 15689 894 15735 932
rect 15689 860 15695 894
rect 15729 860 15735 894
rect 15689 681 15735 860
rect 15821 1029 15827 1063
rect 15861 1029 15867 1063
rect 15821 988 15867 1029
rect 15821 954 15827 988
rect 15861 954 15867 988
rect 15821 913 15867 954
rect 15821 879 15827 913
rect 15861 879 15867 913
rect 15821 839 15867 879
rect 15821 805 15827 839
rect 15861 805 15867 839
rect 15821 765 15867 805
rect 15821 731 15827 765
rect 15861 731 15867 765
rect 15821 691 15867 731
tri 15735 681 15739 685 sw
rect 15566 636 15572 670
rect 15606 636 15612 670
rect 15566 592 15612 636
rect 15566 558 15572 592
rect 15606 558 15612 592
rect 15566 514 15612 558
rect 15566 480 15572 514
rect 15606 480 15612 514
rect 15566 436 15612 480
rect 15566 402 15572 436
rect 15606 402 15612 436
rect 15566 358 15612 402
rect 15566 324 15572 358
rect 15606 324 15612 358
rect 15566 280 15612 324
tri 15687 677 15689 679 se
rect 15689 677 15739 681
rect 15687 671 15739 677
rect 15687 597 15739 619
rect 15687 523 15739 545
rect 15687 448 15739 471
rect 15687 373 15739 396
rect 15821 657 15827 691
rect 15861 657 15867 691
rect 15821 617 15867 657
rect 15821 583 15827 617
rect 15861 583 15867 617
rect 15821 543 15867 583
rect 15821 509 15827 543
rect 15861 509 15867 543
rect 15821 469 15867 509
rect 15821 435 15827 469
rect 15861 435 15867 469
rect 15924 1061 15976 1067
rect 15924 1004 15931 1009
rect 15965 1004 15976 1009
rect 15924 996 15976 1004
rect 15924 932 15931 944
rect 15965 932 15976 944
rect 15924 931 15976 932
rect 15924 866 15931 879
rect 15965 866 15976 879
rect 15924 800 15976 814
rect 15924 653 15976 748
rect 15924 619 15931 653
rect 15965 619 15976 653
rect 15924 581 15976 619
rect 15924 547 15931 581
rect 15965 547 15976 581
rect 15924 509 15976 547
rect 15924 475 15931 509
rect 15965 475 15976 509
rect 15924 463 15976 475
rect 16043 1051 16089 1063
rect 16043 1017 16049 1051
rect 16083 1017 16089 1051
rect 16043 978 16089 1017
rect 16043 944 16049 978
rect 16083 944 16089 978
rect 16043 905 16089 944
rect 16043 871 16049 905
rect 16083 871 16089 905
rect 16043 832 16089 871
rect 16043 798 16049 832
rect 16083 798 16089 832
rect 16043 759 16089 798
rect 16043 725 16049 759
rect 16083 725 16089 759
rect 16043 686 16089 725
rect 16043 652 16049 686
rect 16083 652 16089 686
rect 16043 613 16089 652
rect 16043 579 16049 613
rect 16083 579 16089 613
rect 16043 540 16089 579
rect 16043 506 16049 540
rect 16083 506 16089 540
rect 16043 467 16089 506
rect 15821 428 15867 435
rect 16043 433 16049 467
rect 16083 433 16089 467
tri 15867 428 15869 430 sw
tri 16041 428 16043 430 se
rect 16043 428 16089 433
rect 15821 407 15869 428
tri 15869 407 15890 428 sw
tri 16020 407 16041 428 se
rect 16041 407 16089 428
rect 15821 401 15890 407
tri 15890 401 15896 407 sw
tri 16014 401 16020 407 se
rect 16020 401 16089 407
rect 15821 395 16089 401
rect 15821 361 15899 395
rect 15933 361 15974 395
rect 16008 361 16089 395
rect 15821 355 16089 361
rect 16159 1038 16211 1050
rect 16159 1004 16167 1038
rect 16201 1004 16211 1038
rect 16159 966 16211 1004
rect 16159 932 16167 966
rect 16201 932 16211 966
rect 16159 894 16211 932
rect 16159 860 16167 894
rect 16201 860 16211 894
rect 16159 671 16211 860
rect 16159 597 16211 619
rect 16159 523 16211 545
rect 16159 448 16211 471
rect 16159 373 16211 396
rect 15687 315 15739 321
rect 15687 313 15735 315
tri 15687 311 15689 313 ne
rect 15566 246 15572 280
rect 15606 246 15612 280
rect 15566 202 15612 246
rect 15566 168 15572 202
rect 15606 168 15612 202
tri 15307 103 15309 105 se
rect 15309 103 15357 105
tri 15564 103 15566 105 se
rect 15566 103 15612 168
rect 15689 298 15735 313
tri 15735 311 15739 315 nw
rect 16159 310 16211 321
rect 16346 1039 16352 1073
rect 16386 1039 16392 1073
rect 16346 999 16392 1039
rect 16346 965 16352 999
rect 16386 965 16392 999
rect 16346 925 16392 965
rect 16346 891 16352 925
rect 16386 891 16392 925
rect 16346 851 16392 891
rect 16346 817 16352 851
rect 16386 817 16392 851
rect 16346 777 16392 817
rect 16346 743 16352 777
rect 16386 743 16392 777
rect 16346 703 16392 743
rect 16346 669 16352 703
rect 16386 669 16392 703
rect 16346 629 16392 669
rect 16346 595 16352 629
rect 16386 595 16392 629
rect 16346 555 16392 595
rect 16346 521 16352 555
rect 16386 521 16392 555
rect 16346 481 16392 521
rect 16346 447 16352 481
rect 16386 447 16392 481
rect 16346 407 16392 447
rect 16346 373 16352 407
rect 16386 373 16392 407
rect 16346 333 16392 373
rect 15689 264 15695 298
rect 15729 264 15735 298
rect 16346 299 16352 333
rect 16386 299 16392 333
rect 15689 226 15735 264
rect 15689 192 15695 226
rect 15729 192 15735 226
rect 15895 216 15901 268
rect 15953 216 15971 268
rect 16023 216 16029 268
rect 16085 259 16219 265
tri 16082 225 16085 228 se
rect 16085 225 16097 259
rect 16131 225 16173 259
rect 16207 225 16219 259
tri 16080 223 16082 225 se
rect 16082 223 16219 225
tri 16073 216 16080 223 se
rect 16080 219 16219 223
rect 16346 259 16392 299
rect 16346 225 16352 259
rect 16386 225 16392 259
rect 16080 216 16117 219
tri 16057 200 16073 216 se
rect 16073 200 16117 216
tri 16117 200 16136 219 nw
rect 15689 154 15735 192
tri 16042 185 16057 200 se
rect 16057 185 16102 200
tri 16102 185 16117 200 nw
rect 16346 185 16392 225
tri 16034 177 16042 185 se
rect 16042 177 16094 185
tri 16094 177 16102 185 nw
rect 16034 168 16085 177
tri 16085 168 16094 177 nw
rect 15689 120 15695 154
rect 15729 120 15735 154
rect 15689 108 15735 120
rect 15878 143 15924 155
rect 15878 109 15884 143
rect 15918 109 15924 143
tri 15874 103 15878 107 se
rect 15878 103 15924 109
tri 15303 99 15307 103 se
rect 15307 99 15357 103
tri 15174 77 15196 99 sw
tri 15281 77 15303 99 se
rect 15303 77 15357 99
tri 15357 77 15383 103 sw
tri 15538 77 15564 103 se
rect 15564 77 15612 103
tri 15612 77 15638 103 sw
tri 15848 77 15874 103 se
rect 15874 77 15924 103
rect 15109 75 15196 77
tri 15196 75 15198 77 sw
tri 15279 75 15281 77 se
rect 15281 75 15383 77
tri 15383 75 15385 77 sw
tri 15536 75 15538 77 se
rect 15538 75 15638 77
tri 15638 75 15640 77 sw
tri 15846 75 15848 77 se
rect 15848 75 15924 77
rect 15109 71 15924 75
rect 15109 37 15884 71
rect 15918 37 15924 71
rect 15109 35 15924 37
tri 15109 27 15117 35 ne
rect 15117 27 15924 35
rect 12437 -7 12678 5
rect 12712 3 12737 5
tri 12737 3 12761 27 sw
tri 15117 3 15141 27 ne
rect 15141 3 15924 27
rect 12712 -1 12761 3
tri 12761 -1 12765 3 sw
tri 15846 -1 15850 3 ne
rect 15850 -1 15924 3
rect 12712 -2 12765 -1
tri 12765 -2 12766 -1 sw
tri 15850 -2 15851 -1 ne
rect 15851 -2 15884 -1
rect 12712 -7 12766 -2
rect 12437 -22 12766 -7
rect 12437 -38 12561 -22
rect 12595 -25 12766 -22
tri 12766 -25 12789 -2 sw
tri 15851 -25 15874 -2 ne
rect 15874 -25 15884 -2
rect 12595 -29 12789 -25
tri 12789 -29 12793 -25 sw
tri 15874 -29 15878 -25 ne
rect 12595 -30 12793 -29
tri 12793 -30 12794 -29 sw
rect 12595 -36 15821 -30
rect 12595 -38 13146 -36
rect 12437 -90 12438 -38
rect 12490 -90 12520 -38
rect 12595 -56 12602 -38
rect 12572 -90 12602 -56
rect 12654 -50 12684 -38
rect 12654 -84 12678 -50
rect 12736 -70 13146 -38
rect 13180 -70 13219 -36
rect 13253 -70 13292 -36
rect 13326 -70 13365 -36
rect 13399 -70 13438 -36
rect 13472 -70 13511 -36
rect 13545 -70 13584 -36
rect 13618 -70 13657 -36
rect 13691 -70 13730 -36
rect 13764 -70 13803 -36
rect 13837 -70 13876 -36
rect 13910 -70 13949 -36
rect 13983 -70 14022 -36
rect 14056 -70 14095 -36
rect 14129 -70 14168 -36
rect 14202 -70 14241 -36
rect 14275 -70 14314 -36
rect 14348 -70 14387 -36
rect 14421 -70 14460 -36
rect 14494 -70 14533 -36
rect 14567 -70 14606 -36
rect 14640 -70 14679 -36
rect 14713 -70 14752 -36
rect 14786 -70 14825 -36
rect 14859 -70 14898 -36
rect 14932 -70 14971 -36
rect 15005 -70 15043 -36
rect 15077 -70 15115 -36
rect 15149 -70 15187 -36
rect 15221 -70 15259 -36
rect 15293 -70 15331 -36
rect 15365 -70 15403 -36
rect 15437 -70 15475 -36
rect 15509 -70 15547 -36
rect 15581 -70 15619 -36
rect 15653 -69 15821 -36
rect 15653 -70 15709 -69
rect 12736 -76 15709 -70
rect 12654 -90 12684 -84
rect 12736 -90 12737 -76
rect 12437 -96 12737 -90
tri 12737 -96 12757 -76 nw
tri 15658 -96 15678 -76 ne
rect 15678 -96 15709 -76
tri 15678 -103 15685 -96 ne
rect 15685 -103 15709 -96
rect 15743 -103 15781 -69
rect 15815 -103 15821 -69
tri 15685 -107 15689 -103 ne
rect 15689 -107 15821 -103
tri 15689 -113 15695 -107 ne
rect 15695 -113 15821 -107
tri 15695 -114 15696 -113 ne
rect 15696 -114 15821 -113
tri 15696 -121 15703 -114 ne
tri 2332 -215 2337 -210 sw
rect 2145 -260 2191 -220
tri 2268 -227 2280 -215 se
rect 2280 -219 2337 -215
tri 2337 -219 2341 -215 sw
rect 7418 -219 7808 -167
rect 15703 -142 15821 -114
rect 15703 -176 15709 -142
rect 15743 -176 15781 -142
rect 15815 -176 15821 -142
rect 15703 -215 15821 -176
rect 2280 -227 2341 -219
tri 2341 -227 2349 -219 sw
rect 2145 -294 2151 -260
rect 2185 -294 2191 -260
rect 2221 -279 2227 -227
rect 2279 -279 2291 -227
rect 2343 -279 2349 -227
rect 15703 -249 15709 -215
rect 15743 -249 15781 -215
rect 15815 -249 15821 -215
tri 3355 -279 3366 -268 se
rect 3366 -279 3375 -268
tri 3346 -288 3355 -279 se
rect 3355 -288 3375 -279
tri 3342 -292 3346 -288 se
rect 3346 -292 3375 -288
rect 2145 -322 2191 -294
tri 2191 -322 2221 -292 sw
tri 3312 -322 3342 -292 se
rect 3342 -322 3375 -292
rect 2145 -323 2221 -322
tri 2221 -323 2222 -322 sw
tri 3311 -323 3312 -322 se
rect 3312 -323 3375 -322
rect 2145 -326 2222 -323
tri 2222 -326 2225 -323 sw
tri 3308 -326 3311 -323 se
rect 3311 -326 3375 -323
rect 15703 -288 15821 -249
rect 15703 -322 15709 -288
rect 15743 -322 15781 -288
rect 15815 -322 15821 -288
rect 2145 -332 3366 -326
rect 2145 -366 2227 -332
rect 2261 -366 2303 -332
rect 2337 -366 2379 -332
rect 2413 -366 2455 -332
rect 2489 -366 2531 -332
rect 2565 -366 2607 -332
rect 2641 -366 2683 -332
rect 2717 -366 2759 -332
rect 2793 -366 2835 -332
rect 2869 -366 2911 -332
rect 2945 -366 2987 -332
rect 3021 -366 3063 -332
rect 3097 -366 3140 -332
rect 3174 -366 3217 -332
rect 3251 -366 3294 -332
rect 3328 -366 3366 -332
rect 2145 -372 3366 -366
rect 15703 -361 15821 -322
tri 3308 -395 3331 -372 ne
rect 3331 -395 3375 -372
tri 3331 -412 3348 -395 ne
rect 3348 -412 3375 -395
rect 15703 -395 15709 -361
rect 15743 -395 15781 -361
rect 15815 -395 15821 -361
tri 3348 -413 3349 -412 ne
rect 3349 -413 3375 -412
tri 15702 -413 15703 -412 se
rect 15703 -413 15821 -395
tri 3349 -422 3358 -413 ne
rect 3358 -422 3375 -413
tri 15693 -422 15702 -413 se
rect 15702 -422 15821 -413
rect 2132 -428 2184 -422
tri 3358 -429 3365 -422 ne
rect 3365 -429 3375 -422
tri 15686 -429 15693 -422 se
rect 15693 -429 15821 -422
tri 3365 -430 3366 -429 ne
rect 3366 -430 3375 -429
rect 2132 -492 2184 -480
rect 2132 -1501 2184 -544
rect 15703 -434 15821 -429
rect 15703 -468 15709 -434
rect 15743 -468 15781 -434
rect 15815 -468 15821 -434
rect 15703 -507 15821 -468
rect 15703 -541 15709 -507
rect 15743 -541 15781 -507
rect 15815 -541 15821 -507
rect 15703 -580 15821 -541
rect 15703 -614 15709 -580
rect 15743 -614 15781 -580
rect 15815 -614 15821 -580
rect 15703 -653 15821 -614
rect 15703 -687 15709 -653
rect 15743 -687 15781 -653
rect 15815 -687 15821 -653
rect 15703 -727 15821 -687
rect 15703 -761 15709 -727
rect 15743 -761 15781 -727
rect 15815 -761 15821 -727
rect 15703 -801 15821 -761
rect 15703 -835 15709 -801
rect 15743 -835 15781 -801
rect 15815 -835 15821 -801
rect 15703 -862 15821 -835
rect 15878 -35 15884 -25
rect 15918 -35 15924 -1
rect 15878 -73 15924 -35
rect 15878 -107 15884 -73
rect 15918 -107 15924 -73
rect 15878 -145 15924 -107
rect 15878 -179 15884 -145
rect 15918 -179 15924 -145
rect 15878 -217 15924 -179
rect 15878 -251 15884 -217
rect 15918 -251 15924 -217
rect 15878 -289 15924 -251
rect 15878 -323 15884 -289
rect 15918 -323 15924 -289
rect 15878 -361 15924 -323
rect 15878 -395 15884 -361
rect 15918 -395 15924 -361
rect 15878 -433 15924 -395
rect 15878 -467 15884 -433
rect 15918 -467 15924 -433
rect 15878 -505 15924 -467
rect 15878 -539 15884 -505
rect 15918 -539 15924 -505
rect 15878 -577 15924 -539
rect 15878 -611 15884 -577
rect 15918 -611 15924 -577
rect 15878 -649 15924 -611
rect 15878 -683 15884 -649
rect 15918 -683 15924 -649
rect 15878 -721 15924 -683
rect 15878 -755 15884 -721
rect 15918 -755 15924 -721
rect 15878 -793 15924 -755
rect 15878 -827 15884 -793
rect 15918 -827 15924 -793
rect 15878 -839 15924 -827
rect 16034 143 16080 168
tri 16080 163 16085 168 nw
rect 16034 109 16040 143
rect 16074 109 16080 143
rect 16034 71 16080 109
rect 16034 37 16040 71
rect 16074 37 16080 71
rect 16034 -1 16080 37
rect 16034 -35 16040 -1
rect 16074 -35 16080 -1
rect 16034 -73 16080 -35
rect 16034 -107 16040 -73
rect 16074 -107 16080 -73
rect 16034 -145 16080 -107
rect 16034 -179 16040 -145
rect 16074 -179 16080 -145
rect 16034 -217 16080 -179
rect 16034 -251 16040 -217
rect 16074 -251 16080 -217
rect 16034 -289 16080 -251
rect 16034 -323 16040 -289
rect 16074 -323 16080 -289
rect 16034 -361 16080 -323
rect 16034 -395 16040 -361
rect 16074 -395 16080 -361
rect 16034 -433 16080 -395
rect 16034 -467 16040 -433
rect 16074 -467 16080 -433
rect 16034 -505 16080 -467
rect 16034 -539 16040 -505
rect 16074 -539 16080 -505
rect 16034 -577 16080 -539
rect 16034 -611 16040 -577
rect 16074 -611 16080 -577
rect 16034 -649 16080 -611
rect 16034 -683 16040 -649
rect 16074 -683 16080 -649
rect 16034 -721 16080 -683
rect 16034 -755 16040 -721
rect 16074 -755 16080 -721
rect 16034 -793 16080 -755
rect 16034 -827 16040 -793
rect 16074 -827 16080 -793
tri 16022 -862 16034 -850 se
rect 16034 -862 16080 -827
rect 16187 143 16239 155
rect 16187 129 16196 143
rect 16230 129 16239 143
rect 16187 71 16239 77
rect 16187 56 16196 71
rect 16230 56 16239 71
rect 16187 -1 16239 4
rect 16187 -35 16196 -1
rect 16230 -35 16239 -1
rect 16187 -73 16239 -35
rect 16187 -107 16196 -73
rect 16230 -107 16239 -73
rect 16187 -145 16239 -107
rect 16187 -179 16196 -145
rect 16230 -179 16239 -145
rect 16187 -217 16239 -179
rect 16187 -251 16196 -217
rect 16230 -251 16239 -217
rect 16187 -289 16239 -251
rect 16187 -323 16196 -289
rect 16230 -323 16239 -289
rect 16187 -361 16239 -323
rect 16187 -395 16196 -361
rect 16230 -395 16239 -361
rect 16187 -433 16239 -395
rect 16187 -467 16196 -433
rect 16230 -467 16239 -433
rect 16187 -505 16239 -467
rect 16187 -539 16196 -505
rect 16230 -539 16239 -505
rect 16187 -577 16239 -539
rect 16187 -611 16196 -577
rect 16230 -611 16239 -577
rect 16187 -649 16239 -611
rect 16187 -683 16196 -649
rect 16230 -683 16239 -649
rect 16187 -721 16239 -683
rect 16187 -755 16196 -721
rect 16230 -755 16239 -721
rect 16187 -793 16239 -755
rect 16187 -827 16196 -793
rect 16230 -827 16239 -793
rect 16187 -839 16239 -827
rect 16346 151 16352 185
rect 16386 151 16392 185
rect 16346 111 16392 151
rect 16346 77 16352 111
rect 16386 77 16392 111
rect 16346 37 16392 77
rect 16346 3 16352 37
rect 16386 3 16392 37
rect 16346 -38 16392 3
rect 16346 -72 16352 -38
rect 16386 -72 16392 -38
rect 16346 -113 16392 -72
rect 16346 -147 16352 -113
rect 16386 -147 16392 -113
rect 16346 -188 16392 -147
rect 16346 -222 16352 -188
rect 16386 -222 16392 -188
rect 16346 -263 16392 -222
rect 16346 -297 16352 -263
rect 16386 -297 16392 -263
rect 16346 -338 16392 -297
rect 16346 -372 16352 -338
rect 16386 -372 16392 -338
rect 16346 -413 16392 -372
rect 16346 -447 16352 -413
rect 16386 -447 16392 -413
rect 16346 -488 16392 -447
rect 16346 -522 16352 -488
rect 16386 -522 16392 -488
rect 16346 -563 16392 -522
rect 16346 -597 16352 -563
rect 16386 -597 16392 -563
rect 16346 -638 16392 -597
rect 16346 -672 16352 -638
rect 16386 -672 16392 -638
rect 16346 -713 16392 -672
rect 16346 -747 16352 -713
rect 16386 -747 16392 -713
rect 16346 -788 16392 -747
rect 16346 -822 16352 -788
rect 16386 -822 16392 -788
tri 16345 -850 16346 -849 se
rect 16346 -850 16392 -822
rect 15686 -863 15835 -862
tri 15835 -863 15836 -862 sw
tri 16021 -863 16022 -862 se
rect 16022 -863 16080 -862
tri 16080 -863 16093 -850 sw
tri 16332 -863 16345 -850 se
rect 16345 -863 16392 -850
rect 15686 -867 15836 -863
tri 15836 -867 15840 -863 sw
tri 16017 -867 16021 -863 se
rect 16021 -867 16093 -863
tri 16093 -867 16097 -863 sw
tri 16328 -867 16332 -863 se
rect 16332 -867 16352 -863
rect 15686 -897 15840 -867
tri 15840 -897 15870 -867 sw
tri 15987 -897 16017 -867 se
rect 16017 -897 16097 -867
tri 16097 -897 16127 -867 sw
tri 16298 -897 16328 -867 se
rect 16328 -897 16352 -867
rect 16386 -897 16392 -863
rect 15686 -901 15870 -897
tri 15870 -901 15874 -897 sw
tri 15983 -901 15987 -897 se
rect 15987 -901 16127 -897
tri 16127 -901 16131 -897 sw
tri 16294 -901 16298 -897 se
rect 16298 -901 16392 -897
rect 15686 -935 16392 -901
rect 15686 -969 15917 -935
rect 15951 -969 15990 -935
rect 16024 -969 16063 -935
rect 16097 -969 16136 -935
rect 16170 -969 16208 -935
rect 16242 -969 16280 -935
rect 16314 -969 16392 -935
rect 15686 -1052 16392 -969
rect 16949 -1018 16990 1216
tri 16990 1188 17018 1216 nw
tri 17028 1144 17061 1177 se
rect 17061 1144 18013 1177
tri 17024 1140 17028 1144 se
rect 17028 1140 18013 1144
rect 17024 1125 18013 1140
rect 18065 1125 18077 1177
rect 18129 1125 18135 1177
rect 18857 1150 18903 1216
rect 19967 1344 19973 1378
rect 20007 1344 20013 1378
rect 19967 1300 20013 1344
rect 19967 1266 19973 1300
rect 20007 1266 20013 1300
rect 20246 1433 20347 1550
rect 20246 1399 20252 1433
rect 20286 1399 20347 1433
rect 20246 1325 20347 1399
rect 20246 1291 20252 1325
rect 20286 1291 20347 1325
rect 20246 1274 20347 1291
rect 20505 1544 20868 1551
rect 20505 1492 20519 1544
rect 20571 1492 20592 1544
rect 20644 1492 20665 1544
rect 20717 1492 20738 1544
rect 20790 1492 20810 1544
rect 20862 1492 20868 1544
rect 20505 1474 20868 1492
rect 20505 1422 20519 1474
rect 20571 1422 20592 1474
rect 20644 1422 20665 1474
rect 20717 1422 20738 1474
rect 20790 1422 20810 1474
rect 20862 1422 20868 1474
rect 20505 1404 20868 1422
rect 20505 1352 20519 1404
rect 20571 1352 20592 1404
rect 20644 1352 20665 1404
rect 20717 1352 20738 1404
rect 20790 1352 20810 1404
rect 20862 1352 20868 1404
rect 24462 1352 24664 1888
rect 25297 1828 25427 2023
tri 25427 1994 25456 2023 nw
tri 25944 1888 25972 1916 se
rect 25297 1794 25309 1828
rect 25343 1794 25381 1828
rect 25415 1794 25427 1828
rect 25297 1788 25427 1794
rect 25231 1490 25239 1542
rect 25291 1490 25303 1542
rect 25355 1490 25362 1542
rect 20505 1334 20868 1352
rect 20505 1282 20519 1334
rect 20571 1282 20592 1334
rect 20644 1282 20665 1334
rect 20717 1282 20738 1334
rect 20790 1282 20810 1334
rect 20862 1282 20868 1334
rect 25231 1314 25239 1366
rect 25291 1314 25303 1366
rect 25355 1314 25362 1366
rect 20505 1274 20868 1282
rect 25673 1280 25828 1875
rect 25844 1721 25972 1888
rect 25844 1695 25848 1721
tri 25848 1695 25874 1721 nw
tri 25946 1695 25972 1721 ne
tri 25844 1691 25848 1695 nw
rect 19967 1222 20013 1266
rect 19967 1188 19973 1222
rect 20007 1188 20013 1222
tri 18903 1150 18932 1179 sw
tri 19938 1150 19967 1179 se
rect 19967 1150 20013 1188
rect 18857 1144 20013 1150
rect 17024 1110 17090 1125
tri 17090 1110 17105 1125 nw
rect 18857 1110 18937 1144
rect 18971 1110 19011 1144
rect 19045 1110 19085 1144
rect 19119 1110 19159 1144
rect 19193 1110 19233 1144
rect 19267 1110 19307 1144
rect 19341 1110 19381 1144
rect 19415 1110 19455 1144
rect 19489 1110 19529 1144
rect 19563 1110 19603 1144
rect 19637 1110 19677 1144
rect 19711 1110 19751 1144
rect 19785 1110 19826 1144
rect 19860 1110 19901 1144
rect 19935 1110 20013 1144
rect 17024 -936 17065 1110
tri 17065 1085 17090 1110 nw
rect 18857 1104 20013 1110
rect 18122 1080 18128 1081
tri 17140 1072 17148 1080 se
rect 17148 1072 18128 1080
tri 17118 1050 17140 1072 se
rect 17140 1050 18128 1072
rect 17118 1029 18128 1050
rect 18180 1029 18192 1081
rect 18244 1029 18250 1081
rect 18857 1072 18903 1104
tri 18903 1075 18932 1104 nw
rect 18857 1038 18863 1072
rect 18897 1038 18903 1072
tri 18718 1029 18727 1038 se
rect 17118 -872 17159 1029
tri 17159 998 17190 1029 nw
tri 18687 998 18718 1029 se
rect 18718 998 18727 1029
tri 18684 995 18687 998 se
rect 18687 995 18727 998
tri 18680 991 18684 995 se
rect 18684 991 18727 995
rect 18635 939 18727 991
rect 18857 995 18903 1038
rect 18857 961 18863 995
rect 18897 961 18903 995
rect 18857 918 18903 961
rect 18857 884 18863 918
rect 18897 884 18903 918
rect 18857 842 18903 884
rect 18635 757 18681 809
rect 18857 808 18863 842
rect 18897 808 18903 842
rect 18857 766 18903 808
rect 18857 732 18863 766
rect 18897 732 18903 766
rect 18857 690 18903 732
rect 18857 656 18863 690
rect 18897 656 18903 690
rect 18635 567 18765 619
rect 18857 614 18903 656
rect 18857 580 18863 614
rect 18897 580 18903 614
rect 18857 538 18903 580
rect 18857 504 18863 538
rect 18897 504 18903 538
rect 18857 462 18903 504
rect 18857 428 18863 462
rect 18897 428 18903 462
rect 18370 341 18500 347
rect 18370 307 18382 341
rect 18416 307 18454 341
rect 18488 307 18500 341
rect 18370 301 18500 307
rect 18531 346 18537 398
rect 18589 346 18601 398
rect 18653 346 18659 398
rect 18857 386 18903 428
rect 18857 352 18863 386
rect 18897 352 18903 386
tri 18370 276 18395 301 ne
rect 18395 276 18446 301
tri 18446 276 18471 301 nw
tri 18395 271 18400 276 ne
tri 18395 -170 18400 -165 se
rect 18400 -170 18441 276
tri 18441 271 18446 276 nw
rect 18531 223 18564 346
tri 18564 315 18595 346 nw
rect 18857 310 18903 352
rect 18857 276 18863 310
rect 18897 276 18903 310
rect 18635 257 18765 263
tri 18564 223 18565 224 sw
rect 18635 223 18647 257
rect 18681 223 18719 257
rect 18753 223 18765 257
rect 18531 221 18565 223
tri 18565 221 18567 223 sw
tri 18510 200 18531 221 se
rect 18531 200 18567 221
tri 18567 200 18588 221 sw
tri 18498 188 18510 200 se
rect 18510 188 18588 200
tri 18588 188 18600 200 sw
rect 18470 182 18600 188
rect 18470 148 18482 182
rect 18516 148 18554 182
rect 18588 148 18600 182
rect 18470 142 18600 148
rect 18635 105 18765 223
rect 18857 234 18903 276
rect 18857 200 18863 234
rect 18897 200 18903 234
rect 18857 164 18903 200
rect 19155 282 19354 860
rect 19155 230 19161 282
rect 19213 230 19227 282
rect 19279 230 19354 282
rect 19155 206 19354 230
rect 18857 118 18993 164
rect 18635 71 18647 105
rect 18681 71 18719 105
rect 18753 71 18765 105
rect 18635 65 18765 71
rect 18947 86 18993 118
rect 18635 52 18717 65
tri 18717 52 18730 65 nw
rect 18947 52 18953 86
rect 18987 52 18993 86
rect 18470 26 18600 32
rect 18470 -8 18482 26
rect 18516 -8 18554 26
rect 18588 -8 18600 26
rect 18470 -14 18600 -8
tri 18496 -22 18504 -14 ne
rect 18504 -22 18592 -14
tri 18592 -22 18600 -14 nw
tri 18504 -40 18522 -22 ne
tri 18441 -170 18446 -165 sw
tri 18374 -191 18395 -170 se
rect 18395 -191 18446 -170
tri 18446 -191 18467 -170 sw
rect 18356 -243 18362 -191
rect 18414 -243 18426 -191
rect 18478 -243 18484 -191
rect 18522 -197 18574 -22
tri 18574 -40 18592 -22 nw
rect 18522 -261 18574 -249
rect 18522 -319 18574 -313
tri 18623 -318 18635 -306 se
rect 18635 -318 18696 52
tri 18696 31 18717 52 nw
rect 18947 12 18993 52
rect 18947 -22 18953 12
rect 18987 -22 18993 12
rect 18862 -42 18914 -36
rect 18862 -106 18914 -94
tri 18622 -319 18623 -318 se
rect 18623 -319 18696 -318
tri 18583 -358 18622 -319 se
rect 18622 -346 18696 -319
rect 18622 -358 18684 -346
tri 18684 -358 18696 -346 nw
rect 18751 -120 18803 -114
rect 18751 -184 18803 -172
tri 18581 -360 18583 -358 se
rect 18583 -360 18682 -358
tri 18682 -360 18684 -358 nw
tri 18416 -385 18441 -360 se
rect 18441 -385 18657 -360
tri 18657 -385 18682 -360 nw
rect 18416 -392 18650 -385
tri 18650 -392 18657 -385 nw
rect 18416 -407 18635 -392
tri 18635 -407 18650 -392 nw
rect 18416 -410 18632 -407
tri 18632 -410 18635 -407 nw
rect 18416 -432 18486 -410
tri 18486 -432 18508 -410 nw
rect 18416 -492 18468 -432
tri 18468 -450 18486 -432 nw
tri 17159 -872 17166 -865 sw
rect 17118 -888 17166 -872
tri 17166 -888 17182 -872 sw
tri 17118 -906 17136 -888 ne
rect 17136 -906 17182 -888
tri 17182 -906 17200 -888 sw
tri 17136 -924 17154 -906 ne
rect 17154 -924 17200 -906
tri 17065 -936 17077 -924 sw
tri 17154 -936 17166 -924 ne
rect 17166 -936 17200 -924
tri 17200 -936 17230 -906 sw
rect 17024 -945 17077 -936
tri 17077 -945 17086 -936 sw
tri 17166 -945 17175 -936 ne
rect 17175 -945 17230 -936
tri 17230 -945 17239 -936 sw
rect 17024 -947 17086 -945
tri 17086 -947 17088 -945 sw
tri 17175 -947 17177 -945 ne
rect 17177 -947 17239 -945
tri 17024 -979 17056 -947 ne
rect 17056 -955 17088 -947
tri 17088 -955 17096 -947 sw
tri 17177 -952 17182 -947 ne
rect 17182 -952 17239 -947
tri 17239 -952 17246 -945 sw
tri 17182 -955 17185 -952 ne
rect 17185 -955 17246 -952
rect 17056 -979 17096 -955
tri 17096 -979 17120 -955 sw
tri 17185 -979 17209 -955 ne
rect 17209 -964 17246 -955
tri 17246 -964 17258 -952 sw
rect 17209 -979 17258 -964
tri 17258 -979 17273 -964 sw
tri 17056 -984 17061 -979 ne
rect 17061 -984 17120 -979
tri 17120 -984 17125 -979 sw
tri 17209 -984 17214 -979 ne
rect 17214 -984 17273 -979
tri 17273 -984 17278 -979 sw
tri 17061 -995 17072 -984 ne
rect 17072 -995 17125 -984
tri 16990 -1018 17013 -995 sw
tri 17072 -1011 17088 -995 ne
rect 17088 -1011 17125 -995
tri 17125 -1011 17152 -984 sw
tri 17214 -1011 17241 -984 ne
rect 17241 -1011 17278 -984
tri 17088 -1018 17095 -1011 ne
rect 17095 -1018 17152 -1011
tri 17152 -1018 17159 -1011 sw
tri 17241 -1016 17246 -1011 ne
rect 17246 -1016 17278 -1011
tri 17278 -1016 17310 -984 sw
tri 18250 -1016 18282 -984 se
rect 18282 -1016 18328 -936
tri 17246 -1018 17248 -1016 ne
rect 17248 -1018 17310 -1016
tri 17310 -1018 17312 -1016 sw
tri 18248 -1018 18250 -1016 se
rect 18250 -1018 18328 -1016
rect 16949 -1019 17013 -1018
tri 17013 -1019 17014 -1018 sw
tri 17095 -1019 17096 -1018 ne
rect 17096 -1019 17159 -1018
tri 17159 -1019 17160 -1018 sw
tri 17248 -1019 17249 -1018 ne
rect 17249 -1019 17312 -1018
tri 16392 -1052 16425 -1019 sw
rect 16949 -1021 17014 -1019
tri 17014 -1021 17016 -1019 sw
rect 17096 -1021 17160 -1019
tri 17160 -1021 17162 -1019 sw
tri 17249 -1021 17251 -1019 ne
rect 17251 -1021 17312 -1019
tri 16932 -1038 16949 -1021 se
rect 16949 -1038 17016 -1021
tri 17016 -1038 17033 -1021 sw
rect 15686 -1059 16425 -1052
tri 16425 -1059 16432 -1052 sw
rect 15686 -1060 16758 -1059
tri 15686 -1066 15692 -1060 ne
rect 15692 -1066 16758 -1060
rect 2132 -1580 2184 -1553
rect 2132 -1638 2184 -1632
rect 2225 -1118 2231 -1066
rect 2283 -1118 2295 -1066
rect 2347 -1118 2353 -1066
tri 15692 -1091 15717 -1066 ne
rect 15717 -1091 16758 -1066
tri 16758 -1091 16790 -1059 sw
rect 16905 -1090 16911 -1038
rect 16963 -1090 16975 -1038
rect 17027 -1090 17033 -1038
rect 17096 -1038 17162 -1021
tri 17162 -1038 17179 -1021 sw
tri 17251 -1028 17258 -1021 ne
rect 17258 -1028 17312 -1021
tri 17312 -1028 17322 -1018 sw
tri 18238 -1028 18248 -1018 se
rect 18248 -1028 18328 -1018
rect 17258 -1038 17322 -1028
tri 17322 -1038 17332 -1028 sw
tri 18228 -1038 18238 -1028 se
rect 18238 -1038 18328 -1028
rect 17096 -1090 17102 -1038
rect 17154 -1090 17166 -1038
rect 17218 -1090 17224 -1038
rect 17258 -1090 17264 -1038
rect 17316 -1090 17328 -1038
rect 17380 -1090 17386 -1038
tri 18214 -1052 18228 -1038 se
rect 18228 -1052 18328 -1038
tri 18176 -1090 18214 -1052 se
rect 18214 -1057 18328 -1052
rect 18214 -1081 18304 -1057
tri 18304 -1081 18328 -1057 nw
rect 18214 -1090 18293 -1081
tri 18175 -1091 18176 -1090 se
rect 18176 -1091 18293 -1090
tri 18293 -1091 18303 -1081 nw
tri 15717 -1118 15744 -1091 ne
rect 15744 -1102 16790 -1091
tri 16790 -1102 16801 -1091 sw
tri 18164 -1102 18175 -1091 se
rect 18175 -1102 18282 -1091
tri 18282 -1102 18293 -1091 nw
rect 15744 -1118 16801 -1102
rect 2225 -1125 2317 -1118
tri 2317 -1125 2324 -1118 nw
tri 15744 -1125 15751 -1118 ne
rect 15751 -1125 16801 -1118
tri 16801 -1125 16824 -1102 sw
tri 18141 -1125 18164 -1102 se
rect 18164 -1125 18259 -1102
tri 18259 -1125 18282 -1102 nw
rect 2225 -1134 2308 -1125
tri 2308 -1134 2317 -1125 nw
tri 15751 -1134 15760 -1125 ne
rect 15760 -1134 16824 -1125
tri 16824 -1134 16833 -1125 sw
tri 18132 -1134 18141 -1125 se
rect 18141 -1134 18250 -1125
tri 18250 -1134 18259 -1125 nw
rect 2225 -1740 2281 -1134
tri 2281 -1161 2308 -1134 nw
tri 16726 -1161 16753 -1134 ne
rect 16753 -1161 18220 -1134
tri 16753 -1164 16756 -1161 ne
rect 16756 -1164 18220 -1161
tri 18220 -1164 18250 -1134 nw
tri 16756 -1191 16783 -1164 ne
rect 16783 -1191 18193 -1164
tri 18193 -1191 18220 -1164 nw
rect 17922 -1252 18463 -1226
rect 17922 -1286 17961 -1252
rect 17995 -1286 18037 -1252
rect 18071 -1286 18113 -1252
rect 18147 -1286 18189 -1252
rect 18223 -1286 18265 -1252
rect 18299 -1286 18341 -1252
rect 18375 -1286 18417 -1252
rect 18451 -1286 18463 -1252
rect 17922 -1332 18463 -1286
rect 17922 -1366 17961 -1332
rect 17995 -1366 18037 -1332
rect 18071 -1366 18113 -1332
rect 18147 -1366 18189 -1332
rect 18223 -1366 18265 -1332
rect 18299 -1366 18341 -1332
rect 18375 -1366 18417 -1332
rect 18451 -1366 18463 -1332
rect 17922 -1412 18463 -1366
rect 17922 -1446 17961 -1412
rect 17995 -1446 18037 -1412
rect 18071 -1446 18113 -1412
rect 18147 -1446 18189 -1412
rect 18223 -1446 18265 -1412
rect 18299 -1446 18341 -1412
rect 18375 -1446 18417 -1412
rect 18451 -1446 18463 -1412
rect 17922 -1453 18463 -1446
tri 17922 -1599 18068 -1453 nw
rect 2225 -1792 2227 -1740
rect 2279 -1792 2281 -1740
rect 2225 -1804 2281 -1792
rect 2225 -1856 2227 -1804
rect 2279 -1856 2281 -1804
rect 2225 -1862 2281 -1856
tri 2005 -2670 2011 -2664 se
rect 2011 -2670 2083 -2664
rect 884 -2722 2083 -2670
rect 688 -3231 823 -3225
rect 688 -3265 700 -3231
rect 734 -3265 777 -3231
rect 811 -3265 823 -3231
rect 688 -3432 823 -3265
rect 688 -3484 692 -3432
rect 744 -3484 823 -3432
rect 688 -3496 823 -3484
rect 884 -3369 930 -2722
tri 930 -2748 956 -2722 nw
rect 884 -3403 890 -3369
rect 924 -3403 930 -3369
rect 884 -3441 930 -3403
rect 884 -3475 890 -3441
rect 924 -3475 930 -3441
rect 884 -3487 930 -3475
rect 1033 -3241 1079 -3229
rect 1033 -3275 1039 -3241
rect 1073 -3275 1079 -3241
rect 1033 -3313 1079 -3275
rect 1033 -3347 1039 -3313
rect 1073 -3347 1079 -3313
rect 1033 -3385 1079 -3347
rect 1033 -3419 1039 -3385
rect 1073 -3419 1079 -3385
rect 1033 -3457 1079 -3419
rect 688 -3548 692 -3496
rect 744 -3548 823 -3496
rect 1033 -3491 1039 -3457
rect 1073 -3491 1079 -3457
rect 1033 -3529 1079 -3491
rect 688 -3553 823 -3548
tri 823 -3553 838 -3538 sw
rect 688 -3563 838 -3553
tri 838 -3563 848 -3553 sw
tri 1023 -3563 1033 -3553 se
rect 1033 -3563 1039 -3529
rect 1073 -3563 1079 -3529
rect 688 -3588 848 -3563
tri 848 -3588 873 -3563 sw
tri 998 -3588 1023 -3563 se
rect 1023 -3588 1079 -3563
rect 688 -3601 1079 -3588
rect 688 -3633 1039 -3601
tri 688 -3635 690 -3633 ne
rect 690 -3635 1039 -3633
rect 1073 -3635 1079 -3601
tri 690 -3673 728 -3635 ne
rect 728 -3673 1079 -3635
tri 728 -3707 762 -3673 ne
rect 762 -3707 1039 -3673
rect 1073 -3707 1079 -3673
tri 762 -3745 800 -3707 ne
rect 800 -3745 1079 -3707
tri 800 -3778 833 -3745 ne
rect 833 -3778 1039 -3745
tri 1006 -3779 1007 -3778 ne
rect 1007 -3779 1039 -3778
rect 1073 -3779 1079 -3745
tri 1007 -3805 1033 -3779 ne
rect 1033 -3817 1079 -3779
rect 1033 -3851 1039 -3817
rect 1073 -3851 1079 -3817
rect 1033 -3889 1079 -3851
rect 1033 -3923 1039 -3889
rect 1073 -3923 1079 -3889
rect 1033 -3961 1079 -3923
rect 1033 -3995 1039 -3961
rect 1073 -3995 1079 -3961
rect 1033 -4033 1079 -3995
rect 1033 -4067 1039 -4033
rect 1073 -4067 1079 -4033
rect 1033 -4105 1079 -4067
rect 1033 -4139 1039 -4105
rect 1073 -4139 1079 -4105
rect 1033 -4177 1079 -4139
rect 1033 -4211 1039 -4177
rect 1073 -4211 1079 -4177
tri 1030 -4227 1033 -4224 se
rect 1033 -4227 1079 -4211
tri 1079 -4227 1082 -4224 sw
rect 1030 -4233 1082 -4227
rect 1030 -4299 1082 -4285
rect 1030 -4355 1039 -4351
rect 1073 -4355 1082 -4351
rect 1030 -4365 1082 -4355
rect 1030 -4423 1039 -4417
tri 1030 -4426 1033 -4423 ne
rect 478 -11022 652 -10994
rect 1033 -4427 1039 -4423
rect 1073 -4423 1082 -4417
rect 1691 -4229 1917 -4228
rect 1691 -4281 1697 -4229
rect 1749 -4281 1778 -4229
rect 1830 -4281 1859 -4229
rect 1911 -4281 1917 -4229
rect 1691 -4299 1917 -4281
rect 1691 -4351 1697 -4299
rect 1749 -4351 1778 -4299
rect 1830 -4351 1859 -4299
rect 1911 -4351 1917 -4299
rect 1691 -4369 1917 -4351
rect 1691 -4421 1697 -4369
rect 1749 -4421 1778 -4369
rect 1830 -4421 1859 -4369
rect 1911 -4421 1917 -4369
rect 1691 -4422 1917 -4421
rect 1073 -4427 1079 -4423
tri 1079 -4426 1082 -4423 nw
rect 1033 -4465 1079 -4427
rect 1033 -4499 1039 -4465
rect 1073 -4499 1079 -4465
rect 1033 -4537 1079 -4499
rect 1033 -4571 1039 -4537
rect 1073 -4571 1079 -4537
rect 1033 -4609 1079 -4571
rect 1033 -4643 1039 -4609
rect 1073 -4643 1079 -4609
rect 1033 -4681 1079 -4643
rect 1033 -4715 1039 -4681
rect 1073 -4715 1079 -4681
rect 1033 -4753 1079 -4715
rect 1033 -4787 1039 -4753
rect 1073 -4787 1079 -4753
rect 1033 -4825 1079 -4787
rect 1033 -4859 1039 -4825
rect 1073 -4859 1079 -4825
rect 1033 -4897 1079 -4859
rect 1033 -4931 1039 -4897
rect 1073 -4931 1079 -4897
rect 1033 -4969 1079 -4931
rect 1033 -5003 1039 -4969
rect 1073 -5003 1079 -4969
rect 1033 -5041 1079 -5003
rect 1033 -5075 1039 -5041
rect 1073 -5075 1079 -5041
rect 1033 -5113 1079 -5075
rect 1033 -5147 1039 -5113
rect 1073 -5147 1079 -5113
rect 1033 -5185 1079 -5147
rect 1033 -5219 1039 -5185
rect 1073 -5219 1079 -5185
rect 1033 -5257 1079 -5219
rect 1033 -5291 1039 -5257
rect 1073 -5291 1079 -5257
rect 1033 -5329 1079 -5291
rect 1033 -5363 1039 -5329
rect 1073 -5363 1079 -5329
rect 1033 -5401 1079 -5363
rect 1033 -5435 1039 -5401
rect 1073 -5435 1079 -5401
rect 1033 -5473 1079 -5435
rect 1033 -5507 1039 -5473
rect 1073 -5507 1079 -5473
rect 1033 -5545 1079 -5507
rect 1033 -5579 1039 -5545
rect 1073 -5579 1079 -5545
rect 1033 -5617 1079 -5579
rect 1033 -5651 1039 -5617
rect 1073 -5651 1079 -5617
rect 1033 -5689 1079 -5651
rect 1033 -5723 1039 -5689
rect 1073 -5723 1079 -5689
rect 1033 -5761 1079 -5723
rect 1033 -5795 1039 -5761
rect 1073 -5795 1079 -5761
rect 1033 -5833 1079 -5795
rect 1033 -5867 1039 -5833
rect 1073 -5867 1079 -5833
rect 1033 -5905 1079 -5867
rect 1033 -5939 1039 -5905
rect 1073 -5939 1079 -5905
rect 1033 -5977 1079 -5939
rect 1033 -6011 1039 -5977
rect 1073 -6011 1079 -5977
rect 1033 -6049 1079 -6011
rect 1033 -6083 1039 -6049
rect 1073 -6083 1079 -6049
rect 1033 -6121 1079 -6083
rect 1033 -6155 1039 -6121
rect 1073 -6155 1079 -6121
rect 1033 -6193 1079 -6155
rect 1033 -6227 1039 -6193
rect 1073 -6227 1079 -6193
rect 1033 -6265 1079 -6227
rect 1033 -6299 1039 -6265
rect 1073 -6299 1079 -6265
rect 1033 -6337 1079 -6299
rect 1033 -6371 1039 -6337
rect 1073 -6371 1079 -6337
rect 1033 -6409 1079 -6371
rect 1033 -6443 1039 -6409
rect 1073 -6443 1079 -6409
rect 1033 -6481 1079 -6443
rect 1033 -6515 1039 -6481
rect 1073 -6515 1079 -6481
rect 1033 -6553 1079 -6515
rect 1033 -6587 1039 -6553
rect 1073 -6587 1079 -6553
rect 1033 -6625 1079 -6587
rect 1033 -6659 1039 -6625
rect 1073 -6659 1079 -6625
rect 1033 -6697 1079 -6659
rect 1033 -6731 1039 -6697
rect 1073 -6731 1079 -6697
rect 1033 -6769 1079 -6731
rect 1033 -6803 1039 -6769
rect 1073 -6803 1079 -6769
rect 1033 -6841 1079 -6803
rect 1033 -6875 1039 -6841
rect 1073 -6875 1079 -6841
rect 1033 -6913 1079 -6875
rect 1033 -6947 1039 -6913
rect 1073 -6947 1079 -6913
rect 1033 -6985 1079 -6947
rect 1033 -7019 1039 -6985
rect 1073 -7019 1079 -6985
rect 1033 -7057 1079 -7019
rect 1033 -7091 1039 -7057
rect 1073 -7091 1079 -7057
rect 1033 -7129 1079 -7091
rect 1033 -7163 1039 -7129
rect 1073 -7163 1079 -7129
rect 1033 -7201 1079 -7163
rect 1033 -7235 1039 -7201
rect 1073 -7235 1079 -7201
rect 1033 -7273 1079 -7235
rect 1033 -7307 1039 -7273
rect 1073 -7307 1079 -7273
rect 1033 -7345 1079 -7307
rect 1033 -7379 1039 -7345
rect 1073 -7379 1079 -7345
rect 1033 -7417 1079 -7379
rect 1033 -7451 1039 -7417
rect 1073 -7451 1079 -7417
rect 1033 -7489 1079 -7451
rect 1033 -7523 1039 -7489
rect 1073 -7523 1079 -7489
rect 1033 -7561 1079 -7523
rect 1033 -7595 1039 -7561
rect 1073 -7595 1079 -7561
rect 1033 -7633 1079 -7595
rect 1033 -7667 1039 -7633
rect 1073 -7667 1079 -7633
rect 1033 -7705 1079 -7667
rect 1033 -7739 1039 -7705
rect 1073 -7739 1079 -7705
rect 1033 -7777 1079 -7739
rect 1033 -7811 1039 -7777
rect 1073 -7811 1079 -7777
rect 1033 -7849 1079 -7811
rect 1033 -7883 1039 -7849
rect 1073 -7883 1079 -7849
rect 1033 -7921 1079 -7883
rect 1033 -7955 1039 -7921
rect 1073 -7955 1079 -7921
rect 1033 -7993 1079 -7955
rect 1033 -8027 1039 -7993
rect 1073 -8027 1079 -7993
rect 1033 -8065 1079 -8027
rect 1033 -8099 1039 -8065
rect 1073 -8099 1079 -8065
rect 1033 -8137 1079 -8099
rect 1033 -8171 1039 -8137
rect 1073 -8171 1079 -8137
rect 1033 -8209 1079 -8171
rect 1033 -8243 1039 -8209
rect 1073 -8243 1079 -8209
rect 1033 -8281 1079 -8243
rect 1033 -8315 1039 -8281
rect 1073 -8315 1079 -8281
rect 1033 -8353 1079 -8315
rect 1033 -8387 1039 -8353
rect 1073 -8387 1079 -8353
rect 1033 -8425 1079 -8387
rect 1033 -8459 1039 -8425
rect 1073 -8459 1079 -8425
rect 1033 -8497 1079 -8459
rect 1033 -8531 1039 -8497
rect 1073 -8531 1079 -8497
rect 1033 -8569 1079 -8531
rect 1033 -8603 1039 -8569
rect 1073 -8603 1079 -8569
rect 1033 -8641 1079 -8603
rect 1033 -8675 1039 -8641
rect 1073 -8675 1079 -8641
rect 1033 -8713 1079 -8675
rect 1033 -8747 1039 -8713
rect 1073 -8747 1079 -8713
rect 1033 -8785 1079 -8747
rect 1033 -8819 1039 -8785
rect 1073 -8819 1079 -8785
rect 1033 -8857 1079 -8819
rect 1033 -8891 1039 -8857
rect 1073 -8891 1079 -8857
rect 1033 -8929 1079 -8891
rect 1033 -8963 1039 -8929
rect 1073 -8963 1079 -8929
rect 1033 -9001 1079 -8963
rect 1033 -9035 1039 -9001
rect 1073 -9035 1079 -9001
rect 1033 -9073 1079 -9035
rect 1033 -9107 1039 -9073
rect 1073 -9107 1079 -9073
rect 1033 -9145 1079 -9107
rect 1033 -9179 1039 -9145
rect 1073 -9179 1079 -9145
rect 1033 -9217 1079 -9179
rect 1033 -9251 1039 -9217
rect 1073 -9251 1079 -9217
rect 1033 -9289 1079 -9251
rect 1033 -9323 1039 -9289
rect 1073 -9323 1079 -9289
rect 1033 -9361 1079 -9323
rect 1033 -9395 1039 -9361
rect 1073 -9395 1079 -9361
rect 1033 -9433 1079 -9395
rect 1033 -9467 1039 -9433
rect 1073 -9467 1079 -9433
rect 1033 -9506 1079 -9467
rect 1033 -9540 1039 -9506
rect 1073 -9540 1079 -9506
rect 1033 -9579 1079 -9540
tri 2623 -9572 2665 -9530 se
rect 2665 -9572 2934 -9530
tri 2934 -9572 2976 -9530 sw
tri 2619 -9576 2623 -9572 se
rect 2623 -9576 2976 -9572
rect 1033 -9613 1039 -9579
rect 1073 -9613 1079 -9579
rect 1033 -9652 1079 -9613
rect 1033 -9686 1039 -9652
rect 1073 -9686 1079 -9652
rect 1033 -9725 1079 -9686
rect 1033 -9759 1039 -9725
rect 1073 -9759 1079 -9725
rect 1033 -9798 1079 -9759
rect 1033 -9832 1039 -9798
rect 1073 -9832 1079 -9798
rect 1033 -9871 1079 -9832
rect 1033 -9905 1039 -9871
rect 1073 -9905 1079 -9871
rect 1033 -9944 1079 -9905
rect 1033 -9978 1039 -9944
rect 1073 -9978 1079 -9944
rect 1033 -10017 1079 -9978
rect 1033 -10051 1039 -10017
rect 1073 -10051 1079 -10017
rect 1033 -10090 1079 -10051
rect 1033 -10124 1039 -10090
rect 1073 -10124 1079 -10090
rect 1033 -10163 1079 -10124
rect 1033 -10197 1039 -10163
rect 1073 -10197 1079 -10163
tri 2612 -9583 2619 -9576 se
rect 2619 -9583 2664 -9576
rect 2612 -9624 2664 -9583
tri 2664 -9597 2685 -9576 nw
tri 2914 -9592 2930 -9576 ne
rect 2612 -9625 2624 -9624
rect 2658 -9625 2664 -9624
rect 2612 -9689 2664 -9677
rect 2612 -9772 2664 -9741
rect 2612 -9806 2624 -9772
rect 2658 -9806 2664 -9772
rect 2612 -9846 2664 -9806
rect 2612 -9880 2624 -9846
rect 2658 -9880 2664 -9846
rect 2612 -9920 2664 -9880
rect 2612 -9954 2624 -9920
rect 2658 -9954 2664 -9920
rect 2612 -9994 2664 -9954
rect 2612 -10028 2624 -9994
rect 2658 -10028 2664 -9994
rect 2612 -10068 2664 -10028
rect 2612 -10102 2624 -10068
rect 2658 -10102 2664 -10068
rect 2612 -10142 2664 -10102
rect 2612 -10176 2624 -10142
rect 2658 -10176 2664 -10142
rect 2612 -10188 2664 -10176
rect 2771 -9624 2823 -9612
rect 2771 -9658 2780 -9624
rect 2814 -9658 2823 -9624
rect 2771 -9698 2823 -9658
rect 2771 -9732 2780 -9698
rect 2814 -9732 2823 -9698
rect 2771 -9749 2823 -9732
rect 2771 -9806 2780 -9801
rect 2814 -9806 2823 -9801
rect 2771 -9813 2823 -9806
rect 2771 -9880 2780 -9865
rect 2814 -9880 2823 -9865
rect 2771 -9920 2823 -9880
rect 2771 -9954 2780 -9920
rect 2814 -9954 2823 -9920
rect 2771 -9994 2823 -9954
rect 2771 -10028 2780 -9994
rect 2814 -10028 2823 -9994
rect 2771 -10068 2823 -10028
rect 2771 -10102 2780 -10068
rect 2814 -10102 2823 -10068
rect 2771 -10142 2823 -10102
rect 2771 -10176 2780 -10142
rect 2814 -10176 2823 -10142
rect 2771 -10188 2823 -10176
rect 2930 -9624 2976 -9576
rect 2930 -9658 2936 -9624
rect 2970 -9658 2976 -9624
rect 2930 -9698 2976 -9658
rect 2930 -9732 2936 -9698
rect 2970 -9732 2976 -9698
rect 2930 -9772 2976 -9732
rect 2930 -9806 2936 -9772
rect 2970 -9806 2976 -9772
rect 2930 -9846 2976 -9806
rect 2930 -9880 2936 -9846
rect 2970 -9880 2976 -9846
rect 2930 -9920 2976 -9880
rect 2930 -9954 2936 -9920
rect 2970 -9954 2976 -9920
rect 2930 -9994 2976 -9954
rect 2930 -10028 2936 -9994
rect 2970 -10028 2976 -9994
rect 2930 -10068 2976 -10028
rect 2930 -10102 2936 -10068
rect 2970 -10102 2976 -10068
rect 2930 -10142 2976 -10102
rect 2930 -10176 2936 -10142
rect 2970 -10176 2976 -10142
rect 2930 -10188 2976 -10176
rect 1033 -10236 1079 -10197
rect 1033 -10270 1039 -10236
rect 1073 -10270 1079 -10236
rect 1033 -10309 1079 -10270
rect 2641 -10275 2647 -10223
rect 2699 -10232 2711 -10223
rect 2763 -10226 2769 -10223
rect 2763 -10232 2925 -10226
rect 2763 -10266 2780 -10232
rect 2814 -10266 2879 -10232
rect 2913 -10266 2925 -10232
rect 2699 -10275 2711 -10266
rect 2763 -10272 2925 -10266
rect 2763 -10275 2769 -10272
rect 1033 -10343 1039 -10309
rect 1073 -10343 1079 -10309
rect 1033 -10382 1079 -10343
rect 1033 -10416 1039 -10382
rect 1073 -10416 1079 -10382
rect 1033 -10455 1079 -10416
rect 1033 -10489 1039 -10455
rect 1073 -10489 1079 -10455
rect 1033 -10528 1079 -10489
rect 1033 -10562 1039 -10528
rect 1073 -10562 1079 -10528
rect 1033 -10601 1079 -10562
rect 1033 -10635 1039 -10601
rect 1073 -10635 1079 -10601
rect 1033 -10674 1079 -10635
rect 1033 -10708 1039 -10674
rect 1073 -10708 1079 -10674
rect 1033 -10747 1079 -10708
rect 1033 -10781 1039 -10747
rect 1073 -10781 1079 -10747
rect 1033 -10820 1079 -10781
rect 1033 -10854 1039 -10820
rect 1073 -10854 1079 -10820
rect 1033 -10893 1079 -10854
rect 1033 -10927 1039 -10893
rect 1073 -10927 1079 -10893
rect 1033 -10966 1079 -10927
rect 1033 -11000 1039 -10966
rect 1073 -11000 1079 -10966
rect 2389 -10868 3345 -10862
rect 2441 -10914 3345 -10868
rect 2389 -10932 2441 -10920
rect 2389 -10990 2441 -10984
rect 2473 -10951 3256 -10945
rect 401 -11073 407 -11039
rect 441 -11073 447 -11039
rect 1033 -11039 1079 -11000
tri 447 -11073 449 -11071 sw
tri 1031 -11073 1033 -11071 se
rect 1033 -11073 1039 -11039
rect 1073 -11073 1079 -11039
rect 2525 -10997 3256 -10951
rect 2473 -11015 2525 -11003
rect 2473 -11073 2525 -11067
rect 401 -11105 449 -11073
tri 449 -11105 481 -11073 sw
tri 999 -11105 1031 -11073 se
rect 1031 -11105 1079 -11073
rect 401 -11111 1079 -11105
rect 401 -11145 479 -11111
rect 513 -11145 559 -11111
rect 593 -11145 639 -11111
rect 673 -11145 719 -11111
rect 753 -11145 799 -11111
rect 833 -11145 879 -11111
rect 913 -11145 959 -11111
rect 993 -11145 1079 -11111
rect 401 -11151 1079 -11145
rect 3204 -12013 3256 -10997
rect 3293 -11930 3345 -10914
rect 18751 -11604 18803 -236
rect 18751 -11638 18762 -11604
rect 18796 -11638 18803 -11604
rect 18751 -11692 18803 -11638
rect 18751 -11726 18762 -11692
rect 18796 -11726 18803 -11692
rect 18751 -11740 18803 -11726
rect 3293 -11936 3701 -11930
rect 3293 -11982 3649 -11936
rect 3649 -12000 3701 -11988
rect 3204 -12019 3610 -12013
rect 3204 -12065 3558 -12019
rect 3649 -12058 3701 -12052
rect 3558 -12083 3610 -12071
rect 3558 -12141 3610 -12135
rect 18862 -12797 18914 -158
rect 18947 -62 18993 -22
rect 18947 -96 18953 -62
rect 18987 -96 18993 -62
rect 18947 -136 18993 -96
rect 18947 -170 18953 -136
rect 18987 -170 18993 -136
rect 18947 -210 18993 -170
rect 18947 -244 18953 -210
rect 18987 -244 18993 -210
rect 18947 -284 18993 -244
rect 18947 -318 18953 -284
rect 18987 -318 18993 -284
rect 18947 -358 18993 -318
rect 18947 -392 18953 -358
rect 18987 -392 18993 -358
rect 18947 -432 18993 -392
rect 18947 -466 18953 -432
rect 18987 -466 18993 -432
rect 18947 -506 18993 -466
rect 18947 -540 18953 -506
rect 18987 -540 18993 -506
rect 18947 -580 18993 -540
rect 18947 -614 18953 -580
rect 18987 -614 18993 -580
rect 18947 -653 18993 -614
rect 18947 -687 18953 -653
rect 18987 -687 18993 -653
rect 18947 -726 18993 -687
rect 18947 -760 18953 -726
rect 18987 -760 18993 -726
rect 18947 -799 18993 -760
rect 18947 -833 18953 -799
rect 18987 -833 18993 -799
rect 18947 -872 18993 -833
rect 18947 -906 18953 -872
rect 18987 -906 18993 -872
rect 18947 -945 18993 -906
rect 18947 -979 18953 -945
rect 18987 -979 18993 -945
rect 18947 -1018 18993 -979
rect 18947 -1052 18953 -1018
rect 18987 -1052 18993 -1018
rect 18947 -1091 18993 -1052
rect 18947 -1125 18953 -1091
rect 18987 -1125 18993 -1091
rect 18947 -1164 18993 -1125
rect 18947 -1198 18953 -1164
rect 18987 -1198 18993 -1164
rect 18947 -1237 18993 -1198
rect 18947 -1271 18953 -1237
rect 18987 -1271 18993 -1237
rect 18947 -1310 18993 -1271
rect 18947 -1344 18953 -1310
rect 18987 -1344 18993 -1310
rect 18947 -1383 18993 -1344
rect 18947 -1417 18953 -1383
rect 18987 -1417 18993 -1383
rect 18947 -1455 18993 -1417
rect 19155 154 19161 206
rect 19213 154 19227 206
rect 19279 154 19354 206
rect 19155 -12733 19354 154
rect 22597 -12733 22785 855
rect 18862 -12831 18874 -12797
rect 18908 -12831 18914 -12797
rect 18862 -12940 18914 -12831
rect 18862 -12974 18874 -12940
rect 18908 -12974 18914 -12940
rect 18862 -12986 18914 -12974
tri 3882 -14680 3925 -14637 se
rect 3925 -14680 3980 -14637
rect 3202 -14686 3254 -14680
tri 3824 -14738 3882 -14680 se
rect 3882 -14683 3980 -14680
rect 3882 -14738 3925 -14683
tri 3925 -14738 3980 -14683 nw
rect 3202 -14748 3254 -14738
tri 3814 -14748 3824 -14738 se
rect 3824 -14748 3915 -14738
tri 3915 -14748 3925 -14738 nw
rect 3202 -14750 3855 -14748
rect 3254 -14802 3855 -14750
rect 3202 -14808 3855 -14802
tri 3855 -14808 3915 -14748 nw
rect 3068 -17011 3324 -17005
rect 3068 -17045 3080 -17011
rect 3114 -17045 3179 -17011
rect 3213 -17045 3278 -17011
rect 3312 -17045 3324 -17011
rect 3068 -17051 3324 -17045
rect 3017 -17422 3140 -17416
rect 3017 -17428 3088 -17422
rect 3017 -17462 3023 -17428
rect 3057 -17462 3088 -17428
rect 3017 -17474 3088 -17462
rect 3017 -17488 3140 -17474
rect 3017 -17501 3088 -17488
rect 3017 -17535 3023 -17501
rect 3057 -17535 3088 -17501
rect 3017 -17540 3088 -17535
rect 3017 -17546 3140 -17540
rect 3173 -17425 3225 -17419
rect 3173 -17489 3225 -17477
rect 3017 -17575 3082 -17546
tri 3082 -17575 3111 -17546 nw
rect 3017 -17609 3023 -17575
rect 3057 -17576 3081 -17575
tri 3081 -17576 3082 -17575 nw
rect 3173 -17576 3225 -17541
rect 3057 -17609 3063 -17576
tri 3063 -17594 3081 -17576 nw
rect 3017 -17649 3063 -17609
rect 3017 -17683 3023 -17649
rect 3057 -17683 3063 -17649
rect 3017 -17720 3063 -17683
rect 3173 -17610 3179 -17576
rect 3213 -17610 3225 -17576
rect 3173 -17649 3225 -17610
rect 3173 -17683 3179 -17649
rect 3213 -17683 3225 -17649
rect 3173 -17695 3225 -17683
rect 3329 -17428 3375 -17416
rect 3329 -17462 3335 -17428
rect 3369 -17462 3375 -17428
rect 3329 -17501 3375 -17462
rect 3329 -17535 3335 -17501
rect 3369 -17535 3375 -17501
rect 3329 -17575 3375 -17535
rect 3329 -17609 3335 -17575
rect 3369 -17609 3375 -17575
rect 3329 -17649 3375 -17609
rect 3329 -17683 3335 -17649
rect 3369 -17683 3375 -17649
tri 3063 -17720 3086 -17697 sw
rect 3017 -17734 3086 -17720
tri 3086 -17734 3100 -17720 sw
tri 3315 -17734 3329 -17720 se
rect 3329 -17734 3375 -17683
rect 3017 -17740 3375 -17734
rect 3017 -17752 3363 -17740
tri 3363 -17752 3375 -17740 nw
tri 2951 -17818 3017 -17752 se
rect 3017 -17780 3335 -17752
tri 3335 -17780 3363 -17752 nw
tri 3017 -17818 3055 -17780 nw
tri 2942 -17827 2951 -17818 se
rect 2951 -17827 3008 -17818
tri 3008 -17827 3017 -17818 nw
rect 2625 -17833 2962 -17827
rect 2625 -17867 2637 -17833
rect 2671 -17867 2737 -17833
rect 2771 -17867 2836 -17833
rect 2870 -17867 2962 -17833
rect 2625 -17873 2962 -17867
tri 2962 -17873 3008 -17827 nw
rect 2574 -18114 2932 -18102
rect 2574 -18148 2580 -18114
rect 2614 -18148 2892 -18114
rect 2926 -18148 2932 -18114
rect 2574 -18194 2620 -18148
tri 2620 -18180 2652 -18148 nw
tri 2854 -18180 2886 -18148 ne
rect 2574 -18228 2580 -18194
rect 2614 -18228 2620 -18194
rect 2886 -18187 2932 -18148
rect 2574 -18274 2620 -18228
rect 2574 -18308 2580 -18274
rect 2614 -18308 2620 -18274
rect 2574 -18354 2620 -18308
rect 2574 -18388 2580 -18354
rect 2614 -18388 2620 -18354
rect 2574 -18435 2620 -18388
rect 2574 -18469 2580 -18435
rect 2614 -18469 2620 -18435
rect 2574 -18516 2620 -18469
rect 2574 -18550 2580 -18516
rect 2614 -18550 2620 -18516
rect 2574 -18597 2620 -18550
rect 2574 -18631 2580 -18597
rect 2614 -18631 2620 -18597
rect 2574 -18672 2620 -18631
rect 2492 -18724 2498 -18672
rect 2550 -18724 2562 -18672
rect 2614 -18724 2620 -18672
rect 2730 -18214 2776 -18202
rect 2730 -18248 2736 -18214
rect 2770 -18248 2776 -18214
rect 2730 -18287 2776 -18248
rect 2730 -18321 2736 -18287
rect 2770 -18321 2776 -18287
rect 2730 -18360 2776 -18321
rect 2730 -18394 2736 -18360
rect 2770 -18394 2776 -18360
rect 2730 -18433 2776 -18394
rect 2730 -18467 2736 -18433
rect 2770 -18467 2776 -18433
rect 2730 -18506 2776 -18467
rect 2730 -18540 2736 -18506
rect 2770 -18540 2776 -18506
rect 2730 -18579 2776 -18540
rect 2730 -18613 2736 -18579
rect 2770 -18613 2776 -18579
rect 2730 -18652 2776 -18613
rect 2730 -18686 2736 -18652
rect 2770 -18686 2776 -18652
rect 2730 -18725 2776 -18686
rect 2730 -18759 2736 -18725
rect 2770 -18759 2776 -18725
rect 2730 -18788 2776 -18759
rect 2561 -18794 2776 -18788
rect 2613 -18799 2776 -18794
rect 2613 -18833 2736 -18799
rect 2770 -18833 2776 -18799
rect 2886 -18221 2892 -18187
rect 2926 -18221 2932 -18187
rect 2886 -18260 2932 -18221
rect 2886 -18294 2892 -18260
rect 2926 -18294 2932 -18260
rect 2886 -18333 2932 -18294
rect 2886 -18367 2892 -18333
rect 2926 -18367 2932 -18333
rect 2886 -18406 2932 -18367
rect 2886 -18440 2892 -18406
rect 2926 -18440 2932 -18406
rect 2886 -18479 2932 -18440
rect 2886 -18513 2892 -18479
rect 2926 -18513 2932 -18479
rect 2886 -18552 2932 -18513
rect 2886 -18586 2892 -18552
rect 2926 -18586 2932 -18552
rect 2886 -18625 2932 -18586
rect 2886 -18659 2892 -18625
rect 2926 -18659 2932 -18625
rect 2886 -18699 2932 -18659
rect 2886 -18733 2892 -18699
rect 2926 -18733 2932 -18699
rect 2886 -18773 2932 -18733
rect 2886 -18807 2892 -18773
rect 2926 -18807 2932 -18773
rect 2886 -18819 2932 -18807
rect 2613 -18846 2776 -18833
rect 2561 -18858 2776 -18846
rect 2613 -18873 2776 -18858
rect 2613 -18907 2736 -18873
rect 2770 -18907 2776 -18873
rect 2613 -18910 2776 -18907
rect 2561 -18919 2776 -18910
<< rmetal1 >>
rect 18164 4371 18172 4417
rect 19009 3836 19036 3888
<< via1 >>
rect 454 4942 506 4994
rect 454 4888 467 4912
rect 467 4888 501 4912
rect 501 4888 506 4912
rect 454 4860 506 4888
rect 575 4865 627 4917
rect 639 4865 691 4917
rect 454 4813 467 4830
rect 467 4813 501 4830
rect 501 4813 506 4830
rect 454 4778 506 4813
rect 454 4738 467 4748
rect 467 4738 501 4748
rect 501 4738 506 4748
rect 454 4697 506 4738
rect 454 4696 467 4697
rect 467 4696 501 4697
rect 501 4696 506 4697
rect 454 4663 467 4666
rect 467 4663 501 4666
rect 501 4663 506 4666
rect 454 4622 506 4663
rect 454 4614 467 4622
rect 467 4614 501 4622
rect 501 4614 506 4622
rect 952 4772 1004 4824
rect 1044 4772 1096 4824
rect 1135 4772 1187 4824
rect 1210 4779 1262 4831
rect 1279 4779 1331 4831
rect 1348 4779 1400 4831
rect 1417 4779 1469 4831
rect 1486 4779 1538 4831
rect 1554 4779 1606 4831
rect 1622 4779 1674 4831
rect 1690 4823 1742 4831
rect 1758 4823 1810 4831
rect 1690 4789 1727 4823
rect 1727 4789 1742 4823
rect 1758 4789 1761 4823
rect 1761 4789 1810 4823
rect 1690 4779 1742 4789
rect 1758 4779 1810 4789
rect 1826 4779 1878 4831
rect 1894 4779 1946 4831
rect 1962 4823 2014 4831
rect 1962 4789 1983 4823
rect 1983 4789 2014 4823
rect 1962 4779 2014 4789
rect 952 4692 1004 4744
rect 1044 4692 1096 4744
rect 1135 4692 1187 4744
rect 1210 4701 1262 4753
rect 1279 4701 1331 4753
rect 1348 4701 1400 4753
rect 1417 4701 1469 4753
rect 1486 4701 1538 4753
rect 1554 4701 1606 4753
rect 1622 4701 1674 4753
rect 1690 4751 1742 4753
rect 1758 4751 1810 4753
rect 1690 4717 1727 4751
rect 1727 4717 1742 4751
rect 1758 4717 1761 4751
rect 1761 4717 1810 4751
rect 1690 4701 1742 4717
rect 1758 4701 1810 4717
rect 1826 4701 1878 4753
rect 1894 4701 1946 4753
rect 1962 4751 2014 4753
rect 1962 4717 1983 4751
rect 1983 4717 2014 4751
rect 1962 4701 2014 4717
rect 952 4652 1004 4664
rect 1044 4652 1096 4664
rect 1135 4652 1187 4664
rect 952 4618 962 4652
rect 962 4618 1004 4652
rect 1044 4618 1084 4652
rect 1084 4618 1096 4652
rect 1135 4618 1162 4652
rect 1162 4618 1187 4652
rect 952 4612 1004 4618
rect 1044 4612 1096 4618
rect 1135 4612 1187 4618
rect 2045 4661 2097 4667
rect 2045 4627 2051 4661
rect 2051 4627 2085 4661
rect 2085 4627 2097 4661
rect 2045 4615 2097 4627
rect 2118 4661 2170 4667
rect 2118 4627 2130 4661
rect 2130 4627 2164 4661
rect 2164 4627 2170 4661
rect 2118 4615 2170 4627
rect 2486 4789 2495 4819
rect 2495 4789 2529 4819
rect 2529 4789 2538 4819
rect 2486 4767 2538 4789
rect 2486 4751 2538 4755
rect 2486 4717 2495 4751
rect 2495 4717 2529 4751
rect 2529 4717 2538 4751
rect 2486 4703 2538 4717
rect 2336 4661 2388 4667
rect 2336 4627 2342 4661
rect 2342 4627 2376 4661
rect 2376 4627 2388 4661
rect 2336 4615 2388 4627
rect 2413 4661 2465 4667
rect 2413 4627 2421 4661
rect 2421 4627 2455 4661
rect 2455 4627 2465 4661
rect 2413 4615 2465 4627
rect 2490 4661 2542 4667
rect 2490 4627 2500 4661
rect 2500 4627 2534 4661
rect 2534 4627 2542 4661
rect 2490 4615 2542 4627
rect 2567 4661 2619 4667
rect 2567 4627 2578 4661
rect 2578 4627 2612 4661
rect 2612 4627 2619 4661
rect 2567 4615 2619 4627
rect 2644 4661 2696 4667
rect 2644 4627 2656 4661
rect 2656 4627 2690 4661
rect 2690 4627 2696 4661
rect 2644 4615 2696 4627
rect 2998 4789 3007 4819
rect 3007 4789 3041 4819
rect 3041 4789 3050 4819
rect 2998 4767 3050 4789
rect 2998 4751 3050 4755
rect 2998 4717 3007 4751
rect 3007 4717 3041 4751
rect 3041 4717 3050 4751
rect 2998 4703 3050 4717
rect 3510 4789 3519 4819
rect 3519 4789 3553 4819
rect 3553 4789 3562 4819
rect 3510 4767 3562 4789
rect 3510 4751 3562 4755
rect 3510 4717 3519 4751
rect 3519 4717 3553 4751
rect 3553 4717 3562 4751
rect 2831 4661 2883 4667
rect 2831 4627 2837 4661
rect 2837 4627 2871 4661
rect 2871 4627 2883 4661
rect 2831 4615 2883 4627
rect 2898 4661 2950 4667
rect 2965 4661 3017 4667
rect 3031 4661 3083 4667
rect 3097 4661 3149 4667
rect 2898 4627 2922 4661
rect 2922 4627 2950 4661
rect 2965 4627 3007 4661
rect 3007 4627 3017 4661
rect 3031 4627 3041 4661
rect 3041 4627 3083 4661
rect 3097 4627 3125 4661
rect 3125 4627 3149 4661
rect 2898 4615 2950 4627
rect 2965 4615 3017 4627
rect 3031 4615 3083 4627
rect 3097 4615 3149 4627
rect 3163 4661 3215 4667
rect 3163 4627 3175 4661
rect 3175 4627 3209 4661
rect 3209 4627 3215 4661
rect 3163 4615 3215 4627
rect 3510 4703 3562 4717
rect 3570 4661 3622 4667
rect 3570 4627 3576 4661
rect 3576 4627 3610 4661
rect 3610 4627 3622 4661
rect 3570 4615 3622 4627
rect 3679 4661 3731 4667
rect 3679 4627 3691 4661
rect 3691 4627 3725 4661
rect 3725 4627 3731 4661
rect 3679 4615 3731 4627
rect 454 4547 506 4584
rect 454 4532 467 4547
rect 467 4532 501 4547
rect 501 4532 506 4547
rect 793 4529 845 4581
rect 857 4529 909 4581
rect 4022 4789 4031 4819
rect 4031 4789 4065 4819
rect 4065 4789 4074 4819
rect 4022 4767 4074 4789
rect 4022 4751 4074 4755
rect 4022 4717 4031 4751
rect 4031 4717 4065 4751
rect 4065 4717 4074 4751
rect 4022 4703 4074 4717
rect 3852 4661 3904 4667
rect 3852 4627 3858 4661
rect 3858 4627 3892 4661
rect 3892 4627 3904 4661
rect 3852 4615 3904 4627
rect 3921 4661 3973 4667
rect 3990 4661 4042 4667
rect 4058 4661 4110 4667
rect 4126 4661 4178 4667
rect 3921 4627 3945 4661
rect 3945 4627 3973 4661
rect 3990 4627 4032 4661
rect 4032 4627 4042 4661
rect 4058 4627 4066 4661
rect 4066 4627 4110 4661
rect 4126 4627 4153 4661
rect 4153 4627 4178 4661
rect 3921 4615 3973 4627
rect 3990 4615 4042 4627
rect 4058 4615 4110 4627
rect 4126 4615 4178 4627
rect 4194 4661 4246 4667
rect 4194 4627 4206 4661
rect 4206 4627 4240 4661
rect 4240 4627 4246 4661
rect 4194 4615 4246 4627
rect 4534 4789 4543 4819
rect 4543 4789 4577 4819
rect 4577 4789 4586 4819
rect 4534 4767 4586 4789
rect 4534 4751 4586 4755
rect 4534 4717 4543 4751
rect 4543 4717 4577 4751
rect 4577 4717 4586 4751
rect 4534 4703 4586 4717
rect 4365 4661 4417 4667
rect 4365 4627 4371 4661
rect 4371 4627 4405 4661
rect 4405 4627 4417 4661
rect 4365 4615 4417 4627
rect 4433 4661 4485 4667
rect 4501 4661 4553 4667
rect 4569 4661 4621 4667
rect 4636 4661 4688 4667
rect 4433 4627 4457 4661
rect 4457 4627 4485 4661
rect 4501 4627 4543 4661
rect 4543 4627 4553 4661
rect 4569 4627 4577 4661
rect 4577 4627 4621 4661
rect 4636 4627 4663 4661
rect 4663 4627 4688 4661
rect 4433 4615 4485 4627
rect 4501 4615 4553 4627
rect 4569 4615 4621 4627
rect 4636 4615 4688 4627
rect 4703 4661 4755 4667
rect 4703 4627 4715 4661
rect 4715 4627 4749 4661
rect 4749 4627 4755 4661
rect 4703 4615 4755 4627
rect 5046 4789 5055 4819
rect 5055 4789 5089 4819
rect 5089 4789 5098 4819
rect 5046 4767 5098 4789
rect 5046 4751 5098 4755
rect 5046 4717 5055 4751
rect 5055 4717 5089 4751
rect 5089 4717 5098 4751
rect 5046 4703 5098 4717
rect 5558 4789 5567 4819
rect 5567 4789 5601 4819
rect 5601 4789 5610 4819
rect 5558 4767 5610 4789
rect 5558 4751 5610 4755
rect 5558 4717 5567 4751
rect 5567 4717 5601 4751
rect 5601 4717 5610 4751
rect 5558 4703 5610 4717
rect 6070 4789 6079 4819
rect 6079 4789 6113 4819
rect 6113 4789 6122 4819
rect 6070 4767 6122 4789
rect 6070 4751 6122 4755
rect 6070 4717 6079 4751
rect 6079 4717 6113 4751
rect 6113 4717 6122 4751
rect 6070 4703 6122 4717
rect 6582 4789 6591 4819
rect 6591 4789 6625 4819
rect 6625 4789 6634 4819
rect 6582 4767 6634 4789
rect 6582 4751 6634 4755
rect 6582 4717 6591 4751
rect 6591 4717 6625 4751
rect 6625 4717 6634 4751
rect 6582 4703 6634 4717
rect 6964 4808 7016 4860
rect 7029 4808 7081 4860
rect 7094 4808 7146 4860
rect 7158 4808 7210 4860
rect 7222 4808 7274 4860
rect 7286 4808 7338 4860
rect 7350 4808 7402 4860
rect 7414 4808 7466 4860
rect 7478 4808 7530 4860
rect 7712 4823 7764 4825
rect 7712 4789 7737 4823
rect 7737 4789 7764 4823
rect 7712 4773 7764 4789
rect 7820 4812 7838 4825
rect 7838 4812 7872 4825
rect 7820 4773 7872 4812
rect 6964 4698 7016 4750
rect 7029 4698 7081 4750
rect 7094 4698 7146 4750
rect 7158 4698 7210 4750
rect 7222 4698 7274 4750
rect 7286 4698 7338 4750
rect 7350 4698 7402 4750
rect 7414 4698 7466 4750
rect 7478 4698 7530 4750
rect 7712 4717 7737 4749
rect 7737 4717 7764 4749
rect 7712 4697 7764 4717
rect 7820 4738 7838 4749
rect 7838 4738 7872 4749
rect 7820 4698 7872 4738
rect 7820 4697 7838 4698
rect 7838 4697 7872 4698
rect 4875 4661 4927 4667
rect 4875 4627 4881 4661
rect 4881 4627 4915 4661
rect 4915 4627 4927 4661
rect 4875 4615 4927 4627
rect 4941 4661 4993 4667
rect 4941 4627 4955 4661
rect 4955 4627 4989 4661
rect 4989 4627 4993 4661
rect 4941 4615 4993 4627
rect 5007 4661 5059 4667
rect 5073 4661 5125 4667
rect 5139 4661 5191 4667
rect 5205 4661 5257 4667
rect 5271 4661 5323 4667
rect 5337 4661 5389 4667
rect 5403 4661 5455 4667
rect 5469 4661 5521 4667
rect 5007 4627 5029 4661
rect 5029 4627 5059 4661
rect 5073 4627 5102 4661
rect 5102 4627 5125 4661
rect 5139 4627 5175 4661
rect 5175 4627 5191 4661
rect 5205 4627 5209 4661
rect 5209 4627 5248 4661
rect 5248 4627 5257 4661
rect 5271 4627 5282 4661
rect 5282 4627 5321 4661
rect 5321 4627 5323 4661
rect 5337 4627 5355 4661
rect 5355 4627 5389 4661
rect 5403 4627 5428 4661
rect 5428 4627 5455 4661
rect 5469 4627 5501 4661
rect 5501 4627 5521 4661
rect 5007 4615 5059 4627
rect 5073 4615 5125 4627
rect 5139 4615 5191 4627
rect 5205 4615 5257 4627
rect 5271 4615 5323 4627
rect 5337 4615 5389 4627
rect 5403 4615 5455 4627
rect 5469 4615 5521 4627
rect 5535 4661 5587 4667
rect 5535 4627 5540 4661
rect 5540 4627 5574 4661
rect 5574 4627 5587 4661
rect 5535 4615 5587 4627
rect 5601 4661 5653 4667
rect 5601 4627 5613 4661
rect 5613 4627 5647 4661
rect 5647 4627 5653 4661
rect 5601 4615 5653 4627
rect 5667 4661 5719 4667
rect 5732 4661 5784 4667
rect 5797 4661 5849 4667
rect 5862 4661 5914 4667
rect 5927 4661 5979 4667
rect 5992 4661 6044 4667
rect 6057 4661 6109 4667
rect 5667 4627 5686 4661
rect 5686 4627 5719 4661
rect 5732 4627 5759 4661
rect 5759 4627 5784 4661
rect 5797 4627 5832 4661
rect 5832 4627 5849 4661
rect 5862 4627 5866 4661
rect 5866 4627 5905 4661
rect 5905 4627 5914 4661
rect 5927 4627 5939 4661
rect 5939 4627 5978 4661
rect 5978 4627 5979 4661
rect 5992 4627 6012 4661
rect 6012 4627 6044 4661
rect 6057 4627 6085 4661
rect 6085 4627 6109 4661
rect 5667 4615 5719 4627
rect 5732 4615 5784 4627
rect 5797 4615 5849 4627
rect 5862 4615 5914 4627
rect 5927 4615 5979 4627
rect 5992 4615 6044 4627
rect 6057 4615 6109 4627
rect 6122 4661 6174 4667
rect 6122 4627 6124 4661
rect 6124 4627 6158 4661
rect 6158 4627 6174 4661
rect 6122 4615 6174 4627
rect 6187 4661 6239 4667
rect 6187 4627 6197 4661
rect 6197 4627 6231 4661
rect 6231 4627 6239 4661
rect 6187 4615 6239 4627
rect 6252 4661 6304 4667
rect 6252 4627 6270 4661
rect 6270 4627 6304 4661
rect 6252 4615 6304 4627
rect 6317 4661 6369 4667
rect 6382 4661 6434 4667
rect 6447 4661 6499 4667
rect 6512 4661 6564 4667
rect 6317 4627 6343 4661
rect 6343 4627 6369 4661
rect 6382 4627 6416 4661
rect 6416 4627 6434 4661
rect 6447 4627 6450 4661
rect 6450 4627 6489 4661
rect 6489 4627 6499 4661
rect 6512 4627 6523 4661
rect 6523 4627 6564 4661
rect 6317 4615 6369 4627
rect 6382 4615 6434 4627
rect 6447 4615 6499 4627
rect 6512 4615 6564 4627
rect 6577 4615 6629 4667
rect 6642 4615 6694 4667
rect 6707 4615 6759 4667
rect 6772 4615 6824 4667
rect 8482 4926 8534 4978
rect 8548 4926 8600 4978
rect 8614 4926 8666 4978
rect 8680 4926 8732 4978
rect 8746 4926 8798 4978
rect 8811 4926 8863 4978
rect 8876 4926 8928 4978
rect 8941 4926 8993 4978
rect 9006 4926 9058 4978
rect 9071 4926 9123 4978
rect 9136 4926 9188 4978
rect 9201 4926 9253 4978
rect 9266 4926 9318 4978
rect 9331 4926 9383 4978
rect 9396 4926 9448 4978
rect 9461 4926 9513 4978
rect 9526 4926 9578 4978
rect 9591 4926 9643 4978
rect 9656 4926 9708 4978
rect 9721 4926 9773 4978
rect 9786 4926 9838 4978
rect 9851 4926 9903 4978
rect 9916 4926 9968 4978
rect 9981 4926 10033 4978
rect 10046 4926 10098 4978
rect 10111 4926 10163 4978
rect 10176 4926 10228 4978
rect 10241 4926 10293 4978
rect 10306 4926 10358 4978
rect 10371 4926 10423 4978
rect 10436 4926 10488 4978
rect 10501 4926 10553 4978
rect 10566 4926 10618 4978
rect 10631 4926 10683 4978
rect 10696 4926 10748 4978
rect 10761 4926 10813 4978
rect 10826 4926 10878 4978
rect 10891 4926 10943 4978
rect 10956 4926 11008 4978
rect 11021 4926 11073 4978
rect 11086 4926 11138 4978
rect 11151 4926 11203 4978
rect 11216 4926 11268 4978
rect 11281 4926 11333 4978
rect 11346 4926 11398 4978
rect 11411 4926 11463 4978
rect 11515 4918 11567 4970
rect 11580 4918 11632 4970
rect 11644 4918 11696 4970
rect 19755 4918 19807 4970
rect 19819 4918 19871 4970
rect 19883 4918 19935 4970
rect 19947 4918 19999 4970
rect 8482 4856 8534 4908
rect 8548 4878 8554 4908
rect 8554 4878 8588 4908
rect 8588 4878 8600 4908
rect 8548 4856 8600 4878
rect 8614 4878 8627 4908
rect 8627 4878 8661 4908
rect 8661 4878 8666 4908
rect 8614 4856 8666 4878
rect 8680 4878 8700 4908
rect 8700 4878 8732 4908
rect 8746 4878 8773 4908
rect 8773 4878 8798 4908
rect 8811 4878 8846 4908
rect 8846 4878 8863 4908
rect 8876 4878 8880 4908
rect 8880 4878 8919 4908
rect 8919 4878 8928 4908
rect 8941 4878 8953 4908
rect 8953 4878 8992 4908
rect 8992 4878 8993 4908
rect 9006 4878 9026 4908
rect 9026 4878 9058 4908
rect 9071 4878 9099 4908
rect 9099 4878 9123 4908
rect 8680 4856 8732 4878
rect 8746 4856 8798 4878
rect 8811 4856 8863 4878
rect 8876 4856 8928 4878
rect 8941 4856 8993 4878
rect 9006 4856 9058 4878
rect 9071 4856 9123 4878
rect 9136 4878 9138 4908
rect 9138 4878 9172 4908
rect 9172 4878 9188 4908
rect 9136 4856 9188 4878
rect 9201 4878 9211 4908
rect 9211 4878 9245 4908
rect 9245 4878 9253 4908
rect 9201 4856 9253 4878
rect 9266 4878 9284 4908
rect 9284 4878 9318 4908
rect 9266 4856 9318 4878
rect 9331 4878 9357 4908
rect 9357 4878 9383 4908
rect 9396 4878 9430 4908
rect 9430 4878 9448 4908
rect 9461 4878 9464 4908
rect 9464 4878 9503 4908
rect 9503 4878 9513 4908
rect 9526 4878 9537 4908
rect 9537 4878 9576 4908
rect 9576 4878 9578 4908
rect 9591 4878 9610 4908
rect 9610 4878 9643 4908
rect 9656 4878 9683 4908
rect 9683 4878 9708 4908
rect 9331 4856 9383 4878
rect 9396 4856 9448 4878
rect 9461 4856 9513 4878
rect 9526 4856 9578 4878
rect 9591 4856 9643 4878
rect 9656 4856 9708 4878
rect 9721 4878 9722 4908
rect 9722 4878 9756 4908
rect 9756 4878 9773 4908
rect 9721 4856 9773 4878
rect 9786 4878 9795 4908
rect 9795 4878 9829 4908
rect 9829 4878 9838 4908
rect 9786 4856 9838 4878
rect 9851 4878 9868 4908
rect 9868 4878 9902 4908
rect 9902 4878 9903 4908
rect 9851 4856 9903 4878
rect 9916 4878 9941 4908
rect 9941 4878 9968 4908
rect 9981 4878 10014 4908
rect 10014 4878 10033 4908
rect 10046 4878 10048 4908
rect 10048 4878 10087 4908
rect 10087 4878 10098 4908
rect 10111 4878 10121 4908
rect 10121 4878 10160 4908
rect 10160 4878 10163 4908
rect 10176 4878 10194 4908
rect 10194 4878 10228 4908
rect 10241 4878 10267 4908
rect 10267 4878 10293 4908
rect 9916 4856 9968 4878
rect 9981 4856 10033 4878
rect 10046 4856 10098 4878
rect 10111 4856 10163 4878
rect 10176 4856 10228 4878
rect 10241 4856 10293 4878
rect 10306 4878 10340 4908
rect 10340 4878 10358 4908
rect 10306 4856 10358 4878
rect 10371 4878 10379 4908
rect 10379 4878 10413 4908
rect 10413 4878 10423 4908
rect 10371 4856 10423 4878
rect 10436 4878 10452 4908
rect 10452 4878 10486 4908
rect 10486 4878 10488 4908
rect 10436 4856 10488 4878
rect 10501 4878 10525 4908
rect 10525 4878 10553 4908
rect 10566 4878 10598 4908
rect 10598 4878 10618 4908
rect 10631 4878 10632 4908
rect 10632 4878 10671 4908
rect 10671 4878 10683 4908
rect 10696 4878 10705 4908
rect 10705 4878 10744 4908
rect 10744 4878 10748 4908
rect 10761 4878 10778 4908
rect 10778 4878 10813 4908
rect 10826 4878 10851 4908
rect 10851 4878 10878 4908
rect 10891 4878 10924 4908
rect 10924 4878 10943 4908
rect 10501 4856 10553 4878
rect 10566 4856 10618 4878
rect 10631 4856 10683 4878
rect 10696 4856 10748 4878
rect 10761 4856 10813 4878
rect 10826 4856 10878 4878
rect 10891 4856 10943 4878
rect 10956 4878 10963 4908
rect 10963 4878 10997 4908
rect 10997 4878 11008 4908
rect 10956 4856 11008 4878
rect 11021 4878 11036 4908
rect 11036 4878 11070 4908
rect 11070 4878 11073 4908
rect 11021 4856 11073 4878
rect 11086 4878 11109 4908
rect 11109 4878 11138 4908
rect 11151 4878 11182 4908
rect 11182 4878 11203 4908
rect 11216 4878 11255 4908
rect 11255 4878 11268 4908
rect 11281 4878 11289 4908
rect 11289 4878 11328 4908
rect 11328 4878 11333 4908
rect 11346 4878 11362 4908
rect 11362 4878 11398 4908
rect 11411 4878 11435 4908
rect 11435 4878 11463 4908
rect 19755 4878 19757 4879
rect 19757 4878 19791 4879
rect 19791 4878 19807 4879
rect 11086 4856 11138 4878
rect 11151 4856 11203 4878
rect 11216 4856 11268 4878
rect 11281 4856 11333 4878
rect 11346 4856 11398 4878
rect 11411 4856 11463 4878
rect 8473 4804 8482 4806
rect 8482 4804 8516 4806
rect 8516 4804 8525 4806
rect 8473 4764 8525 4804
rect 8473 4754 8482 4764
rect 8482 4754 8516 4764
rect 8516 4754 8525 4764
rect 8473 4690 8525 4723
rect 8473 4671 8482 4690
rect 8482 4671 8516 4690
rect 8516 4671 8525 4690
rect 8861 4774 8870 4806
rect 8870 4774 8904 4806
rect 8904 4774 8913 4806
rect 8861 4754 8913 4774
rect 8861 4702 8870 4723
rect 8870 4702 8904 4723
rect 8904 4702 8913 4723
rect 8861 4671 8913 4702
rect 454 4472 506 4502
rect 454 4450 467 4472
rect 467 4450 501 4472
rect 501 4450 506 4472
rect 454 4397 506 4420
rect 454 4368 467 4397
rect 467 4368 501 4397
rect 501 4368 506 4397
rect 454 4322 506 4338
rect 454 4288 467 4322
rect 467 4288 501 4322
rect 501 4288 506 4322
rect 454 4286 506 4288
rect 952 4492 1004 4497
rect 1044 4492 1096 4497
rect 1135 4492 1187 4497
rect 952 4458 962 4492
rect 962 4458 1004 4492
rect 1044 4458 1084 4492
rect 1084 4458 1096 4492
rect 1135 4458 1162 4492
rect 1162 4458 1187 4492
rect 952 4445 1004 4458
rect 1044 4445 1096 4458
rect 1135 4445 1187 4458
rect 1783 4486 1835 4498
rect 1783 4452 1789 4486
rect 1789 4452 1823 4486
rect 1823 4452 1835 4486
rect 1783 4446 1835 4452
rect 1850 4486 1902 4498
rect 1850 4452 1865 4486
rect 1865 4452 1899 4486
rect 1899 4452 1902 4486
rect 1850 4446 1902 4452
rect 1917 4486 1969 4498
rect 1983 4486 2035 4498
rect 2049 4486 2101 4498
rect 2115 4486 2167 4498
rect 2181 4486 2233 4498
rect 2247 4486 2299 4498
rect 1917 4452 1941 4486
rect 1941 4452 1969 4486
rect 1983 4452 2017 4486
rect 2017 4452 2035 4486
rect 2049 4452 2051 4486
rect 2051 4452 2093 4486
rect 2093 4452 2101 4486
rect 2115 4452 2127 4486
rect 2127 4452 2167 4486
rect 2181 4452 2203 4486
rect 2203 4452 2233 4486
rect 2247 4452 2278 4486
rect 2278 4452 2299 4486
rect 1917 4446 1969 4452
rect 1983 4446 2035 4452
rect 2049 4446 2101 4452
rect 2115 4446 2167 4452
rect 2181 4446 2233 4452
rect 2247 4446 2299 4452
rect 2313 4486 2365 4498
rect 2313 4452 2319 4486
rect 2319 4452 2353 4486
rect 2353 4452 2365 4486
rect 2313 4446 2365 4452
rect 2379 4486 2431 4498
rect 2379 4452 2394 4486
rect 2394 4452 2428 4486
rect 2428 4452 2431 4486
rect 2379 4446 2431 4452
rect 2445 4486 2497 4498
rect 2511 4486 2563 4498
rect 2577 4486 2629 4498
rect 2643 4486 2695 4498
rect 2709 4486 2761 4498
rect 2775 4486 2827 4498
rect 2445 4452 2469 4486
rect 2469 4452 2497 4486
rect 2511 4452 2544 4486
rect 2544 4452 2563 4486
rect 2577 4452 2578 4486
rect 2578 4452 2619 4486
rect 2619 4452 2629 4486
rect 2643 4452 2653 4486
rect 2653 4452 2694 4486
rect 2694 4452 2695 4486
rect 2709 4452 2728 4486
rect 2728 4452 2761 4486
rect 2775 4452 2803 4486
rect 2803 4452 2827 4486
rect 2445 4446 2497 4452
rect 2511 4446 2563 4452
rect 2577 4446 2629 4452
rect 2643 4446 2695 4452
rect 2709 4446 2761 4452
rect 2775 4446 2827 4452
rect 2841 4486 2893 4498
rect 2841 4452 2844 4486
rect 2844 4452 2878 4486
rect 2878 4452 2893 4486
rect 2841 4446 2893 4452
rect 2907 4486 2959 4498
rect 2907 4452 2919 4486
rect 2919 4452 2953 4486
rect 2953 4452 2959 4486
rect 2907 4446 2959 4452
rect 952 4365 1004 4417
rect 1044 4365 1096 4417
rect 1135 4365 1187 4417
rect 1665 4361 1717 4413
rect 1746 4393 1798 4413
rect 1746 4361 1761 4393
rect 1761 4361 1798 4393
rect 952 4285 1004 4337
rect 1044 4285 1096 4337
rect 1135 4285 1187 4337
rect 1665 4285 1717 4337
rect 1746 4321 1798 4337
rect 1746 4287 1761 4321
rect 1761 4287 1798 4321
rect 1746 4285 1798 4287
rect 454 4247 506 4256
rect 454 4213 467 4247
rect 467 4213 501 4247
rect 501 4213 506 4247
rect 454 4204 506 4213
rect 2230 4393 2282 4407
rect 2230 4359 2239 4393
rect 2239 4359 2273 4393
rect 2273 4359 2282 4393
rect 2230 4355 2282 4359
rect 2230 4321 2282 4343
rect 2230 4291 2239 4321
rect 2239 4291 2273 4321
rect 2273 4291 2282 4321
rect 2742 4393 2794 4407
rect 2742 4359 2751 4393
rect 2751 4359 2785 4393
rect 2785 4359 2794 4393
rect 2742 4355 2794 4359
rect 2742 4321 2794 4343
rect 2742 4291 2751 4321
rect 2751 4291 2785 4321
rect 2785 4291 2794 4321
rect 3089 4486 3141 4498
rect 3089 4452 3095 4486
rect 3095 4452 3129 4486
rect 3129 4452 3141 4486
rect 3089 4446 3141 4452
rect 3158 4486 3210 4498
rect 3158 4452 3173 4486
rect 3173 4452 3207 4486
rect 3207 4452 3210 4486
rect 3158 4446 3210 4452
rect 3227 4486 3279 4498
rect 3296 4486 3348 4498
rect 3365 4486 3417 4498
rect 3434 4486 3486 4498
rect 3502 4486 3554 4498
rect 3570 4486 3622 4498
rect 3227 4452 3251 4486
rect 3251 4452 3279 4486
rect 3296 4452 3329 4486
rect 3329 4452 3348 4486
rect 3365 4452 3407 4486
rect 3407 4452 3417 4486
rect 3434 4452 3441 4486
rect 3441 4452 3485 4486
rect 3485 4452 3486 4486
rect 3502 4452 3519 4486
rect 3519 4452 3554 4486
rect 3570 4452 3597 4486
rect 3597 4452 3622 4486
rect 3227 4446 3279 4452
rect 3296 4446 3348 4452
rect 3365 4446 3417 4452
rect 3434 4446 3486 4452
rect 3502 4446 3554 4452
rect 3570 4446 3622 4452
rect 3638 4486 3690 4498
rect 3638 4452 3641 4486
rect 3641 4452 3675 4486
rect 3675 4452 3690 4486
rect 3638 4446 3690 4452
rect 3706 4486 3758 4498
rect 3706 4452 3718 4486
rect 3718 4452 3752 4486
rect 3752 4452 3758 4486
rect 3706 4446 3758 4452
rect 3254 4393 3306 4407
rect 3254 4359 3263 4393
rect 3263 4359 3297 4393
rect 3297 4359 3306 4393
rect 3254 4355 3306 4359
rect 3254 4321 3306 4343
rect 3254 4291 3263 4321
rect 3263 4291 3297 4321
rect 3297 4291 3306 4321
rect 3766 4393 3818 4407
rect 3766 4359 3775 4393
rect 3775 4359 3809 4393
rect 3809 4359 3818 4393
rect 3766 4355 3818 4359
rect 3766 4321 3818 4343
rect 3766 4291 3775 4321
rect 3775 4291 3809 4321
rect 3809 4291 3818 4321
rect 3889 4355 3941 4407
rect 3889 4291 3941 4343
rect 4127 4486 4179 4498
rect 4127 4452 4133 4486
rect 4133 4452 4167 4486
rect 4167 4452 4179 4486
rect 4127 4446 4179 4452
rect 4218 4486 4270 4498
rect 4218 4452 4230 4486
rect 4230 4452 4264 4486
rect 4264 4452 4270 4486
rect 4218 4446 4270 4452
rect 4594 4486 4646 4498
rect 4594 4452 4600 4486
rect 4600 4452 4634 4486
rect 4634 4452 4646 4486
rect 4594 4446 4646 4452
rect 4659 4486 4711 4498
rect 4659 4452 4675 4486
rect 4675 4452 4709 4486
rect 4709 4452 4711 4486
rect 4659 4446 4711 4452
rect 4724 4486 4776 4498
rect 4789 4486 4841 4498
rect 4853 4486 4905 4498
rect 4917 4486 4969 4498
rect 4981 4486 5033 4498
rect 4724 4452 4750 4486
rect 4750 4452 4776 4486
rect 4789 4452 4825 4486
rect 4825 4452 4841 4486
rect 4853 4452 4859 4486
rect 4859 4452 4900 4486
rect 4900 4452 4905 4486
rect 4917 4452 4934 4486
rect 4934 4452 4969 4486
rect 4981 4452 5009 4486
rect 5009 4452 5033 4486
rect 4724 4446 4776 4452
rect 4789 4446 4841 4452
rect 4853 4446 4905 4452
rect 4917 4446 4969 4452
rect 4981 4446 5033 4452
rect 5045 4486 5097 4498
rect 5045 4452 5050 4486
rect 5050 4452 5084 4486
rect 5084 4452 5097 4486
rect 5045 4446 5097 4452
rect 5109 4486 5161 4498
rect 5109 4452 5125 4486
rect 5125 4452 5159 4486
rect 5159 4452 5161 4486
rect 5109 4446 5161 4452
rect 5173 4486 5225 4498
rect 5237 4486 5289 4498
rect 5301 4486 5353 4498
rect 5365 4486 5417 4498
rect 5429 4486 5481 4498
rect 5173 4452 5199 4486
rect 5199 4452 5225 4486
rect 5237 4452 5273 4486
rect 5273 4452 5289 4486
rect 5301 4452 5307 4486
rect 5307 4452 5347 4486
rect 5347 4452 5353 4486
rect 5365 4452 5381 4486
rect 5381 4452 5417 4486
rect 5429 4452 5455 4486
rect 5455 4452 5481 4486
rect 5173 4446 5225 4452
rect 5237 4446 5289 4452
rect 5301 4446 5353 4452
rect 5365 4446 5417 4452
rect 5429 4446 5481 4452
rect 5493 4486 5545 4498
rect 5493 4452 5495 4486
rect 5495 4452 5529 4486
rect 5529 4452 5545 4486
rect 5493 4446 5545 4452
rect 5557 4486 5609 4498
rect 5557 4452 5569 4486
rect 5569 4452 5603 4486
rect 5603 4452 5609 4486
rect 5557 4446 5609 4452
rect 5621 4486 5673 4498
rect 5685 4486 5737 4498
rect 5749 4486 5801 4498
rect 5813 4486 5865 4498
rect 5877 4486 5929 4498
rect 5941 4486 5993 4498
rect 5621 4452 5643 4486
rect 5643 4452 5673 4486
rect 5685 4452 5717 4486
rect 5717 4452 5737 4486
rect 5749 4452 5751 4486
rect 5751 4452 5791 4486
rect 5791 4452 5801 4486
rect 5813 4452 5825 4486
rect 5825 4452 5865 4486
rect 5877 4452 5899 4486
rect 5899 4452 5929 4486
rect 5941 4452 5973 4486
rect 5973 4452 5993 4486
rect 5621 4446 5673 4452
rect 5685 4446 5737 4452
rect 5749 4446 5801 4452
rect 5813 4446 5865 4452
rect 5877 4446 5929 4452
rect 5941 4446 5993 4452
rect 6005 4486 6057 4498
rect 6005 4452 6013 4486
rect 6013 4452 6047 4486
rect 6047 4452 6057 4486
rect 6005 4446 6057 4452
rect 6069 4486 6121 4498
rect 6069 4452 6087 4486
rect 6087 4452 6121 4486
rect 6069 4446 6121 4452
rect 6133 4486 6185 4498
rect 6197 4486 6249 4498
rect 6261 4486 6313 4498
rect 6325 4486 6377 4498
rect 6389 4486 6441 4498
rect 6133 4452 6161 4486
rect 6161 4452 6185 4486
rect 6197 4452 6235 4486
rect 6235 4452 6249 4486
rect 6261 4452 6269 4486
rect 6269 4452 6309 4486
rect 6309 4452 6313 4486
rect 6325 4452 6343 4486
rect 6343 4452 6377 4486
rect 6389 4452 6417 4486
rect 6417 4452 6441 4486
rect 6133 4446 6185 4452
rect 6197 4446 6249 4452
rect 6261 4446 6313 4452
rect 6325 4446 6377 4452
rect 6389 4446 6441 4452
rect 6453 4486 6505 4498
rect 6453 4452 6457 4486
rect 6457 4452 6491 4486
rect 6491 4452 6505 4486
rect 6453 4446 6505 4452
rect 6517 4486 6569 4498
rect 6517 4452 6531 4486
rect 6531 4452 6565 4486
rect 6565 4452 6569 4486
rect 6517 4446 6569 4452
rect 6674 4446 6726 4498
rect 6743 4446 6795 4498
rect 4278 4393 4330 4407
rect 4278 4359 4287 4393
rect 4287 4359 4321 4393
rect 4321 4359 4330 4393
rect 4278 4355 4330 4359
rect 4278 4321 4330 4343
rect 4278 4291 4287 4321
rect 4287 4291 4321 4321
rect 4321 4291 4330 4321
rect 4401 4355 4453 4407
rect 4401 4291 4453 4343
rect 4790 4393 4842 4407
rect 4790 4359 4799 4393
rect 4799 4359 4833 4393
rect 4833 4359 4842 4393
rect 4790 4355 4842 4359
rect 4790 4321 4842 4343
rect 4790 4291 4799 4321
rect 4799 4291 4833 4321
rect 4833 4291 4842 4321
rect 5302 4393 5354 4407
rect 5302 4359 5311 4393
rect 5311 4359 5345 4393
rect 5345 4359 5354 4393
rect 5302 4355 5354 4359
rect 5302 4321 5354 4343
rect 5302 4291 5311 4321
rect 5311 4291 5345 4321
rect 5345 4291 5354 4321
rect 3007 4195 3059 4247
rect 3071 4195 3123 4247
rect 3519 4195 3571 4247
rect 3583 4195 3635 4247
rect 4365 4195 4417 4247
rect 4429 4195 4481 4247
rect 4973 4195 5025 4247
rect 5037 4195 5089 4247
rect 5814 4393 5866 4407
rect 5814 4359 5823 4393
rect 5823 4359 5857 4393
rect 5857 4359 5866 4393
rect 5814 4355 5866 4359
rect 5814 4321 5866 4343
rect 5814 4291 5823 4321
rect 5823 4291 5857 4321
rect 5857 4291 5866 4321
rect 6326 4393 6378 4407
rect 6326 4359 6335 4393
rect 6335 4359 6369 4393
rect 6369 4359 6378 4393
rect 6326 4355 6378 4359
rect 6326 4321 6378 4343
rect 6326 4291 6335 4321
rect 6335 4291 6369 4321
rect 6369 4291 6378 4321
rect 454 4172 506 4174
rect 454 4138 467 4172
rect 467 4138 501 4172
rect 501 4138 506 4172
rect 454 4122 506 4138
rect 454 4063 467 4092
rect 467 4063 501 4092
rect 501 4063 506 4092
rect 454 4040 506 4063
rect 699 4109 751 4161
rect 2454 4119 2506 4171
rect 2518 4119 2570 4171
rect 5908 4115 5960 4167
rect 5972 4115 6024 4167
rect 6847 4393 6899 4413
rect 6847 4361 6881 4393
rect 6881 4361 6899 4393
rect 6953 4361 7005 4413
rect 7058 4361 7110 4413
rect 7163 4361 7215 4413
rect 7268 4361 7320 4413
rect 7373 4361 7425 4413
rect 7478 4361 7530 4413
rect 7597 4361 7649 4413
rect 7705 4393 7757 4413
rect 7705 4361 7737 4393
rect 7737 4361 7757 4393
rect 6847 4321 6899 4337
rect 6847 4287 6881 4321
rect 6881 4287 6899 4321
rect 6847 4285 6899 4287
rect 6953 4285 7005 4337
rect 7058 4285 7110 4337
rect 7163 4285 7215 4337
rect 7268 4285 7320 4337
rect 7373 4285 7425 4337
rect 7478 4285 7530 4337
rect 7597 4285 7649 4337
rect 7705 4321 7757 4337
rect 7705 4287 7737 4321
rect 7737 4287 7757 4321
rect 7705 4285 7757 4287
rect 8103 4562 8155 4614
rect 8103 4498 8155 4550
rect 6674 4198 6726 4250
rect 6743 4198 6795 4250
rect 454 3988 467 4010
rect 467 3988 501 4010
rect 501 3988 506 4010
rect 454 3958 506 3988
rect 617 4005 669 4057
rect 699 4045 751 4097
rect 1264 4027 1316 4079
rect 1328 4027 1380 4079
rect 3519 4027 3571 4079
rect 3583 4027 3635 4079
rect 4973 4027 5025 4079
rect 5037 4027 5089 4079
rect 617 3941 669 3993
rect 3007 3935 3059 3987
rect 3071 3935 3123 3987
rect 454 3913 467 3928
rect 467 3913 501 3928
rect 501 3913 506 3928
rect 454 3876 506 3913
rect 454 3838 467 3846
rect 467 3838 501 3846
rect 501 3838 506 3846
rect 454 3797 506 3838
rect 454 3794 467 3797
rect 467 3794 501 3797
rect 501 3794 506 3797
rect 2454 3851 2506 3903
rect 2518 3851 2570 3903
rect 454 3763 467 3764
rect 467 3763 501 3764
rect 501 3763 506 3764
rect 454 3722 506 3763
rect 454 3712 467 3722
rect 467 3712 501 3722
rect 501 3712 506 3722
rect 454 3647 506 3681
rect 454 3629 467 3647
rect 467 3629 501 3647
rect 501 3629 506 3647
rect 952 3763 1004 3815
rect 1044 3763 1096 3815
rect 1135 3763 1187 3815
rect 1624 3763 1676 3815
rect 1709 3813 1761 3815
rect 1709 3779 1727 3813
rect 1727 3779 1761 3813
rect 1709 3763 1761 3779
rect 952 3683 1004 3735
rect 1044 3683 1096 3735
rect 1135 3683 1187 3735
rect 1624 3687 1676 3739
rect 1709 3707 1727 3739
rect 1727 3707 1761 3739
rect 1709 3687 1761 3707
rect 2230 3779 2239 3809
rect 2239 3779 2273 3809
rect 2273 3779 2282 3809
rect 2230 3757 2282 3779
rect 2230 3741 2282 3745
rect 2230 3707 2239 3741
rect 2239 3707 2273 3741
rect 2273 3707 2282 3741
rect 2230 3693 2282 3707
rect 2742 3779 2751 3809
rect 2751 3779 2785 3809
rect 2785 3779 2794 3809
rect 2742 3757 2794 3779
rect 2742 3741 2794 3745
rect 2742 3707 2751 3741
rect 2751 3707 2785 3741
rect 2785 3707 2794 3741
rect 2742 3693 2794 3707
rect 3519 3853 3571 3905
rect 3583 3853 3635 3905
rect 4365 3853 4417 3905
rect 4429 3853 4481 3905
rect 4973 3853 5025 3905
rect 5037 3853 5089 3905
rect 3254 3779 3263 3809
rect 3263 3779 3297 3809
rect 3297 3779 3306 3809
rect 3254 3757 3306 3779
rect 3254 3741 3306 3745
rect 3254 3707 3263 3741
rect 3263 3707 3297 3741
rect 3297 3707 3306 3741
rect 3254 3693 3306 3707
rect 3766 3779 3775 3809
rect 3775 3779 3809 3809
rect 3809 3779 3818 3809
rect 3766 3757 3818 3779
rect 3766 3741 3818 3745
rect 3766 3707 3775 3741
rect 3775 3707 3809 3741
rect 3809 3707 3818 3741
rect 3766 3693 3818 3707
rect 4145 3757 4197 3809
rect 4145 3693 4197 3745
rect 454 3572 506 3598
rect 454 3546 467 3572
rect 467 3546 501 3572
rect 501 3546 506 3572
rect 454 3498 506 3515
rect 454 3464 467 3498
rect 467 3464 501 3498
rect 501 3464 506 3498
rect 454 3463 506 3464
rect 535 3565 587 3617
rect 952 3642 1004 3655
rect 1044 3642 1096 3655
rect 1135 3642 1187 3655
rect 4278 3779 4287 3809
rect 4287 3779 4321 3809
rect 4321 3779 4330 3809
rect 4278 3757 4330 3779
rect 4278 3741 4330 3745
rect 4278 3707 4287 3741
rect 4287 3707 4321 3741
rect 4321 3707 4330 3741
rect 4278 3693 4330 3707
rect 952 3608 962 3642
rect 962 3608 1004 3642
rect 1044 3608 1084 3642
rect 1084 3608 1096 3642
rect 1135 3608 1162 3642
rect 1162 3608 1187 3642
rect 952 3603 1004 3608
rect 1044 3603 1096 3608
rect 1135 3603 1187 3608
rect 2553 3645 2605 3653
rect 2553 3611 2557 3645
rect 2557 3611 2591 3645
rect 2591 3611 2605 3645
rect 2553 3601 2605 3611
rect 2618 3645 2670 3653
rect 2618 3611 2633 3645
rect 2633 3611 2667 3645
rect 2667 3611 2670 3645
rect 2618 3601 2670 3611
rect 2682 3645 2734 3653
rect 2746 3645 2798 3653
rect 2810 3645 2862 3653
rect 2874 3645 2926 3653
rect 2938 3645 2990 3653
rect 2682 3611 2709 3645
rect 2709 3611 2734 3645
rect 2746 3611 2785 3645
rect 2785 3611 2798 3645
rect 2810 3611 2819 3645
rect 2819 3611 2861 3645
rect 2861 3611 2862 3645
rect 2874 3611 2895 3645
rect 2895 3611 2926 3645
rect 2938 3611 2970 3645
rect 2970 3611 2990 3645
rect 2682 3601 2734 3611
rect 2746 3601 2798 3611
rect 2810 3601 2862 3611
rect 2874 3601 2926 3611
rect 2938 3601 2990 3611
rect 3002 3645 3054 3653
rect 3002 3611 3011 3645
rect 3011 3611 3045 3645
rect 3045 3611 3054 3645
rect 3002 3601 3054 3611
rect 3066 3645 3118 3653
rect 3130 3645 3182 3653
rect 3194 3645 3246 3653
rect 3258 3645 3310 3653
rect 3322 3645 3374 3653
rect 3066 3611 3086 3645
rect 3086 3611 3118 3645
rect 3130 3611 3161 3645
rect 3161 3611 3182 3645
rect 3194 3611 3195 3645
rect 3195 3611 3236 3645
rect 3236 3611 3246 3645
rect 3258 3611 3270 3645
rect 3270 3611 3310 3645
rect 3322 3611 3345 3645
rect 3345 3611 3374 3645
rect 3066 3601 3118 3611
rect 3130 3601 3182 3611
rect 3194 3601 3246 3611
rect 3258 3601 3310 3611
rect 3322 3601 3374 3611
rect 3386 3645 3438 3653
rect 3386 3611 3420 3645
rect 3420 3611 3438 3645
rect 3386 3601 3438 3611
rect 3450 3645 3502 3653
rect 3450 3611 3461 3645
rect 3461 3611 3495 3645
rect 3495 3611 3502 3645
rect 3450 3601 3502 3611
rect 3514 3645 3566 3653
rect 3578 3645 3630 3653
rect 3642 3645 3694 3653
rect 3706 3645 3758 3653
rect 3770 3645 3822 3653
rect 3514 3611 3536 3645
rect 3536 3611 3566 3645
rect 3578 3611 3611 3645
rect 3611 3611 3630 3645
rect 3642 3611 3645 3645
rect 3645 3611 3686 3645
rect 3686 3611 3694 3645
rect 3706 3611 3720 3645
rect 3720 3611 3758 3645
rect 3770 3611 3795 3645
rect 3795 3611 3822 3645
rect 3514 3601 3566 3611
rect 3578 3601 3630 3611
rect 3642 3601 3694 3611
rect 3706 3601 3758 3611
rect 3770 3601 3822 3611
rect 3834 3645 3886 3653
rect 3834 3611 3836 3645
rect 3836 3611 3870 3645
rect 3870 3611 3886 3645
rect 3834 3601 3886 3611
rect 3898 3645 3950 3653
rect 3898 3611 3911 3645
rect 3911 3611 3945 3645
rect 3945 3611 3950 3645
rect 3898 3601 3950 3611
rect 3962 3645 4014 3653
rect 3962 3611 3986 3645
rect 3986 3611 4014 3645
rect 3962 3601 4014 3611
rect 4338 3645 4390 3653
rect 4338 3611 4366 3645
rect 4366 3611 4390 3645
rect 4338 3601 4390 3611
rect 4433 3645 4485 3653
rect 4433 3611 4445 3645
rect 4445 3611 4479 3645
rect 4479 3611 4485 3645
rect 4433 3601 4485 3611
rect 4657 3757 4709 3809
rect 4657 3693 4709 3745
rect 4790 3779 4799 3809
rect 4799 3779 4833 3809
rect 4833 3779 4842 3809
rect 4790 3757 4842 3779
rect 4790 3741 4842 3745
rect 4790 3707 4799 3741
rect 4799 3707 4833 3741
rect 4833 3707 4842 3741
rect 4790 3693 4842 3707
rect 5302 3779 5311 3809
rect 5311 3779 5345 3809
rect 5345 3779 5354 3809
rect 5302 3757 5354 3779
rect 5302 3741 5354 3745
rect 5302 3707 5311 3741
rect 5311 3707 5345 3741
rect 5345 3707 5354 3741
rect 5302 3693 5354 3707
rect 5908 3853 5960 3905
rect 5972 3853 6024 3905
rect 5814 3779 5823 3809
rect 5823 3779 5857 3809
rect 5857 3779 5866 3809
rect 5814 3757 5866 3779
rect 5814 3741 5866 3745
rect 5814 3707 5823 3741
rect 5823 3707 5857 3741
rect 5857 3707 5866 3741
rect 5814 3693 5866 3707
rect 6326 3779 6335 3809
rect 6335 3779 6369 3809
rect 6369 3779 6378 3809
rect 6326 3757 6378 3779
rect 6326 3741 6378 3745
rect 6326 3707 6335 3741
rect 6335 3707 6369 3741
rect 6369 3707 6378 3741
rect 6326 3693 6378 3707
rect 7826 4141 7838 4170
rect 7838 4141 7872 4170
rect 7872 4141 7878 4170
rect 7826 4118 7878 4141
rect 7826 4100 7878 4106
rect 7826 4066 7838 4100
rect 7838 4066 7872 4100
rect 7872 4066 7878 4100
rect 7826 4054 7878 4066
rect 6847 3813 6899 3815
rect 6847 3779 6881 3813
rect 6881 3779 6899 3813
rect 6847 3763 6899 3779
rect 6954 3763 7006 3815
rect 7061 3763 7113 3815
rect 7168 3763 7220 3815
rect 7275 3763 7327 3815
rect 7382 3763 7434 3815
rect 6847 3707 6881 3739
rect 6881 3707 6899 3739
rect 6847 3687 6899 3707
rect 6954 3687 7006 3739
rect 7061 3687 7113 3739
rect 7168 3687 7220 3739
rect 7275 3687 7327 3739
rect 7382 3687 7434 3739
rect 4850 3645 4902 3653
rect 4921 3645 4973 3653
rect 4992 3645 5044 3653
rect 5062 3645 5114 3653
rect 4850 3611 4878 3645
rect 4878 3611 4902 3645
rect 4921 3611 4950 3645
rect 4950 3611 4973 3645
rect 4992 3611 5022 3645
rect 5022 3611 5044 3645
rect 5062 3611 5094 3645
rect 5094 3611 5114 3645
rect 4850 3601 4902 3611
rect 4921 3601 4973 3611
rect 4992 3601 5044 3611
rect 5062 3601 5114 3611
rect 5132 3645 5184 3653
rect 5132 3611 5166 3645
rect 5166 3611 5184 3645
rect 5132 3601 5184 3611
rect 5202 3645 5254 3653
rect 5202 3611 5204 3645
rect 5204 3611 5238 3645
rect 5238 3611 5254 3645
rect 5202 3601 5254 3611
rect 5272 3645 5324 3653
rect 5272 3611 5276 3645
rect 5276 3611 5310 3645
rect 5310 3611 5324 3645
rect 5272 3601 5324 3611
rect 5342 3645 5394 3653
rect 5342 3611 5348 3645
rect 5348 3611 5382 3645
rect 5382 3611 5394 3645
rect 5342 3601 5394 3611
rect 5412 3645 5464 3653
rect 5412 3611 5420 3645
rect 5420 3611 5454 3645
rect 5454 3611 5464 3645
rect 5412 3601 5464 3611
rect 5482 3645 5534 3653
rect 5482 3611 5492 3645
rect 5492 3611 5526 3645
rect 5526 3611 5534 3645
rect 5482 3601 5534 3611
rect 5552 3645 5604 3653
rect 5552 3611 5564 3645
rect 5564 3611 5598 3645
rect 5598 3611 5604 3645
rect 5552 3601 5604 3611
rect 5649 3645 5701 3653
rect 5649 3611 5655 3645
rect 5655 3611 5689 3645
rect 5689 3611 5701 3645
rect 5649 3601 5701 3611
rect 5715 3645 5767 3653
rect 5715 3611 5729 3645
rect 5729 3611 5763 3645
rect 5763 3611 5767 3645
rect 5715 3601 5767 3611
rect 5780 3645 5832 3653
rect 5845 3645 5897 3653
rect 5910 3645 5962 3653
rect 5975 3645 6027 3653
rect 6040 3645 6092 3653
rect 6105 3645 6157 3653
rect 5780 3611 5803 3645
rect 5803 3611 5832 3645
rect 5845 3611 5877 3645
rect 5877 3611 5897 3645
rect 5910 3611 5911 3645
rect 5911 3611 5951 3645
rect 5951 3611 5962 3645
rect 5975 3611 5985 3645
rect 5985 3611 6025 3645
rect 6025 3611 6027 3645
rect 6040 3611 6059 3645
rect 6059 3611 6092 3645
rect 6105 3611 6133 3645
rect 6133 3611 6157 3645
rect 5780 3601 5832 3611
rect 5845 3601 5897 3611
rect 5910 3601 5962 3611
rect 5975 3601 6027 3611
rect 6040 3601 6092 3611
rect 6105 3601 6157 3611
rect 6170 3645 6222 3653
rect 6170 3611 6173 3645
rect 6173 3611 6207 3645
rect 6207 3611 6222 3645
rect 6170 3601 6222 3611
rect 6235 3645 6287 3653
rect 6235 3611 6247 3645
rect 6247 3611 6281 3645
rect 6281 3611 6287 3645
rect 6235 3601 6287 3611
rect 6410 3645 6462 3653
rect 6410 3611 6416 3645
rect 6416 3611 6450 3645
rect 6450 3611 6462 3645
rect 6410 3601 6462 3611
rect 6523 3645 6575 3653
rect 6523 3611 6535 3645
rect 6535 3611 6569 3645
rect 6569 3611 6575 3645
rect 6523 3601 6575 3611
rect 6674 3601 6726 3653
rect 6743 3601 6795 3653
rect 535 3501 587 3553
rect 454 3424 506 3432
rect 454 3390 467 3424
rect 467 3390 501 3424
rect 501 3390 506 3424
rect 454 3380 506 3390
rect 454 3316 467 3349
rect 467 3316 501 3349
rect 501 3316 506 3349
rect 454 3297 506 3316
rect 454 3242 467 3266
rect 467 3242 501 3266
rect 501 3242 506 3266
rect 454 3214 506 3242
rect 952 3482 1004 3489
rect 1044 3482 1096 3489
rect 1135 3482 1187 3489
rect 952 3448 962 3482
rect 962 3448 1004 3482
rect 1044 3448 1084 3482
rect 1084 3448 1096 3482
rect 1135 3448 1162 3482
rect 1162 3448 1187 3482
rect 952 3437 1004 3448
rect 1044 3437 1096 3448
rect 1135 3437 1187 3448
rect 1778 3476 1830 3485
rect 1778 3442 1785 3476
rect 1785 3442 1819 3476
rect 1819 3442 1830 3476
rect 1778 3433 1830 3442
rect 1844 3476 1896 3485
rect 1844 3442 1859 3476
rect 1859 3442 1893 3476
rect 1893 3442 1896 3476
rect 1844 3433 1896 3442
rect 1910 3476 1962 3485
rect 1976 3476 2028 3485
rect 2042 3476 2094 3485
rect 2108 3476 2160 3485
rect 2174 3476 2226 3485
rect 2240 3476 2292 3485
rect 2306 3476 2358 3485
rect 2372 3476 2424 3485
rect 1910 3442 1932 3476
rect 1932 3442 1962 3476
rect 1976 3442 2005 3476
rect 2005 3442 2028 3476
rect 2042 3442 2078 3476
rect 2078 3442 2094 3476
rect 2108 3442 2112 3476
rect 2112 3442 2151 3476
rect 2151 3442 2160 3476
rect 2174 3442 2185 3476
rect 2185 3442 2224 3476
rect 2224 3442 2226 3476
rect 2240 3442 2258 3476
rect 2258 3442 2292 3476
rect 2306 3442 2331 3476
rect 2331 3442 2358 3476
rect 2372 3442 2404 3476
rect 2404 3442 2424 3476
rect 1910 3433 1962 3442
rect 1976 3433 2028 3442
rect 2042 3433 2094 3442
rect 2108 3433 2160 3442
rect 2174 3433 2226 3442
rect 2240 3433 2292 3442
rect 2306 3433 2358 3442
rect 2372 3433 2424 3442
rect 2437 3476 2489 3485
rect 2437 3442 2443 3476
rect 2443 3442 2477 3476
rect 2477 3442 2489 3476
rect 2437 3433 2489 3442
rect 2502 3476 2554 3485
rect 2502 3442 2516 3476
rect 2516 3442 2550 3476
rect 2550 3442 2554 3476
rect 2502 3433 2554 3442
rect 2567 3476 2619 3485
rect 2632 3476 2684 3485
rect 2697 3476 2749 3485
rect 2762 3476 2814 3485
rect 2827 3476 2879 3485
rect 2892 3476 2944 3485
rect 2957 3476 3009 3485
rect 2567 3442 2589 3476
rect 2589 3442 2619 3476
rect 2632 3442 2662 3476
rect 2662 3442 2684 3476
rect 2697 3442 2735 3476
rect 2735 3442 2749 3476
rect 2762 3442 2769 3476
rect 2769 3442 2808 3476
rect 2808 3442 2814 3476
rect 2827 3442 2842 3476
rect 2842 3442 2879 3476
rect 2892 3442 2915 3476
rect 2915 3442 2944 3476
rect 2957 3442 2988 3476
rect 2988 3442 3009 3476
rect 2567 3433 2619 3442
rect 2632 3433 2684 3442
rect 2697 3433 2749 3442
rect 2762 3433 2814 3442
rect 2827 3433 2879 3442
rect 2892 3433 2944 3442
rect 2957 3433 3009 3442
rect 3022 3476 3074 3485
rect 3022 3442 3027 3476
rect 3027 3442 3061 3476
rect 3061 3442 3074 3476
rect 3022 3433 3074 3442
rect 3087 3476 3139 3485
rect 3087 3442 3100 3476
rect 3100 3442 3134 3476
rect 3134 3442 3139 3476
rect 3087 3433 3139 3442
rect 3152 3476 3204 3485
rect 3217 3476 3269 3485
rect 3282 3476 3334 3485
rect 3347 3476 3399 3485
rect 3412 3476 3464 3485
rect 3477 3476 3529 3485
rect 3542 3476 3594 3485
rect 3152 3442 3173 3476
rect 3173 3442 3204 3476
rect 3217 3442 3246 3476
rect 3246 3442 3269 3476
rect 3282 3442 3319 3476
rect 3319 3442 3334 3476
rect 3347 3442 3353 3476
rect 3353 3442 3392 3476
rect 3392 3442 3399 3476
rect 3412 3442 3426 3476
rect 3426 3442 3464 3476
rect 3477 3442 3499 3476
rect 3499 3442 3529 3476
rect 3542 3442 3572 3476
rect 3572 3442 3594 3476
rect 3152 3433 3204 3442
rect 3217 3433 3269 3442
rect 3282 3433 3334 3442
rect 3347 3433 3399 3442
rect 3412 3433 3464 3442
rect 3477 3433 3529 3442
rect 3542 3433 3594 3442
rect 3607 3476 3659 3485
rect 3607 3442 3611 3476
rect 3611 3442 3645 3476
rect 3645 3442 3659 3476
rect 3607 3433 3659 3442
rect 3672 3476 3724 3485
rect 3672 3442 3684 3476
rect 3684 3442 3718 3476
rect 3718 3442 3724 3476
rect 3672 3433 3724 3442
rect 952 3373 1004 3425
rect 1044 3373 1096 3425
rect 1135 3373 1187 3425
rect 1581 3351 1633 3403
rect 1581 3275 1633 3327
rect 1974 3383 2026 3397
rect 1974 3349 1983 3383
rect 1983 3349 2017 3383
rect 2017 3349 2026 3383
rect 1974 3345 2026 3349
rect 1974 3311 2026 3333
rect 1974 3281 1983 3311
rect 1983 3281 2017 3311
rect 2017 3281 2026 3311
rect 2486 3383 2538 3397
rect 2486 3349 2495 3383
rect 2495 3349 2529 3383
rect 2529 3349 2538 3383
rect 2486 3345 2538 3349
rect 2486 3311 2538 3333
rect 2486 3281 2495 3311
rect 2495 3281 2529 3311
rect 2529 3281 2538 3311
rect 2998 3383 3050 3397
rect 2998 3349 3007 3383
rect 3007 3349 3041 3383
rect 3041 3349 3050 3383
rect 2998 3345 3050 3349
rect 2998 3311 3050 3333
rect 2998 3281 3007 3311
rect 3007 3281 3041 3311
rect 3041 3281 3050 3311
rect 3510 3383 3562 3397
rect 3510 3349 3519 3383
rect 3519 3349 3553 3383
rect 3553 3349 3562 3383
rect 3510 3345 3562 3349
rect 3510 3311 3562 3333
rect 3510 3281 3519 3311
rect 3519 3281 3553 3311
rect 3553 3281 3562 3311
rect 3855 3476 3907 3485
rect 3855 3442 3861 3476
rect 3861 3442 3895 3476
rect 3895 3442 3907 3476
rect 3855 3433 3907 3442
rect 3922 3476 3974 3485
rect 3989 3476 4041 3485
rect 4056 3476 4108 3485
rect 4123 3476 4175 3485
rect 3922 3442 3946 3476
rect 3946 3442 3974 3476
rect 3989 3442 4031 3476
rect 4031 3442 4041 3476
rect 4056 3442 4065 3476
rect 4065 3442 4108 3476
rect 4123 3442 4150 3476
rect 4150 3442 4175 3476
rect 3922 3433 3974 3442
rect 3989 3433 4041 3442
rect 4056 3433 4108 3442
rect 4123 3433 4175 3442
rect 4189 3476 4241 3485
rect 4189 3442 4201 3476
rect 4201 3442 4235 3476
rect 4235 3442 4241 3476
rect 4189 3433 4241 3442
rect 4022 3383 4074 3397
rect 4022 3349 4031 3383
rect 4031 3349 4065 3383
rect 4065 3349 4074 3383
rect 4022 3345 4074 3349
rect 4022 3311 4074 3333
rect 4022 3281 4031 3311
rect 4031 3281 4065 3311
rect 4065 3281 4074 3311
rect 4367 3476 4419 3485
rect 4367 3442 4373 3476
rect 4373 3442 4407 3476
rect 4407 3442 4419 3476
rect 4367 3433 4419 3442
rect 4434 3476 4486 3485
rect 4501 3476 4553 3485
rect 4568 3476 4620 3485
rect 4635 3476 4687 3485
rect 4434 3442 4458 3476
rect 4458 3442 4486 3476
rect 4501 3442 4543 3476
rect 4543 3442 4553 3476
rect 4568 3442 4577 3476
rect 4577 3442 4620 3476
rect 4635 3442 4662 3476
rect 4662 3442 4687 3476
rect 4434 3433 4486 3442
rect 4501 3433 4553 3442
rect 4568 3433 4620 3442
rect 4635 3433 4687 3442
rect 4701 3476 4753 3485
rect 4701 3442 4713 3476
rect 4713 3442 4747 3476
rect 4747 3442 4753 3476
rect 4701 3433 4753 3442
rect 4534 3383 4586 3397
rect 4534 3349 4543 3383
rect 4543 3349 4577 3383
rect 4577 3349 4586 3383
rect 4534 3345 4586 3349
rect 4534 3311 4586 3333
rect 4534 3281 4543 3311
rect 4543 3281 4577 3311
rect 4577 3281 4586 3311
rect 4879 3476 4931 3485
rect 4879 3442 4885 3476
rect 4885 3442 4919 3476
rect 4919 3442 4931 3476
rect 4879 3433 4931 3442
rect 4986 3476 5038 3485
rect 4986 3442 4998 3476
rect 4998 3442 5032 3476
rect 5032 3442 5038 3476
rect 4986 3433 5038 3442
rect 5618 3476 5670 3485
rect 5618 3442 5624 3476
rect 5624 3442 5658 3476
rect 5658 3442 5670 3476
rect 5618 3433 5670 3442
rect 5684 3476 5736 3485
rect 5684 3442 5700 3476
rect 5700 3442 5734 3476
rect 5734 3442 5736 3476
rect 5684 3433 5736 3442
rect 5750 3476 5802 3485
rect 5816 3476 5868 3485
rect 5882 3476 5934 3485
rect 5948 3476 6000 3485
rect 6014 3476 6066 3485
rect 5750 3442 5776 3476
rect 5776 3442 5802 3476
rect 5816 3442 5852 3476
rect 5852 3442 5868 3476
rect 5882 3442 5886 3476
rect 5886 3442 5928 3476
rect 5928 3442 5934 3476
rect 5948 3442 5962 3476
rect 5962 3442 6000 3476
rect 6014 3442 6038 3476
rect 6038 3442 6066 3476
rect 5750 3433 5802 3442
rect 5816 3433 5868 3442
rect 5882 3433 5934 3442
rect 5948 3433 6000 3442
rect 6014 3433 6066 3442
rect 6079 3476 6131 3485
rect 6079 3442 6080 3476
rect 6080 3442 6114 3476
rect 6114 3442 6131 3476
rect 6079 3433 6131 3442
rect 6144 3476 6196 3485
rect 6144 3442 6156 3476
rect 6156 3442 6190 3476
rect 6190 3442 6196 3476
rect 6144 3433 6196 3442
rect 6209 3476 6261 3485
rect 6274 3476 6326 3485
rect 6339 3476 6391 3485
rect 6404 3476 6456 3485
rect 6469 3476 6521 3485
rect 6209 3442 6232 3476
rect 6232 3442 6261 3476
rect 6274 3442 6308 3476
rect 6308 3442 6326 3476
rect 6339 3442 6342 3476
rect 6342 3442 6384 3476
rect 6384 3442 6391 3476
rect 6404 3442 6418 3476
rect 6418 3442 6456 3476
rect 6469 3442 6493 3476
rect 6493 3442 6521 3476
rect 6209 3433 6261 3442
rect 6274 3433 6326 3442
rect 6339 3433 6391 3442
rect 6404 3433 6456 3442
rect 6469 3433 6521 3442
rect 6534 3476 6586 3485
rect 6534 3442 6568 3476
rect 6568 3442 6586 3476
rect 6534 3433 6586 3442
rect 6674 3433 6726 3485
rect 6743 3433 6795 3485
rect 5046 3383 5098 3397
rect 5302 3383 5354 3397
rect 5558 3383 5610 3397
rect 5046 3349 5055 3383
rect 5055 3349 5089 3383
rect 5089 3349 5098 3383
rect 5046 3345 5098 3349
rect 5046 3311 5098 3333
rect 5046 3281 5055 3311
rect 5055 3281 5089 3311
rect 5089 3281 5098 3311
rect 5302 3349 5311 3383
rect 5311 3349 5345 3383
rect 5345 3349 5354 3383
rect 5302 3345 5354 3349
rect 5302 3311 5354 3333
rect 5302 3281 5311 3311
rect 5311 3281 5345 3311
rect 5345 3281 5354 3311
rect 5558 3349 5567 3383
rect 5567 3349 5601 3383
rect 5601 3349 5610 3383
rect 5558 3345 5610 3349
rect 5558 3311 5610 3333
rect 5558 3281 5567 3311
rect 5567 3281 5601 3311
rect 5601 3281 5610 3311
rect 6070 3383 6122 3397
rect 6070 3349 6079 3383
rect 6079 3349 6113 3383
rect 6113 3349 6122 3383
rect 6070 3345 6122 3349
rect 6070 3311 6122 3333
rect 6070 3281 6079 3311
rect 6079 3281 6113 3311
rect 6113 3281 6122 3311
rect 6582 3383 6634 3397
rect 6582 3349 6591 3383
rect 6591 3349 6625 3383
rect 6625 3349 6634 3383
rect 6582 3345 6634 3349
rect 6582 3311 6634 3333
rect 6582 3281 6591 3311
rect 6591 3281 6625 3311
rect 6625 3281 6634 3311
rect 6986 3351 7038 3403
rect 7085 3351 7137 3403
rect 7184 3351 7236 3403
rect 7283 3351 7335 3403
rect 7382 3351 7434 3403
rect 7712 3383 7764 3403
rect 7712 3351 7737 3383
rect 7737 3351 7764 3383
rect 7820 3391 7838 3403
rect 7838 3391 7872 3403
rect 7820 3351 7872 3391
rect 6986 3275 7038 3327
rect 7085 3275 7137 3327
rect 7184 3275 7236 3327
rect 7283 3275 7335 3327
rect 7382 3275 7434 3327
rect 7712 3311 7764 3327
rect 7712 3277 7737 3311
rect 7737 3277 7764 3311
rect 7712 3275 7764 3277
rect 7820 3316 7838 3327
rect 7838 3316 7872 3327
rect 7820 3275 7872 3316
rect 454 3168 467 3183
rect 467 3168 501 3183
rect 501 3168 506 3183
rect 454 3131 506 3168
rect 781 3177 833 3229
rect 6289 3183 6341 3235
rect 6353 3183 6405 3235
rect 454 3094 482 3100
rect 482 3094 506 3100
rect 781 3113 833 3165
rect 454 3048 506 3094
rect 863 3091 915 3143
rect 5035 3128 5087 3134
rect 5102 3128 5154 3134
rect 5169 3128 5221 3134
rect 5236 3128 5288 3134
rect 5303 3128 5355 3134
rect 5371 3128 5423 3134
rect 1582 3111 1634 3117
rect 863 3027 915 3079
rect 1582 3077 1584 3111
rect 1584 3077 1618 3111
rect 1618 3077 1634 3111
rect 1582 3065 1634 3077
rect 1646 3111 1698 3117
rect 1964 3111 2016 3117
rect 2028 3111 2080 3117
rect 1646 3077 1656 3111
rect 1656 3077 1690 3111
rect 1690 3077 1698 3111
rect 1964 3077 1978 3111
rect 1978 3077 2016 3111
rect 2028 3077 2050 3111
rect 2050 3077 2080 3111
rect 5035 3094 5064 3128
rect 5064 3094 5087 3128
rect 5102 3094 5137 3128
rect 5137 3094 5154 3128
rect 5169 3094 5171 3128
rect 5171 3094 5210 3128
rect 5210 3094 5221 3128
rect 5236 3094 5244 3128
rect 5244 3094 5283 3128
rect 5283 3094 5288 3128
rect 5303 3094 5317 3128
rect 5317 3094 5355 3128
rect 5371 3094 5390 3128
rect 5390 3094 5423 3128
rect 1646 3065 1698 3077
rect 1964 3065 2016 3077
rect 2028 3065 2080 3077
rect 5035 3082 5087 3094
rect 5102 3082 5154 3094
rect 5169 3082 5221 3094
rect 5236 3082 5288 3094
rect 5303 3082 5355 3094
rect 5371 3082 5423 3094
rect 7936 4092 7988 4144
rect 7936 4028 7988 4080
rect 8020 4020 8072 4072
rect 8020 3956 8072 4008
rect 1751 2989 1803 3041
rect 1815 2989 1867 3041
rect 5166 2989 5218 3041
rect 5230 2989 5282 3041
rect 1017 2843 1069 2895
rect 1116 2859 1232 2975
rect 8215 4573 8267 4625
rect 8279 4573 8331 4625
rect 1017 2779 1069 2831
rect 8269 4412 8321 4464
rect 8333 4412 8385 4464
rect 863 2687 915 2739
rect 8348 3949 8400 4001
rect 8348 3885 8400 3937
rect 9609 4774 9618 4806
rect 9618 4774 9652 4806
rect 9652 4774 9661 4806
rect 9609 4754 9661 4774
rect 9609 4702 9618 4723
rect 9618 4702 9652 4723
rect 9652 4702 9661 4723
rect 9609 4671 9661 4702
rect 9889 4774 9898 4806
rect 9898 4774 9932 4806
rect 9932 4774 9941 4806
rect 9889 4754 9941 4774
rect 9889 4702 9898 4723
rect 9898 4702 9932 4723
rect 9932 4702 9941 4723
rect 9889 4671 9941 4702
rect 10322 4774 10331 4806
rect 10331 4774 10365 4806
rect 10365 4774 10374 4806
rect 10322 4754 10374 4774
rect 10322 4702 10331 4723
rect 10331 4702 10365 4723
rect 10365 4702 10374 4723
rect 10322 4671 10374 4702
rect 10634 4774 10643 4806
rect 10643 4774 10677 4806
rect 10677 4774 10686 4806
rect 10634 4754 10686 4774
rect 10634 4702 10643 4723
rect 10643 4702 10677 4723
rect 10677 4702 10686 4723
rect 10634 4671 10686 4702
rect 10946 4774 10955 4806
rect 10955 4774 10989 4806
rect 10989 4774 10998 4806
rect 10946 4754 10998 4774
rect 10946 4702 10955 4723
rect 10955 4702 10989 4723
rect 10989 4702 10998 4723
rect 10946 4671 10998 4702
rect 9712 4304 9764 4322
rect 9712 4270 9742 4304
rect 9742 4270 9764 4304
rect 9776 4270 9828 4322
rect 9454 3982 9462 4007
rect 9462 3982 9496 4007
rect 9496 3982 9506 4007
rect 9454 3955 9506 3982
rect 9518 3955 9570 4007
rect 8655 3886 8707 3938
rect 8719 3910 8748 3938
rect 8748 3910 8771 3938
rect 8719 3886 8771 3910
rect 8978 3910 9026 3938
rect 9026 3910 9030 3938
rect 9042 3910 9060 3938
rect 9060 3910 9094 3938
rect 8978 3886 9030 3910
rect 9042 3886 9094 3910
rect 9296 3910 9338 3938
rect 9338 3910 9348 3938
rect 9360 3910 9372 3938
rect 9372 3910 9412 3938
rect 9296 3886 9348 3910
rect 9360 3886 9412 3910
rect 10045 4342 10054 4374
rect 10054 4342 10088 4374
rect 10088 4342 10097 4374
rect 10045 4322 10097 4342
rect 10045 4304 10097 4310
rect 10045 4270 10054 4304
rect 10054 4270 10088 4304
rect 10088 4270 10097 4304
rect 10045 4258 10097 4270
rect 10478 4160 10530 4170
rect 10478 4126 10487 4160
rect 10487 4126 10521 4160
rect 10521 4126 10530 4160
rect 10478 4118 10530 4126
rect 10478 4088 10530 4104
rect 10478 4054 10487 4088
rect 10487 4054 10521 4088
rect 10521 4054 10530 4088
rect 10478 4052 10530 4054
rect 10787 4160 10839 4170
rect 10787 4126 10799 4160
rect 10799 4126 10833 4160
rect 10833 4126 10839 4160
rect 10787 4118 10839 4126
rect 10787 4088 10839 4104
rect 10787 4054 10799 4088
rect 10799 4054 10833 4088
rect 10833 4054 10839 4088
rect 10787 4052 10839 4054
rect 10867 4127 10919 4179
rect 10867 4061 10919 4113
rect 11184 4757 11236 4809
rect 11184 4671 11236 4723
rect 11103 3910 11111 3921
rect 11111 3910 11145 3921
rect 11145 3910 11155 3921
rect 11103 3872 11155 3910
rect 11103 3869 11111 3872
rect 11111 3869 11145 3872
rect 11145 3869 11155 3872
rect 11103 3838 11111 3855
rect 11111 3838 11145 3855
rect 11145 3838 11155 3855
rect 11103 3803 11155 3838
rect 8646 3650 8657 3667
rect 8657 3650 8691 3667
rect 8691 3650 8698 3667
rect 8646 3615 8698 3650
rect 9019 3617 9071 3669
rect 9083 3617 9135 3669
rect 9192 3617 9244 3669
rect 9256 3617 9308 3669
rect 9648 3617 9700 3669
rect 9712 3617 9764 3669
rect 10077 3612 10129 3664
rect 10141 3612 10193 3664
rect 8646 3551 8698 3603
rect 9731 3509 9783 3518
rect 9799 3509 9851 3518
rect 9731 3475 9753 3509
rect 9753 3475 9783 3509
rect 9799 3475 9825 3509
rect 9825 3475 9851 3509
rect 10723 3504 10775 3556
rect 10787 3504 10839 3556
rect 11515 4824 11567 4876
rect 11580 4824 11632 4876
rect 11644 4824 11696 4876
rect 11290 4806 11298 4807
rect 11298 4806 11332 4807
rect 11332 4806 11342 4807
rect 11290 4766 11342 4806
rect 11290 4755 11298 4766
rect 11298 4755 11332 4766
rect 11332 4755 11342 4766
rect 11515 4730 11567 4782
rect 11580 4730 11632 4782
rect 11644 4730 11696 4782
rect 19755 4827 19807 4878
rect 19819 4878 19829 4879
rect 19829 4878 19863 4879
rect 19863 4878 19871 4879
rect 19819 4827 19871 4878
rect 19883 4878 19901 4879
rect 19901 4878 19935 4879
rect 19883 4827 19935 4878
rect 19947 4840 19999 4879
rect 19947 4827 19973 4840
rect 19973 4827 19999 4840
rect 11290 4692 11342 4721
rect 11290 4669 11298 4692
rect 11298 4669 11332 4692
rect 11332 4669 11342 4692
rect 19755 4736 19807 4788
rect 19819 4736 19871 4788
rect 19883 4736 19935 4788
rect 19947 4767 19999 4788
rect 19947 4736 19973 4767
rect 19973 4736 19999 4767
rect 11671 4593 11723 4645
rect 11735 4593 11787 4645
rect 17057 4590 17109 4642
rect 17121 4590 17173 4642
rect 17529 4620 17581 4672
rect 17593 4620 17645 4672
rect 19964 4660 19973 4686
rect 19973 4660 20007 4686
rect 20007 4660 20016 4686
rect 14443 4516 14495 4568
rect 14507 4516 14559 4568
rect 18726 4601 18778 4653
rect 18790 4601 18842 4653
rect 19964 4634 20016 4660
rect 19964 4587 19973 4621
rect 19973 4587 20007 4621
rect 20007 4587 20016 4621
rect 9731 3466 9783 3475
rect 9799 3466 9851 3475
rect 9350 3389 9402 3441
rect 9414 3389 9466 3441
rect 11097 3412 11149 3464
rect 11161 3412 11213 3464
rect 8470 2988 8522 3008
rect 8470 2956 8482 2988
rect 8482 2956 8516 2988
rect 8516 2956 8522 2988
rect 8470 2914 8522 2944
rect 8470 2892 8482 2914
rect 8482 2892 8516 2914
rect 8516 2892 8522 2914
rect 863 2623 915 2675
rect 8348 2677 8400 2729
rect 1734 2594 1786 2646
rect 1734 2530 1786 2582
rect 454 2441 506 2450
rect 454 2407 466 2441
rect 466 2407 500 2441
rect 500 2407 506 2441
rect 454 2398 506 2407
rect 1334 2433 1386 2436
rect 1334 2399 1362 2433
rect 1362 2399 1386 2433
rect 454 2369 506 2370
rect 454 2335 466 2369
rect 466 2335 500 2369
rect 500 2335 506 2369
rect 454 2318 506 2335
rect 1334 2384 1386 2399
rect 1334 2320 1386 2372
rect 454 2263 466 2290
rect 466 2263 500 2290
rect 500 2263 506 2290
rect 1487 2306 1539 2358
rect 454 2238 506 2263
rect 1487 2277 1539 2294
rect 1487 2243 1506 2277
rect 1506 2243 1539 2277
rect 1487 2242 1539 2243
rect 1616 2222 1668 2274
rect 454 2191 466 2210
rect 466 2191 500 2210
rect 500 2191 506 2210
rect 454 2158 506 2191
rect 454 2119 466 2130
rect 466 2119 500 2130
rect 500 2119 506 2130
rect 1616 2158 1668 2210
rect 454 2081 506 2119
rect 454 2078 466 2081
rect 466 2078 500 2081
rect 500 2078 506 2081
rect 1664 2070 1716 2122
rect 1728 2070 1780 2122
rect 454 2047 466 2050
rect 466 2047 500 2050
rect 500 2047 506 2050
rect 454 2009 506 2047
rect 454 1998 466 2009
rect 466 1998 500 2009
rect 500 1998 506 2009
rect 454 1937 506 1970
rect 454 1918 466 1937
rect 466 1918 500 1937
rect 500 1918 506 1937
rect 454 1865 506 1890
rect 454 1838 466 1865
rect 466 1838 500 1865
rect 500 1838 506 1865
rect 454 1793 506 1810
rect 1283 1841 1335 1850
rect 1283 1807 1290 1841
rect 1290 1807 1324 1841
rect 1324 1807 1335 1841
rect 1283 1798 1335 1807
rect 1347 1841 1399 1850
rect 1347 1807 1362 1841
rect 1362 1807 1396 1841
rect 1396 1807 1399 1841
rect 1347 1798 1399 1807
rect 454 1759 466 1793
rect 466 1759 500 1793
rect 500 1759 506 1793
rect 454 1758 506 1759
rect 454 1721 506 1730
rect 1108 1764 1160 1773
rect 1108 1730 1114 1764
rect 1114 1730 1148 1764
rect 1148 1730 1160 1764
rect 1108 1721 1160 1730
rect 1174 1764 1226 1773
rect 1174 1730 1186 1764
rect 1186 1730 1220 1764
rect 1220 1730 1226 1764
rect 1174 1721 1226 1730
rect 454 1687 466 1721
rect 466 1687 500 1721
rect 500 1687 506 1721
rect 454 1678 506 1687
rect 454 1649 506 1650
rect 454 1615 466 1649
rect 466 1615 500 1649
rect 500 1615 506 1649
rect 1610 1677 1662 1729
rect 454 1598 506 1615
rect 454 1543 466 1570
rect 466 1543 500 1570
rect 500 1543 506 1570
rect 1108 1607 1160 1615
rect 1108 1573 1114 1607
rect 1114 1573 1148 1607
rect 1148 1573 1160 1607
rect 1108 1563 1160 1573
rect 1174 1607 1226 1615
rect 1174 1573 1186 1607
rect 1186 1573 1220 1607
rect 1220 1573 1226 1607
rect 1174 1563 1226 1573
rect 1610 1613 1662 1665
rect 454 1518 506 1543
rect 454 1471 466 1490
rect 466 1471 500 1490
rect 500 1471 506 1490
rect 1283 1529 1335 1538
rect 1283 1495 1290 1529
rect 1290 1495 1324 1529
rect 1324 1495 1335 1529
rect 1283 1486 1335 1495
rect 1347 1529 1399 1538
rect 1347 1495 1362 1529
rect 1362 1495 1396 1529
rect 1396 1495 1399 1529
rect 1347 1486 1399 1495
rect 454 1438 506 1471
rect 454 1399 466 1410
rect 466 1399 500 1410
rect 500 1399 506 1410
rect 454 1361 506 1399
rect 1734 1404 1786 1456
rect 454 1358 466 1361
rect 466 1358 500 1361
rect 500 1358 506 1361
rect 454 1327 466 1330
rect 466 1327 500 1330
rect 500 1327 506 1330
rect 454 1289 506 1327
rect 1734 1325 1786 1377
rect 1821 2594 1873 2646
rect 1821 2530 1873 2582
rect 1821 2222 1873 2274
rect 1821 2158 1873 2210
rect 454 1278 466 1289
rect 466 1278 500 1289
rect 500 1278 506 1289
rect 454 1217 506 1250
rect 1262 1279 1314 1291
rect 1326 1279 1378 1291
rect 1262 1245 1290 1279
rect 1290 1245 1314 1279
rect 1326 1245 1362 1279
rect 1362 1245 1378 1279
rect 1901 2594 1953 2646
rect 1901 2530 1953 2582
rect 1901 1677 1953 1729
rect 1901 1608 1953 1660
rect 1901 1539 1953 1591
rect 1901 1470 1953 1522
rect 1901 1400 1953 1452
rect 1262 1239 1314 1245
rect 1326 1239 1378 1245
rect 8093 2613 8145 2665
rect 8157 2613 8209 2665
rect 8348 2613 8400 2665
rect 454 1198 466 1217
rect 466 1198 500 1217
rect 500 1198 506 1217
rect 454 1145 506 1170
rect 454 1118 466 1145
rect 466 1118 500 1145
rect 500 1118 506 1145
rect 454 1073 506 1090
rect 781 1123 833 1167
rect 781 1115 786 1123
rect 786 1115 820 1123
rect 820 1115 833 1123
rect 781 1089 786 1097
rect 786 1089 820 1097
rect 820 1089 833 1097
rect 454 1039 466 1073
rect 466 1039 500 1073
rect 500 1039 506 1073
rect 781 1045 833 1089
rect 454 1038 506 1039
rect 454 1001 506 1010
rect 454 967 466 1001
rect 466 967 500 1001
rect 500 967 506 1001
rect 454 958 506 967
rect 454 929 506 930
rect 1262 967 1314 976
rect 1326 967 1378 976
rect 1262 933 1290 967
rect 1290 933 1314 967
rect 1326 933 1362 967
rect 1362 933 1378 967
rect 454 895 466 929
rect 466 895 500 929
rect 500 895 506 929
rect 1262 924 1314 933
rect 1326 924 1378 933
rect 454 878 506 895
rect 454 823 466 850
rect 466 823 500 850
rect 500 823 506 850
rect 454 798 506 823
rect 1174 777 1180 811
rect 1180 777 1218 811
rect 1218 777 1226 811
rect 454 751 466 770
rect 466 751 500 770
rect 500 751 506 770
rect 454 718 506 751
rect 1174 759 1226 777
rect 454 679 466 690
rect 466 679 500 690
rect 500 679 506 690
rect 454 641 506 679
rect 454 638 466 641
rect 466 638 500 641
rect 500 638 506 641
rect 699 655 751 699
rect 1174 695 1226 747
rect 699 647 714 655
rect 714 647 748 655
rect 748 647 751 655
rect 699 621 714 629
rect 714 621 748 629
rect 748 621 751 629
rect 454 607 466 610
rect 466 607 500 610
rect 500 607 506 610
rect 454 569 506 607
rect 699 577 751 621
rect 454 558 466 569
rect 466 558 500 569
rect 500 558 506 569
rect 454 497 506 530
rect 1174 529 1226 581
rect 454 478 466 497
rect 466 478 500 497
rect 500 478 506 497
rect 1174 499 1226 517
rect 1174 465 1180 499
rect 1180 465 1218 499
rect 1218 465 1226 499
rect 454 425 506 450
rect 454 398 466 425
rect 466 398 500 425
rect 500 398 506 425
rect 454 353 506 370
rect 454 319 466 353
rect 466 319 500 353
rect 500 319 506 353
rect 454 318 506 319
rect 707 343 759 352
rect 707 309 714 343
rect 714 309 748 343
rect 748 309 759 343
rect 707 300 759 309
rect 771 343 823 352
rect 771 309 786 343
rect 786 309 820 343
rect 820 309 823 343
rect 771 300 823 309
rect 454 281 506 290
rect 454 247 466 281
rect 466 247 500 281
rect 500 247 506 281
rect 454 238 506 247
rect 454 209 506 210
rect 454 175 466 209
rect 466 175 500 209
rect 500 175 506 209
rect 454 158 506 175
rect 617 187 669 230
rect 617 178 642 187
rect 642 178 669 187
rect 617 153 642 160
rect 642 153 669 160
rect 454 103 466 130
rect 466 103 500 130
rect 500 103 506 130
rect 454 78 506 103
rect 617 108 669 153
rect 454 31 466 50
rect 466 31 500 50
rect 500 31 506 50
rect 454 -2 506 31
rect 707 31 759 40
rect 707 -3 714 31
rect 714 -3 748 31
rect 748 -3 759 31
rect 707 -12 759 -3
rect 771 31 823 40
rect 771 -3 786 31
rect 786 -3 820 31
rect 820 -3 823 31
rect 771 -12 823 -3
rect 454 -41 466 -30
rect 466 -41 500 -30
rect 500 -41 506 -30
rect 454 -79 506 -41
rect 454 -82 466 -79
rect 466 -82 500 -79
rect 500 -82 506 -79
rect 454 -113 466 -110
rect 466 -113 500 -110
rect 500 -113 506 -110
rect 454 -151 506 -113
rect 454 -162 466 -151
rect 466 -162 500 -151
rect 500 -162 506 -151
rect 693 -159 714 -125
rect 714 -159 745 -125
rect 693 -177 745 -159
rect 454 -223 506 -190
rect 454 -242 466 -223
rect 466 -242 500 -223
rect 500 -242 506 -223
rect 454 -295 506 -270
rect 454 -322 466 -295
rect 466 -322 500 -295
rect 500 -322 506 -295
rect 454 -368 506 -350
rect 535 -281 587 -237
rect 693 -241 745 -189
rect 535 -289 570 -281
rect 570 -289 587 -281
rect 535 -315 570 -307
rect 570 -315 587 -307
rect 535 -359 587 -315
rect 454 -402 466 -368
rect 466 -402 500 -368
rect 500 -402 506 -368
rect 693 -410 745 -358
rect 1866 160 1918 212
rect 1866 92 1918 144
rect 1866 24 1918 76
rect 6269 2533 6321 2585
rect 6349 2533 6401 2585
rect 6455 2533 6507 2585
rect 6519 2533 6571 2585
rect 7303 2533 7355 2585
rect 7367 2533 7419 2585
rect 7664 2533 7716 2585
rect 7728 2533 7780 2585
rect 8096 2499 8148 2508
rect 2065 169 2117 221
rect 2065 105 2117 157
rect 8096 2465 8112 2499
rect 8112 2465 8146 2499
rect 8146 2465 8148 2499
rect 8096 2456 8148 2465
rect 8160 2499 8212 2508
rect 8160 2465 8184 2499
rect 8184 2465 8212 2499
rect 8160 2456 8212 2465
rect 1866 -44 1918 8
rect 1866 -112 1918 -60
rect 1866 -180 1918 -128
rect 1866 -248 1918 -196
rect 1866 -317 1918 -265
rect 1866 -386 1918 -334
rect 1948 -105 2000 -53
rect 1948 -169 2000 -117
rect 454 -441 506 -430
rect 454 -475 466 -441
rect 466 -475 500 -441
rect 500 -475 506 -441
rect 693 -437 745 -422
rect 693 -471 714 -437
rect 714 -471 745 -437
rect 693 -474 745 -471
rect 454 -482 506 -475
rect 454 -514 506 -510
rect 454 -548 466 -514
rect 466 -548 500 -514
rect 500 -548 506 -514
rect 454 -562 506 -548
rect 454 -621 466 -590
rect 466 -621 500 -590
rect 500 -621 506 -590
rect 454 -642 506 -621
rect 1098 -627 1108 -593
rect 1108 -627 1146 -593
rect 1146 -627 1150 -593
rect 1098 -645 1150 -627
rect 454 -694 466 -670
rect 466 -694 500 -670
rect 500 -694 506 -670
rect 454 -722 506 -694
rect 937 -719 989 -667
rect 1098 -709 1150 -657
rect 454 -767 466 -750
rect 466 -767 500 -750
rect 500 -767 506 -750
rect 454 -802 506 -767
rect 454 -840 466 -830
rect 466 -840 500 -830
rect 500 -840 506 -830
rect 454 -879 506 -840
rect 617 -779 669 -727
rect 937 -749 989 -731
rect 937 -783 945 -749
rect 945 -783 986 -749
rect 986 -783 989 -749
rect 617 -843 669 -791
rect 1610 -818 1662 -766
rect 454 -882 466 -879
rect 466 -882 500 -879
rect 500 -882 506 -879
rect 454 -913 466 -910
rect 466 -913 500 -910
rect 500 -913 506 -910
rect 454 -952 506 -913
rect 1610 -882 1662 -830
rect 454 -962 466 -952
rect 466 -962 500 -952
rect 500 -962 506 -952
rect 454 -1025 506 -990
rect 541 -1009 593 -957
rect 605 -1009 657 -957
rect 1628 -993 1680 -941
rect 454 -1042 466 -1025
rect 466 -1042 500 -1025
rect 500 -1042 506 -1025
rect 454 -1098 506 -1070
rect 1343 -1034 1395 -1024
rect 1343 -1068 1377 -1034
rect 1377 -1068 1395 -1034
rect 1343 -1076 1395 -1068
rect 1415 -1034 1467 -1024
rect 1415 -1068 1423 -1034
rect 1423 -1068 1457 -1034
rect 1457 -1068 1467 -1034
rect 1415 -1076 1467 -1068
rect 1487 -1034 1539 -1024
rect 1487 -1068 1503 -1034
rect 1503 -1068 1537 -1034
rect 1537 -1068 1539 -1034
rect 1487 -1076 1539 -1068
rect 1628 -1057 1680 -1005
rect 454 -1122 466 -1098
rect 466 -1122 500 -1098
rect 500 -1122 506 -1098
rect 454 -1171 506 -1150
rect 947 -1156 999 -1104
rect 1011 -1156 1063 -1104
rect 454 -1202 466 -1171
rect 466 -1202 500 -1171
rect 500 -1202 506 -1171
rect 1256 -1224 1290 -1190
rect 1290 -1224 1308 -1190
rect 454 -1244 506 -1230
rect 454 -1278 466 -1244
rect 466 -1278 500 -1244
rect 500 -1278 506 -1244
rect 1256 -1242 1308 -1224
rect 454 -1282 506 -1278
rect 454 -1317 506 -1310
rect 1256 -1306 1308 -1254
rect 454 -1351 466 -1317
rect 466 -1351 500 -1317
rect 500 -1351 506 -1317
rect 454 -1362 506 -1351
rect 1343 -1346 1395 -1337
rect 1415 -1346 1467 -1337
rect 1487 -1346 1539 -1337
rect 1343 -1380 1362 -1346
rect 1362 -1380 1395 -1346
rect 1415 -1380 1434 -1346
rect 1434 -1380 1467 -1346
rect 1487 -1380 1506 -1346
rect 1506 -1380 1539 -1346
rect 1343 -1389 1395 -1380
rect 1415 -1389 1467 -1380
rect 1487 -1389 1539 -1380
rect 1609 -1371 1661 -1319
rect 454 -1424 466 -1390
rect 466 -1424 500 -1390
rect 500 -1424 506 -1390
rect 454 -1442 506 -1424
rect 956 -1468 1008 -1416
rect 1035 -1468 1087 -1416
rect 1609 -1450 1661 -1398
rect 454 -1497 466 -1470
rect 466 -1497 500 -1470
rect 500 -1497 506 -1470
rect 454 -1522 506 -1497
rect 1141 -1502 1193 -1490
rect 1141 -1536 1146 -1502
rect 1146 -1536 1180 -1502
rect 1180 -1536 1193 -1502
rect 1141 -1542 1193 -1536
rect 1205 -1502 1257 -1490
rect 1205 -1536 1218 -1502
rect 1218 -1536 1252 -1502
rect 1252 -1536 1257 -1502
rect 1205 -1542 1257 -1536
rect 1613 -1507 1665 -1501
rect 1613 -1541 1622 -1507
rect 1622 -1541 1656 -1507
rect 1656 -1541 1665 -1507
rect 454 -1570 466 -1550
rect 466 -1570 500 -1550
rect 500 -1570 506 -1550
rect 454 -1602 506 -1570
rect 454 -1643 466 -1630
rect 466 -1643 500 -1630
rect 500 -1643 506 -1630
rect 1613 -1553 1665 -1541
rect 1613 -1592 1665 -1580
rect 1613 -1626 1622 -1592
rect 1622 -1626 1656 -1592
rect 1656 -1626 1665 -1592
rect 1613 -1632 1665 -1626
rect 454 -1682 506 -1643
rect 1343 -1658 1395 -1646
rect 1415 -1658 1467 -1646
rect 1487 -1658 1539 -1646
rect 1343 -1692 1362 -1658
rect 1362 -1692 1395 -1658
rect 1415 -1692 1434 -1658
rect 1434 -1692 1467 -1658
rect 1487 -1692 1506 -1658
rect 1506 -1692 1539 -1658
rect 1343 -1698 1395 -1692
rect 1415 -1698 1467 -1692
rect 1487 -1698 1539 -1692
rect 454 -1716 466 -1710
rect 466 -1716 500 -1710
rect 500 -1716 506 -1710
rect 454 -1755 506 -1716
rect 454 -1762 466 -1755
rect 466 -1762 500 -1755
rect 500 -1762 506 -1755
rect 454 -1828 506 -1790
rect 454 -1842 466 -1828
rect 466 -1842 500 -1828
rect 500 -1842 506 -1828
rect 777 -1814 829 -1769
rect 777 -1821 786 -1814
rect 786 -1821 820 -1814
rect 820 -1821 829 -1814
rect 777 -1848 786 -1833
rect 786 -1848 820 -1833
rect 820 -1848 829 -1833
rect 1501 -1848 1506 -1814
rect 1506 -1848 1540 -1814
rect 1540 -1848 1553 -1814
rect 454 -1901 506 -1870
rect 777 -1885 829 -1848
rect 1501 -1866 1553 -1848
rect 454 -1922 466 -1901
rect 466 -1922 500 -1901
rect 500 -1922 506 -1901
rect 1501 -1930 1553 -1878
rect 1779 -853 1831 -801
rect 1779 -917 1831 -865
rect 454 -1974 506 -1950
rect 454 -2002 466 -1974
rect 466 -2002 500 -1974
rect 500 -2002 506 -1974
rect 1117 -1970 1169 -1958
rect 1189 -1970 1241 -1958
rect 1261 -1970 1313 -1958
rect 1117 -2004 1146 -1970
rect 1146 -2004 1169 -1970
rect 1189 -2004 1218 -1970
rect 1218 -2004 1241 -1970
rect 1261 -2004 1290 -1970
rect 1290 -2004 1313 -1970
rect 1117 -2010 1169 -2004
rect 1189 -2010 1241 -2004
rect 1261 -2010 1313 -2004
rect 454 -2047 506 -2031
rect 454 -2081 466 -2047
rect 466 -2081 500 -2047
rect 500 -2081 506 -2047
rect 454 -2083 506 -2081
rect 454 -2120 506 -2112
rect 454 -2154 466 -2120
rect 466 -2154 500 -2120
rect 500 -2154 506 -2120
rect 454 -2164 506 -2154
rect 693 -2126 745 -2085
rect 865 -2092 917 -2040
rect 929 -2092 981 -2040
rect 693 -2137 718 -2126
rect 718 -2137 745 -2126
rect 693 -2160 718 -2149
rect 718 -2160 745 -2149
rect 693 -2201 745 -2160
rect 1110 -2202 1162 -2150
rect 1185 -2202 1237 -2150
rect 1260 -2202 1312 -2150
rect 1860 -948 1912 -896
rect 1860 -1012 1912 -960
rect 395 -3462 447 -3432
rect 395 -3484 407 -3462
rect 407 -3484 441 -3462
rect 441 -3484 447 -3462
rect 395 -3535 447 -3496
rect 395 -3548 407 -3535
rect 407 -3548 441 -3535
rect 441 -3548 447 -3535
rect 398 -4265 450 -4233
rect 398 -4285 407 -4265
rect 407 -4285 441 -4265
rect 441 -4285 450 -4265
rect 398 -4338 450 -4299
rect 398 -4351 407 -4338
rect 407 -4351 441 -4338
rect 441 -4351 450 -4338
rect 398 -4372 407 -4365
rect 407 -4372 441 -4365
rect 441 -4372 450 -4365
rect 398 -4411 450 -4372
rect 398 -4417 407 -4411
rect 407 -4417 441 -4411
rect 441 -4417 450 -4411
rect 1949 -1039 2001 -987
rect 1949 -1103 2001 -1051
rect 2221 -105 2273 -53
rect 2221 -169 2273 -117
rect 7465 2256 7517 2308
rect 7529 2256 7581 2308
rect 4392 2231 4444 2241
rect 4476 2231 4528 2241
rect 4560 2231 4612 2241
rect 4644 2231 4696 2241
rect 4392 2197 4413 2231
rect 4413 2197 4444 2231
rect 4476 2197 4486 2231
rect 4486 2197 4525 2231
rect 4525 2197 4528 2231
rect 4560 2197 4598 2231
rect 4598 2197 4612 2231
rect 4644 2197 4671 2231
rect 4671 2197 4696 2231
rect 4392 2189 4444 2197
rect 4476 2189 4528 2197
rect 4560 2189 4612 2197
rect 4644 2189 4696 2197
rect 7147 2188 7199 2240
rect 7211 2188 7263 2240
rect 7664 2237 7716 2246
rect 7664 2203 7667 2237
rect 7667 2203 7701 2237
rect 7701 2203 7716 2237
rect 7664 2194 7716 2203
rect 7728 2237 7780 2246
rect 8601 2245 8653 2272
rect 7728 2203 7744 2237
rect 7744 2203 7778 2237
rect 7778 2203 7780 2237
rect 7728 2194 7780 2203
rect 3044 2137 3096 2145
rect 3115 2137 3167 2145
rect 3186 2137 3238 2145
rect 3256 2137 3308 2145
rect 3044 2103 3068 2137
rect 3068 2103 3096 2137
rect 3115 2103 3140 2137
rect 3140 2103 3167 2137
rect 3186 2103 3212 2137
rect 3212 2103 3238 2137
rect 3256 2103 3284 2137
rect 3284 2103 3308 2137
rect 3044 2093 3096 2103
rect 3115 2093 3167 2103
rect 3186 2093 3238 2103
rect 3256 2093 3308 2103
rect 6054 2137 6106 2146
rect 6054 2103 6056 2137
rect 6056 2103 6090 2137
rect 6090 2103 6106 2137
rect 6054 2094 6106 2103
rect 6118 2137 6170 2146
rect 6118 2103 6128 2137
rect 6128 2103 6162 2137
rect 6162 2103 6170 2137
rect 6118 2094 6170 2103
rect 4463 2082 4515 2088
rect 4463 2048 4472 2082
rect 4472 2048 4506 2082
rect 4506 2048 4515 2082
rect 4463 2036 4515 2048
rect 4463 2005 4515 2022
rect 4463 1971 4472 2005
rect 4472 1971 4506 2005
rect 4506 1971 4515 2005
rect 4463 1970 4515 1971
rect 4463 1928 4515 1955
rect 2422 1901 2474 1910
rect 2493 1901 2545 1910
rect 2422 1867 2454 1901
rect 2454 1867 2474 1901
rect 2493 1867 2526 1901
rect 2526 1867 2545 1901
rect 2422 1858 2474 1867
rect 2493 1858 2545 1867
rect 2564 1901 2616 1910
rect 2564 1867 2598 1901
rect 2598 1867 2616 1901
rect 2564 1858 2616 1867
rect 2634 1901 2686 1910
rect 3869 1901 3921 1910
rect 3940 1901 3992 1910
rect 4011 1901 4063 1910
rect 4081 1901 4133 1910
rect 2634 1867 2636 1901
rect 2636 1867 2670 1901
rect 2670 1867 2686 1901
rect 3869 1867 3894 1901
rect 3894 1867 3921 1901
rect 3940 1867 3966 1901
rect 3966 1867 3992 1901
rect 4011 1867 4038 1901
rect 4038 1867 4063 1901
rect 4081 1867 4110 1901
rect 4110 1867 4133 1901
rect 2634 1858 2686 1867
rect 3869 1858 3921 1867
rect 3940 1858 3992 1867
rect 4011 1858 4063 1867
rect 4081 1858 4133 1867
rect 4463 1903 4472 1928
rect 4472 1903 4506 1928
rect 4506 1903 4515 1928
rect 4463 1851 4515 1888
rect 4463 1836 4472 1851
rect 4472 1836 4506 1851
rect 4506 1836 4515 1851
rect 4463 1817 4472 1821
rect 4472 1817 4506 1821
rect 4506 1817 4515 1821
rect 4463 1774 4515 1817
rect 4463 1769 4472 1774
rect 4472 1769 4506 1774
rect 4506 1769 4515 1774
rect 4463 1740 4472 1754
rect 4472 1740 4506 1754
rect 4506 1740 4515 1754
rect 4463 1702 4515 1740
rect 3044 1665 3096 1674
rect 3115 1665 3167 1674
rect 3186 1665 3238 1674
rect 3256 1665 3308 1674
rect 3044 1631 3068 1665
rect 3068 1631 3096 1665
rect 3115 1631 3140 1665
rect 3140 1631 3167 1665
rect 3186 1631 3212 1665
rect 3212 1631 3238 1665
rect 3256 1631 3284 1665
rect 3284 1631 3308 1665
rect 3044 1622 3096 1631
rect 3115 1622 3167 1631
rect 3186 1622 3238 1631
rect 3256 1622 3308 1631
rect 4463 1663 4472 1687
rect 4472 1663 4506 1687
rect 4506 1663 4515 1687
rect 4568 2077 4620 2088
rect 8601 2220 8613 2245
rect 8613 2220 8647 2245
rect 8647 2220 8653 2245
rect 8601 2173 8653 2208
rect 8601 2156 8613 2173
rect 8613 2156 8647 2173
rect 8647 2156 8653 2173
rect 4568 2043 4580 2077
rect 4580 2043 4614 2077
rect 4614 2043 4620 2077
rect 4568 2036 4620 2043
rect 4568 1989 4620 2018
rect 4568 1966 4580 1989
rect 4580 1966 4614 1989
rect 4614 1966 4620 1989
rect 4568 1900 4620 1947
rect 4568 1895 4580 1900
rect 4580 1895 4614 1900
rect 4614 1895 4620 1900
rect 4568 1866 4580 1876
rect 4580 1866 4614 1876
rect 4614 1866 4620 1876
rect 4568 1824 4620 1866
rect 6659 1901 6711 1910
rect 6659 1867 6666 1901
rect 6666 1867 6711 1901
rect 6659 1858 6711 1867
rect 6723 1858 6775 1910
rect 4568 1777 4580 1805
rect 4580 1777 4614 1805
rect 4614 1777 4620 1805
rect 4568 1753 4620 1777
rect 4568 1722 4620 1734
rect 4568 1688 4580 1722
rect 4580 1688 4614 1722
rect 4614 1688 4620 1722
rect 4568 1682 4620 1688
rect 4463 1635 4515 1663
rect 6054 1665 6106 1674
rect 6054 1631 6056 1665
rect 6056 1631 6090 1665
rect 6090 1631 6106 1665
rect 6054 1622 6106 1631
rect 6118 1665 6170 1674
rect 6118 1631 6128 1665
rect 6128 1631 6162 1665
rect 6162 1631 6170 1665
rect 6118 1622 6170 1631
rect 7303 1919 7355 1971
rect 7367 1919 7419 1971
rect 8143 1919 8195 1971
rect 8207 1919 8259 1971
rect 7896 1823 7948 1835
rect 7977 1823 8029 1835
rect 7896 1789 7910 1823
rect 7910 1789 7948 1823
rect 7977 1789 7985 1823
rect 7985 1789 8026 1823
rect 8026 1789 8029 1823
rect 7896 1783 7948 1789
rect 7977 1783 8029 1789
rect 7007 1663 7059 1715
rect 7105 1663 7157 1715
rect 7202 1663 7254 1715
rect 8598 1722 8650 1774
rect 8598 1658 8650 1710
rect 9572 3197 9624 3209
rect 9640 3197 9692 3209
rect 10797 3214 10849 3220
rect 10869 3214 10921 3220
rect 10941 3214 10993 3220
rect 11012 3214 11064 3220
rect 11083 3214 11135 3220
rect 9572 3163 9609 3197
rect 9609 3163 9624 3197
rect 9640 3163 9643 3197
rect 9643 3163 9681 3197
rect 9681 3163 9692 3197
rect 9572 3157 9624 3163
rect 9640 3157 9692 3163
rect 8881 3075 8933 3127
rect 8945 3075 8997 3127
rect 9893 3075 9945 3127
rect 9957 3075 10009 3127
rect 10797 3180 10834 3214
rect 10834 3180 10849 3214
rect 10869 3180 10906 3214
rect 10906 3180 10921 3214
rect 10941 3180 10978 3214
rect 10978 3180 10993 3214
rect 11012 3180 11050 3214
rect 11050 3180 11064 3214
rect 11083 3180 11084 3214
rect 11084 3180 11122 3214
rect 11122 3180 11135 3214
rect 10797 3168 10849 3180
rect 10869 3168 10921 3180
rect 10941 3168 10993 3180
rect 11012 3168 11064 3180
rect 11083 3168 11135 3180
rect 10070 3055 10122 3107
rect 10134 3055 10186 3107
rect 11591 4439 11643 4491
rect 11656 4439 11708 4491
rect 19964 4569 20016 4587
rect 19964 4548 20016 4556
rect 19964 4514 19973 4548
rect 19973 4514 20007 4548
rect 20007 4514 20016 4548
rect 19964 4504 20016 4514
rect 19964 4475 20016 4491
rect 19964 4441 19973 4475
rect 19973 4441 20007 4475
rect 20007 4441 20016 4475
rect 19964 4439 20016 4441
rect 11636 4359 11688 4411
rect 11700 4359 11752 4411
rect 19964 4402 20016 4426
rect 19964 4374 19973 4402
rect 19973 4374 20007 4402
rect 20007 4374 20016 4402
rect 19964 4329 20016 4361
rect 19964 4309 19973 4329
rect 19973 4309 20007 4329
rect 20007 4309 20016 4329
rect 19964 4295 19973 4296
rect 19973 4295 20007 4296
rect 20007 4295 20016 4296
rect 13247 4254 13299 4263
rect 13247 4220 13250 4254
rect 13250 4220 13284 4254
rect 13284 4220 13299 4254
rect 13247 4211 13299 4220
rect 13311 4254 13363 4263
rect 13311 4220 13322 4254
rect 13322 4220 13356 4254
rect 13356 4220 13363 4254
rect 13311 4211 13363 4220
rect 19964 4256 20016 4295
rect 19964 4244 19973 4256
rect 19973 4244 20007 4256
rect 20007 4244 20016 4256
rect 19964 4222 19973 4231
rect 19973 4222 20007 4231
rect 20007 4222 20016 4231
rect 12394 4123 12400 4151
rect 12400 4123 12434 4151
rect 12434 4123 12446 4151
rect 12394 4099 12446 4123
rect 12460 4123 12472 4151
rect 12472 4123 12506 4151
rect 12506 4123 12512 4151
rect 12460 4099 12512 4123
rect 13083 4114 13135 4120
rect 13083 4080 13089 4114
rect 13089 4080 13123 4114
rect 13123 4080 13135 4114
rect 13083 4068 13135 4080
rect 13147 4114 13199 4120
rect 13147 4080 13161 4114
rect 13161 4080 13195 4114
rect 13195 4080 13199 4114
rect 13147 4068 13199 4080
rect 16316 4121 16368 4127
rect 16316 4087 16317 4121
rect 16317 4087 16351 4121
rect 16351 4087 16368 4121
rect 16316 4075 16368 4087
rect 16380 4121 16432 4127
rect 16380 4087 16389 4121
rect 16389 4087 16423 4121
rect 16423 4087 16432 4121
rect 16380 4075 16432 4087
rect 16837 4115 16889 4121
rect 16837 4081 16843 4115
rect 16843 4081 16877 4115
rect 16877 4081 16889 4115
rect 16837 4069 16889 4081
rect 16996 4119 17048 4129
rect 16996 4085 17015 4119
rect 17015 4085 17048 4119
rect 16996 4077 17048 4085
rect 17062 4077 17114 4129
rect 12442 4058 12494 4067
rect 12442 4024 12448 4058
rect 12448 4024 12482 4058
rect 12482 4024 12494 4058
rect 12442 4015 12494 4024
rect 12506 4058 12558 4067
rect 12506 4024 12520 4058
rect 12520 4024 12554 4058
rect 12554 4024 12558 4058
rect 12506 4015 12558 4024
rect 16837 4043 16889 4055
rect 16837 4009 16843 4043
rect 16843 4009 16877 4043
rect 16877 4009 16889 4043
rect 16837 4003 16889 4009
rect 17675 4010 17727 4062
rect 17765 4073 17817 4082
rect 17765 4039 17779 4073
rect 17779 4039 17813 4073
rect 17813 4039 17817 4073
rect 17765 4030 17817 4039
rect 17839 4073 17891 4082
rect 17839 4039 17855 4073
rect 17855 4039 17889 4073
rect 17889 4039 17891 4073
rect 17839 4030 17891 4039
rect 17912 4073 17964 4082
rect 17912 4039 17931 4073
rect 17931 4039 17964 4073
rect 19259 4090 19311 4098
rect 19259 4056 19268 4090
rect 19268 4056 19302 4090
rect 19302 4056 19311 4090
rect 19964 4183 20016 4222
rect 19964 4179 19973 4183
rect 19973 4179 20007 4183
rect 20007 4179 20016 4183
rect 19964 4149 19973 4166
rect 19973 4149 20007 4166
rect 20007 4149 20016 4166
rect 19964 4114 20016 4149
rect 19964 4076 19973 4100
rect 19973 4076 20007 4100
rect 20007 4076 20016 4100
rect 17912 4030 17964 4039
rect 19259 4046 19311 4056
rect 19259 4018 19311 4034
rect 11638 3942 11690 3994
rect 11702 3942 11754 3994
rect 17675 3946 17727 3998
rect 18588 3961 18640 4013
rect 18652 3961 18704 4013
rect 19259 3984 19268 4018
rect 19268 3984 19302 4018
rect 19302 3984 19311 4018
rect 19259 3982 19311 3984
rect 17107 3926 17159 3932
rect 11783 3852 11835 3904
rect 11847 3852 11899 3904
rect 17107 3892 17116 3926
rect 17116 3892 17150 3926
rect 17150 3892 17159 3926
rect 19964 4048 20016 4076
rect 19964 4003 19973 4034
rect 19973 4003 20007 4034
rect 20007 4003 20016 4034
rect 19964 3982 20016 4003
rect 19964 3964 20016 3968
rect 19964 3930 19973 3964
rect 19973 3930 20007 3964
rect 20007 3930 20016 3964
rect 19964 3916 20016 3930
rect 17107 3880 17159 3892
rect 19964 3891 20016 3902
rect 17107 3854 17159 3866
rect 17107 3820 17116 3854
rect 17116 3820 17150 3854
rect 17150 3820 17159 3854
rect 18766 3836 18818 3888
rect 18833 3836 18885 3888
rect 19964 3857 19973 3891
rect 19973 3857 20007 3891
rect 20007 3857 20016 3891
rect 19964 3850 20016 3857
rect 17107 3814 17159 3820
rect 19964 3818 20016 3836
rect 19964 3784 19973 3818
rect 19973 3784 20007 3818
rect 20007 3784 20016 3818
rect 19088 3719 19140 3771
rect 19165 3719 19217 3771
rect 19242 3719 19294 3771
rect 19088 3649 19140 3701
rect 19165 3649 19217 3701
rect 19242 3649 19294 3701
rect 19088 3579 19140 3631
rect 19165 3579 19217 3631
rect 19242 3579 19294 3631
rect 19964 3745 20016 3770
rect 19964 3718 19973 3745
rect 19973 3718 20007 3745
rect 20007 3718 20016 3745
rect 19964 3672 20016 3704
rect 19964 3652 19973 3672
rect 19973 3652 20007 3672
rect 20007 3652 20016 3672
rect 19964 3599 20016 3638
rect 19964 3586 19973 3599
rect 19973 3586 20007 3599
rect 20007 3586 20016 3599
rect 19964 3565 19973 3572
rect 19973 3565 20007 3572
rect 20007 3565 20016 3572
rect 19964 3526 20016 3565
rect 19964 3520 19973 3526
rect 19973 3520 20007 3526
rect 20007 3520 20016 3526
rect 11580 3412 11632 3464
rect 11644 3412 11696 3464
rect 13083 3412 13135 3464
rect 13147 3412 13199 3464
rect 13247 3412 13299 3464
rect 13311 3412 13363 3464
rect 18767 3412 18819 3464
rect 18833 3412 18885 3464
rect 19964 3492 19973 3506
rect 19973 3492 20007 3506
rect 20007 3492 20016 3506
rect 19964 3454 20016 3492
rect 19964 3420 19973 3440
rect 19973 3420 20007 3440
rect 20007 3420 20016 3440
rect 19964 3388 20016 3420
rect 17298 3377 17350 3382
rect 17298 3343 17331 3377
rect 17331 3343 17350 3377
rect 17298 3330 17350 3343
rect 17362 3377 17414 3382
rect 17362 3343 17369 3377
rect 17369 3343 17403 3377
rect 17403 3343 17414 3377
rect 17362 3330 17414 3343
rect 8851 3002 8903 3014
rect 8851 2968 8867 3002
rect 8867 2968 8901 3002
rect 8901 2968 8903 3002
rect 8851 2962 8903 2968
rect 8915 3002 8967 3014
rect 8915 2968 8942 3002
rect 8942 2968 8967 3002
rect 17765 3248 17817 3300
rect 17839 3248 17891 3300
rect 8915 2962 8967 2968
rect 9195 2866 9247 2918
rect 9259 2866 9311 2918
rect 10775 2856 10827 2868
rect 10839 2856 10891 2868
rect 10775 2822 10805 2856
rect 10805 2822 10827 2856
rect 10839 2822 10884 2856
rect 10884 2822 10891 2856
rect 10775 2816 10827 2822
rect 10839 2816 10891 2822
rect 11477 2728 11529 2780
rect 8868 2658 8920 2710
rect 8932 2658 8984 2710
rect 11477 2664 11529 2716
rect 8865 2578 8917 2630
rect 8929 2578 8981 2630
rect 10098 2578 10150 2630
rect 10206 2578 10258 2630
rect 10314 2578 10366 2630
rect 10602 2618 10654 2630
rect 10602 2584 10613 2618
rect 10613 2584 10647 2618
rect 10647 2584 10654 2618
rect 10602 2578 10654 2584
rect 10673 2618 10725 2630
rect 10673 2584 10685 2618
rect 10685 2584 10719 2618
rect 10719 2584 10725 2618
rect 10673 2578 10725 2584
rect 16930 3166 16982 3218
rect 16994 3166 17046 3218
rect 17298 3216 17350 3222
rect 17362 3216 17414 3222
rect 17298 3182 17307 3216
rect 17307 3182 17350 3216
rect 17362 3182 17391 3216
rect 17391 3182 17414 3216
rect 17298 3170 17350 3182
rect 17362 3170 17414 3182
rect 4463 1619 4515 1620
rect 4463 1585 4472 1619
rect 4472 1585 4506 1619
rect 4506 1585 4515 1619
rect 4463 1568 4515 1585
rect 15831 3084 15883 3136
rect 15895 3084 15947 3136
rect 16316 3084 16368 3136
rect 16380 3084 16432 3136
rect 17451 3071 17503 3123
rect 4463 1541 4515 1553
rect 4463 1507 4472 1541
rect 4472 1507 4506 1541
rect 4506 1507 4515 1541
rect 4463 1501 4515 1507
rect 17037 3002 17089 3054
rect 17101 3002 17153 3054
rect 17451 3047 17503 3059
rect 17451 3013 17457 3047
rect 17457 3013 17491 3047
rect 17491 3013 17503 3047
rect 17451 3007 17503 3013
rect 17613 3096 17619 3128
rect 17619 3096 17653 3128
rect 17653 3096 17665 3128
rect 17613 3076 17665 3096
rect 17613 3012 17665 3064
rect 18104 3148 18156 3154
rect 18104 3114 18110 3148
rect 18110 3114 18144 3148
rect 18144 3114 18156 3148
rect 18104 3102 18156 3114
rect 18104 3076 18156 3088
rect 18104 3042 18110 3076
rect 18110 3042 18144 3076
rect 18144 3042 18156 3076
rect 18104 3036 18156 3042
rect 18273 3148 18325 3154
rect 18273 3114 18282 3148
rect 18282 3114 18316 3148
rect 18316 3114 18325 3148
rect 18273 3102 18325 3114
rect 18273 3076 18325 3088
rect 18273 3042 18282 3076
rect 18282 3042 18316 3076
rect 18316 3042 18325 3076
rect 18273 3036 18325 3042
rect 18583 3148 18635 3154
rect 18583 3114 18594 3148
rect 18594 3114 18628 3148
rect 18628 3114 18635 3148
rect 18583 3102 18635 3114
rect 18583 3076 18635 3088
rect 18583 3042 18594 3076
rect 18594 3042 18628 3076
rect 18628 3042 18635 3076
rect 18583 3036 18635 3042
rect 18733 3148 18785 3154
rect 18733 3114 18744 3148
rect 18744 3114 18778 3148
rect 18778 3114 18785 3148
rect 18733 3102 18785 3114
rect 18733 3076 18785 3088
rect 18733 3042 18744 3076
rect 18744 3042 18778 3076
rect 18778 3042 18785 3076
rect 18733 3036 18785 3042
rect 18821 3101 18873 3153
rect 18821 3035 18873 3087
rect 2422 1429 2474 1439
rect 2493 1429 2545 1439
rect 2422 1395 2454 1429
rect 2454 1395 2474 1429
rect 2493 1395 2526 1429
rect 2526 1395 2545 1429
rect 2422 1387 2474 1395
rect 2493 1387 2545 1395
rect 2564 1429 2616 1439
rect 2564 1395 2598 1429
rect 2598 1395 2616 1429
rect 2564 1387 2616 1395
rect 2634 1429 2686 1439
rect 3869 1429 3921 1439
rect 3940 1429 3992 1439
rect 4011 1429 4063 1439
rect 4081 1429 4133 1439
rect 2634 1395 2636 1429
rect 2636 1395 2670 1429
rect 2670 1395 2686 1429
rect 3869 1395 3894 1429
rect 3894 1395 3921 1429
rect 3940 1395 3966 1429
rect 3966 1395 3992 1429
rect 4011 1395 4038 1429
rect 4038 1395 4063 1429
rect 4081 1395 4110 1429
rect 4110 1395 4133 1429
rect 2634 1387 2686 1395
rect 3869 1387 3921 1395
rect 3940 1387 3992 1395
rect 4011 1387 4063 1395
rect 4081 1387 4133 1395
rect 4467 1321 4486 1355
rect 4486 1321 4519 1355
rect 4467 1303 4519 1321
rect 4467 1273 4519 1291
rect 4467 1239 4486 1273
rect 4486 1239 4519 1273
rect 6204 1297 6256 1349
rect 7142 1381 7194 1433
rect 7208 1381 7260 1433
rect 6204 1233 6256 1285
rect 6996 1271 7048 1323
rect 6996 1207 7048 1259
rect 3044 1193 3096 1202
rect 3115 1193 3167 1202
rect 3186 1193 3238 1202
rect 3256 1193 3308 1202
rect 3044 1159 3068 1193
rect 3068 1159 3096 1193
rect 3115 1159 3140 1193
rect 3140 1159 3167 1193
rect 3186 1159 3212 1193
rect 3212 1159 3238 1193
rect 3256 1159 3284 1193
rect 3284 1159 3308 1193
rect 3044 1150 3096 1159
rect 3115 1150 3167 1159
rect 3186 1150 3238 1159
rect 3256 1150 3308 1159
rect 6808 1153 6860 1205
rect 6872 1153 6924 1205
rect 3867 1098 3919 1117
rect 3867 1065 3876 1098
rect 3876 1065 3919 1098
rect 3931 1098 3983 1117
rect 3931 1065 3933 1098
rect 3933 1065 3967 1098
rect 3967 1065 3983 1098
rect 5518 1066 5570 1118
rect 5582 1066 5634 1118
rect 5739 1098 5791 1125
rect 5739 1073 5764 1098
rect 5764 1073 5791 1098
rect 5803 1098 5855 1125
rect 5803 1073 5807 1098
rect 5807 1073 5841 1098
rect 5841 1073 5855 1098
rect 6054 1071 6106 1123
rect 6118 1071 6170 1123
rect 2377 478 2429 515
rect 2377 463 2406 478
rect 2406 463 2429 478
rect 2441 463 2493 515
rect 3177 660 3186 668
rect 3186 660 3220 668
rect 3220 660 3229 668
rect 3177 622 3229 660
rect 3177 616 3186 622
rect 3186 616 3220 622
rect 3220 616 3229 622
rect 3177 588 3186 604
rect 3186 588 3220 604
rect 3220 588 3229 604
rect 3177 552 3229 588
rect 2718 478 2770 515
rect 2718 463 2752 478
rect 2752 463 2770 478
rect 2782 463 2834 515
rect 2994 478 3046 515
rect 3058 478 3110 515
rect 2994 463 3030 478
rect 3030 463 3046 478
rect 3058 463 3064 478
rect 3064 463 3110 478
rect 2630 260 2682 312
rect 2630 196 2682 248
rect 2553 118 2605 154
rect 2553 102 2562 118
rect 2562 102 2596 118
rect 2596 102 2605 118
rect 2553 84 2562 89
rect 2562 84 2596 89
rect 2596 84 2605 89
rect 2553 46 2605 84
rect 2553 37 2562 46
rect 2562 37 2596 46
rect 2596 37 2605 46
rect 2553 12 2562 24
rect 2562 12 2596 24
rect 2596 12 2605 24
rect 2553 -28 2605 12
rect 2865 118 2917 154
rect 2865 102 2874 118
rect 2874 102 2908 118
rect 2908 102 2917 118
rect 2865 84 2874 89
rect 2874 84 2908 89
rect 2908 84 2917 89
rect 2865 46 2917 84
rect 2865 37 2874 46
rect 2874 37 2908 46
rect 2908 37 2917 46
rect 2865 12 2874 24
rect 2874 12 2908 24
rect 2908 12 2917 24
rect 2865 -28 2917 12
rect 3489 660 3498 668
rect 3498 660 3532 668
rect 3532 660 3541 668
rect 3489 622 3541 660
rect 3489 616 3498 622
rect 3498 616 3532 622
rect 3532 616 3541 622
rect 3489 588 3498 604
rect 3498 588 3532 604
rect 3532 588 3541 604
rect 3489 552 3541 588
rect 3342 478 3394 515
rect 3342 463 3376 478
rect 3376 463 3394 478
rect 3406 463 3458 515
rect 3618 478 3670 515
rect 3682 478 3734 515
rect 3618 463 3654 478
rect 3654 463 3670 478
rect 3682 463 3688 478
rect 3688 463 3734 478
rect 3925 660 3934 668
rect 3934 660 3968 668
rect 3968 660 3977 668
rect 3925 622 3977 660
rect 3925 616 3934 622
rect 3934 616 3968 622
rect 3968 616 3977 622
rect 3925 588 3934 604
rect 3934 588 3968 604
rect 3968 588 3977 604
rect 3925 552 3977 588
rect 3254 342 3306 394
rect 3254 278 3306 330
rect 3846 424 3898 476
rect 3846 360 3898 412
rect 4004 424 4056 476
rect 4004 360 4056 412
rect 3769 118 3821 154
rect 3769 102 3778 118
rect 3778 102 3812 118
rect 3812 102 3821 118
rect 3769 84 3778 89
rect 3778 84 3812 89
rect 3812 84 3821 89
rect 3769 46 3821 84
rect 3769 37 3778 46
rect 3778 37 3812 46
rect 3812 37 3821 46
rect 3769 12 3778 24
rect 3778 12 3812 24
rect 3812 12 3821 24
rect 3769 -28 3821 12
rect 4237 948 4246 971
rect 4246 948 4280 971
rect 4280 948 4289 971
rect 4237 919 4289 948
rect 4237 876 4246 907
rect 4246 876 4280 907
rect 4280 876 4289 907
rect 4237 855 4289 876
rect 4081 118 4133 154
rect 4081 102 4090 118
rect 4090 102 4124 118
rect 4124 102 4133 118
rect 4081 84 4090 89
rect 4090 84 4124 89
rect 4124 84 4133 89
rect 4081 46 4133 84
rect 4081 37 4090 46
rect 4090 37 4124 46
rect 4124 37 4133 46
rect 4081 12 4090 24
rect 4090 12 4124 24
rect 4124 12 4133 24
rect 4081 -28 4133 12
rect 4393 118 4445 154
rect 4393 102 4402 118
rect 4402 102 4436 118
rect 4436 102 4445 118
rect 4393 84 4402 89
rect 4402 84 4436 89
rect 4436 84 4445 89
rect 4393 46 4445 84
rect 4393 37 4402 46
rect 4402 37 4436 46
rect 4436 37 4445 46
rect 4393 12 4402 24
rect 4402 12 4436 24
rect 4436 12 4445 24
rect 4393 -28 4445 12
rect 4709 478 4761 507
rect 4709 455 4714 478
rect 4714 455 4748 478
rect 4748 455 4761 478
rect 4773 455 4825 507
rect 4549 118 4601 154
rect 4549 102 4558 118
rect 4558 102 4592 118
rect 4592 102 4601 118
rect 4549 84 4558 89
rect 4558 84 4592 89
rect 4592 84 4601 89
rect 4549 46 4601 84
rect 4549 37 4558 46
rect 4558 37 4592 46
rect 4592 37 4601 46
rect 4549 12 4558 24
rect 4558 12 4592 24
rect 4592 12 4601 24
rect 4549 -28 4601 12
rect 5173 948 5182 971
rect 5182 948 5216 971
rect 5216 948 5225 971
rect 5173 919 5225 948
rect 5173 876 5182 907
rect 5182 876 5216 907
rect 5216 876 5225 907
rect 5173 855 5225 876
rect 4861 118 4913 154
rect 4861 102 4870 118
rect 4870 102 4904 118
rect 4904 102 4913 118
rect 4861 84 4870 89
rect 4870 84 4904 89
rect 4904 84 4913 89
rect 4861 46 4913 84
rect 4861 37 4870 46
rect 4870 37 4904 46
rect 4904 37 4913 46
rect 4861 12 4870 24
rect 4870 12 4904 24
rect 4904 12 4913 24
rect 4861 -28 4913 12
rect 5017 118 5069 154
rect 5017 102 5026 118
rect 5026 102 5060 118
rect 5060 102 5069 118
rect 5017 84 5026 89
rect 5026 84 5060 89
rect 5060 84 5069 89
rect 5017 46 5069 84
rect 5017 37 5026 46
rect 5026 37 5060 46
rect 5060 37 5069 46
rect 5017 12 5026 24
rect 5026 12 5060 24
rect 5060 12 5069 24
rect 5017 -28 5069 12
rect 5483 948 5494 971
rect 5494 948 5528 971
rect 5528 948 5535 971
rect 5483 919 5535 948
rect 5483 876 5494 907
rect 5494 876 5528 907
rect 5528 876 5535 907
rect 5483 855 5535 876
rect 5662 732 5668 754
rect 5668 732 5702 754
rect 5702 732 5714 754
rect 5662 702 5714 732
rect 5729 702 5781 754
rect 5567 506 5619 558
rect 5567 442 5619 494
rect 5329 118 5381 154
rect 5329 102 5338 118
rect 5338 102 5372 118
rect 5372 102 5381 118
rect 5329 84 5338 89
rect 5338 84 5372 89
rect 5372 84 5381 89
rect 5329 46 5381 84
rect 5329 37 5338 46
rect 5338 37 5372 46
rect 5372 37 5381 46
rect 5329 12 5338 24
rect 5338 12 5372 24
rect 5372 12 5381 24
rect 5329 -28 5381 12
rect 6204 1098 6256 1110
rect 6204 1064 6226 1098
rect 6226 1064 6256 1098
rect 6204 1058 6256 1064
rect 6455 1096 6507 1108
rect 6519 1096 6571 1108
rect 6455 1062 6476 1096
rect 6476 1062 6507 1096
rect 6519 1062 6550 1096
rect 6550 1062 6571 1096
rect 6455 1056 6507 1062
rect 6519 1056 6571 1062
rect 6204 994 6256 1046
rect 6285 982 6337 1016
rect 6285 964 6292 982
rect 6292 964 6326 982
rect 6326 964 6337 982
rect 6285 948 6292 952
rect 6292 948 6326 952
rect 6326 948 6337 952
rect 6285 910 6337 948
rect 6285 900 6292 910
rect 6292 900 6326 910
rect 6326 900 6337 910
rect 5902 603 5954 655
rect 5969 622 6021 655
rect 5969 603 5980 622
rect 5980 603 6014 622
rect 6014 603 6021 622
rect 6085 478 6137 490
rect 6149 478 6201 490
rect 6085 444 6136 478
rect 6136 444 6137 478
rect 6149 444 6170 478
rect 6170 444 6201 478
rect 6085 438 6137 444
rect 6149 438 6201 444
rect 5814 118 5866 154
rect 5814 102 5824 118
rect 5824 102 5858 118
rect 5858 102 5866 118
rect 5814 84 5824 89
rect 5824 84 5858 89
rect 5858 84 5866 89
rect 5814 46 5866 84
rect 5814 37 5824 46
rect 5824 37 5858 46
rect 5858 37 5866 46
rect 5814 12 5824 24
rect 5824 12 5858 24
rect 5858 12 5866 24
rect 5814 -28 5866 12
rect 6687 982 6739 1017
rect 6687 965 6696 982
rect 6696 965 6730 982
rect 6730 965 6739 982
rect 6687 948 6696 953
rect 6696 948 6730 953
rect 6730 948 6739 953
rect 6687 910 6739 948
rect 6687 901 6696 910
rect 6696 901 6730 910
rect 6730 901 6739 910
rect 6563 622 6615 647
rect 6563 595 6572 622
rect 6572 595 6606 622
rect 6606 595 6615 622
rect 6563 550 6615 583
rect 6563 531 6572 550
rect 6572 531 6606 550
rect 6606 531 6615 550
rect 6407 118 6459 154
rect 6407 102 6416 118
rect 6416 102 6450 118
rect 6450 102 6459 118
rect 6407 84 6416 89
rect 6416 84 6450 89
rect 6450 84 6459 89
rect 6407 46 6459 84
rect 6407 37 6416 46
rect 6416 37 6450 46
rect 6450 37 6459 46
rect 6407 12 6416 24
rect 6416 12 6450 24
rect 6450 12 6459 24
rect 6407 -28 6459 12
rect 6843 118 6895 154
rect 6843 102 6852 118
rect 6852 102 6886 118
rect 6886 102 6895 118
rect 6843 84 6852 89
rect 6852 84 6886 89
rect 6886 84 6895 89
rect 6843 46 6895 84
rect 6843 37 6852 46
rect 6852 37 6886 46
rect 6886 37 6895 46
rect 6843 12 6852 24
rect 6852 12 6886 24
rect 6886 12 6895 24
rect 6843 -28 6895 12
rect 7142 1312 7194 1364
rect 7208 1312 7260 1364
rect 7142 1242 7194 1294
rect 7208 1242 7260 1294
rect 7142 1172 7194 1224
rect 7208 1172 7260 1224
rect 12862 2910 12914 2962
rect 12926 2910 12978 2962
rect 16301 2909 16353 2961
rect 16365 2909 16417 2961
rect 16772 2920 16824 2972
rect 16836 2920 16888 2972
rect 17795 2930 17847 2982
rect 17859 2976 17911 2982
rect 17859 2942 17889 2976
rect 17889 2942 17911 2976
rect 17859 2930 17911 2942
rect 18953 2883 19005 2895
rect 19044 2883 19096 2895
rect 7325 595 7377 647
rect 7501 1283 7510 1293
rect 7510 1283 7544 1293
rect 7544 1283 7553 1293
rect 7501 1245 7553 1283
rect 7501 1241 7510 1245
rect 7510 1241 7544 1245
rect 7544 1241 7553 1245
rect 7501 1211 7510 1229
rect 7510 1211 7544 1229
rect 7544 1211 7553 1229
rect 7501 1177 7553 1211
rect 7325 531 7377 583
rect 7414 597 7466 604
rect 7414 563 7424 597
rect 7424 563 7458 597
rect 7458 563 7466 597
rect 7414 552 7466 563
rect 7414 525 7466 540
rect 7414 491 7424 525
rect 7424 491 7458 525
rect 7458 491 7466 525
rect 7414 488 7466 491
rect 7142 102 7194 154
rect 7208 102 7260 154
rect 7142 32 7194 84
rect 7208 32 7260 84
rect 7142 -39 7194 13
rect 7208 -39 7260 13
rect 2748 -58 2800 -46
rect 2813 -58 2865 -46
rect 2878 -58 2930 -46
rect 2943 -58 2995 -46
rect 3008 -58 3060 -46
rect 3073 -58 3125 -46
rect 2748 -92 2775 -58
rect 2775 -92 2800 -58
rect 2813 -92 2848 -58
rect 2848 -92 2865 -58
rect 2878 -92 2882 -58
rect 2882 -92 2921 -58
rect 2921 -92 2930 -58
rect 2943 -92 2955 -58
rect 2955 -92 2994 -58
rect 2994 -92 2995 -58
rect 3008 -92 3028 -58
rect 3028 -92 3060 -58
rect 3073 -92 3101 -58
rect 3101 -92 3125 -58
rect 2748 -98 2800 -92
rect 2813 -98 2865 -92
rect 2878 -98 2930 -92
rect 2943 -98 2995 -92
rect 3008 -98 3060 -92
rect 3073 -98 3125 -92
rect 3138 -58 3190 -46
rect 3138 -92 3140 -58
rect 3140 -92 3174 -58
rect 3174 -92 3190 -58
rect 3138 -98 3190 -92
rect 3203 -58 3255 -46
rect 3203 -92 3213 -58
rect 3213 -92 3247 -58
rect 3247 -92 3255 -58
rect 3203 -98 3255 -92
rect 3268 -58 3320 -46
rect 3268 -92 3286 -58
rect 3286 -92 3320 -58
rect 3268 -98 3320 -92
rect 3333 -58 3385 -46
rect 3398 -58 3450 -46
rect 3463 -58 3515 -46
rect 3528 -58 3580 -46
rect 3593 -58 3645 -46
rect 3658 -58 3710 -46
rect 3333 -92 3359 -58
rect 3359 -92 3385 -58
rect 3398 -92 3432 -58
rect 3432 -92 3450 -58
rect 3463 -92 3466 -58
rect 3466 -92 3505 -58
rect 3505 -92 3515 -58
rect 3528 -92 3539 -58
rect 3539 -92 3578 -58
rect 3578 -92 3580 -58
rect 3593 -92 3612 -58
rect 3612 -92 3645 -58
rect 3658 -92 3685 -58
rect 3685 -92 3710 -58
rect 3333 -98 3385 -92
rect 3398 -98 3450 -92
rect 3463 -98 3515 -92
rect 3528 -98 3580 -92
rect 3593 -98 3645 -92
rect 3658 -98 3710 -92
rect 3723 -58 3775 -46
rect 3723 -92 3724 -58
rect 3724 -92 3758 -58
rect 3758 -92 3775 -58
rect 3723 -98 3775 -92
rect 3788 -58 3840 -46
rect 3788 -92 3797 -58
rect 3797 -92 3831 -58
rect 3831 -92 3840 -58
rect 3788 -98 3840 -92
rect 3853 -58 3905 -46
rect 3853 -92 3870 -58
rect 3870 -92 3904 -58
rect 3904 -92 3905 -58
rect 3853 -98 3905 -92
rect 3918 -58 3970 -46
rect 3983 -58 4035 -46
rect 4048 -58 4100 -46
rect 4113 -58 4165 -46
rect 4178 -58 4230 -46
rect 4243 -58 4295 -46
rect 4308 -58 4360 -46
rect 3918 -92 3943 -58
rect 3943 -92 3970 -58
rect 3983 -92 4016 -58
rect 4016 -92 4035 -58
rect 4048 -92 4050 -58
rect 4050 -92 4089 -58
rect 4089 -92 4100 -58
rect 4113 -92 4123 -58
rect 4123 -92 4161 -58
rect 4161 -92 4165 -58
rect 4178 -92 4195 -58
rect 4195 -92 4230 -58
rect 4243 -92 4267 -58
rect 4267 -92 4295 -58
rect 4308 -92 4339 -58
rect 4339 -92 4360 -58
rect 3918 -98 3970 -92
rect 3983 -98 4035 -92
rect 4048 -98 4100 -92
rect 4113 -98 4165 -92
rect 4178 -98 4230 -92
rect 4243 -98 4295 -92
rect 4308 -98 4360 -92
rect 4373 -58 4425 -46
rect 4373 -92 4377 -58
rect 4377 -92 4411 -58
rect 4411 -92 4425 -58
rect 4373 -98 4425 -92
rect 4438 -58 4490 -46
rect 4438 -92 4449 -58
rect 4449 -92 4483 -58
rect 4483 -92 4490 -58
rect 4438 -98 4490 -92
rect 4503 -58 4555 -46
rect 4503 -92 4521 -58
rect 4521 -92 4555 -58
rect 4503 -98 4555 -92
rect 4568 -58 4620 -46
rect 4632 -58 4684 -46
rect 4696 -58 4748 -46
rect 4760 -58 4812 -46
rect 4824 -58 4876 -46
rect 4888 -58 4940 -46
rect 4568 -92 4593 -58
rect 4593 -92 4620 -58
rect 4632 -92 4665 -58
rect 4665 -92 4684 -58
rect 4696 -92 4699 -58
rect 4699 -92 4737 -58
rect 4737 -92 4748 -58
rect 4760 -92 4771 -58
rect 4771 -92 4809 -58
rect 4809 -92 4812 -58
rect 4824 -92 4843 -58
rect 4843 -92 4876 -58
rect 4888 -92 4915 -58
rect 4915 -92 4940 -58
rect 4568 -98 4620 -92
rect 4632 -98 4684 -92
rect 4696 -98 4748 -92
rect 4760 -98 4812 -92
rect 4824 -98 4876 -92
rect 4888 -98 4940 -92
rect 4952 -58 5004 -46
rect 4952 -92 4953 -58
rect 4953 -92 4987 -58
rect 4987 -92 5004 -58
rect 4952 -98 5004 -92
rect 5016 -58 5068 -46
rect 5016 -92 5025 -58
rect 5025 -92 5059 -58
rect 5059 -92 5068 -58
rect 5016 -98 5068 -92
rect 5080 -58 5132 -46
rect 5080 -92 5097 -58
rect 5097 -92 5131 -58
rect 5131 -92 5132 -58
rect 5080 -98 5132 -92
rect 5144 -58 5196 -46
rect 5208 -58 5260 -46
rect 5272 -58 5324 -46
rect 5336 -58 5388 -46
rect 5400 -58 5452 -46
rect 5464 -58 5516 -46
rect 5144 -92 5169 -58
rect 5169 -92 5196 -58
rect 5208 -92 5241 -58
rect 5241 -92 5260 -58
rect 5272 -92 5275 -58
rect 5275 -92 5313 -58
rect 5313 -92 5324 -58
rect 5336 -92 5347 -58
rect 5347 -92 5385 -58
rect 5385 -92 5388 -58
rect 5400 -92 5419 -58
rect 5419 -92 5452 -58
rect 5464 -92 5491 -58
rect 5491 -92 5516 -58
rect 5144 -98 5196 -92
rect 5208 -98 5260 -92
rect 5272 -98 5324 -92
rect 5336 -98 5388 -92
rect 5400 -98 5452 -92
rect 5464 -98 5516 -92
rect 5528 -58 5580 -46
rect 5528 -92 5529 -58
rect 5529 -92 5563 -58
rect 5563 -92 5580 -58
rect 5528 -98 5580 -92
rect 5592 -58 5644 -46
rect 5592 -92 5601 -58
rect 5601 -92 5635 -58
rect 5635 -92 5644 -58
rect 5592 -98 5644 -92
rect 5680 -58 5732 -46
rect 5680 -92 5686 -58
rect 5686 -92 5720 -58
rect 5720 -92 5732 -58
rect 5680 -98 5732 -92
rect 5745 -58 5797 -46
rect 5745 -92 5760 -58
rect 5760 -92 5794 -58
rect 5794 -92 5797 -58
rect 5745 -98 5797 -92
rect 5810 -58 5862 -46
rect 5875 -58 5927 -46
rect 5940 -58 5992 -46
rect 6005 -58 6057 -46
rect 6070 -58 6122 -46
rect 6135 -58 6187 -46
rect 5810 -92 5834 -58
rect 5834 -92 5862 -58
rect 5875 -92 5908 -58
rect 5908 -92 5927 -58
rect 5940 -92 5942 -58
rect 5942 -92 5982 -58
rect 5982 -92 5992 -58
rect 6005 -92 6016 -58
rect 6016 -92 6056 -58
rect 6056 -92 6057 -58
rect 6070 -92 6090 -58
rect 6090 -92 6122 -58
rect 6135 -92 6163 -58
rect 6163 -92 6187 -58
rect 5810 -98 5862 -92
rect 5875 -98 5927 -92
rect 5940 -98 5992 -92
rect 6005 -98 6057 -92
rect 6070 -98 6122 -92
rect 6135 -98 6187 -92
rect 6200 -58 6252 -46
rect 6200 -92 6202 -58
rect 6202 -92 6236 -58
rect 6236 -92 6252 -58
rect 6200 -98 6252 -92
rect 6265 -58 6317 -46
rect 6265 -92 6275 -58
rect 6275 -92 6309 -58
rect 6309 -92 6317 -58
rect 6265 -98 6317 -92
rect 6330 -58 6382 -46
rect 6330 -92 6348 -58
rect 6348 -92 6382 -58
rect 6330 -98 6382 -92
rect 6395 -58 6447 -46
rect 6460 -58 6512 -46
rect 6525 -58 6577 -46
rect 6590 -58 6642 -46
rect 6655 -58 6707 -46
rect 6720 -58 6772 -46
rect 6395 -92 6421 -58
rect 6421 -92 6447 -58
rect 6460 -92 6494 -58
rect 6494 -92 6512 -58
rect 6525 -92 6528 -58
rect 6528 -92 6567 -58
rect 6567 -92 6577 -58
rect 6590 -92 6601 -58
rect 6601 -92 6640 -58
rect 6640 -92 6642 -58
rect 6655 -92 6674 -58
rect 6674 -92 6707 -58
rect 6720 -92 6747 -58
rect 6747 -92 6772 -58
rect 6395 -98 6447 -92
rect 6460 -98 6512 -92
rect 6525 -98 6577 -92
rect 6590 -98 6642 -92
rect 6655 -98 6707 -92
rect 6720 -98 6772 -92
rect 6785 -58 6837 -46
rect 6785 -92 6786 -58
rect 6786 -92 6820 -58
rect 6820 -92 6837 -58
rect 6785 -98 6837 -92
rect 6850 -58 6902 -46
rect 6850 -92 6859 -58
rect 6859 -92 6893 -58
rect 6893 -92 6902 -58
rect 6850 -98 6902 -92
rect 7142 -110 7194 -58
rect 7208 -110 7260 -58
rect 7673 1283 7682 1293
rect 7682 1283 7716 1293
rect 7716 1283 7725 1293
rect 7673 1245 7725 1283
rect 7673 1241 7682 1245
rect 7682 1241 7716 1245
rect 7716 1241 7725 1245
rect 7673 1211 7682 1229
rect 7682 1211 7716 1229
rect 7716 1211 7725 1229
rect 7673 1177 7725 1211
rect 7845 1283 7854 1293
rect 7854 1283 7888 1293
rect 7888 1283 7897 1293
rect 7845 1245 7897 1283
rect 7845 1241 7854 1245
rect 7854 1241 7888 1245
rect 7888 1241 7897 1245
rect 7845 1211 7854 1229
rect 7854 1211 7888 1229
rect 7888 1211 7897 1229
rect 7845 1177 7897 1211
rect 7586 597 7638 604
rect 7586 563 7596 597
rect 7596 563 7630 597
rect 7630 563 7638 597
rect 7586 552 7638 563
rect 7586 525 7638 540
rect 7586 491 7596 525
rect 7596 491 7630 525
rect 7630 491 7638 525
rect 7586 488 7638 491
rect 7758 707 7768 714
rect 7768 707 7802 714
rect 7802 707 7810 714
rect 7758 669 7810 707
rect 7758 662 7768 669
rect 7768 662 7802 669
rect 7802 662 7810 669
rect 7758 635 7768 650
rect 7768 635 7802 650
rect 7802 635 7810 650
rect 7758 598 7810 635
rect 7929 478 7981 530
rect 7929 414 7981 466
rect 10607 2213 10659 2222
rect 10607 2179 10613 2213
rect 10613 2179 10647 2213
rect 10647 2179 10659 2213
rect 10607 2170 10659 2179
rect 10671 2213 10723 2222
rect 10671 2179 10685 2213
rect 10685 2179 10719 2213
rect 10719 2179 10723 2213
rect 10671 2170 10723 2179
rect 16764 2831 16816 2883
rect 16828 2831 16880 2883
rect 18066 2831 18118 2883
rect 18132 2831 18184 2883
rect 18953 2849 18977 2883
rect 18977 2849 19005 2883
rect 19044 2849 19056 2883
rect 19056 2849 19090 2883
rect 19090 2849 19096 2883
rect 18953 2843 19005 2849
rect 19044 2843 19096 2849
rect 17132 2737 17184 2789
rect 17196 2737 17248 2789
rect 16773 2640 16825 2692
rect 16837 2640 16889 2692
rect 18218 2640 18270 2692
rect 18282 2640 18334 2692
rect 18401 2727 18453 2739
rect 18492 2727 18544 2739
rect 18401 2693 18430 2727
rect 18430 2693 18453 2727
rect 18492 2693 18509 2727
rect 18509 2693 18543 2727
rect 18543 2693 18544 2727
rect 18401 2687 18453 2693
rect 18492 2687 18544 2693
rect 17298 2560 17350 2612
rect 17362 2560 17414 2612
rect 8010 394 8062 446
rect 8010 330 8062 382
rect 9929 2086 9981 2138
rect 9993 2086 10045 2138
rect 10775 2047 10827 2052
rect 9201 1932 9253 1984
rect 9201 1868 9253 1920
rect 9401 1987 9453 2013
rect 9401 1961 9411 1987
rect 9411 1961 9445 1987
rect 9445 1961 9453 1987
rect 10775 2013 10792 2047
rect 10792 2013 10826 2047
rect 10826 2013 10827 2047
rect 10775 2000 10827 2013
rect 10839 2047 10891 2052
rect 10927 2047 10979 2052
rect 10839 2013 10865 2047
rect 10865 2013 10891 2047
rect 10927 2013 10938 2047
rect 10938 2013 10972 2047
rect 10972 2013 10979 2047
rect 10839 2000 10891 2013
rect 10927 2000 10979 2013
rect 10992 2047 11044 2052
rect 10992 2013 11010 2047
rect 11010 2013 11044 2047
rect 10992 2000 11044 2013
rect 11057 2047 11109 2052
rect 11122 2047 11174 2052
rect 11187 2047 11239 2052
rect 11252 2047 11304 2052
rect 11317 2047 11369 2052
rect 11382 2047 11434 2052
rect 11447 2047 11499 2052
rect 11057 2013 11082 2047
rect 11082 2013 11109 2047
rect 11122 2013 11154 2047
rect 11154 2013 11174 2047
rect 11187 2013 11188 2047
rect 11188 2013 11226 2047
rect 11226 2013 11239 2047
rect 11252 2013 11260 2047
rect 11260 2013 11298 2047
rect 11298 2013 11304 2047
rect 11317 2013 11332 2047
rect 11332 2013 11369 2047
rect 11382 2013 11404 2047
rect 11404 2013 11434 2047
rect 11447 2013 11476 2047
rect 11476 2013 11499 2047
rect 11057 2000 11109 2013
rect 11122 2000 11174 2013
rect 11187 2000 11239 2013
rect 11252 2000 11304 2013
rect 11317 2000 11369 2013
rect 11382 2000 11434 2013
rect 11447 2000 11499 2013
rect 11512 2047 11564 2052
rect 11512 2013 11514 2047
rect 11514 2013 11548 2047
rect 11548 2013 11564 2047
rect 11512 2000 11564 2013
rect 11577 2047 11629 2052
rect 11577 2013 11586 2047
rect 11586 2013 11620 2047
rect 11620 2013 11629 2047
rect 11577 2000 11629 2013
rect 11642 2047 11694 2052
rect 11642 2013 11658 2047
rect 11658 2013 11692 2047
rect 11692 2013 11694 2047
rect 11642 2000 11694 2013
rect 11707 2047 11759 2052
rect 11772 2047 11824 2052
rect 11837 2047 11889 2052
rect 11901 2047 11953 2052
rect 11965 2047 12017 2052
rect 12029 2047 12081 2052
rect 12093 2047 12145 2052
rect 11707 2013 11730 2047
rect 11730 2013 11759 2047
rect 11772 2013 11802 2047
rect 11802 2013 11824 2047
rect 11837 2013 11874 2047
rect 11874 2013 11889 2047
rect 11901 2013 11908 2047
rect 11908 2013 11946 2047
rect 11946 2013 11953 2047
rect 11965 2013 11980 2047
rect 11980 2013 12017 2047
rect 12029 2013 12052 2047
rect 12052 2013 12081 2047
rect 12093 2013 12124 2047
rect 12124 2013 12145 2047
rect 11707 2000 11759 2013
rect 11772 2000 11824 2013
rect 11837 2000 11889 2013
rect 11901 2000 11953 2013
rect 11965 2000 12017 2013
rect 12029 2000 12081 2013
rect 12093 2000 12145 2013
rect 12157 2047 12209 2052
rect 12157 2013 12162 2047
rect 12162 2013 12196 2047
rect 12196 2013 12209 2047
rect 12157 2000 12209 2013
rect 12221 2047 12273 2052
rect 12221 2013 12234 2047
rect 12234 2013 12268 2047
rect 12268 2013 12273 2047
rect 12221 2000 12273 2013
rect 12285 2047 12337 2052
rect 12349 2047 12401 2052
rect 12413 2047 12465 2052
rect 12477 2047 12529 2052
rect 12541 2047 12593 2052
rect 12605 2047 12657 2052
rect 12669 2047 12721 2052
rect 12285 2013 12306 2047
rect 12306 2013 12337 2047
rect 12349 2013 12378 2047
rect 12378 2013 12401 2047
rect 12413 2013 12450 2047
rect 12450 2013 12465 2047
rect 12477 2013 12484 2047
rect 12484 2013 12522 2047
rect 12522 2013 12529 2047
rect 12541 2013 12556 2047
rect 12556 2013 12593 2047
rect 12605 2013 12628 2047
rect 12628 2013 12657 2047
rect 12669 2013 12700 2047
rect 12700 2013 12721 2047
rect 12285 2000 12337 2013
rect 12349 2000 12401 2013
rect 12413 2000 12465 2013
rect 12477 2000 12529 2013
rect 12541 2000 12593 2013
rect 12605 2000 12657 2013
rect 12669 2000 12721 2013
rect 12733 2047 12785 2052
rect 12733 2013 12738 2047
rect 12738 2013 12772 2047
rect 12772 2013 12785 2047
rect 12733 2000 12785 2013
rect 12797 2047 12849 2052
rect 12797 2013 12810 2047
rect 12810 2013 12844 2047
rect 12844 2013 12849 2047
rect 12797 2000 12849 2013
rect 12861 2047 12913 2052
rect 12925 2047 12977 2052
rect 12989 2047 13041 2052
rect 13053 2047 13105 2052
rect 13117 2047 13169 2052
rect 13181 2047 13233 2052
rect 13245 2047 13297 2052
rect 12861 2013 12882 2047
rect 12882 2013 12913 2047
rect 12925 2013 12954 2047
rect 12954 2013 12977 2047
rect 12989 2013 13026 2047
rect 13026 2013 13041 2047
rect 13053 2013 13060 2047
rect 13060 2013 13098 2047
rect 13098 2013 13105 2047
rect 13117 2013 13132 2047
rect 13132 2013 13169 2047
rect 13181 2013 13204 2047
rect 13204 2013 13233 2047
rect 13245 2013 13276 2047
rect 13276 2013 13297 2047
rect 12861 2000 12913 2013
rect 12925 2000 12977 2013
rect 12989 2000 13041 2013
rect 13053 2000 13105 2013
rect 13117 2000 13169 2013
rect 13181 2000 13233 2013
rect 13245 2000 13297 2013
rect 13309 2047 13361 2052
rect 13309 2013 13314 2047
rect 13314 2013 13348 2047
rect 13348 2013 13361 2047
rect 13309 2000 13361 2013
rect 13373 2047 13425 2052
rect 13373 2013 13386 2047
rect 13386 2013 13420 2047
rect 13420 2013 13425 2047
rect 13373 2000 13425 2013
rect 13437 2047 13489 2052
rect 13437 2013 13458 2047
rect 13458 2013 13489 2047
rect 13437 2000 13489 2013
rect 25334 2023 25386 2075
rect 25398 2023 25450 2075
rect 9401 1908 9453 1932
rect 9401 1880 9411 1908
rect 9411 1880 9445 1908
rect 9445 1880 9453 1908
rect 9401 1829 9453 1850
rect 9401 1798 9411 1829
rect 9411 1798 9445 1829
rect 9445 1798 9453 1829
rect 9203 1722 9255 1774
rect 9203 1658 9255 1710
rect 10762 1884 10765 1885
rect 10765 1884 10799 1885
rect 10799 1884 10814 1885
rect 10762 1836 10814 1884
rect 10762 1833 10765 1836
rect 10765 1833 10799 1836
rect 10799 1833 10814 1836
rect 10829 1884 10838 1885
rect 10838 1884 10872 1885
rect 10872 1884 10881 1885
rect 10829 1836 10881 1884
rect 10829 1833 10838 1836
rect 10838 1833 10872 1836
rect 10872 1833 10881 1836
rect 10896 1884 10911 1885
rect 10911 1884 10945 1885
rect 10945 1884 10948 1885
rect 10896 1836 10948 1884
rect 10896 1833 10911 1836
rect 10911 1833 10945 1836
rect 10945 1833 10948 1836
rect 10963 1884 10984 1885
rect 10984 1884 11015 1885
rect 11030 1884 11057 1885
rect 11057 1884 11082 1885
rect 11097 1884 11130 1885
rect 11130 1884 11149 1885
rect 11164 1884 11203 1885
rect 11203 1884 11216 1885
rect 11231 1884 11237 1885
rect 11237 1884 11276 1885
rect 11276 1884 11283 1885
rect 11298 1884 11310 1885
rect 11310 1884 11349 1885
rect 11349 1884 11350 1885
rect 11365 1884 11383 1885
rect 11383 1884 11417 1885
rect 11432 1884 11456 1885
rect 11456 1884 11484 1885
rect 11499 1884 11529 1885
rect 11529 1884 11551 1885
rect 10963 1836 11015 1884
rect 11030 1836 11082 1884
rect 11097 1836 11149 1884
rect 11164 1836 11216 1884
rect 11231 1836 11283 1884
rect 11298 1836 11350 1884
rect 11365 1836 11417 1884
rect 11432 1836 11484 1884
rect 11499 1836 11551 1884
rect 10963 1833 10984 1836
rect 10984 1833 11015 1836
rect 11030 1833 11057 1836
rect 11057 1833 11082 1836
rect 11097 1833 11130 1836
rect 11130 1833 11149 1836
rect 11164 1833 11203 1836
rect 11203 1833 11216 1836
rect 11231 1833 11237 1836
rect 11237 1833 11276 1836
rect 11276 1833 11283 1836
rect 11298 1833 11310 1836
rect 11310 1833 11349 1836
rect 11349 1833 11350 1836
rect 11365 1833 11383 1836
rect 11383 1833 11417 1836
rect 11432 1833 11456 1836
rect 11456 1833 11484 1836
rect 11499 1833 11529 1836
rect 11529 1833 11551 1836
rect 11566 1884 11568 1885
rect 11568 1884 11602 1885
rect 11602 1884 11618 1885
rect 11566 1836 11618 1884
rect 11566 1833 11568 1836
rect 11568 1833 11602 1836
rect 11602 1833 11618 1836
rect 11633 1884 11641 1885
rect 11641 1884 11675 1885
rect 11675 1884 11685 1885
rect 11633 1836 11685 1884
rect 11633 1833 11641 1836
rect 11641 1833 11675 1836
rect 11675 1833 11685 1836
rect 11699 1884 11714 1885
rect 11714 1884 11748 1885
rect 11748 1884 11751 1885
rect 11699 1836 11751 1884
rect 11699 1833 11714 1836
rect 11714 1833 11748 1836
rect 11748 1833 11751 1836
rect 11765 1884 11787 1885
rect 11787 1884 11817 1885
rect 11831 1884 11860 1885
rect 11860 1884 11883 1885
rect 11897 1884 11933 1885
rect 11933 1884 11949 1885
rect 11963 1884 11967 1885
rect 11967 1884 12006 1885
rect 12006 1884 12015 1885
rect 12029 1884 12040 1885
rect 12040 1884 12079 1885
rect 12079 1884 12081 1885
rect 12095 1884 12113 1885
rect 12113 1884 12147 1885
rect 12161 1884 12186 1885
rect 12186 1884 12213 1885
rect 12227 1884 12259 1885
rect 12259 1884 12279 1885
rect 11765 1836 11817 1884
rect 11831 1836 11883 1884
rect 11897 1836 11949 1884
rect 11963 1836 12015 1884
rect 12029 1836 12081 1884
rect 12095 1836 12147 1884
rect 12161 1836 12213 1884
rect 12227 1836 12279 1884
rect 11765 1833 11787 1836
rect 11787 1833 11817 1836
rect 11831 1833 11860 1836
rect 11860 1833 11883 1836
rect 11897 1833 11933 1836
rect 11933 1833 11949 1836
rect 11963 1833 11967 1836
rect 11967 1833 12006 1836
rect 12006 1833 12015 1836
rect 12029 1833 12040 1836
rect 12040 1833 12079 1836
rect 12079 1833 12081 1836
rect 12095 1833 12113 1836
rect 12113 1833 12147 1836
rect 12161 1833 12186 1836
rect 12186 1833 12213 1836
rect 12227 1833 12259 1836
rect 12259 1833 12279 1836
rect 12293 1884 12298 1885
rect 12298 1884 12332 1885
rect 12332 1884 12345 1885
rect 12293 1836 12345 1884
rect 12293 1833 12298 1836
rect 12298 1833 12332 1836
rect 12332 1833 12345 1836
rect 12359 1884 12371 1885
rect 12371 1884 12405 1885
rect 12405 1884 12411 1885
rect 12359 1836 12411 1884
rect 12359 1833 12371 1836
rect 12371 1833 12405 1836
rect 12405 1833 12411 1836
rect 10762 1802 10765 1805
rect 10765 1802 10799 1805
rect 10799 1802 10814 1805
rect 10762 1754 10814 1802
rect 10762 1753 10765 1754
rect 10765 1753 10799 1754
rect 10799 1753 10814 1754
rect 10829 1802 10838 1805
rect 10838 1802 10872 1805
rect 10872 1802 10881 1805
rect 10829 1754 10881 1802
rect 10829 1753 10838 1754
rect 10838 1753 10872 1754
rect 10872 1753 10881 1754
rect 10896 1802 10911 1805
rect 10911 1802 10945 1805
rect 10945 1802 10948 1805
rect 10896 1754 10948 1802
rect 10896 1753 10911 1754
rect 10911 1753 10945 1754
rect 10945 1753 10948 1754
rect 10963 1802 10984 1805
rect 10984 1802 11015 1805
rect 11030 1802 11057 1805
rect 11057 1802 11082 1805
rect 11097 1802 11130 1805
rect 11130 1802 11149 1805
rect 11164 1802 11203 1805
rect 11203 1802 11216 1805
rect 11231 1802 11237 1805
rect 11237 1802 11276 1805
rect 11276 1802 11283 1805
rect 11298 1802 11310 1805
rect 11310 1802 11349 1805
rect 11349 1802 11350 1805
rect 11365 1802 11383 1805
rect 11383 1802 11417 1805
rect 11432 1802 11456 1805
rect 11456 1802 11484 1805
rect 11499 1802 11529 1805
rect 11529 1802 11551 1805
rect 10963 1754 11015 1802
rect 11030 1754 11082 1802
rect 11097 1754 11149 1802
rect 11164 1754 11216 1802
rect 11231 1754 11283 1802
rect 11298 1754 11350 1802
rect 11365 1754 11417 1802
rect 11432 1754 11484 1802
rect 11499 1754 11551 1802
rect 10963 1753 10984 1754
rect 10984 1753 11015 1754
rect 11030 1753 11057 1754
rect 11057 1753 11082 1754
rect 11097 1753 11130 1754
rect 11130 1753 11149 1754
rect 11164 1753 11203 1754
rect 11203 1753 11216 1754
rect 11231 1753 11237 1754
rect 11237 1753 11276 1754
rect 11276 1753 11283 1754
rect 11298 1753 11310 1754
rect 11310 1753 11349 1754
rect 11349 1753 11350 1754
rect 11365 1753 11383 1754
rect 11383 1753 11417 1754
rect 11432 1753 11456 1754
rect 11456 1753 11484 1754
rect 11499 1753 11529 1754
rect 11529 1753 11551 1754
rect 11566 1802 11568 1805
rect 11568 1802 11602 1805
rect 11602 1802 11618 1805
rect 11566 1754 11618 1802
rect 11566 1753 11568 1754
rect 11568 1753 11602 1754
rect 11602 1753 11618 1754
rect 11633 1802 11641 1805
rect 11641 1802 11675 1805
rect 11675 1802 11685 1805
rect 11633 1754 11685 1802
rect 11633 1753 11641 1754
rect 11641 1753 11675 1754
rect 11675 1753 11685 1754
rect 11699 1802 11714 1805
rect 11714 1802 11748 1805
rect 11748 1802 11751 1805
rect 11699 1754 11751 1802
rect 11699 1753 11714 1754
rect 11714 1753 11748 1754
rect 11748 1753 11751 1754
rect 11765 1802 11787 1805
rect 11787 1802 11817 1805
rect 11831 1802 11860 1805
rect 11860 1802 11883 1805
rect 11897 1802 11933 1805
rect 11933 1802 11949 1805
rect 11963 1802 11967 1805
rect 11967 1802 12006 1805
rect 12006 1802 12015 1805
rect 12029 1802 12040 1805
rect 12040 1802 12079 1805
rect 12079 1802 12081 1805
rect 12095 1802 12113 1805
rect 12113 1802 12147 1805
rect 12161 1802 12186 1805
rect 12186 1802 12213 1805
rect 12227 1802 12259 1805
rect 12259 1802 12279 1805
rect 11765 1754 11817 1802
rect 11831 1754 11883 1802
rect 11897 1754 11949 1802
rect 11963 1754 12015 1802
rect 12029 1754 12081 1802
rect 12095 1754 12147 1802
rect 12161 1754 12213 1802
rect 12227 1754 12279 1802
rect 11765 1753 11787 1754
rect 11787 1753 11817 1754
rect 11831 1753 11860 1754
rect 11860 1753 11883 1754
rect 11897 1753 11933 1754
rect 11933 1753 11949 1754
rect 11963 1753 11967 1754
rect 11967 1753 12006 1754
rect 12006 1753 12015 1754
rect 12029 1753 12040 1754
rect 12040 1753 12079 1754
rect 12079 1753 12081 1754
rect 12095 1753 12113 1754
rect 12113 1753 12147 1754
rect 12161 1753 12186 1754
rect 12186 1753 12213 1754
rect 12227 1753 12259 1754
rect 12259 1753 12279 1754
rect 12293 1802 12298 1805
rect 12298 1802 12332 1805
rect 12332 1802 12345 1805
rect 12293 1754 12345 1802
rect 12293 1753 12298 1754
rect 12298 1753 12332 1754
rect 12332 1753 12345 1754
rect 12359 1802 12371 1805
rect 12371 1802 12405 1805
rect 12405 1802 12411 1805
rect 12359 1754 12411 1802
rect 12359 1753 12371 1754
rect 12371 1753 12405 1754
rect 12405 1753 12411 1754
rect 10762 1720 10765 1725
rect 10765 1720 10799 1725
rect 10799 1720 10814 1725
rect 10762 1673 10814 1720
rect 10829 1720 10838 1725
rect 10838 1720 10872 1725
rect 10872 1720 10881 1725
rect 10829 1673 10881 1720
rect 10896 1720 10911 1725
rect 10911 1720 10945 1725
rect 10945 1720 10948 1725
rect 10896 1673 10948 1720
rect 10963 1720 10984 1725
rect 10984 1720 11015 1725
rect 11030 1720 11057 1725
rect 11057 1720 11082 1725
rect 11097 1720 11130 1725
rect 11130 1720 11149 1725
rect 11164 1720 11203 1725
rect 11203 1720 11216 1725
rect 11231 1720 11237 1725
rect 11237 1720 11276 1725
rect 11276 1720 11283 1725
rect 11298 1720 11310 1725
rect 11310 1720 11349 1725
rect 11349 1720 11350 1725
rect 11365 1720 11383 1725
rect 11383 1720 11417 1725
rect 11432 1720 11456 1725
rect 11456 1720 11484 1725
rect 11499 1720 11529 1725
rect 11529 1720 11551 1725
rect 10963 1673 11015 1720
rect 11030 1673 11082 1720
rect 11097 1673 11149 1720
rect 11164 1673 11216 1720
rect 11231 1673 11283 1720
rect 11298 1673 11350 1720
rect 11365 1673 11417 1720
rect 11432 1673 11484 1720
rect 11499 1673 11551 1720
rect 11566 1720 11568 1725
rect 11568 1720 11602 1725
rect 11602 1720 11618 1725
rect 11566 1673 11618 1720
rect 11633 1720 11641 1725
rect 11641 1720 11675 1725
rect 11675 1720 11685 1725
rect 11633 1673 11685 1720
rect 11699 1720 11714 1725
rect 11714 1720 11748 1725
rect 11748 1720 11751 1725
rect 11699 1673 11751 1720
rect 11765 1720 11787 1725
rect 11787 1720 11817 1725
rect 11831 1720 11860 1725
rect 11860 1720 11883 1725
rect 11897 1720 11933 1725
rect 11933 1720 11949 1725
rect 11963 1720 11967 1725
rect 11967 1720 12006 1725
rect 12006 1720 12015 1725
rect 12029 1720 12040 1725
rect 12040 1720 12079 1725
rect 12079 1720 12081 1725
rect 12095 1720 12113 1725
rect 12113 1720 12147 1725
rect 12161 1720 12186 1725
rect 12186 1720 12213 1725
rect 12227 1720 12259 1725
rect 12259 1720 12279 1725
rect 11765 1673 11817 1720
rect 11831 1673 11883 1720
rect 11897 1673 11949 1720
rect 11963 1673 12015 1720
rect 12029 1673 12081 1720
rect 12095 1673 12147 1720
rect 12161 1673 12213 1720
rect 12227 1673 12279 1720
rect 12293 1720 12298 1725
rect 12298 1720 12332 1725
rect 12332 1720 12345 1725
rect 12293 1673 12345 1720
rect 12359 1720 12371 1725
rect 12371 1720 12405 1725
rect 12405 1720 12411 1725
rect 12359 1673 12411 1720
rect 16535 1708 16587 1760
rect 16611 1708 16663 1760
rect 16687 1708 16739 1760
rect 10762 1638 10765 1645
rect 10765 1638 10799 1645
rect 10799 1638 10814 1645
rect 10762 1593 10814 1638
rect 10829 1638 10838 1645
rect 10838 1638 10872 1645
rect 10872 1638 10881 1645
rect 10829 1593 10881 1638
rect 10896 1638 10911 1645
rect 10911 1638 10945 1645
rect 10945 1638 10948 1645
rect 10896 1593 10948 1638
rect 10963 1638 10984 1645
rect 10984 1638 11015 1645
rect 11030 1638 11057 1645
rect 11057 1638 11082 1645
rect 11097 1638 11130 1645
rect 11130 1638 11149 1645
rect 11164 1638 11203 1645
rect 11203 1638 11216 1645
rect 11231 1638 11237 1645
rect 11237 1638 11276 1645
rect 11276 1638 11283 1645
rect 11298 1638 11310 1645
rect 11310 1638 11349 1645
rect 11349 1638 11350 1645
rect 11365 1638 11383 1645
rect 11383 1638 11417 1645
rect 11432 1638 11456 1645
rect 11456 1638 11484 1645
rect 11499 1638 11529 1645
rect 11529 1638 11551 1645
rect 10963 1593 11015 1638
rect 11030 1593 11082 1638
rect 11097 1593 11149 1638
rect 11164 1593 11216 1638
rect 11231 1593 11283 1638
rect 11298 1593 11350 1638
rect 11365 1593 11417 1638
rect 11432 1593 11484 1638
rect 11499 1593 11551 1638
rect 11566 1638 11568 1645
rect 11568 1638 11602 1645
rect 11602 1638 11618 1645
rect 11566 1593 11618 1638
rect 11633 1638 11641 1645
rect 11641 1638 11675 1645
rect 11675 1638 11685 1645
rect 11633 1593 11685 1638
rect 11699 1638 11714 1645
rect 11714 1638 11748 1645
rect 11748 1638 11751 1645
rect 11699 1593 11751 1638
rect 11765 1638 11787 1645
rect 11787 1638 11817 1645
rect 11831 1638 11860 1645
rect 11860 1638 11883 1645
rect 11897 1638 11933 1645
rect 11933 1638 11949 1645
rect 11963 1638 11967 1645
rect 11967 1638 12006 1645
rect 12006 1638 12015 1645
rect 12029 1638 12040 1645
rect 12040 1638 12079 1645
rect 12079 1638 12081 1645
rect 12095 1638 12113 1645
rect 12113 1638 12147 1645
rect 12161 1638 12186 1645
rect 12186 1638 12213 1645
rect 12227 1638 12259 1645
rect 12259 1638 12279 1645
rect 11765 1593 11817 1638
rect 11831 1593 11883 1638
rect 11897 1593 11949 1638
rect 11963 1593 12015 1638
rect 12029 1593 12081 1638
rect 12095 1593 12147 1638
rect 12161 1593 12213 1638
rect 12227 1593 12279 1638
rect 12293 1638 12298 1645
rect 12298 1638 12332 1645
rect 12332 1638 12345 1645
rect 12293 1593 12345 1638
rect 12359 1638 12371 1645
rect 12371 1638 12405 1645
rect 12405 1638 12411 1645
rect 12359 1593 12411 1638
rect 16535 1629 16587 1681
rect 16611 1629 16663 1681
rect 16687 1629 16739 1681
rect 18875 1730 18927 1755
rect 18941 1730 18993 1755
rect 18875 1703 18897 1730
rect 18897 1703 18927 1730
rect 18941 1703 18969 1730
rect 18969 1703 18993 1730
rect 19007 1730 19059 1755
rect 19007 1703 19041 1730
rect 19041 1703 19059 1730
rect 19073 1730 19125 1755
rect 19073 1703 19079 1730
rect 19079 1703 19113 1730
rect 19113 1703 19125 1730
rect 19139 1730 19191 1755
rect 19139 1703 19151 1730
rect 19151 1703 19185 1730
rect 19185 1703 19191 1730
rect 18875 1644 18927 1655
rect 18941 1644 18993 1655
rect 18875 1610 18897 1644
rect 18897 1610 18927 1644
rect 18941 1610 18969 1644
rect 18969 1610 18993 1644
rect 18875 1603 18927 1610
rect 18941 1603 18993 1610
rect 19007 1644 19059 1655
rect 19007 1610 19041 1644
rect 19041 1610 19059 1644
rect 19007 1603 19059 1610
rect 19073 1644 19125 1655
rect 19073 1610 19079 1644
rect 19079 1610 19113 1644
rect 19113 1610 19125 1644
rect 19073 1603 19125 1610
rect 19139 1644 19191 1655
rect 19139 1610 19151 1644
rect 19151 1610 19185 1644
rect 19185 1610 19191 1644
rect 19139 1603 19191 1610
rect 16535 1550 16587 1602
rect 16611 1550 16663 1602
rect 16687 1550 16739 1602
rect 14443 1462 14495 1514
rect 14507 1462 14559 1514
rect 17619 1485 17671 1537
rect 17683 1485 17735 1537
rect 12264 1355 12316 1367
rect 12328 1355 12380 1367
rect 12264 1321 12282 1355
rect 12282 1321 12316 1355
rect 12328 1321 12354 1355
rect 12354 1321 12380 1355
rect 12264 1315 12316 1321
rect 12328 1315 12380 1321
rect 8431 1164 8483 1216
rect 8509 1164 8561 1216
rect 8587 1164 8639 1216
rect 8665 1164 8717 1216
rect 8743 1164 8795 1216
rect 8090 260 8142 312
rect 8090 196 8142 248
rect 8431 770 8483 808
rect 8431 756 8440 770
rect 8440 756 8474 770
rect 8474 756 8483 770
rect 8431 736 8440 744
rect 8440 736 8474 744
rect 8474 736 8483 744
rect 8431 698 8483 736
rect 8431 692 8440 698
rect 8440 692 8474 698
rect 8474 692 8483 698
rect 8171 148 8223 154
rect 8171 114 8177 148
rect 8177 114 8211 148
rect 8211 114 8223 148
rect 8171 102 8223 114
rect 8275 122 8327 154
rect 8275 102 8284 122
rect 8284 102 8318 122
rect 8318 102 8327 122
rect 8171 71 8223 72
rect 8171 37 8177 71
rect 8177 37 8211 71
rect 8211 37 8223 71
rect 8171 20 8223 37
rect 8275 50 8327 72
rect 8275 20 8284 50
rect 8284 20 8318 50
rect 8318 20 8327 50
rect 8171 -40 8177 -11
rect 8177 -40 8211 -11
rect 8211 -40 8223 -11
rect 8171 -63 8223 -40
rect 8275 -22 8327 -11
rect 8275 -56 8284 -22
rect 8284 -56 8318 -22
rect 8318 -56 8327 -22
rect 8275 -63 8327 -56
rect 8743 770 8795 808
rect 8743 756 8752 770
rect 8752 756 8786 770
rect 8786 756 8795 770
rect 8743 736 8752 744
rect 8752 736 8786 744
rect 8786 736 8795 744
rect 8743 698 8795 736
rect 8743 692 8752 698
rect 8752 692 8786 698
rect 8786 692 8795 698
rect 8587 122 8639 154
rect 8587 102 8596 122
rect 8596 102 8630 122
rect 8630 102 8639 122
rect 8587 50 8639 72
rect 8587 20 8596 50
rect 8596 20 8630 50
rect 8630 20 8639 50
rect 8587 -22 8639 -11
rect 8587 -56 8596 -22
rect 8596 -56 8630 -22
rect 8630 -56 8639 -22
rect 8587 -63 8639 -56
rect 9055 592 9064 618
rect 9064 592 9098 618
rect 9098 592 9107 618
rect 9055 566 9107 592
rect 9055 520 9064 554
rect 9064 520 9098 554
rect 9098 520 9107 554
rect 9055 502 9107 520
rect 8899 122 8951 154
rect 8899 102 8908 122
rect 8908 102 8942 122
rect 8942 102 8951 122
rect 8899 50 8951 72
rect 8899 20 8908 50
rect 8908 20 8942 50
rect 8942 20 8951 50
rect 8899 -22 8951 -11
rect 8899 -56 8908 -22
rect 8908 -56 8942 -22
rect 8942 -56 8951 -22
rect 8899 -63 8951 -56
rect 9367 592 9376 618
rect 9376 592 9410 618
rect 9410 592 9419 618
rect 9367 566 9419 592
rect 9367 520 9376 554
rect 9376 520 9410 554
rect 9410 520 9419 554
rect 9367 502 9419 520
rect 9211 122 9263 154
rect 9211 102 9220 122
rect 9220 102 9254 122
rect 9254 102 9263 122
rect 9211 50 9263 72
rect 9211 20 9220 50
rect 9220 20 9254 50
rect 9254 20 9263 50
rect 9211 -22 9263 -11
rect 9211 -56 9220 -22
rect 9220 -56 9254 -22
rect 9254 -56 9263 -22
rect 9211 -63 9263 -56
rect 9679 592 9688 618
rect 9688 592 9722 618
rect 9722 592 9731 618
rect 9679 566 9731 592
rect 9679 520 9688 554
rect 9688 520 9722 554
rect 9722 520 9731 554
rect 9679 502 9731 520
rect 9991 592 10000 618
rect 10000 592 10034 618
rect 10034 592 10043 618
rect 9991 566 10043 592
rect 9991 520 10000 554
rect 10000 520 10034 554
rect 10034 520 10043 554
rect 9991 502 10043 520
rect 9834 410 9886 420
rect 9834 376 9844 410
rect 9844 376 9878 410
rect 9878 376 9886 410
rect 9834 368 9886 376
rect 9834 338 9886 350
rect 9834 304 9844 338
rect 9844 304 9878 338
rect 9878 304 9886 338
rect 9834 298 9886 304
rect 9523 122 9575 154
rect 9523 102 9532 122
rect 9532 102 9566 122
rect 9566 102 9575 122
rect 9523 50 9575 72
rect 9523 20 9532 50
rect 9532 20 9566 50
rect 9566 20 9575 50
rect 9523 -22 9575 -11
rect 9523 -56 9532 -22
rect 9532 -56 9566 -22
rect 9566 -56 9575 -22
rect 9523 -63 9575 -56
rect 10303 592 10312 618
rect 10312 592 10346 618
rect 10346 592 10355 618
rect 10303 566 10355 592
rect 10303 520 10312 554
rect 10312 520 10346 554
rect 10346 520 10355 554
rect 10303 502 10355 520
rect 10146 410 10198 420
rect 10146 376 10156 410
rect 10156 376 10190 410
rect 10190 376 10198 410
rect 10146 368 10198 376
rect 10146 338 10198 350
rect 10146 304 10156 338
rect 10156 304 10190 338
rect 10190 304 10198 338
rect 10146 298 10198 304
rect 10458 410 10510 420
rect 10458 376 10468 410
rect 10468 376 10502 410
rect 10502 376 10510 410
rect 10458 368 10510 376
rect 10458 338 10510 350
rect 10458 304 10468 338
rect 10468 304 10502 338
rect 10502 304 10510 338
rect 10458 298 10510 304
rect 15831 1391 15883 1443
rect 15895 1391 15947 1443
rect 17381 1391 17433 1443
rect 17445 1391 17497 1443
rect 10595 144 10604 151
rect 10604 144 10638 151
rect 10638 144 10647 151
rect 10595 102 10647 144
rect 10595 99 10604 102
rect 10604 99 10638 102
rect 10638 99 10647 102
rect 10595 26 10647 57
rect 10595 5 10604 26
rect 10604 5 10638 26
rect 10638 5 10647 26
rect 10595 -50 10647 -38
rect 10595 -84 10604 -50
rect 10604 -84 10638 -50
rect 10638 -84 10647 -50
rect 10595 -90 10647 -84
rect 10728 122 10780 151
rect 10728 99 10737 122
rect 10737 99 10771 122
rect 10771 99 10780 122
rect 10728 50 10780 57
rect 10728 16 10737 50
rect 10737 16 10771 50
rect 10771 16 10780 50
rect 10728 5 10780 16
rect 10728 -56 10737 -38
rect 10737 -56 10771 -38
rect 10771 -56 10780 -38
rect 10728 -90 10780 -56
rect 11184 122 11236 151
rect 11184 99 11193 122
rect 11193 99 11227 122
rect 11227 99 11236 122
rect 11184 50 11236 57
rect 11184 16 11193 50
rect 11193 16 11227 50
rect 11227 16 11236 50
rect 11184 5 11236 16
rect 11184 -56 11193 -38
rect 11193 -56 11227 -38
rect 11227 -56 11236 -38
rect 11184 -90 11236 -56
rect 11640 122 11692 151
rect 11640 99 11649 122
rect 11649 99 11683 122
rect 11683 99 11692 122
rect 11640 50 11692 57
rect 11640 16 11649 50
rect 11649 16 11683 50
rect 11683 16 11692 50
rect 11640 5 11692 16
rect 11640 -56 11649 -38
rect 11649 -56 11683 -38
rect 11683 -56 11692 -38
rect 11640 -90 11692 -56
rect 13501 1355 13553 1367
rect 13565 1355 13617 1367
rect 13501 1321 13526 1355
rect 13526 1321 13553 1355
rect 13565 1321 13599 1355
rect 13599 1321 13617 1355
rect 13501 1315 13553 1321
rect 13565 1315 13617 1321
rect 17939 1223 17991 1275
rect 18003 1223 18055 1275
rect 13805 1069 13857 1079
rect 13873 1069 13925 1079
rect 13941 1069 13993 1079
rect 13805 1035 13826 1069
rect 13826 1035 13857 1069
rect 13873 1035 13898 1069
rect 13898 1035 13925 1069
rect 13941 1035 13970 1069
rect 13970 1035 13993 1069
rect 13805 1027 13857 1035
rect 13873 1027 13925 1035
rect 13941 1027 13993 1035
rect 14008 1069 14060 1079
rect 14008 1035 14042 1069
rect 14042 1035 14060 1069
rect 14008 1027 14060 1035
rect 14075 1069 14127 1079
rect 14075 1035 14080 1069
rect 14080 1035 14114 1069
rect 14114 1035 14127 1069
rect 14075 1027 14127 1035
rect 14142 1069 14194 1079
rect 14142 1035 14152 1069
rect 14152 1035 14186 1069
rect 14186 1035 14194 1069
rect 14142 1027 14194 1035
rect 14209 1069 14261 1079
rect 14209 1035 14224 1069
rect 14224 1035 14258 1069
rect 14258 1035 14261 1069
rect 14209 1027 14261 1035
rect 14276 1069 14328 1079
rect 14343 1069 14395 1079
rect 14410 1069 14462 1079
rect 14477 1069 14529 1079
rect 14544 1069 14596 1079
rect 14611 1069 14663 1079
rect 14678 1069 14730 1079
rect 14745 1069 14797 1079
rect 14812 1069 14864 1079
rect 14879 1069 14931 1079
rect 14946 1069 14998 1079
rect 14276 1035 14296 1069
rect 14296 1035 14328 1069
rect 14343 1035 14368 1069
rect 14368 1035 14395 1069
rect 14410 1035 14440 1069
rect 14440 1035 14462 1069
rect 14477 1035 14512 1069
rect 14512 1035 14529 1069
rect 14544 1035 14546 1069
rect 14546 1035 14584 1069
rect 14584 1035 14596 1069
rect 14611 1035 14618 1069
rect 14618 1035 14656 1069
rect 14656 1035 14663 1069
rect 14678 1035 14690 1069
rect 14690 1035 14728 1069
rect 14728 1035 14730 1069
rect 14745 1035 14762 1069
rect 14762 1035 14797 1069
rect 14812 1035 14834 1069
rect 14834 1035 14864 1069
rect 14879 1035 14906 1069
rect 14906 1035 14931 1069
rect 14946 1035 14978 1069
rect 14978 1035 14998 1069
rect 14276 1027 14328 1035
rect 14343 1027 14395 1035
rect 14410 1027 14462 1035
rect 14477 1027 14529 1035
rect 14544 1027 14596 1035
rect 14611 1027 14663 1035
rect 14678 1027 14730 1035
rect 14745 1027 14797 1035
rect 14812 1027 14864 1035
rect 14879 1027 14931 1035
rect 14946 1027 14998 1035
rect 13289 833 13341 842
rect 13289 799 13322 833
rect 13322 799 13341 833
rect 13289 790 13341 799
rect 13354 833 13406 842
rect 13354 799 13360 833
rect 13360 799 13394 833
rect 13394 799 13406 833
rect 13354 790 13406 799
rect 13419 833 13471 842
rect 13419 799 13432 833
rect 13432 799 13466 833
rect 13466 799 13471 833
rect 13419 790 13471 799
rect 13484 833 13536 842
rect 13549 833 13601 842
rect 13614 833 13666 842
rect 13678 833 13730 842
rect 14484 833 14536 842
rect 14555 833 14607 842
rect 14626 833 14678 842
rect 14697 833 14749 842
rect 14768 833 14820 842
rect 14838 833 14890 842
rect 14908 833 14960 842
rect 13484 799 13504 833
rect 13504 799 13536 833
rect 13549 799 13576 833
rect 13576 799 13601 833
rect 13614 799 13648 833
rect 13648 799 13666 833
rect 13678 799 13682 833
rect 13682 799 13720 833
rect 13720 799 13730 833
rect 14484 799 14512 833
rect 14512 799 14536 833
rect 14555 799 14584 833
rect 14584 799 14607 833
rect 14626 799 14656 833
rect 14656 799 14678 833
rect 14697 799 14728 833
rect 14728 799 14749 833
rect 14768 799 14800 833
rect 14800 799 14820 833
rect 14838 799 14872 833
rect 14872 799 14890 833
rect 14908 799 14944 833
rect 14944 799 14960 833
rect 13484 790 13536 799
rect 13549 790 13601 799
rect 13614 790 13666 799
rect 13678 790 13730 799
rect 14484 790 14536 799
rect 14555 790 14607 799
rect 14626 790 14678 799
rect 14697 790 14749 799
rect 14768 790 14820 799
rect 14838 790 14890 799
rect 14908 790 14960 799
rect 13805 597 13857 606
rect 13876 597 13928 606
rect 13947 597 13999 606
rect 14018 597 14070 606
rect 14089 597 14141 606
rect 14159 597 14211 606
rect 14229 597 14281 606
rect 14299 597 14351 606
rect 13805 563 13826 597
rect 13826 563 13857 597
rect 13876 563 13898 597
rect 13898 563 13928 597
rect 13947 563 13970 597
rect 13970 563 13999 597
rect 14018 563 14042 597
rect 14042 563 14070 597
rect 14089 563 14114 597
rect 14114 563 14141 597
rect 14159 563 14186 597
rect 14186 563 14211 597
rect 14229 563 14258 597
rect 14258 563 14281 597
rect 14299 563 14330 597
rect 14330 563 14351 597
rect 13805 554 13857 563
rect 13876 554 13928 563
rect 13947 554 13999 563
rect 14018 554 14070 563
rect 14089 554 14141 563
rect 14159 554 14211 563
rect 14229 554 14281 563
rect 14299 554 14351 563
rect 15214 653 15266 671
rect 15214 619 15223 653
rect 15223 619 15257 653
rect 15257 619 15266 653
rect 15214 581 15266 597
rect 15214 547 15223 581
rect 15223 547 15257 581
rect 15257 547 15266 581
rect 15214 545 15266 547
rect 12758 464 12810 516
rect 12758 381 12810 433
rect 13289 361 13341 369
rect 12758 298 12810 350
rect 13289 327 13322 361
rect 13322 327 13341 361
rect 13289 317 13341 327
rect 13354 361 13406 369
rect 13354 327 13360 361
rect 13360 327 13394 361
rect 13394 327 13406 361
rect 13354 317 13406 327
rect 13419 361 13471 369
rect 13419 327 13432 361
rect 13432 327 13466 361
rect 13466 327 13471 361
rect 13419 317 13471 327
rect 13484 361 13536 369
rect 13549 361 13601 369
rect 13614 361 13666 369
rect 13678 361 13730 369
rect 14484 361 14536 369
rect 14555 361 14607 369
rect 14626 361 14678 369
rect 14697 361 14749 369
rect 14768 361 14820 369
rect 14838 361 14890 369
rect 14908 361 14960 369
rect 13484 327 13504 361
rect 13504 327 13536 361
rect 13549 327 13576 361
rect 13576 327 13601 361
rect 13614 327 13648 361
rect 13648 327 13666 361
rect 13678 327 13682 361
rect 13682 327 13720 361
rect 13720 327 13730 361
rect 14484 327 14512 361
rect 14512 327 14536 361
rect 14555 327 14584 361
rect 14584 327 14607 361
rect 14626 327 14656 361
rect 14656 327 14678 361
rect 14697 327 14728 361
rect 14728 327 14749 361
rect 14768 327 14800 361
rect 14800 327 14820 361
rect 14838 327 14872 361
rect 14872 327 14890 361
rect 14908 327 14944 361
rect 14944 327 14960 361
rect 13484 317 13536 327
rect 13549 317 13601 327
rect 13614 317 13666 327
rect 13678 317 13730 327
rect 14484 317 14536 327
rect 14555 317 14607 327
rect 14626 317 14678 327
rect 14697 317 14749 327
rect 14768 317 14820 327
rect 14838 317 14890 327
rect 14908 317 14960 327
rect 12097 122 12149 151
rect 12097 99 12105 122
rect 12105 99 12139 122
rect 12139 99 12149 122
rect 12097 50 12149 57
rect 12097 16 12105 50
rect 12105 16 12139 50
rect 12139 16 12149 50
rect 12097 5 12149 16
rect 12097 -56 12105 -38
rect 12105 -56 12139 -38
rect 12139 -56 12149 -38
rect 12097 -90 12149 -56
rect 13805 176 13857 228
rect 13876 176 13928 228
rect 13947 176 13999 228
rect 14018 176 14070 228
rect 14089 176 14141 228
rect 14159 176 14211 228
rect 14229 176 14281 228
rect 14299 176 14351 228
rect 12438 99 12490 151
rect 12520 122 12572 151
rect 12520 99 12561 122
rect 12561 99 12572 122
rect 12602 99 12654 151
rect 12684 146 12712 151
rect 12712 146 12736 151
rect 12684 104 12736 146
rect 12684 99 12712 104
rect 12712 99 12736 104
rect 12438 5 12490 57
rect 12520 50 12572 57
rect 12520 16 12561 50
rect 12561 16 12572 50
rect 12520 5 12572 16
rect 12602 5 12654 57
rect 12684 27 12736 57
rect 12684 5 12712 27
rect 12712 5 12736 27
rect 15214 509 15266 523
rect 15214 475 15223 509
rect 15223 475 15257 509
rect 15257 475 15266 509
rect 15214 471 15266 475
rect 15214 396 15266 448
rect 15214 321 15266 373
rect 15452 1038 15504 1061
rect 15452 1009 15459 1038
rect 15459 1009 15493 1038
rect 15493 1009 15504 1038
rect 15452 966 15504 996
rect 15452 944 15459 966
rect 15459 944 15493 966
rect 15493 944 15504 966
rect 15452 894 15504 931
rect 15452 879 15459 894
rect 15459 879 15493 894
rect 15493 879 15504 894
rect 15452 860 15459 866
rect 15459 860 15493 866
rect 15493 860 15504 866
rect 15452 814 15504 860
rect 15452 748 15504 800
rect 15687 653 15739 671
rect 15687 619 15695 653
rect 15695 619 15729 653
rect 15729 619 15739 653
rect 15687 581 15739 597
rect 15687 547 15695 581
rect 15695 547 15729 581
rect 15729 547 15739 581
rect 15687 545 15739 547
rect 15687 509 15739 523
rect 15687 475 15695 509
rect 15695 475 15729 509
rect 15729 475 15739 509
rect 15687 471 15739 475
rect 15687 396 15739 448
rect 15687 321 15739 373
rect 15924 1038 15976 1061
rect 15924 1009 15931 1038
rect 15931 1009 15965 1038
rect 15965 1009 15976 1038
rect 15924 966 15976 996
rect 15924 944 15931 966
rect 15931 944 15965 966
rect 15965 944 15976 966
rect 15924 894 15976 931
rect 15924 879 15931 894
rect 15931 879 15965 894
rect 15965 879 15976 894
rect 15924 860 15931 866
rect 15931 860 15965 866
rect 15965 860 15976 866
rect 15924 814 15976 860
rect 15924 748 15976 800
rect 16159 653 16211 671
rect 16159 619 16167 653
rect 16167 619 16201 653
rect 16201 619 16211 653
rect 16159 581 16211 597
rect 16159 547 16167 581
rect 16167 547 16201 581
rect 16201 547 16211 581
rect 16159 545 16211 547
rect 16159 509 16211 523
rect 16159 475 16167 509
rect 16167 475 16201 509
rect 16201 475 16211 509
rect 16159 471 16211 475
rect 16159 396 16211 448
rect 16159 321 16211 373
rect 15901 259 15953 268
rect 15901 225 15911 259
rect 15911 225 15945 259
rect 15945 225 15953 259
rect 15901 216 15953 225
rect 15971 259 16023 268
rect 15971 225 15983 259
rect 15983 225 16017 259
rect 16017 225 16023 259
rect 15971 216 16023 225
rect 12438 -90 12490 -38
rect 12520 -56 12561 -38
rect 12561 -56 12572 -38
rect 12520 -90 12572 -56
rect 12602 -90 12654 -38
rect 12684 -50 12736 -38
rect 12684 -84 12712 -50
rect 12712 -84 12736 -50
rect 12684 -90 12736 -84
rect 2227 -279 2279 -227
rect 2291 -279 2343 -227
rect 2132 -480 2184 -428
rect 2132 -544 2184 -492
rect 16187 109 16196 129
rect 16196 109 16230 129
rect 16230 109 16239 129
rect 16187 77 16239 109
rect 16187 37 16196 56
rect 16196 37 16230 56
rect 16230 37 16239 56
rect 16187 4 16239 37
rect 18013 1125 18065 1177
rect 18077 1125 18129 1177
rect 20519 1492 20571 1544
rect 20592 1492 20644 1544
rect 20665 1492 20717 1544
rect 20738 1492 20790 1544
rect 20810 1492 20862 1544
rect 20519 1422 20571 1474
rect 20592 1422 20644 1474
rect 20665 1422 20717 1474
rect 20738 1422 20790 1474
rect 20810 1422 20862 1474
rect 20519 1352 20571 1404
rect 20592 1352 20644 1404
rect 20665 1352 20717 1404
rect 20738 1352 20790 1404
rect 20810 1352 20862 1404
rect 25239 1530 25291 1542
rect 25239 1496 25243 1530
rect 25243 1496 25277 1530
rect 25277 1496 25291 1530
rect 25239 1490 25291 1496
rect 25303 1530 25355 1542
rect 25303 1496 25315 1530
rect 25315 1496 25349 1530
rect 25349 1496 25355 1530
rect 25303 1490 25355 1496
rect 20519 1282 20571 1334
rect 20592 1282 20644 1334
rect 20665 1282 20717 1334
rect 20738 1282 20790 1334
rect 20810 1282 20862 1334
rect 25239 1354 25291 1366
rect 25239 1320 25243 1354
rect 25243 1320 25277 1354
rect 25277 1320 25291 1354
rect 25239 1314 25291 1320
rect 25303 1354 25355 1366
rect 25303 1320 25315 1354
rect 25315 1320 25349 1354
rect 25349 1320 25355 1354
rect 25303 1314 25355 1320
rect 18128 1029 18180 1081
rect 18192 1029 18244 1081
rect 18537 346 18589 398
rect 18601 346 18653 398
rect 19161 230 19213 282
rect 19227 230 19279 282
rect 18362 -243 18414 -191
rect 18426 -243 18478 -191
rect 18522 -249 18574 -197
rect 18522 -313 18574 -261
rect 18862 -94 18914 -42
rect 18751 -172 18803 -120
rect 18751 -236 18803 -184
rect 2132 -1553 2184 -1501
rect 2132 -1632 2184 -1580
rect 2231 -1118 2283 -1066
rect 2295 -1118 2347 -1066
rect 16911 -1090 16963 -1038
rect 16975 -1090 17027 -1038
rect 17102 -1090 17154 -1038
rect 17166 -1090 17218 -1038
rect 17264 -1090 17316 -1038
rect 17328 -1090 17380 -1038
rect 2227 -1792 2279 -1740
rect 2227 -1856 2279 -1804
rect 692 -3484 744 -3432
rect 692 -3548 744 -3496
rect 1030 -4249 1082 -4233
rect 1030 -4283 1039 -4249
rect 1039 -4283 1073 -4249
rect 1073 -4283 1082 -4249
rect 1030 -4285 1082 -4283
rect 1030 -4321 1082 -4299
rect 1030 -4351 1039 -4321
rect 1039 -4351 1073 -4321
rect 1073 -4351 1082 -4321
rect 1030 -4393 1082 -4365
rect 1030 -4417 1039 -4393
rect 1039 -4417 1073 -4393
rect 1073 -4417 1082 -4393
rect 1697 -4281 1749 -4229
rect 1778 -4281 1830 -4229
rect 1859 -4281 1911 -4229
rect 1697 -4351 1749 -4299
rect 1778 -4351 1830 -4299
rect 1859 -4351 1911 -4299
rect 1697 -4421 1749 -4369
rect 1778 -4421 1830 -4369
rect 1859 -4421 1911 -4369
rect 2612 -9658 2624 -9625
rect 2624 -9658 2658 -9625
rect 2658 -9658 2664 -9625
rect 2612 -9677 2664 -9658
rect 2612 -9698 2664 -9689
rect 2612 -9732 2624 -9698
rect 2624 -9732 2658 -9698
rect 2658 -9732 2664 -9698
rect 2612 -9741 2664 -9732
rect 2771 -9772 2823 -9749
rect 2771 -9801 2780 -9772
rect 2780 -9801 2814 -9772
rect 2814 -9801 2823 -9772
rect 2771 -9846 2823 -9813
rect 2771 -9865 2780 -9846
rect 2780 -9865 2814 -9846
rect 2814 -9865 2823 -9846
rect 2647 -10232 2699 -10223
rect 2711 -10232 2763 -10223
rect 2647 -10266 2681 -10232
rect 2681 -10266 2699 -10232
rect 2711 -10266 2715 -10232
rect 2715 -10266 2763 -10232
rect 2647 -10275 2699 -10266
rect 2711 -10275 2763 -10266
rect 2389 -10920 2441 -10868
rect 2389 -10984 2441 -10932
rect 2473 -11003 2525 -10951
rect 2473 -11067 2525 -11015
rect 18862 -158 18914 -106
rect 3649 -11988 3701 -11936
rect 3558 -12071 3610 -12019
rect 3649 -12052 3701 -12000
rect 3558 -12135 3610 -12083
rect 19161 154 19213 206
rect 19227 154 19279 206
rect 3202 -14738 3254 -14686
rect 3202 -14802 3254 -14750
rect 3088 -17474 3140 -17422
rect 3088 -17540 3140 -17488
rect 3173 -17431 3225 -17425
rect 3173 -17465 3179 -17431
rect 3179 -17465 3213 -17431
rect 3213 -17465 3225 -17431
rect 3173 -17477 3225 -17465
rect 3173 -17503 3225 -17489
rect 3173 -17537 3179 -17503
rect 3179 -17537 3213 -17503
rect 3213 -17537 3225 -17503
rect 3173 -17541 3225 -17537
rect 2498 -18724 2550 -18672
rect 2562 -18678 2614 -18672
rect 2562 -18712 2580 -18678
rect 2580 -18712 2614 -18678
rect 2562 -18724 2614 -18712
rect 2561 -18846 2613 -18794
rect 2561 -18910 2613 -18858
<< metal2 >>
rect 357 4994 506 5029
rect 357 4942 454 4994
rect 357 4912 506 4942
rect 946 4926 8482 4978
rect 8534 4926 8548 4978
rect 8600 4926 8614 4978
rect 8666 4926 8680 4978
rect 8732 4926 8746 4978
rect 8798 4926 8811 4978
rect 8863 4926 8876 4978
rect 8928 4926 8941 4978
rect 8993 4926 9006 4978
rect 9058 4926 9071 4978
rect 9123 4926 9136 4978
rect 9188 4926 9201 4978
rect 9253 4926 9266 4978
rect 9318 4926 9331 4978
rect 9383 4926 9396 4978
rect 9448 4926 9461 4978
rect 9513 4926 9526 4978
rect 9578 4926 9591 4978
rect 9643 4926 9656 4978
rect 9708 4926 9721 4978
rect 9773 4926 9786 4978
rect 9838 4926 9851 4978
rect 9903 4926 9916 4978
rect 9968 4926 9981 4978
rect 10033 4926 10046 4978
rect 10098 4926 10111 4978
rect 10163 4926 10176 4978
rect 10228 4926 10241 4978
rect 10293 4926 10306 4978
rect 10358 4926 10371 4978
rect 10423 4926 10436 4978
rect 10488 4926 10501 4978
rect 10553 4926 10566 4978
rect 10618 4926 10631 4978
rect 10683 4926 10696 4978
rect 10748 4926 10761 4978
rect 10813 4926 10826 4978
rect 10878 4926 10891 4978
rect 10943 4926 10956 4978
rect 11008 4926 11021 4978
rect 11073 4926 11086 4978
rect 11138 4926 11151 4978
rect 11203 4926 11216 4978
rect 11268 4926 11281 4978
rect 11333 4926 11346 4978
rect 11398 4926 11411 4978
rect 11463 4970 11707 4978
rect 11463 4926 11515 4970
rect 946 4918 11515 4926
rect 11567 4918 11580 4970
rect 11632 4918 11644 4970
rect 11696 4918 11707 4970
rect 357 4860 454 4912
rect 569 4865 575 4917
rect 627 4865 639 4917
rect 691 4865 697 4917
tri 577 4860 582 4865 ne
rect 582 4860 692 4865
tri 692 4860 697 4865 nw
rect 946 4908 11707 4918
rect 19753 4970 20024 4978
rect 19753 4918 19755 4970
rect 19807 4918 19819 4970
rect 19871 4918 19883 4970
rect 19935 4918 19947 4970
rect 19999 4918 20024 4970
rect 946 4860 8482 4908
rect 357 4830 506 4860
tri 582 4831 611 4860 ne
rect 357 4778 454 4830
rect 357 4748 506 4778
rect 357 4696 454 4748
rect 357 4666 506 4696
rect 357 4614 454 4666
rect 357 4584 506 4614
rect 357 4532 454 4584
rect 357 4502 506 4532
rect 357 4450 454 4502
rect 357 4420 506 4450
rect 357 4368 454 4420
rect 357 4338 506 4368
rect 611 4389 663 4860
tri 663 4831 692 4860 nw
rect 946 4831 6964 4860
rect 946 4824 1210 4831
rect 946 4772 952 4824
rect 1004 4772 1044 4824
rect 1096 4772 1135 4824
rect 1187 4779 1210 4824
rect 1262 4779 1279 4831
rect 1331 4779 1348 4831
rect 1400 4779 1417 4831
rect 1469 4779 1486 4831
rect 1538 4779 1554 4831
rect 1606 4779 1622 4831
rect 1674 4779 1690 4831
rect 1742 4779 1758 4831
rect 1810 4779 1826 4831
rect 1878 4779 1894 4831
rect 1946 4779 1962 4831
rect 2014 4819 6964 4831
rect 2014 4779 2486 4819
rect 1187 4772 2486 4779
rect 946 4767 2486 4772
rect 2538 4767 2998 4819
rect 3050 4767 3510 4819
rect 3562 4767 4022 4819
rect 4074 4767 4534 4819
rect 4586 4767 5046 4819
rect 5098 4767 5558 4819
rect 5610 4767 6070 4819
rect 6122 4767 6582 4819
rect 6634 4808 6964 4819
rect 7016 4808 7029 4860
rect 7081 4808 7094 4860
rect 7146 4808 7158 4860
rect 7210 4808 7222 4860
rect 7274 4808 7286 4860
rect 7338 4808 7350 4860
rect 7402 4808 7414 4860
rect 7466 4808 7478 4860
rect 7530 4856 8482 4860
rect 8534 4856 8548 4908
rect 8600 4856 8614 4908
rect 8666 4856 8680 4908
rect 8732 4856 8746 4908
rect 8798 4856 8811 4908
rect 8863 4856 8876 4908
rect 8928 4856 8941 4908
rect 8993 4856 9006 4908
rect 9058 4856 9071 4908
rect 9123 4856 9136 4908
rect 9188 4856 9201 4908
rect 9253 4856 9266 4908
rect 9318 4856 9331 4908
rect 9383 4856 9396 4908
rect 9448 4856 9461 4908
rect 9513 4856 9526 4908
rect 9578 4856 9591 4908
rect 9643 4856 9656 4908
rect 9708 4856 9721 4908
rect 9773 4856 9786 4908
rect 9838 4856 9851 4908
rect 9903 4856 9916 4908
rect 9968 4856 9981 4908
rect 10033 4856 10046 4908
rect 10098 4856 10111 4908
rect 10163 4856 10176 4908
rect 10228 4856 10241 4908
rect 10293 4856 10306 4908
rect 10358 4856 10371 4908
rect 10423 4856 10436 4908
rect 10488 4856 10501 4908
rect 10553 4856 10566 4908
rect 10618 4856 10631 4908
rect 10683 4856 10696 4908
rect 10748 4856 10761 4908
rect 10813 4856 10826 4908
rect 10878 4856 10891 4908
rect 10943 4856 10956 4908
rect 11008 4856 11021 4908
rect 11073 4856 11086 4908
rect 11138 4856 11151 4908
rect 11203 4856 11216 4908
rect 11268 4856 11281 4908
rect 11333 4856 11346 4908
rect 11398 4856 11411 4908
rect 11463 4876 11707 4908
rect 11463 4856 11515 4876
rect 7530 4825 11515 4856
rect 7530 4808 7712 4825
rect 6634 4773 7712 4808
rect 7764 4773 7820 4825
rect 7872 4824 11515 4825
rect 11567 4824 11580 4876
rect 11632 4824 11644 4876
rect 11696 4824 11707 4876
rect 18720 4852 18729 4908
rect 18785 4852 18809 4908
rect 18865 4852 18874 4908
tri 14379 4827 14381 4829 se
rect 14381 4827 16586 4829
tri 16586 4827 16588 4829 sw
rect 18720 4827 18849 4852
tri 18849 4827 18874 4852 nw
rect 19753 4879 20024 4918
rect 19753 4827 19755 4879
rect 19807 4827 19819 4879
rect 19871 4827 19883 4879
rect 19935 4827 19947 4879
rect 19999 4827 20024 4879
rect 7872 4809 11707 4824
tri 14373 4821 14379 4827 se
rect 14379 4821 16588 4827
tri 16588 4821 16594 4827 sw
rect 7872 4806 11184 4809
rect 7872 4773 8473 4806
rect 6634 4767 8473 4773
rect 946 4755 8473 4767
rect 946 4753 2486 4755
rect 946 4744 1210 4753
rect 946 4692 952 4744
rect 1004 4692 1044 4744
rect 1096 4692 1135 4744
rect 1187 4701 1210 4744
rect 1262 4701 1279 4753
rect 1331 4701 1348 4753
rect 1400 4701 1417 4753
rect 1469 4701 1486 4753
rect 1538 4701 1554 4753
rect 1606 4701 1622 4753
rect 1674 4701 1690 4753
rect 1742 4701 1758 4753
rect 1810 4701 1826 4753
rect 1878 4701 1894 4753
rect 1946 4701 1962 4753
rect 2014 4703 2486 4753
rect 2538 4703 2998 4755
rect 3050 4703 3510 4755
rect 3562 4703 4022 4755
rect 4074 4703 4534 4755
rect 4586 4703 5046 4755
rect 5098 4703 5558 4755
rect 5610 4703 6070 4755
rect 6122 4703 6582 4755
rect 6634 4754 8473 4755
rect 8525 4754 8861 4806
rect 8913 4754 9609 4806
rect 9661 4754 9889 4806
rect 9941 4754 10322 4806
rect 10374 4754 10634 4806
rect 10686 4754 10946 4806
rect 10998 4757 11184 4806
rect 11236 4807 11707 4809
rect 11236 4757 11290 4807
rect 10998 4755 11290 4757
rect 11342 4782 11707 4807
tri 14340 4788 14373 4821 se
rect 14373 4793 16594 4821
rect 14373 4788 14392 4793
tri 14392 4788 14397 4793 nw
tri 16570 4788 16575 4793 ne
rect 16575 4788 16594 4793
tri 16594 4788 16627 4821 sw
rect 11342 4755 11515 4782
rect 10998 4754 11515 4755
rect 6634 4750 11515 4754
rect 6634 4703 6964 4750
rect 2014 4701 6964 4703
rect 1187 4698 6964 4701
rect 7016 4698 7029 4750
rect 7081 4698 7094 4750
rect 7146 4698 7158 4750
rect 7210 4698 7222 4750
rect 7274 4698 7286 4750
rect 7338 4698 7350 4750
rect 7402 4698 7414 4750
rect 7466 4698 7478 4750
rect 7530 4749 11515 4750
rect 7530 4698 7712 4749
rect 1187 4697 7712 4698
rect 7764 4697 7820 4749
rect 7872 4730 11515 4749
rect 11567 4730 11580 4782
rect 11632 4730 11644 4782
rect 11696 4730 11707 4782
tri 14329 4777 14340 4788 se
rect 14340 4777 14381 4788
tri 14381 4777 14392 4788 nw
tri 16575 4777 16586 4788 ne
rect 16586 4777 16627 4788
tri 14321 4769 14329 4777 se
rect 14329 4769 14373 4777
tri 14373 4769 14381 4777 nw
tri 16586 4769 16594 4777 ne
rect 16594 4769 16627 4777
tri 16627 4769 16646 4788 sw
tri 14313 4761 14321 4769 se
rect 14321 4761 14365 4769
tri 14365 4761 14373 4769 nw
tri 16594 4761 16602 4769 ne
rect 16602 4761 16646 4769
tri 16646 4761 16654 4769 sw
tri 14291 4739 14313 4761 se
rect 14313 4739 14343 4761
tri 14343 4739 14365 4761 nw
tri 14389 4739 14411 4761 se
rect 14411 4739 16556 4761
tri 16556 4739 16578 4761 sw
tri 16602 4739 16624 4761 ne
rect 16624 4739 16654 4761
tri 16654 4739 16676 4761 sw
tri 14288 4736 14291 4739 se
rect 14291 4736 14340 4739
tri 14340 4736 14343 4739 nw
tri 14386 4736 14389 4739 se
rect 14389 4736 16578 4739
tri 16578 4736 16581 4739 sw
tri 16624 4736 16627 4739 ne
rect 16627 4736 16676 4739
tri 16676 4736 16679 4739 sw
tri 14282 4730 14288 4736 se
rect 14288 4731 14335 4736
tri 14335 4731 14340 4736 nw
tri 14381 4731 14386 4736 se
rect 14386 4731 16581 4736
rect 14288 4730 14334 4731
tri 14334 4730 14335 4731 nw
tri 14380 4730 14381 4731 se
rect 14381 4730 16581 4731
tri 16581 4730 16587 4736 sw
tri 16627 4730 16633 4736 ne
rect 16633 4730 16679 4736
tri 16679 4730 16685 4736 sw
rect 7872 4723 11707 4730
tri 14277 4725 14282 4730 se
rect 14282 4725 14329 4730
tri 14329 4725 14334 4730 nw
tri 14375 4725 14380 4730 se
rect 14380 4725 16587 4730
rect 7872 4697 8473 4723
rect 1187 4692 1235 4697
rect 946 4671 1235 4692
tri 1235 4671 1261 4697 nw
tri 1382 4671 1408 4697 ne
rect 1408 4671 1452 4697
tri 1452 4671 1478 4697 nw
tri 7927 4671 7953 4697 ne
rect 7953 4671 8473 4697
rect 8525 4671 8861 4723
rect 8913 4671 9609 4723
rect 9661 4671 9889 4723
rect 9941 4671 10322 4723
rect 10374 4671 10634 4723
rect 10686 4671 10946 4723
rect 10998 4671 11184 4723
rect 11236 4721 11707 4723
rect 11236 4671 11290 4721
rect 946 4669 1233 4671
tri 1233 4669 1235 4671 nw
tri 1408 4669 1410 4671 ne
rect 1410 4669 1450 4671
tri 1450 4669 1452 4671 nw
tri 7953 4669 7955 4671 ne
rect 7955 4669 11290 4671
rect 11342 4720 11707 4721
tri 14272 4720 14277 4725 se
rect 14277 4720 14313 4725
rect 11342 4709 11405 4720
tri 11405 4709 11416 4720 nw
tri 14261 4709 14272 4720 se
rect 14272 4709 14313 4720
tri 14313 4709 14329 4725 nw
tri 14359 4709 14375 4725 se
rect 14375 4709 14411 4725
tri 14411 4709 14427 4725 nw
tri 16540 4709 16556 4725 ne
rect 16556 4723 16587 4725
tri 16587 4723 16594 4730 sw
tri 16633 4723 16640 4730 ne
rect 16640 4723 16685 4730
rect 16556 4717 16594 4723
tri 16594 4717 16600 4723 sw
tri 16640 4717 16646 4723 ne
rect 16646 4717 16685 4723
tri 16685 4717 16698 4730 sw
rect 16556 4709 16600 4717
rect 11342 4693 11389 4709
tri 11389 4693 11405 4709 nw
tri 14245 4693 14261 4709 se
rect 14261 4693 14297 4709
tri 14297 4693 14313 4709 nw
tri 14343 4693 14359 4709 se
rect 14359 4693 14395 4709
tri 14395 4693 14411 4709 nw
tri 16556 4693 16572 4709 ne
rect 16572 4693 16600 4709
tri 16600 4693 16624 4717 sw
tri 16646 4693 16670 4717 ne
rect 16670 4693 16698 4717
tri 16698 4693 16722 4717 sw
rect 11342 4686 11382 4693
tri 11382 4686 11389 4693 nw
tri 14238 4686 14245 4693 se
rect 14245 4686 14290 4693
tri 14290 4686 14297 4693 nw
tri 14336 4686 14343 4693 se
rect 14343 4686 14388 4693
tri 14388 4686 14395 4693 nw
tri 14434 4686 14441 4693 se
rect 14441 4692 16526 4693
tri 16526 4692 16527 4693 sw
tri 16572 4692 16573 4693 ne
rect 16573 4692 16624 4693
tri 16624 4692 16625 4693 sw
tri 16670 4692 16671 4693 ne
rect 16671 4692 16722 4693
tri 16722 4692 16723 4693 sw
rect 14441 4687 16527 4692
tri 16527 4687 16532 4692 sw
tri 16573 4687 16578 4692 ne
rect 16578 4687 16625 4692
tri 16625 4687 16630 4692 sw
tri 16671 4687 16676 4692 ne
rect 16676 4687 16723 4692
tri 16723 4687 16728 4692 sw
rect 14441 4686 16532 4687
tri 16532 4686 16533 4687 sw
tri 16578 4686 16579 4687 ne
rect 16579 4686 16630 4687
tri 16630 4686 16631 4687 sw
tri 16676 4686 16677 4687 ne
rect 16677 4686 16728 4687
tri 16728 4686 16729 4687 sw
rect 11342 4673 11369 4686
tri 11369 4673 11382 4686 nw
tri 14225 4673 14238 4686 se
rect 14238 4679 14283 4686
tri 14283 4679 14290 4686 nw
tri 14329 4679 14336 4686 se
rect 14336 4679 14374 4686
rect 14238 4673 14277 4679
tri 14277 4673 14283 4679 nw
tri 14323 4673 14329 4679 se
rect 14329 4673 14374 4679
rect 11342 4672 11368 4673
tri 11368 4672 11369 4673 nw
tri 14224 4672 14225 4673 se
rect 14225 4672 14276 4673
tri 14276 4672 14277 4673 nw
tri 14322 4672 14323 4673 se
rect 14323 4672 14374 4673
tri 14374 4672 14388 4686 nw
tri 14420 4672 14434 4686 se
rect 14434 4672 16533 4686
tri 16533 4672 16547 4686 sw
tri 16579 4672 16593 4686 ne
rect 16593 4672 16631 4686
tri 16631 4672 16645 4686 sw
tri 16677 4672 16691 4686 ne
rect 16691 4672 16729 4686
tri 16729 4672 16743 4686 sw
rect 11342 4669 11359 4672
rect 946 4667 1231 4669
tri 1231 4667 1233 4669 nw
tri 1410 4667 1412 4669 ne
rect 1412 4667 1448 4669
tri 1448 4667 1450 4669 nw
tri 7955 4667 7957 4669 ne
rect 7957 4667 11359 4669
rect 946 4664 1193 4667
rect 946 4612 952 4664
rect 1004 4612 1044 4664
rect 1096 4612 1135 4664
rect 1187 4612 1193 4664
tri 1193 4629 1231 4667 nw
tri 1412 4663 1416 4667 ne
rect 787 4529 793 4581
rect 845 4529 857 4581
rect 909 4529 915 4581
tri 829 4498 860 4529 ne
rect 860 4498 915 4529
tri 860 4497 861 4498 ne
rect 861 4497 915 4498
tri 861 4495 863 4497 ne
tri 663 4389 669 4395 sw
rect 611 4365 669 4389
tri 669 4365 693 4389 sw
tri 611 4361 615 4365 ne
rect 615 4361 693 4365
tri 693 4361 697 4365 sw
tri 615 4355 621 4361 ne
rect 621 4355 697 4361
tri 697 4355 703 4361 sw
tri 621 4343 633 4355 ne
rect 633 4343 703 4355
tri 703 4343 715 4355 sw
rect 357 4286 454 4338
tri 633 4337 639 4343 ne
rect 639 4337 715 4343
tri 715 4337 721 4343 sw
tri 639 4307 669 4337 ne
rect 669 4307 721 4337
tri 721 4307 751 4337 sw
rect 357 4256 506 4286
tri 669 4285 691 4307 ne
rect 691 4285 751 4307
tri 751 4285 773 4307 sw
tri 691 4270 706 4285 ne
rect 706 4270 773 4285
tri 773 4270 788 4285 sw
tri 706 4258 718 4270 ne
rect 718 4258 788 4270
tri 788 4258 800 4270 sw
rect 357 4204 454 4256
tri 718 4250 726 4258 ne
rect 726 4250 800 4258
tri 800 4250 808 4258 sw
tri 726 4247 729 4250 ne
rect 729 4247 808 4250
tri 808 4247 811 4250 sw
tri 729 4225 751 4247 ne
rect 751 4225 811 4247
tri 811 4225 833 4247 sw
rect 357 4174 506 4204
tri 751 4195 781 4225 ne
rect 357 4122 454 4174
rect 357 4092 506 4122
rect 357 4040 454 4092
rect 699 4161 751 4167
rect 699 4097 751 4109
rect 357 4010 506 4040
rect 357 3958 454 4010
rect 357 3928 506 3958
rect 357 3876 454 3928
rect 357 3846 506 3876
rect 357 3794 454 3846
rect 357 3764 506 3794
rect 357 3712 454 3764
rect 357 3681 506 3712
rect 357 3629 454 3681
rect 357 3598 506 3629
rect 617 4057 669 4063
rect 617 3993 669 4005
rect 357 3546 454 3598
rect 357 3515 506 3546
rect 357 3463 454 3515
rect 357 3432 506 3463
rect 357 3380 454 3432
rect 357 3349 506 3380
rect 357 3297 454 3349
rect 357 3266 506 3297
rect 357 3214 454 3266
rect 357 3183 506 3214
rect 357 3131 454 3183
rect 357 3100 506 3131
rect 357 3048 454 3100
rect 357 2450 506 3048
rect 357 2398 454 2450
rect 357 2370 506 2398
rect 357 2318 454 2370
rect 357 2290 506 2318
rect 357 2238 454 2290
rect 357 2210 506 2238
rect 357 2158 454 2210
rect 357 2130 506 2158
rect 357 2078 454 2130
rect 357 2050 506 2078
rect 357 1998 454 2050
rect 357 1970 506 1998
rect 357 1918 454 1970
rect 357 1890 506 1918
rect 357 1838 454 1890
rect 357 1810 506 1838
rect 357 1758 454 1810
rect 357 1730 506 1758
rect 357 1678 454 1730
rect 357 1650 506 1678
rect 357 1598 454 1650
rect 357 1570 506 1598
rect 357 1518 454 1570
rect 357 1490 506 1518
rect 357 1438 454 1490
rect 357 1410 506 1438
rect 357 1358 454 1410
rect 357 1330 506 1358
rect 357 1278 454 1330
rect 357 1250 506 1278
rect 357 1198 454 1250
rect 357 1170 506 1198
rect 357 1118 454 1170
rect 357 1090 506 1118
rect 357 1038 454 1090
rect 357 1010 506 1038
rect 357 958 454 1010
rect 357 930 506 958
rect 357 878 454 930
rect 357 850 506 878
rect 357 798 454 850
rect 357 770 506 798
rect 357 718 454 770
rect 357 690 506 718
rect 357 638 454 690
rect 357 610 506 638
rect 357 558 454 610
rect 357 530 506 558
rect 357 478 454 530
rect 357 450 506 478
rect 357 398 454 450
rect 357 370 506 398
rect 357 318 454 370
rect 357 290 506 318
rect 357 238 454 290
rect 357 210 506 238
rect 357 158 454 210
rect 357 130 506 158
rect 357 78 454 130
rect 357 50 506 78
rect 357 -2 454 50
rect 357 -30 506 -2
rect 357 -82 454 -30
rect 357 -110 506 -82
rect 357 -162 454 -110
rect 357 -190 506 -162
rect 357 -242 454 -190
rect 357 -270 506 -242
rect 357 -322 454 -270
rect 357 -350 506 -322
rect 357 -402 454 -350
rect 357 -430 506 -402
rect 357 -482 454 -430
rect 357 -510 506 -482
rect 357 -562 454 -510
rect 357 -590 506 -562
rect 357 -642 454 -590
rect 357 -670 506 -642
rect 357 -722 454 -670
rect 357 -750 506 -722
rect 357 -802 454 -750
rect 357 -830 506 -802
rect 357 -882 454 -830
rect 357 -910 506 -882
rect 357 -962 454 -910
rect 357 -990 506 -962
rect 357 -1042 454 -990
rect 535 3617 587 3623
rect 535 3553 587 3565
rect 535 -237 587 3501
rect 535 -307 587 -289
rect 535 -917 587 -359
rect 617 230 669 3941
rect 699 699 751 4045
rect 699 629 751 647
rect 699 571 751 577
rect 781 3229 833 4225
rect 781 3165 833 3177
rect 781 1167 833 3113
rect 863 3143 915 4497
rect 946 4497 1193 4612
rect 946 4445 952 4497
rect 1004 4445 1044 4497
rect 1096 4445 1135 4497
rect 1187 4445 1193 4497
rect 946 4417 1193 4445
rect 946 4365 952 4417
rect 1004 4365 1044 4417
rect 1096 4365 1135 4417
rect 1187 4365 1193 4417
rect 946 4337 1193 4365
rect 946 4285 952 4337
rect 1004 4285 1044 4337
rect 1096 4285 1135 4337
rect 1187 4285 1193 4337
rect 946 3815 1193 4285
rect 1258 4027 1264 4079
rect 1316 4027 1328 4079
rect 1380 4027 1386 4079
tri 1258 4022 1263 4027 ne
rect 946 3763 952 3815
rect 1004 3763 1044 3815
rect 1096 3763 1135 3815
rect 1187 3763 1193 3815
rect 946 3735 1193 3763
rect 946 3683 952 3735
rect 1004 3683 1044 3735
rect 1096 3683 1135 3735
rect 1187 3683 1193 3735
rect 946 3655 1193 3683
rect 946 3603 952 3655
rect 1004 3603 1044 3655
rect 1096 3603 1135 3655
rect 1187 3603 1193 3655
rect 946 3489 1193 3603
rect 1263 3604 1386 4027
tri 1263 3601 1266 3604 ne
rect 1266 3601 1386 3604
tri 1266 3551 1316 3601 ne
rect 1316 3551 1386 3601
tri 1316 3533 1334 3551 ne
rect 946 3437 952 3489
rect 1004 3437 1044 3489
rect 1096 3437 1135 3489
rect 1187 3437 1193 3489
rect 946 3425 1193 3437
rect 946 3373 952 3425
rect 1004 3373 1044 3425
rect 1096 3373 1135 3425
rect 1187 3373 1193 3425
rect 863 3079 915 3091
rect 863 2901 915 3027
rect 1102 2975 1232 2981
tri 915 2901 940 2926 sw
tri 863 2895 869 2901 ne
rect 869 2895 940 2901
tri 940 2895 946 2901 sw
rect 1017 2895 1069 2901
tri 869 2856 908 2895 ne
rect 908 2856 946 2895
tri 946 2856 985 2895 sw
tri 908 2849 915 2856 ne
rect 915 2849 985 2856
tri 915 2843 921 2849 ne
rect 921 2843 985 2849
tri 921 2831 933 2843 ne
rect 933 2831 985 2843
tri 933 2819 945 2831 ne
rect 781 1097 833 1115
tri 777 540 781 544 se
rect 781 540 833 1045
rect 777 531 833 540
rect 777 451 833 475
rect 777 386 833 395
rect 863 2739 915 2745
rect 863 2675 915 2687
rect 863 2617 915 2623
rect 617 160 669 178
rect 617 -93 669 108
rect 701 300 707 352
rect 759 300 771 352
rect 823 300 829 352
rect 701 40 829 300
rect 701 -12 707 40
rect 759 -12 771 40
rect 823 -12 829 40
rect 701 -28 829 -12
tri 741 -44 757 -28 ne
rect 757 -44 829 -28
tri 757 -46 759 -44 ne
rect 759 -46 829 -44
tri 759 -53 766 -46 ne
rect 766 -53 829 -46
tri 766 -60 773 -53 ne
rect 773 -60 829 -53
tri 773 -64 777 -60 ne
rect 617 -719 663 -93
tri 663 -99 669 -93 nw
rect 693 -125 745 -119
rect 693 -189 745 -177
rect 693 -358 745 -241
rect 693 -422 745 -410
rect 693 -682 745 -474
tri 693 -688 699 -682 ne
tri 663 -719 667 -715 sw
rect 617 -721 667 -719
tri 667 -721 669 -719 sw
rect 617 -727 669 -721
rect 617 -791 669 -779
rect 617 -849 669 -843
tri 693 -896 699 -890 se
rect 699 -896 745 -682
tri 587 -917 593 -911 sw
rect 535 -941 593 -917
tri 593 -941 617 -917 sw
rect 535 -957 617 -941
tri 617 -957 633 -941 sw
rect 535 -1009 541 -957
rect 593 -1009 605 -957
rect 657 -1009 663 -957
rect 357 -1070 506 -1042
rect 357 -1122 454 -1070
rect 357 -1150 506 -1122
rect 357 -1202 454 -1150
rect 357 -1230 506 -1202
rect 357 -1282 454 -1230
rect 357 -1310 506 -1282
rect 357 -1362 454 -1310
rect 357 -1390 506 -1362
rect 357 -1442 454 -1390
rect 357 -1470 506 -1442
rect 357 -1522 454 -1470
rect 357 -1550 506 -1522
rect 357 -1602 454 -1550
rect 357 -1630 506 -1602
rect 357 -1682 454 -1630
rect 357 -1710 506 -1682
rect 357 -1762 454 -1710
rect 357 -1790 506 -1762
rect 357 -1842 454 -1790
rect 357 -1870 506 -1842
rect 357 -1922 454 -1870
rect 357 -1950 506 -1922
rect 357 -2002 454 -1950
rect 357 -2031 506 -2002
rect 357 -2083 454 -2031
rect 357 -2112 506 -2083
rect 357 -2164 454 -2112
rect 357 -2170 506 -2164
rect 693 -2085 745 -896
rect 777 -1769 829 -60
rect 777 -1833 829 -1821
rect 777 -1891 829 -1885
tri 859 256 863 260 se
rect 863 256 911 2617
tri 911 2613 915 2617 nw
rect 859 232 911 256
rect 859 -2010 907 232
tri 907 228 911 232 nw
tri 941 -657 945 -653 se
rect 945 -657 985 2831
rect 1017 2831 1069 2843
tri 937 -661 941 -657 se
rect 941 -661 985 -657
tri 985 -661 989 -657 sw
rect 937 -667 989 -661
rect 937 -731 989 -719
rect 937 -789 989 -783
tri 1011 -1076 1017 -1070 se
rect 1017 -1076 1069 2779
rect 1102 2859 1116 2975
rect 1102 2530 1232 2859
tri 1232 2530 1233 2531 sw
rect 1102 2508 1233 2530
tri 1233 2508 1255 2530 sw
rect 1102 2507 1255 2508
tri 1255 2507 1256 2508 sw
rect 1102 2451 1111 2507
rect 1167 2451 1191 2507
rect 1247 2451 1256 2507
rect 1102 2436 1241 2451
tri 1241 2436 1256 2451 nw
rect 1334 2436 1386 3551
rect 1416 2468 1444 4667
tri 1444 4663 1448 4667 nw
tri 1492 4663 1496 4667 se
rect 1496 4663 2045 4667
tri 1475 4646 1492 4663 se
rect 1492 4646 2045 4663
rect 1475 4615 2045 4646
rect 2097 4615 2118 4667
rect 2170 4615 2336 4667
rect 2388 4615 2413 4667
rect 2465 4615 2490 4667
rect 2542 4615 2567 4667
rect 2619 4615 2644 4667
rect 2696 4615 2831 4667
rect 2883 4615 2898 4667
rect 2950 4615 2965 4667
rect 3017 4615 3031 4667
rect 3083 4615 3097 4667
rect 3149 4615 3163 4667
rect 3215 4615 3570 4667
rect 3622 4615 3679 4667
rect 3731 4615 3852 4667
rect 3904 4615 3921 4667
rect 3973 4615 3990 4667
rect 4042 4615 4058 4667
rect 4110 4615 4126 4667
rect 4178 4615 4194 4667
rect 4246 4615 4365 4667
rect 4417 4615 4433 4667
rect 4485 4615 4501 4667
rect 4553 4615 4569 4667
rect 4621 4615 4636 4667
rect 4688 4615 4703 4667
rect 4755 4615 4875 4667
rect 4927 4615 4941 4667
rect 4993 4615 5007 4667
rect 5059 4615 5073 4667
rect 5125 4615 5139 4667
rect 5191 4615 5205 4667
rect 5257 4615 5271 4667
rect 5323 4615 5337 4667
rect 5389 4615 5403 4667
rect 5455 4615 5469 4667
rect 5521 4615 5535 4667
rect 5587 4615 5601 4667
rect 5653 4615 5667 4667
rect 5719 4615 5732 4667
rect 5784 4615 5797 4667
rect 5849 4615 5862 4667
rect 5914 4615 5927 4667
rect 5979 4615 5992 4667
rect 6044 4615 6057 4667
rect 6109 4615 6122 4667
rect 6174 4615 6187 4667
rect 6239 4615 6252 4667
rect 6304 4615 6317 4667
rect 6369 4615 6382 4667
rect 6434 4615 6447 4667
rect 6499 4615 6512 4667
rect 6564 4615 6577 4667
rect 6629 4615 6642 4667
rect 6694 4615 6707 4667
rect 6759 4615 6772 4667
rect 6824 4615 6830 4667
tri 7957 4665 7959 4667 ne
rect 7959 4665 11359 4667
tri 11288 4663 11290 4665 ne
rect 11290 4663 11359 4665
tri 11359 4663 11368 4672 nw
tri 14215 4663 14224 4672 se
rect 14224 4663 14267 4672
tri 14267 4663 14276 4672 nw
tri 14313 4663 14322 4672 se
rect 14322 4663 14365 4672
tri 14365 4663 14374 4672 nw
tri 14411 4663 14420 4672 se
rect 14420 4663 16547 4672
tri 16547 4663 16556 4672 sw
tri 16593 4663 16602 4672 ne
rect 16602 4671 16645 4672
tri 16645 4671 16646 4672 sw
tri 16691 4671 16692 4672 ne
rect 16692 4671 16743 4672
rect 16602 4665 16646 4671
tri 16646 4665 16652 4671 sw
tri 16692 4665 16698 4671 ne
rect 16698 4665 16743 4671
tri 16743 4665 16750 4672 sw
rect 16602 4663 16652 4665
tri 16652 4663 16654 4665 sw
tri 16698 4663 16700 4665 ne
rect 16700 4663 16750 4665
tri 16750 4663 16752 4665 sw
tri 14209 4657 14215 4663 se
rect 14215 4657 14261 4663
tri 14261 4657 14267 4663 nw
tri 14307 4657 14313 4663 se
rect 14313 4657 14359 4663
tri 14359 4657 14365 4663 nw
tri 14405 4657 14411 4663 se
rect 14411 4657 16556 4663
tri 16556 4657 16562 4663 sw
tri 16602 4657 16608 4663 ne
rect 16608 4657 16654 4663
tri 16654 4657 16660 4663 sw
tri 16700 4657 16706 4663 ne
rect 16706 4657 16752 4663
tri 16752 4657 16758 4663 sw
tri 14197 4645 14209 4657 se
rect 14209 4645 14249 4657
tri 14249 4645 14261 4657 nw
tri 14295 4645 14307 4657 se
rect 14307 4645 14347 4657
tri 14347 4645 14359 4657 nw
tri 14393 4645 14405 4657 se
rect 14405 4645 14442 4657
tri 11597 4625 11617 4645 se
rect 11617 4625 11671 4645
rect 1475 4614 1551 4615
tri 1551 4614 1552 4615 nw
rect 8103 4614 8155 4620
rect 1475 4498 1527 4614
tri 1527 4590 1551 4614 nw
rect 8209 4573 8215 4625
rect 8267 4573 8279 4625
rect 8331 4593 11671 4625
rect 11723 4593 11735 4645
rect 11787 4593 11793 4645
tri 13027 4642 13030 4645 se
rect 13030 4642 14246 4645
tri 14246 4642 14249 4645 nw
tri 14292 4642 14295 4645 se
rect 14295 4642 14344 4645
tri 14344 4642 14347 4645 nw
tri 14390 4642 14393 4645 se
rect 14393 4642 14442 4645
tri 14442 4642 14457 4657 nw
tri 16510 4642 16525 4657 ne
rect 16525 4645 16562 4657
tri 16562 4645 16574 4657 sw
tri 16608 4645 16620 4657 ne
rect 16620 4645 16660 4657
tri 16660 4645 16672 4657 sw
tri 16706 4645 16718 4657 ne
rect 16718 4645 16758 4657
tri 16758 4645 16770 4657 sw
rect 16525 4642 16574 4645
tri 16574 4642 16577 4645 sw
tri 16620 4642 16623 4645 ne
rect 16623 4642 16672 4645
tri 16672 4642 16675 4645 sw
tri 16718 4642 16721 4645 ne
rect 16721 4642 16770 4645
tri 16770 4642 16773 4645 sw
tri 13026 4641 13027 4642 se
rect 13027 4641 14245 4642
tri 14245 4641 14246 4642 nw
tri 14291 4641 14292 4642 se
rect 14292 4641 14343 4642
tri 14343 4641 14344 4642 nw
tri 14389 4641 14390 4642 se
rect 14390 4641 14441 4642
tri 14441 4641 14442 4642 nw
tri 16525 4641 16526 4642 ne
rect 16526 4641 16577 4642
tri 16577 4641 16578 4642 sw
tri 16623 4641 16624 4642 ne
rect 16624 4641 16675 4642
tri 12990 4605 13026 4641 se
rect 13026 4609 14213 4641
tri 14213 4609 14245 4641 nw
tri 14259 4609 14291 4641 se
rect 14291 4611 14313 4641
tri 14313 4611 14343 4641 nw
tri 14359 4611 14389 4641 se
rect 14389 4611 14405 4641
rect 14291 4609 14307 4611
rect 13026 4605 13042 4609
tri 13042 4605 13046 4609 nw
tri 14255 4605 14259 4609 se
rect 14259 4605 14307 4609
tri 14307 4605 14313 4611 nw
tri 14353 4605 14359 4611 se
rect 14359 4605 14405 4611
tri 14405 4605 14441 4641 nw
tri 16526 4605 16562 4641 ne
rect 16562 4635 16578 4641
tri 16578 4635 16584 4641 sw
tri 16624 4635 16630 4641 ne
rect 16630 4635 16675 4641
tri 16675 4635 16682 4642 sw
tri 16721 4635 16728 4642 ne
rect 16728 4635 16773 4642
tri 16773 4635 16780 4642 sw
rect 16562 4620 16584 4635
tri 16584 4620 16599 4635 sw
tri 16630 4620 16645 4635 ne
rect 16645 4620 16682 4635
tri 16682 4620 16697 4635 sw
tri 16728 4620 16743 4635 ne
rect 16743 4620 16780 4635
tri 16780 4620 16795 4635 sw
rect 16562 4605 16599 4620
tri 16599 4605 16614 4620 sw
tri 16645 4605 16660 4620 ne
rect 16660 4619 16697 4620
tri 16697 4619 16698 4620 sw
tri 16743 4619 16744 4620 ne
rect 16744 4619 16795 4620
rect 16660 4613 16698 4619
tri 16698 4613 16704 4619 sw
tri 16744 4613 16750 4619 ne
rect 16750 4613 16795 4619
tri 16795 4613 16802 4620 sw
rect 16660 4605 16704 4613
tri 16704 4605 16712 4613 sw
tri 16750 4605 16758 4613 ne
rect 16758 4605 16802 4613
tri 12978 4593 12990 4605 se
rect 12990 4593 13030 4605
tri 13030 4593 13042 4605 nw
tri 14243 4593 14255 4605 se
rect 14255 4593 14295 4605
tri 14295 4593 14307 4605 nw
tri 14341 4593 14353 4605 se
rect 14353 4593 14390 4605
rect 8331 4590 11636 4593
tri 11636 4590 11639 4593 nw
tri 12975 4590 12978 4593 se
rect 12978 4590 13027 4593
tri 13027 4590 13030 4593 nw
tri 14240 4590 14243 4593 se
rect 14243 4590 14292 4593
tri 14292 4590 14295 4593 nw
tri 14338 4590 14341 4593 se
rect 14341 4590 14390 4593
tri 14390 4590 14405 4605 nw
tri 16562 4590 16577 4605 ne
rect 16577 4593 16614 4605
tri 16614 4593 16626 4605 sw
tri 16660 4593 16672 4605 ne
rect 16672 4593 16712 4605
tri 16712 4593 16724 4605 sw
tri 16758 4597 16766 4605 ne
rect 16577 4590 16626 4593
tri 16626 4590 16629 4593 sw
tri 16672 4590 16675 4593 ne
rect 16675 4590 16724 4593
tri 16724 4590 16727 4593 sw
rect 8331 4573 11619 4590
tri 11619 4573 11636 4590 nw
tri 12974 4589 12975 4590 se
rect 12975 4589 13026 4590
tri 13026 4589 13027 4590 nw
tri 14239 4589 14240 4590 se
rect 14240 4589 14291 4590
tri 14291 4589 14292 4590 nw
tri 14337 4589 14338 4590 se
rect 14338 4589 14389 4590
tri 14389 4589 14390 4590 nw
tri 16577 4589 16578 4590 ne
rect 16578 4589 16629 4590
tri 16629 4589 16630 4590 sw
tri 16675 4589 16676 4590 ne
rect 16676 4589 16727 4590
tri 12962 4577 12974 4589 se
rect 12974 4577 13014 4589
tri 13014 4577 13026 4589 nw
tri 14227 4577 14239 4589 se
rect 14239 4577 14279 4589
tri 14279 4577 14291 4589 nw
tri 14325 4577 14337 4589 se
rect 14337 4577 14369 4589
tri 12958 4573 12962 4577 se
rect 12962 4573 13010 4577
tri 13010 4573 13014 4577 nw
tri 13056 4573 13060 4577 se
rect 13060 4573 14275 4577
tri 14275 4573 14279 4577 nw
tri 14321 4573 14325 4577 se
rect 14325 4573 14369 4577
tri 12954 4569 12958 4573 se
rect 12958 4569 13006 4573
tri 13006 4569 13010 4573 nw
tri 13052 4569 13056 4573 se
rect 13056 4569 14271 4573
tri 14271 4569 14275 4573 nw
tri 14317 4569 14321 4573 se
rect 14321 4569 14369 4573
tri 14369 4569 14389 4589 nw
tri 16578 4569 16598 4589 ne
rect 16598 4583 16630 4589
tri 16630 4583 16636 4589 sw
tri 16676 4583 16682 4589 ne
rect 16682 4583 16727 4589
tri 16727 4583 16734 4590 sw
rect 16598 4573 16636 4583
tri 16636 4573 16646 4583 sw
tri 16682 4573 16692 4583 ne
rect 16692 4573 16734 4583
rect 16598 4569 16646 4573
tri 16646 4569 16650 4573 sw
tri 16692 4569 16696 4573 ne
rect 16696 4569 16734 4573
tri 8155 4568 8156 4569 sw
tri 12953 4568 12954 4569 se
rect 12954 4568 13005 4569
tri 13005 4568 13006 4569 nw
tri 13051 4568 13052 4569 se
rect 13052 4568 14270 4569
tri 14270 4568 14271 4569 nw
tri 14316 4568 14317 4569 se
rect 14317 4568 14368 4569
tri 14368 4568 14369 4569 nw
tri 16598 4568 16599 4569 ne
rect 16599 4568 16650 4569
tri 16650 4568 16651 4569 sw
tri 16696 4568 16697 4569 ne
rect 16697 4568 16734 4569
rect 8155 4562 8156 4568
rect 8103 4550 8156 4562
tri 1527 4498 1552 4523 sw
rect 8155 4544 8156 4550
tri 8156 4544 8180 4568 sw
tri 12929 4544 12953 4568 se
rect 12953 4547 12984 4568
tri 12984 4547 13005 4568 nw
tri 13030 4547 13051 4568 se
rect 13051 4547 14243 4568
rect 12953 4544 12978 4547
rect 8155 4541 11407 4544
tri 11407 4541 11410 4544 sw
tri 12926 4541 12929 4544 se
rect 12929 4541 12978 4544
tri 12978 4541 12984 4547 nw
tri 13024 4541 13030 4547 se
rect 13030 4541 14243 4547
tri 14243 4541 14270 4568 nw
tri 14289 4541 14316 4568 se
rect 14316 4541 14337 4568
rect 8155 4537 11410 4541
tri 11410 4537 11414 4541 sw
tri 12922 4537 12926 4541 se
rect 12926 4537 12974 4541
tri 12974 4537 12978 4541 nw
tri 13020 4537 13024 4541 se
rect 13024 4537 13072 4541
tri 13072 4537 13076 4541 nw
tri 14285 4537 14289 4541 se
rect 14289 4537 14337 4541
tri 14337 4537 14368 4568 nw
rect 8155 4525 11414 4537
tri 11414 4525 11426 4537 sw
tri 12910 4525 12922 4537 se
rect 12922 4525 12962 4537
tri 12962 4525 12974 4537 nw
tri 13008 4525 13020 4537 se
rect 13020 4525 13060 4537
tri 13060 4525 13072 4537 nw
tri 14273 4525 14285 4537 se
rect 14285 4525 14316 4537
rect 8155 4516 11426 4525
tri 11426 4516 11435 4525 sw
tri 12901 4516 12910 4525 se
rect 12910 4516 12953 4525
tri 12953 4516 12962 4525 nw
tri 12999 4516 13008 4525 se
rect 13008 4516 13051 4525
tri 13051 4516 13060 4525 nw
tri 14264 4516 14273 4525 se
rect 14273 4516 14316 4525
tri 14316 4516 14337 4537 nw
rect 14437 4516 14443 4568
rect 14495 4516 14507 4568
rect 14559 4516 14565 4568
tri 16599 4556 16611 4568 ne
rect 16611 4556 16651 4568
tri 16651 4556 16663 4568 sw
tri 16697 4567 16698 4568 ne
tri 16611 4553 16614 4556 ne
rect 16614 4553 16663 4556
tri 16663 4553 16666 4556 sw
tri 16614 4537 16630 4553 ne
rect 8155 4509 11435 4516
tri 11435 4509 11442 4516 sw
tri 12894 4509 12901 4516 se
rect 12901 4509 12946 4516
tri 12946 4509 12953 4516 nw
tri 12992 4509 12999 4516 se
rect 12999 4509 13044 4516
tri 13044 4509 13051 4516 nw
tri 14257 4509 14264 4516 se
rect 14264 4509 14309 4516
tri 14309 4509 14316 4516 nw
rect 8155 4504 11442 4509
tri 11442 4504 11447 4509 sw
tri 12889 4504 12894 4509 se
rect 12894 4504 12941 4509
tri 12941 4504 12946 4509 nw
tri 12987 4504 12992 4509 se
rect 12992 4504 13039 4509
tri 13039 4504 13044 4509 nw
tri 13085 4504 13090 4509 se
rect 13090 4504 14304 4509
tri 14304 4504 14309 4509 nw
rect 8155 4498 11447 4504
rect 1475 4446 1783 4498
rect 1835 4446 1850 4498
rect 1902 4446 1917 4498
rect 1969 4446 1983 4498
rect 2035 4446 2049 4498
rect 2101 4446 2115 4498
rect 2167 4446 2181 4498
rect 2233 4446 2247 4498
rect 2299 4446 2313 4498
rect 2365 4446 2379 4498
rect 2431 4446 2445 4498
rect 2497 4446 2511 4498
rect 2563 4446 2577 4498
rect 2629 4446 2643 4498
rect 2695 4446 2709 4498
rect 2761 4446 2775 4498
rect 2827 4446 2841 4498
rect 2893 4446 2907 4498
rect 2959 4446 3089 4498
rect 3141 4446 3158 4498
rect 3210 4446 3227 4498
rect 3279 4446 3296 4498
rect 3348 4446 3365 4498
rect 3417 4446 3434 4498
rect 3486 4446 3502 4498
rect 3554 4446 3570 4498
rect 3622 4446 3638 4498
rect 3690 4446 3706 4498
rect 3758 4446 4127 4498
rect 4179 4446 4218 4498
rect 4270 4446 4594 4498
rect 4646 4446 4659 4498
rect 4711 4446 4724 4498
rect 4776 4446 4789 4498
rect 4841 4446 4853 4498
rect 4905 4446 4917 4498
rect 4969 4446 4981 4498
rect 5033 4446 5045 4498
rect 5097 4446 5109 4498
rect 5161 4446 5173 4498
rect 5225 4446 5237 4498
rect 5289 4446 5301 4498
rect 5353 4446 5365 4498
rect 5417 4446 5429 4498
rect 5481 4446 5493 4498
rect 5545 4446 5557 4498
rect 5609 4446 5621 4498
rect 5673 4446 5685 4498
rect 5737 4446 5749 4498
rect 5801 4446 5813 4498
rect 5865 4446 5877 4498
rect 5929 4446 5941 4498
rect 5993 4446 6005 4498
rect 6057 4446 6069 4498
rect 6121 4446 6133 4498
rect 6185 4446 6197 4498
rect 6249 4446 6261 4498
rect 6313 4446 6325 4498
rect 6377 4446 6389 4498
rect 6441 4446 6453 4498
rect 6505 4446 6517 4498
rect 6569 4446 6674 4498
rect 6726 4446 6743 4498
rect 6795 4446 6801 4498
rect 8103 4492 11447 4498
tri 11447 4492 11459 4504 sw
tri 12877 4492 12889 4504 se
rect 12889 4495 12932 4504
tri 12932 4495 12941 4504 nw
tri 12978 4495 12987 4504 se
rect 12987 4495 13027 4504
rect 12889 4492 12929 4495
tri 12929 4492 12932 4495 nw
tri 12975 4492 12978 4495 se
rect 12978 4492 13027 4495
tri 13027 4492 13039 4504 nw
tri 13073 4492 13085 4504 se
rect 13085 4492 14291 4504
tri 11393 4491 11394 4492 ne
rect 11394 4491 11459 4492
tri 11459 4491 11460 4492 sw
tri 12876 4491 12877 4492 se
rect 12877 4491 12928 4492
tri 12928 4491 12929 4492 nw
tri 12974 4491 12975 4492 se
rect 12975 4491 13026 4492
tri 13026 4491 13027 4492 nw
tri 13072 4491 13073 4492 se
rect 13073 4491 14291 4492
tri 14291 4491 14304 4504 nw
tri 11394 4478 11407 4491 ne
rect 11407 4478 11591 4491
tri 11407 4464 11421 4478 ne
rect 11421 4464 11591 4478
rect 1475 3676 1527 4446
tri 1527 4421 1552 4446 nw
rect 1618 4361 1665 4413
rect 1717 4361 1746 4413
rect 1798 4407 6847 4413
rect 1798 4361 2230 4407
rect 1618 4355 2230 4361
rect 2282 4379 2742 4407
rect 2794 4379 3254 4407
rect 3306 4379 3766 4407
rect 2282 4355 2689 4379
rect 1618 4343 2689 4355
rect 2745 4343 2771 4355
rect 1618 4337 2230 4343
rect 1618 4285 1665 4337
rect 1717 4285 1746 4337
rect 1798 4291 2230 4337
rect 2282 4323 2689 4343
rect 2827 4323 2853 4379
rect 2909 4323 2935 4379
rect 2991 4323 3017 4379
rect 3073 4323 3099 4379
rect 3155 4323 3180 4379
rect 3236 4355 3254 4379
rect 3236 4343 3261 4355
rect 3236 4323 3254 4343
rect 3317 4323 3342 4379
rect 3398 4323 3423 4379
rect 3479 4323 3504 4379
rect 3560 4355 3766 4379
rect 3818 4355 3889 4407
rect 3941 4355 4278 4407
rect 4330 4355 4401 4407
rect 4453 4355 4790 4407
rect 4842 4355 5302 4407
rect 5354 4355 5814 4407
rect 5866 4355 6326 4407
rect 6378 4361 6847 4407
rect 6899 4361 6953 4413
rect 7005 4361 7058 4413
rect 7110 4361 7163 4413
rect 7215 4361 7268 4413
rect 7320 4361 7373 4413
rect 7425 4361 7478 4413
rect 7530 4361 7597 4413
rect 7649 4361 7705 4413
rect 7757 4393 7763 4413
rect 8263 4412 8269 4464
rect 8321 4412 8333 4464
rect 8385 4446 11365 4464
tri 11365 4446 11383 4464 sw
tri 11421 4446 11439 4464 ne
rect 11439 4446 11591 4464
rect 8385 4439 11383 4446
tri 11383 4439 11390 4446 sw
tri 11439 4439 11446 4446 ne
rect 11446 4439 11591 4446
rect 11643 4439 11656 4491
rect 11708 4439 11714 4491
tri 12874 4489 12876 4491 se
rect 12876 4489 12926 4491
tri 12926 4489 12928 4491 nw
tri 12972 4489 12974 4491 se
rect 12974 4489 13014 4491
tri 12858 4473 12874 4489 se
rect 12874 4473 12910 4489
tri 12910 4473 12926 4489 nw
tri 12956 4473 12972 4489 se
rect 12972 4479 13014 4489
tri 13014 4479 13026 4491 nw
tri 13060 4479 13072 4491 se
rect 13072 4479 14273 4491
rect 12972 4473 13008 4479
tri 13008 4473 13014 4479 nw
tri 13054 4473 13060 4479 se
rect 13060 4473 14273 4479
tri 14273 4473 14291 4491 nw
tri 12842 4457 12858 4473 se
rect 12858 4457 12894 4473
tri 12894 4457 12910 4473 nw
tri 12940 4457 12956 4473 se
rect 12956 4457 12992 4473
tri 12992 4457 13008 4473 nw
tri 13038 4457 13054 4473 se
rect 13054 4457 13090 4473
tri 13090 4457 13106 4473 nw
tri 12824 4439 12842 4457 se
rect 12842 4443 12880 4457
tri 12880 4443 12894 4457 nw
tri 12926 4443 12940 4457 se
rect 12940 4443 12974 4457
rect 12842 4439 12876 4443
tri 12876 4439 12880 4443 nw
tri 12922 4439 12926 4443 se
rect 12926 4439 12974 4443
tri 12974 4439 12992 4457 nw
tri 13020 4439 13038 4457 se
rect 13038 4439 13072 4457
tri 13072 4439 13090 4457 nw
rect 8385 4426 11390 4439
tri 11390 4426 11403 4439 sw
tri 12822 4437 12824 4439 se
rect 12824 4437 12874 4439
tri 12874 4437 12876 4439 nw
tri 12920 4437 12922 4439 se
rect 12922 4437 12962 4439
tri 12811 4426 12822 4437 se
rect 12822 4426 12863 4437
tri 12863 4426 12874 4437 nw
tri 12909 4426 12920 4437 se
rect 12920 4427 12962 4437
tri 12962 4427 12974 4439 nw
tri 13008 4427 13020 4439 se
rect 13020 4427 13059 4439
rect 12920 4426 12961 4427
tri 12961 4426 12962 4427 nw
tri 13007 4426 13008 4427 se
rect 13008 4426 13059 4427
tri 13059 4426 13072 4439 nw
rect 8385 4419 11403 4426
rect 8385 4413 10261 4419
tri 10261 4413 10267 4419 nw
tri 11339 4413 11345 4419 ne
rect 11345 4413 11403 4419
tri 11403 4413 11416 4426 sw
tri 12806 4421 12811 4426 se
rect 12811 4421 12858 4426
tri 12858 4421 12863 4426 nw
tri 12904 4421 12909 4426 se
rect 12909 4421 12956 4426
tri 12956 4421 12961 4426 nw
tri 13002 4421 13007 4426 se
rect 13007 4421 13038 4426
tri 12798 4413 12806 4421 se
rect 12806 4413 12850 4421
tri 12850 4413 12858 4421 nw
tri 12896 4413 12904 4421 se
rect 12904 4413 12948 4421
tri 12948 4413 12956 4421 nw
tri 12994 4413 13002 4421 se
rect 13002 4413 13038 4421
rect 8385 4412 10260 4413
tri 10260 4412 10261 4413 nw
tri 11345 4412 11346 4413 ne
rect 11346 4412 11416 4413
tri 11346 4411 11347 4412 ne
rect 11347 4411 11416 4412
tri 11416 4411 11418 4413 sw
tri 12796 4411 12798 4413 se
rect 12798 4411 12848 4413
tri 12848 4411 12850 4413 nw
tri 12894 4411 12896 4413 se
rect 12896 4411 12946 4413
tri 12946 4411 12948 4413 nw
tri 12992 4411 12994 4413 se
rect 12994 4411 13038 4413
tri 11347 4407 11351 4411 ne
rect 11351 4407 11636 4411
tri 7763 4393 7777 4407 sw
tri 11351 4393 11365 4407 ne
rect 11365 4393 11636 4407
rect 7757 4380 7777 4393
tri 7777 4380 7790 4393 sw
tri 11365 4390 11368 4393 ne
rect 11368 4390 11636 4393
tri 10296 4387 10299 4390 se
rect 10299 4387 11319 4390
tri 11319 4387 11322 4390 sw
tri 11368 4387 11371 4390 ne
rect 11371 4387 11636 4390
tri 10289 4380 10296 4387 se
rect 10296 4380 11322 4387
tri 11322 4380 11329 4387 sw
tri 11371 4380 11378 4387 ne
rect 11378 4380 11636 4387
rect 7757 4379 7790 4380
tri 7790 4379 7791 4380 sw
rect 7757 4361 9908 4379
rect 6378 4355 9908 4361
rect 3560 4351 9908 4355
rect 3560 4343 7763 4351
rect 3560 4323 3766 4343
rect 2282 4291 2742 4323
rect 2794 4291 3254 4323
rect 3306 4291 3766 4323
rect 3818 4291 3889 4343
rect 3941 4291 4278 4343
rect 4330 4291 4401 4343
rect 4453 4291 4790 4343
rect 4842 4291 5302 4343
rect 5354 4291 5814 4343
rect 5866 4291 6326 4343
rect 6378 4337 7763 4343
rect 6378 4291 6847 4337
rect 1798 4285 6847 4291
rect 6899 4285 6953 4337
rect 7005 4285 7058 4337
rect 7110 4285 7163 4337
rect 7215 4285 7268 4337
rect 7320 4285 7373 4337
rect 7425 4285 7478 4337
rect 7530 4285 7597 4337
rect 7649 4285 7705 4337
rect 7757 4285 7763 4337
tri 7763 4323 7791 4351 nw
tri 9852 4323 9880 4351 ne
tri 9701 4320 9703 4322 se
rect 9703 4320 9712 4322
tri 7810 4285 7845 4320 se
rect 7845 4285 9712 4320
rect 1618 4270 1764 4285
tri 1764 4270 1779 4285 nw
tri 7795 4270 7810 4285 se
rect 7810 4275 9712 4285
rect 7810 4270 7870 4275
tri 7870 4270 7875 4275 nw
tri 9701 4270 9706 4275 ne
rect 9706 4270 9712 4275
rect 9764 4270 9776 4322
rect 9828 4270 9834 4322
rect 1618 4258 1752 4270
tri 1752 4258 1764 4270 nw
tri 7783 4258 7795 4270 se
rect 7795 4258 7858 4270
tri 7858 4258 7870 4270 nw
tri 9868 4258 9880 4270 se
rect 9880 4258 9908 4351
rect 10045 4374 10097 4380
tri 10268 4359 10289 4380 se
rect 10289 4359 11329 4380
tri 11329 4359 11350 4380 sw
tri 11378 4359 11399 4380 ne
rect 11399 4359 11636 4380
rect 11688 4359 11700 4411
rect 11752 4359 11758 4411
tri 12790 4405 12796 4411 se
rect 12796 4405 12842 4411
tri 12842 4405 12848 4411 nw
tri 12888 4405 12894 4411 se
rect 12894 4405 12940 4411
tri 12940 4405 12946 4411 nw
tri 12986 4405 12992 4411 se
rect 12992 4405 13038 4411
tri 13038 4405 13059 4426 nw
tri 12770 4385 12790 4405 se
rect 12790 4391 12828 4405
tri 12828 4391 12842 4405 nw
tri 12874 4391 12888 4405 se
rect 12888 4391 12910 4405
rect 12790 4385 12822 4391
tri 12822 4385 12828 4391 nw
tri 12868 4385 12874 4391 se
rect 12874 4385 12910 4391
tri 12759 4374 12770 4385 se
rect 12770 4374 12811 4385
tri 12811 4374 12822 4385 nw
tri 12857 4374 12868 4385 se
rect 12868 4375 12910 4385
tri 12910 4375 12940 4405 nw
tri 12956 4375 12986 4405 se
rect 12986 4375 13007 4405
rect 12868 4374 12909 4375
tri 12909 4374 12910 4375 nw
tri 12955 4374 12956 4375 se
rect 12956 4374 13007 4375
tri 13007 4374 13038 4405 nw
tri 12754 4369 12759 4374 se
rect 12759 4369 12806 4374
tri 12806 4369 12811 4374 nw
tri 12852 4369 12857 4374 se
rect 12857 4369 12904 4374
tri 12904 4369 12909 4374 nw
tri 12950 4369 12955 4374 se
rect 12955 4369 12994 4374
tri 12746 4361 12754 4369 se
rect 12754 4361 12798 4369
tri 12798 4361 12806 4369 nw
tri 12844 4361 12852 4369 se
rect 12852 4361 12896 4369
tri 12896 4361 12904 4369 nw
tri 12942 4361 12950 4369 se
rect 12950 4361 12994 4369
tri 12994 4361 13007 4374 nw
tri 12744 4359 12746 4361 se
rect 12746 4359 12796 4361
tri 12796 4359 12798 4361 nw
tri 12842 4359 12844 4361 se
rect 12844 4359 12894 4361
tri 12894 4359 12896 4361 nw
tri 12940 4359 12942 4361 se
rect 12942 4359 12986 4361
tri 10253 4344 10268 4359 se
rect 10268 4358 11350 4359
rect 10268 4344 10299 4358
tri 10299 4344 10313 4358 nw
tri 11295 4344 11309 4358 ne
rect 11309 4353 11350 4358
tri 11350 4353 11356 4359 sw
tri 12738 4353 12744 4359 se
rect 12744 4353 12790 4359
tri 12790 4353 12796 4359 nw
tri 12836 4353 12842 4359 se
rect 12842 4353 12888 4359
tri 12888 4353 12894 4359 nw
tri 12934 4353 12940 4359 se
rect 12940 4353 12986 4359
tri 12986 4353 12994 4361 nw
rect 11309 4344 11356 4353
tri 10240 4331 10253 4344 se
rect 10253 4331 10286 4344
tri 10286 4331 10299 4344 nw
tri 11309 4331 11322 4344 ne
rect 11322 4333 11356 4344
tri 11356 4333 11376 4353 sw
tri 12718 4333 12738 4353 se
rect 12738 4339 12776 4353
tri 12776 4339 12790 4353 nw
tri 12822 4339 12836 4353 se
rect 12836 4339 12858 4353
rect 12738 4333 12770 4339
tri 12770 4333 12776 4339 nw
tri 12816 4333 12822 4339 se
rect 12822 4333 12858 4339
rect 11322 4331 11376 4333
tri 11376 4331 11378 4333 sw
tri 12716 4331 12718 4333 se
rect 12718 4331 12768 4333
tri 12768 4331 12770 4333 nw
tri 12814 4331 12816 4333 se
rect 12816 4331 12858 4333
tri 10238 4329 10240 4331 se
rect 10240 4329 10284 4331
tri 10284 4329 10286 4331 nw
tri 11322 4329 11324 4331 ne
rect 11324 4329 12754 4331
tri 10236 4327 10238 4329 se
rect 10238 4327 10282 4329
tri 10282 4327 10284 4329 nw
tri 10322 4327 10324 4329 se
rect 10324 4327 11271 4329
tri 11271 4327 11273 4329 sw
tri 11324 4327 11326 4329 ne
rect 11326 4327 12754 4329
rect 10045 4310 10097 4322
tri 10019 4270 10045 4296 se
tri 10007 4258 10019 4270 se
rect 10019 4258 10045 4270
tri 10218 4309 10236 4327 se
rect 10236 4309 10264 4327
tri 10264 4309 10282 4327 nw
tri 10304 4309 10322 4327 se
rect 10322 4317 11273 4327
tri 11273 4317 11283 4327 sw
tri 11326 4317 11336 4327 ne
rect 11336 4317 12754 4327
tri 12754 4317 12768 4331 nw
tri 12800 4317 12814 4331 se
rect 12814 4323 12858 4331
tri 12858 4323 12888 4353 nw
tri 12904 4323 12934 4353 se
rect 12934 4323 12942 4353
rect 12814 4317 12852 4323
tri 12852 4317 12858 4323 nw
tri 12898 4317 12904 4323 se
rect 12904 4317 12942 4323
rect 10322 4309 11283 4317
tri 11283 4309 11291 4317 sw
tri 11336 4309 11344 4317 ne
rect 11344 4309 12746 4317
tri 12746 4309 12754 4317 nw
tri 12792 4309 12800 4317 se
rect 12800 4309 12844 4317
tri 12844 4309 12852 4317 nw
tri 12890 4309 12898 4317 se
rect 12898 4309 12942 4317
tri 12942 4309 12986 4353 nw
tri 10207 4298 10218 4309 se
rect 10218 4304 10259 4309
tri 10259 4304 10264 4309 nw
tri 10299 4304 10304 4309 se
rect 10304 4304 11291 4309
rect 10218 4298 10253 4304
tri 10253 4298 10259 4304 nw
tri 10293 4298 10299 4304 se
rect 10299 4301 11291 4304
tri 11291 4301 11299 4309 sw
tri 11344 4301 11352 4309 ne
rect 11352 4301 12738 4309
tri 12738 4301 12746 4309 nw
tri 12784 4301 12792 4309 se
rect 12792 4301 12836 4309
tri 12836 4301 12844 4309 nw
tri 12882 4301 12890 4309 se
rect 12890 4301 12934 4309
tri 12934 4301 12942 4309 nw
rect 10299 4299 11299 4301
tri 11299 4299 11301 4301 sw
tri 11352 4299 11354 4301 ne
rect 11354 4299 12736 4301
tri 12736 4299 12738 4301 nw
tri 12782 4299 12784 4301 se
rect 12784 4299 12831 4301
rect 10299 4298 11301 4299
tri 10205 4296 10207 4298 se
rect 10207 4296 10251 4298
tri 10251 4296 10253 4298 nw
tri 10291 4296 10293 4298 se
rect 10293 4297 11301 4298
rect 10293 4296 10337 4297
tri 10337 4296 10338 4297 nw
tri 11247 4296 11248 4297 ne
rect 11248 4296 11301 4297
tri 11301 4296 11304 4299 sw
tri 12779 4296 12782 4299 se
rect 12782 4296 12831 4299
tri 12831 4296 12836 4301 nw
tri 12877 4296 12882 4301 se
rect 12882 4296 12929 4301
tri 12929 4296 12934 4301 nw
tri 10192 4283 10205 4296 se
rect 10205 4283 10238 4296
tri 10238 4283 10251 4296 nw
tri 10278 4283 10291 4296 se
rect 10291 4283 10324 4296
tri 10324 4283 10337 4296 nw
tri 11248 4283 11261 4296 ne
rect 11261 4283 11304 4296
tri 10180 4271 10192 4283 se
rect 10192 4271 10226 4283
tri 10226 4271 10238 4283 nw
tri 10266 4271 10278 4283 se
rect 10278 4271 10312 4283
tri 10312 4271 10324 4283 nw
tri 11261 4271 11273 4283 ne
rect 11273 4271 11304 4283
tri 11304 4271 11329 4296 sw
tri 12754 4271 12779 4296 se
rect 12779 4271 12806 4296
tri 12806 4271 12831 4296 nw
tri 12852 4271 12877 4296 se
rect 12877 4271 12896 4296
tri 10177 4268 10180 4271 se
rect 10180 4268 10223 4271
tri 10223 4268 10226 4271 nw
tri 10263 4268 10266 4271 se
rect 10266 4268 10309 4271
tri 10309 4268 10312 4271 nw
tri 11273 4268 11276 4271 ne
rect 11276 4268 12798 4271
tri 10176 4267 10177 4268 se
rect 10177 4267 10222 4268
tri 10222 4267 10223 4268 nw
tri 10262 4267 10263 4268 se
rect 10263 4267 10308 4268
tri 10308 4267 10309 4268 nw
tri 10348 4267 10349 4268 se
rect 10349 4267 11228 4268
tri 11228 4267 11229 4268 sw
tri 11276 4267 11277 4268 ne
rect 11277 4267 12798 4268
tri 10172 4263 10176 4267 se
rect 10176 4263 10218 4267
tri 10218 4263 10222 4267 nw
tri 10258 4263 10262 4267 se
rect 10262 4263 10304 4267
tri 10304 4263 10308 4267 nw
tri 10344 4263 10348 4267 se
rect 10348 4263 11229 4267
tri 11229 4263 11233 4267 sw
tri 11277 4263 11281 4267 ne
rect 11281 4263 12798 4267
tri 12798 4263 12806 4271 nw
tri 12844 4263 12852 4271 se
rect 12852 4263 12896 4271
tri 12896 4263 12929 4296 nw
rect 1618 4250 1744 4258
tri 1744 4250 1752 4258 nw
tri 7778 4253 7783 4258 se
rect 7783 4253 7853 4258
tri 7853 4253 7858 4258 nw
tri 9863 4253 9868 4258 se
rect 9868 4253 9908 4258
tri 10002 4253 10007 4258 se
rect 10007 4253 10097 4258
tri 7777 4252 7778 4253 se
rect 7778 4252 7852 4253
tri 7852 4252 7853 4253 nw
tri 9862 4252 9863 4253 se
rect 9863 4252 9908 4253
tri 10001 4252 10002 4253 se
rect 10002 4252 10097 4253
tri 10161 4252 10172 4263 se
rect 10172 4258 10213 4263
tri 10213 4258 10218 4263 nw
tri 10253 4258 10258 4263 se
rect 10258 4258 10293 4263
rect 10172 4252 10207 4258
tri 10207 4252 10213 4258 nw
tri 10247 4252 10253 4258 se
rect 10253 4252 10293 4258
tri 10293 4252 10304 4263 nw
tri 10333 4252 10344 4263 se
rect 10344 4252 11233 4263
tri 11233 4252 11244 4263 sw
tri 11281 4252 11292 4263 ne
rect 11292 4252 12787 4263
tri 12787 4252 12798 4263 nw
tri 12833 4252 12844 4263 se
rect 12844 4252 12882 4263
tri 7775 4250 7777 4252 se
rect 7777 4250 7850 4252
tri 7850 4250 7852 4252 nw
tri 9860 4250 9862 4252 se
rect 9862 4250 9908 4252
rect 1618 4247 1741 4250
tri 1741 4247 1744 4250 nw
rect 1618 3851 1708 4247
tri 1708 4214 1741 4247 nw
rect 3001 4195 3007 4247
rect 3059 4195 3071 4247
rect 3123 4195 3129 4247
rect 2448 4119 2454 4171
rect 2506 4119 2518 4171
rect 2570 4119 2576 4171
rect 2448 3903 2576 4119
rect 3001 3987 3129 4195
rect 3001 3935 3007 3987
rect 3059 3935 3071 3987
rect 3123 3935 3129 3987
rect 3513 4195 3519 4247
rect 3571 4195 3583 4247
rect 3635 4195 3641 4247
rect 3513 4079 3641 4195
rect 3513 4027 3519 4079
rect 3571 4027 3583 4079
rect 3635 4027 3641 4079
tri 1708 3851 1743 3886 sw
rect 2448 3851 2454 3903
rect 2506 3851 2518 3903
rect 2570 3851 2576 3903
rect 3513 3905 3641 4027
rect 3513 3853 3519 3905
rect 3571 3853 3583 3905
rect 3635 3853 3641 3905
rect 4359 4195 4365 4247
rect 4417 4195 4429 4247
rect 4481 4195 4487 4247
rect 4359 3905 4487 4195
rect 4359 3853 4365 3905
rect 4417 3853 4429 3905
rect 4481 3853 4487 3905
rect 4967 4195 4973 4247
rect 5025 4195 5037 4247
rect 5089 4230 6145 4247
tri 6145 4230 6162 4247 sw
rect 5089 4198 6162 4230
tri 6162 4198 6194 4230 sw
rect 6668 4198 6674 4250
rect 6726 4198 6743 4250
rect 6795 4247 7847 4250
tri 7847 4247 7850 4250 nw
tri 9857 4247 9860 4250 se
rect 9860 4247 9908 4250
tri 9996 4247 10001 4252 se
rect 10001 4247 10019 4252
rect 6795 4242 7842 4247
tri 7842 4242 7847 4247 nw
tri 9852 4242 9857 4247 se
rect 9857 4242 9908 4247
rect 6795 4240 7840 4242
tri 7840 4240 7842 4242 nw
tri 7890 4240 7892 4242 se
rect 7892 4240 9685 4242
tri 9685 4240 9687 4242 sw
tri 9847 4240 9849 4242 se
rect 9849 4240 9908 4242
rect 6795 4211 7811 4240
tri 7811 4211 7840 4240 nw
tri 7861 4211 7890 4240 se
rect 7890 4211 9908 4240
tri 9960 4211 9996 4247 se
rect 9996 4211 10019 4247
tri 10019 4211 10060 4252 nw
tri 10146 4237 10161 4252 se
rect 10161 4237 10192 4252
tri 10192 4237 10207 4252 nw
tri 10232 4237 10247 4252 se
rect 10247 4243 10284 4252
tri 10284 4243 10293 4252 nw
tri 10324 4243 10333 4252 se
rect 10333 4249 11244 4252
tri 11244 4249 11247 4252 sw
tri 11292 4249 11295 4252 ne
rect 11295 4249 12784 4252
tri 12784 4249 12787 4252 nw
tri 12830 4249 12833 4252 se
rect 12833 4249 12882 4252
tri 12882 4249 12896 4263 nw
rect 10333 4243 11247 4249
rect 10247 4237 10278 4243
tri 10278 4237 10284 4243 nw
tri 10318 4237 10324 4243 se
rect 10324 4239 11247 4243
tri 11247 4239 11257 4249 sw
tri 11295 4239 11305 4249 ne
rect 11305 4239 12774 4249
tri 12774 4239 12784 4249 nw
tri 12820 4239 12830 4249 se
rect 12830 4239 12844 4249
rect 10324 4237 11257 4239
tri 10131 4222 10146 4237 se
rect 10146 4222 10177 4237
tri 10177 4222 10192 4237 nw
tri 10217 4222 10232 4237 se
rect 10232 4222 10263 4237
tri 10263 4222 10278 4237 nw
tri 10303 4222 10318 4237 se
rect 10318 4236 11257 4237
rect 10318 4222 10349 4236
tri 10349 4222 10363 4236 nw
tri 11204 4222 11218 4236 ne
rect 11218 4222 11257 4236
tri 10120 4211 10131 4222 se
rect 10131 4212 10167 4222
tri 10167 4212 10177 4222 nw
tri 10207 4212 10217 4222 se
rect 10217 4212 10252 4222
rect 10131 4211 10166 4212
tri 10166 4211 10167 4212 nw
tri 10206 4211 10207 4212 se
rect 10207 4211 10252 4212
tri 10252 4211 10263 4222 nw
tri 10292 4211 10303 4222 se
rect 10303 4211 10338 4222
tri 10338 4211 10349 4222 nw
tri 11218 4211 11229 4222 ne
rect 11229 4211 11257 4222
tri 11257 4211 11285 4239 sw
tri 12792 4211 12820 4239 se
rect 12820 4211 12844 4239
tri 12844 4211 12882 4249 nw
rect 13241 4211 13247 4263
rect 13299 4211 13311 4263
rect 13363 4211 13369 4263
rect 6795 4206 7806 4211
tri 7806 4206 7811 4211 nw
tri 7856 4206 7861 4211 se
rect 7861 4209 9908 4211
tri 9958 4209 9960 4211 se
rect 9960 4209 10002 4211
rect 7861 4206 7892 4209
rect 6795 4198 6801 4206
tri 6801 4198 6809 4206 nw
tri 7848 4198 7856 4206 se
rect 7856 4198 7892 4206
rect 5089 4195 6194 4198
rect 4967 4179 5132 4195
tri 5132 4179 5148 4195 nw
tri 6116 4179 6132 4195 ne
rect 6132 4194 6194 4195
tri 6194 4194 6198 4198 sw
tri 7844 4194 7848 4198 se
rect 7848 4194 7892 4198
tri 7892 4194 7907 4209 nw
tri 9943 4194 9958 4209 se
rect 9958 4194 10002 4209
tri 10002 4194 10019 4211 nw
tri 10115 4206 10120 4211 se
rect 10120 4206 10161 4211
tri 10161 4206 10166 4211 nw
tri 10201 4206 10206 4211 se
rect 10206 4206 10238 4211
tri 10103 4194 10115 4206 se
rect 10115 4194 10149 4206
tri 10149 4194 10161 4206 nw
tri 10189 4194 10201 4206 se
rect 10201 4197 10238 4206
tri 10238 4197 10252 4211 nw
tri 10278 4197 10292 4211 se
rect 10292 4197 10312 4211
rect 10201 4194 10235 4197
tri 10235 4194 10238 4197 nw
tri 10275 4194 10278 4197 se
rect 10278 4194 10312 4197
rect 6132 4179 6198 4194
tri 6198 4179 6213 4194 sw
tri 7829 4179 7844 4194 se
rect 7844 4179 7878 4194
tri 7878 4180 7892 4194 nw
tri 9929 4180 9943 4194 se
rect 9943 4180 9987 4194
tri 9928 4179 9929 4180 se
rect 9929 4179 9987 4180
tri 9987 4179 10002 4194 nw
tri 10100 4191 10103 4194 se
rect 10103 4191 10146 4194
tri 10146 4191 10149 4194 nw
tri 10186 4191 10189 4194 se
rect 10189 4191 10232 4194
tri 10232 4191 10235 4194 nw
tri 10272 4191 10275 4194 se
rect 10275 4191 10312 4194
tri 10094 4185 10100 4191 se
rect 10100 4185 10140 4191
tri 10140 4185 10146 4191 nw
tri 10180 4185 10186 4191 se
rect 10186 4185 10226 4191
tri 10226 4185 10232 4191 nw
tri 10266 4185 10272 4191 se
rect 10272 4185 10312 4191
tri 10312 4185 10338 4211 nw
tri 11229 4185 11255 4211 ne
rect 11255 4185 12812 4211
tri 10088 4179 10094 4185 se
rect 10094 4179 10134 4185
tri 10134 4179 10140 4185 nw
tri 10174 4179 10180 4185 se
rect 10180 4179 10220 4185
tri 10220 4179 10226 4185 nw
tri 10260 4179 10266 4185 se
rect 10266 4179 10306 4185
tri 10306 4179 10312 4185 nw
rect 10867 4179 10919 4185
tri 10919 4179 10925 4185 sw
tri 11255 4179 11261 4185 ne
rect 11261 4179 12812 4185
tri 12812 4179 12844 4211 nw
rect 4967 4170 5123 4179
tri 5123 4170 5132 4179 nw
tri 6132 4170 6141 4179 ne
rect 6141 4170 6213 4179
tri 6213 4170 6222 4179 sw
tri 7826 4176 7829 4179 se
rect 7829 4176 7878 4179
rect 7826 4170 7878 4176
tri 9923 4174 9928 4179 se
rect 9928 4174 9982 4179
tri 9982 4174 9987 4179 nw
tri 10085 4176 10088 4179 se
rect 10088 4176 10131 4179
tri 10131 4176 10134 4179 nw
tri 10171 4176 10174 4179 se
rect 10174 4176 10217 4179
tri 10217 4176 10220 4179 nw
tri 10257 4176 10260 4179 se
rect 10260 4176 10303 4179
tri 10303 4176 10306 4179 nw
tri 10083 4174 10085 4176 se
rect 10085 4174 10129 4176
tri 10129 4174 10131 4176 nw
tri 10169 4174 10171 4176 se
rect 10171 4174 10215 4176
tri 10215 4174 10217 4176 nw
tri 10255 4174 10257 4176 se
rect 10257 4174 10301 4176
tri 10301 4174 10303 4176 nw
tri 10381 4174 10383 4176 se
rect 10383 4174 10839 4176
tri 7956 4170 7960 4174 se
rect 7960 4170 9978 4174
tri 9978 4170 9982 4174 nw
tri 10079 4170 10083 4174 se
rect 10083 4170 10125 4174
tri 10125 4170 10129 4174 nw
tri 10165 4170 10169 4174 se
rect 10169 4170 10211 4174
tri 10211 4170 10215 4174 nw
tri 10251 4170 10255 4174 se
rect 10255 4170 10297 4174
tri 10297 4170 10301 4174 nw
tri 10377 4170 10381 4174 se
rect 10381 4170 10839 4174
rect 4967 4167 5120 4170
tri 5120 4167 5123 4170 nw
tri 6141 4167 6144 4170 ne
rect 6144 4167 6222 4170
tri 6222 4167 6225 4170 sw
rect 4967 4079 5095 4167
tri 5095 4142 5120 4167 nw
rect 4967 4027 4973 4079
rect 5025 4027 5037 4079
rect 5089 4027 5095 4079
rect 4967 3905 5095 4027
rect 4967 3853 4973 3905
rect 5025 3853 5037 3905
rect 5089 3853 5095 3905
rect 5902 4115 5908 4167
rect 5960 4115 5972 4167
rect 6024 4115 6030 4167
tri 6144 4149 6162 4167 ne
rect 6162 4149 6225 4167
tri 6225 4149 6243 4167 sw
tri 6162 4118 6193 4149 ne
rect 6193 4118 7672 4149
rect 5902 4054 6030 4115
tri 6193 4106 6205 4118 ne
rect 6205 4106 7672 4118
tri 6205 4097 6214 4106 ne
rect 6214 4097 7672 4106
tri 7592 4065 7624 4097 ne
tri 6030 4054 6034 4058 sw
rect 5902 4048 6034 4054
tri 6034 4048 6040 4054 sw
rect 5902 4028 6040 4048
tri 6040 4028 6060 4048 sw
rect 5902 3956 7552 4028
rect 5902 3949 6055 3956
tri 6055 3949 6062 3956 nw
tri 7442 3949 7449 3956 ne
rect 7449 3949 7552 3956
rect 5902 3942 6048 3949
tri 6048 3942 6055 3949 nw
tri 7449 3942 7456 3949 ne
rect 7456 3942 7552 3949
rect 5902 3938 6044 3942
tri 6044 3938 6048 3942 nw
tri 7456 3938 7460 3942 ne
rect 7460 3938 7552 3942
rect 5902 3937 6043 3938
tri 6043 3937 6044 3938 nw
tri 7460 3937 7461 3938 ne
rect 7461 3937 7552 3938
rect 5902 3905 6030 3937
tri 6030 3924 6043 3937 nw
tri 7461 3924 7474 3937 ne
rect 7474 3924 7552 3937
tri 7474 3905 7493 3924 ne
rect 7493 3905 7552 3924
rect 5902 3853 5908 3905
rect 5960 3853 5972 3905
rect 6024 3853 6030 3905
tri 7493 3898 7500 3905 ne
rect 1618 3815 1743 3851
tri 1743 3815 1779 3851 sw
rect 1618 3763 1624 3815
rect 1676 3763 1709 3815
rect 1761 3809 6847 3815
rect 1761 3763 2230 3809
rect 1618 3757 2230 3763
rect 2282 3777 2742 3809
rect 2794 3777 3254 3809
rect 3306 3777 3766 3809
rect 2282 3757 2689 3777
rect 1618 3745 2689 3757
rect 2745 3745 2771 3757
rect 1618 3739 2230 3745
rect 1618 3687 1624 3739
rect 1676 3687 1709 3739
rect 1761 3693 2230 3739
rect 2282 3721 2689 3745
rect 2827 3721 2853 3777
rect 2909 3721 2935 3777
rect 2991 3721 3017 3777
rect 3073 3721 3099 3777
rect 3155 3721 3180 3777
rect 3236 3757 3254 3777
rect 3236 3745 3261 3757
rect 3236 3721 3254 3745
rect 3317 3721 3342 3777
rect 3398 3721 3423 3777
rect 3479 3721 3504 3777
rect 3560 3757 3766 3777
rect 3818 3757 4145 3809
rect 4197 3757 4278 3809
rect 4330 3757 4657 3809
rect 4709 3757 4790 3809
rect 4842 3757 5302 3809
rect 5354 3757 5814 3809
rect 5866 3757 6326 3809
rect 6378 3763 6847 3809
rect 6899 3763 6954 3815
rect 7006 3763 7061 3815
rect 7113 3763 7168 3815
rect 7220 3763 7275 3815
rect 7327 3763 7382 3815
rect 7434 3763 7462 3815
rect 6378 3757 7462 3763
rect 3560 3745 7462 3757
rect 3560 3721 3766 3745
rect 2282 3693 2742 3721
rect 2794 3693 3254 3721
rect 3306 3693 3766 3721
rect 3818 3693 4145 3745
rect 4197 3693 4278 3745
rect 4330 3693 4657 3745
rect 4709 3693 4790 3745
rect 4842 3693 5302 3745
rect 5354 3693 5814 3745
rect 5866 3693 6326 3745
rect 6378 3739 7462 3745
rect 6378 3693 6847 3739
rect 1761 3687 6847 3693
rect 6899 3687 6954 3739
rect 7006 3687 7061 3739
rect 7113 3687 7168 3739
rect 7220 3687 7275 3739
rect 7327 3687 7382 3739
rect 7434 3687 7462 3739
rect 7500 3784 7552 3905
rect 7624 3856 7672 4097
tri 7953 4167 7956 4170 se
rect 7956 4167 9958 4170
rect 7826 4106 7878 4118
rect 7826 4048 7878 4054
tri 7936 4150 7953 4167 se
rect 7953 4150 9958 4167
tri 9958 4150 9978 4170 nw
tri 10069 4160 10079 4170 se
rect 10079 4166 10121 4170
tri 10121 4166 10125 4170 nw
tri 10161 4166 10165 4170 se
rect 10165 4166 10192 4170
rect 10079 4160 10115 4166
tri 10115 4160 10121 4166 nw
tri 10155 4160 10161 4166 se
rect 10161 4160 10192 4166
tri 10059 4150 10069 4160 se
rect 10069 4150 10105 4160
tri 10105 4150 10115 4160 nw
tri 10145 4150 10155 4160 se
rect 10155 4151 10192 4160
tri 10192 4151 10211 4170 nw
tri 10232 4151 10251 4170 se
rect 10251 4151 10277 4170
rect 10155 4150 10191 4151
tri 10191 4150 10192 4151 nw
tri 10231 4150 10232 4151 se
rect 10232 4150 10277 4151
tri 10277 4150 10297 4170 nw
tri 10357 4150 10377 4170 se
rect 10377 4150 10478 4170
rect 7936 4144 9937 4150
rect 7988 4129 9937 4144
tri 9937 4129 9958 4150 nw
tri 10054 4145 10059 4150 se
rect 10059 4145 10100 4150
tri 10100 4145 10105 4150 nw
tri 10140 4145 10145 4150 se
rect 10145 4145 10186 4150
tri 10186 4145 10191 4150 nw
tri 10226 4145 10231 4150 se
rect 10231 4145 10257 4150
tri 10039 4130 10054 4145 se
rect 10054 4130 10085 4145
tri 10085 4130 10100 4145 nw
tri 10125 4130 10140 4145 se
rect 10140 4130 10171 4145
tri 10171 4130 10186 4145 nw
tri 10211 4130 10226 4145 se
rect 10226 4130 10257 4145
tri 10257 4130 10277 4150 nw
tri 10337 4130 10357 4150 se
rect 10357 4130 10478 4150
tri 10038 4129 10039 4130 se
rect 10039 4129 10084 4130
tri 10084 4129 10085 4130 nw
tri 10124 4129 10125 4130 se
rect 10125 4129 10170 4130
tri 10170 4129 10171 4130 nw
tri 10210 4129 10211 4130 se
rect 10211 4129 10256 4130
tri 10256 4129 10257 4130 nw
tri 10336 4129 10337 4130 se
rect 10337 4129 10478 4130
rect 7988 4127 9935 4129
tri 9935 4127 9937 4129 nw
tri 10036 4127 10038 4129 se
rect 10038 4127 10082 4129
tri 10082 4127 10084 4129 nw
tri 10122 4127 10124 4129 se
rect 10124 4127 10168 4129
tri 10168 4127 10170 4129 nw
tri 10208 4127 10210 4129 se
rect 10210 4127 10254 4129
tri 10254 4127 10256 4129 nw
tri 10334 4127 10336 4129 se
rect 10336 4127 10478 4129
rect 7988 4122 9930 4127
tri 9930 4122 9935 4127 nw
tri 10031 4122 10036 4127 se
rect 10036 4122 10077 4127
tri 10077 4122 10082 4127 nw
tri 10117 4122 10122 4127 se
rect 10122 4122 10163 4127
tri 10163 4122 10168 4127 nw
tri 10203 4122 10208 4127 se
rect 10208 4122 10249 4127
tri 10249 4122 10254 4127 nw
tri 10329 4122 10334 4127 se
rect 10334 4122 10478 4127
rect 7988 4118 8009 4122
tri 8009 4118 8013 4122 nw
tri 10027 4118 10031 4122 se
rect 10031 4120 10075 4122
tri 10075 4120 10077 4122 nw
tri 10115 4120 10117 4122 se
rect 10117 4120 10159 4122
rect 10031 4118 10073 4120
tri 10073 4118 10075 4120 nw
tri 10113 4118 10115 4120 se
rect 10115 4118 10159 4120
tri 10159 4118 10163 4122 nw
tri 10199 4118 10203 4122 se
rect 10203 4118 10245 4122
tri 10245 4118 10249 4122 nw
tri 10325 4118 10329 4122 se
rect 10329 4118 10478 4122
rect 10530 4118 10787 4170
rect 7988 4113 8004 4118
tri 8004 4113 8009 4118 nw
tri 10023 4114 10027 4118 se
rect 10027 4114 10069 4118
tri 10069 4114 10073 4118 nw
tri 10109 4114 10113 4118 se
rect 10113 4114 10154 4118
tri 10022 4113 10023 4114 se
rect 10023 4113 10068 4114
tri 10068 4113 10069 4114 nw
tri 10108 4113 10109 4114 se
rect 10109 4113 10154 4114
tri 10154 4113 10159 4118 nw
tri 10194 4113 10199 4118 se
rect 10199 4113 10240 4118
tri 10240 4113 10245 4118 nw
tri 10320 4113 10325 4118 se
rect 10325 4113 10839 4118
rect 7988 4104 7995 4113
tri 7995 4104 8004 4113 nw
tri 10013 4104 10022 4113 se
rect 10022 4104 10059 4113
tri 10059 4104 10068 4113 nw
tri 10099 4104 10108 4113 se
rect 10108 4105 10146 4113
tri 10146 4105 10154 4113 nw
tri 10186 4105 10194 4113 se
rect 10194 4105 10231 4113
rect 10108 4104 10145 4105
tri 10145 4104 10146 4105 nw
tri 10185 4104 10186 4105 se
rect 10186 4104 10231 4105
tri 10231 4104 10240 4113 nw
tri 10311 4104 10320 4113 se
rect 10320 4104 10839 4113
tri 7988 4097 7995 4104 nw
tri 10008 4099 10013 4104 se
rect 10013 4099 10054 4104
tri 10054 4099 10059 4104 nw
tri 10094 4099 10099 4104 se
rect 10099 4099 10140 4104
tri 10140 4099 10145 4104 nw
tri 10180 4099 10185 4104 se
rect 10185 4099 10224 4104
tri 10006 4097 10008 4099 se
rect 10008 4097 10052 4099
tri 10052 4097 10054 4099 nw
tri 10092 4097 10094 4099 se
rect 10094 4097 10138 4099
tri 10138 4097 10140 4099 nw
tri 10178 4097 10180 4099 se
rect 10180 4097 10224 4099
tri 10224 4097 10231 4104 nw
tri 10304 4097 10311 4104 se
rect 10311 4097 10478 4104
rect 7936 4080 7988 4092
tri 9999 4090 10006 4097 se
rect 10006 4090 10039 4097
tri 8026 4084 8032 4090 se
rect 8032 4084 9847 4090
tri 9993 4084 9999 4090 se
rect 9999 4084 10039 4090
tri 10039 4084 10052 4097 nw
tri 10079 4084 10092 4097 se
rect 10092 4084 10125 4097
tri 10125 4084 10138 4097 nw
tri 10165 4084 10178 4097 se
rect 10178 4084 10211 4097
tri 10211 4084 10224 4097 nw
tri 10291 4084 10304 4097 se
rect 10304 4084 10478 4097
rect 7936 4022 7988 4028
tri 8020 4078 8026 4084 se
rect 8026 4078 9847 4084
rect 8020 4072 9847 4078
rect 8072 4038 9847 4072
tri 9977 4068 9993 4084 se
rect 9993 4074 10029 4084
tri 10029 4074 10039 4084 nw
tri 10069 4074 10079 4084 se
rect 10079 4074 10100 4084
rect 9993 4068 10023 4074
tri 10023 4068 10029 4074 nw
tri 10063 4068 10069 4074 se
rect 10069 4068 10100 4074
tri 9962 4053 9977 4068 se
rect 9977 4053 10008 4068
tri 10008 4053 10023 4068 nw
tri 10048 4053 10063 4068 se
rect 10063 4059 10100 4068
tri 10100 4059 10125 4084 nw
tri 10140 4059 10165 4084 se
rect 10165 4059 10179 4084
rect 10063 4053 10094 4059
tri 10094 4053 10100 4059 nw
tri 10134 4053 10140 4059 se
rect 10140 4053 10179 4059
tri 9961 4052 9962 4053 se
rect 9962 4052 10007 4053
tri 10007 4052 10008 4053 nw
tri 10047 4052 10048 4053 se
rect 10048 4052 10093 4053
tri 10093 4052 10094 4053 nw
tri 10133 4052 10134 4053 se
rect 10134 4052 10179 4053
tri 10179 4052 10211 4084 nw
tri 10259 4052 10291 4084 se
rect 10291 4052 10478 4084
rect 10530 4052 10787 4104
rect 10919 4166 10925 4179
tri 10925 4166 10938 4179 sw
rect 10919 4151 10938 4166
tri 10938 4151 10953 4166 sw
rect 10919 4127 12394 4151
rect 10867 4113 12394 4127
rect 10919 4099 12394 4113
rect 12446 4099 12460 4151
rect 12512 4099 12984 4151
tri 10919 4079 10939 4099 nw
tri 12822 4079 12842 4099 ne
rect 12842 4079 12984 4099
tri 12842 4068 12853 4079 ne
rect 12853 4068 12984 4079
tri 12853 4067 12854 4068 ne
rect 12854 4067 12984 4068
rect 10867 4055 10919 4061
tri 12190 4055 12202 4067 se
rect 12202 4055 12442 4067
tri 9955 4046 9961 4052 se
rect 9961 4046 10001 4052
tri 10001 4046 10007 4052 nw
tri 10041 4046 10047 4052 se
rect 10047 4046 10087 4052
tri 10087 4046 10093 4052 nw
tri 10127 4046 10133 4052 se
rect 10133 4046 10173 4052
tri 10173 4046 10179 4052 nw
tri 10253 4046 10259 4052 se
rect 10259 4046 10839 4052
tri 12181 4046 12190 4055 se
rect 12190 4046 12442 4055
tri 9947 4038 9955 4046 se
rect 9955 4038 9993 4046
tri 9993 4038 10001 4046 nw
tri 10033 4038 10041 4046 se
rect 10041 4038 10079 4046
tri 10079 4038 10087 4046 nw
tri 10119 4038 10127 4046 se
rect 10127 4038 10165 4046
tri 10165 4038 10173 4046 nw
tri 10245 4038 10253 4046 se
rect 10253 4038 10319 4046
rect 8072 4022 8092 4038
tri 8092 4022 8108 4038 nw
tri 9931 4022 9947 4038 se
rect 9947 4028 9983 4038
tri 9983 4028 9993 4038 nw
tri 10023 4028 10033 4038 se
rect 10033 4028 10063 4038
rect 9947 4022 9977 4028
tri 9977 4022 9983 4028 nw
tri 10017 4022 10023 4028 se
rect 10023 4022 10063 4028
tri 10063 4022 10079 4038 nw
tri 10103 4022 10119 4038 se
rect 10119 4022 10149 4038
tri 10149 4022 10165 4038 nw
tri 10229 4022 10245 4038 se
rect 10245 4022 10319 4038
tri 10319 4022 10343 4046 nw
tri 12157 4022 12181 4046 se
rect 12181 4022 12442 4046
rect 8072 4020 8085 4022
rect 8020 4015 8085 4020
tri 8085 4015 8092 4022 nw
tri 9924 4015 9931 4022 se
rect 9931 4015 9970 4022
tri 9970 4015 9977 4022 nw
tri 10010 4015 10017 4022 se
rect 10017 4015 10056 4022
tri 10056 4015 10063 4022 nw
tri 10096 4015 10103 4022 se
rect 10103 4015 10142 4022
tri 10142 4015 10149 4022 nw
tri 10222 4015 10229 4022 se
rect 10229 4015 10312 4022
tri 10312 4015 10319 4022 nw
tri 12150 4015 12157 4022 se
rect 12157 4015 12442 4022
rect 12494 4015 12506 4067
rect 12558 4015 12564 4067
tri 12854 4065 12856 4067 ne
rect 8020 4008 8077 4015
rect 8072 4007 8077 4008
tri 8077 4007 8085 4015 nw
tri 9916 4007 9924 4015 se
rect 9924 4007 9962 4015
tri 9962 4007 9970 4015 nw
tri 10002 4007 10010 4015 se
rect 10010 4013 10054 4015
tri 10054 4013 10056 4015 nw
tri 10094 4013 10096 4015 se
rect 10096 4013 10134 4015
rect 10010 4007 10048 4013
tri 10048 4007 10054 4013 nw
tri 10088 4007 10094 4013 se
rect 10094 4007 10134 4013
tri 10134 4007 10142 4015 nw
tri 10214 4007 10222 4015 se
rect 10222 4007 10304 4015
tri 10304 4007 10312 4015 nw
tri 12148 4013 12150 4015 se
rect 12150 4013 12216 4015
tri 10557 4007 10563 4013 se
rect 10563 4007 11760 4013
tri 12142 4007 12148 4013 se
rect 12148 4007 12216 4013
tri 12216 4007 12224 4015 nw
tri 8072 4002 8077 4007 nw
rect 8020 3950 8072 3956
rect 8348 4001 9454 4007
rect 8400 3968 9454 4001
rect 8400 3955 8440 3968
tri 8440 3955 8453 3968 nw
tri 9435 3955 9448 3968 ne
rect 9448 3955 9454 3968
rect 9506 3955 9518 4007
rect 9570 3955 9576 4007
tri 9912 4003 9916 4007 se
rect 9916 4003 9958 4007
tri 9958 4003 9962 4007 nw
tri 9998 4003 10002 4007 se
rect 10002 4003 10044 4007
tri 10044 4003 10048 4007 nw
tri 10084 4003 10088 4007 se
rect 10088 4003 10130 4007
tri 10130 4003 10134 4007 nw
tri 10210 4003 10214 4007 se
rect 10214 4003 10300 4007
tri 10300 4003 10304 4007 nw
tri 10553 4003 10557 4007 se
rect 10557 4003 11760 4007
tri 12138 4003 12142 4007 se
rect 12142 4003 12212 4007
tri 12212 4003 12216 4007 nw
tri 9907 3998 9912 4003 se
rect 9912 3998 9953 4003
tri 9953 3998 9958 4003 nw
tri 9993 3998 9998 4003 se
rect 9998 3998 10039 4003
tri 10039 3998 10044 4003 nw
tri 10079 3998 10084 4003 se
rect 10084 3998 10125 4003
tri 10125 3998 10130 4003 nw
tri 10205 3998 10210 4003 se
rect 10210 3998 10295 4003
tri 10295 3998 10300 4003 nw
tri 10548 3998 10553 4003 se
rect 10553 3998 11760 4003
tri 12133 3998 12138 4003 se
rect 12138 3998 12207 4003
tri 12207 3998 12212 4003 nw
tri 9903 3994 9907 3998 se
rect 9907 3994 9949 3998
tri 9949 3994 9953 3998 nw
tri 9989 3994 9993 3998 se
rect 9993 3994 10035 3998
tri 10035 3994 10039 3998 nw
tri 10075 3994 10079 3998 se
rect 10079 3994 10121 3998
tri 10121 3994 10125 3998 nw
tri 10201 3994 10205 3998 se
rect 10205 3994 10291 3998
tri 10291 3994 10295 3998 nw
tri 10544 3994 10548 3998 se
rect 10548 3994 11760 3998
tri 9901 3992 9903 3994 se
rect 9903 3992 9947 3994
tri 9947 3992 9949 3994 nw
tri 9987 3992 9989 3994 se
rect 9989 3992 10033 3994
tri 10033 3992 10035 3994 nw
tri 10073 3992 10075 3994 se
rect 10075 3992 10119 3994
tri 10119 3992 10121 3994 nw
tri 10199 3992 10201 3994 se
rect 10201 3992 10253 3994
tri 9885 3976 9901 3992 se
rect 9901 3982 9937 3992
tri 9937 3982 9947 3992 nw
tri 9977 3982 9987 3992 se
rect 9987 3982 10008 3992
rect 9901 3976 9931 3982
tri 9931 3976 9937 3982 nw
tri 9971 3976 9977 3982 se
rect 9977 3976 10008 3982
tri 9870 3961 9885 3976 se
rect 9885 3961 9916 3976
tri 9916 3961 9931 3976 nw
tri 9956 3961 9971 3976 se
rect 9971 3967 10008 3976
tri 10008 3967 10033 3992 nw
tri 10048 3967 10073 3992 se
rect 10073 3967 10083 3992
rect 9971 3961 10002 3967
tri 10002 3961 10008 3967 nw
tri 10042 3961 10048 3967 se
rect 10048 3961 10083 3967
tri 9865 3956 9870 3961 se
rect 9870 3956 9911 3961
tri 9911 3956 9916 3961 nw
tri 9951 3956 9956 3961 se
rect 9956 3956 9997 3961
tri 9997 3956 10002 3961 nw
tri 10037 3956 10042 3961 se
rect 10042 3956 10083 3961
tri 10083 3956 10119 3992 nw
tri 10163 3956 10199 3992 se
rect 10199 3956 10253 3992
tri 10253 3956 10291 3994 nw
tri 10506 3956 10544 3994 se
rect 10544 3961 11638 3994
rect 10544 3956 10566 3961
tri 9864 3955 9865 3956 se
rect 9865 3955 9910 3956
tri 9910 3955 9911 3956 nw
tri 9950 3955 9951 3956 se
rect 9951 3955 9996 3956
tri 9996 3955 9997 3956 nw
tri 10036 3955 10037 3956 se
rect 10037 3955 10082 3956
tri 10082 3955 10083 3956 nw
tri 10162 3955 10163 3956 se
rect 10163 3955 10239 3956
rect 8400 3949 8427 3955
rect 8348 3942 8427 3949
tri 8427 3942 8440 3955 nw
tri 9855 3946 9864 3955 se
rect 9864 3946 9901 3955
tri 9901 3946 9910 3955 nw
tri 9941 3946 9950 3955 se
rect 9950 3946 9987 3955
tri 9987 3946 9996 3955 nw
tri 10027 3946 10036 3955 se
rect 10036 3946 10073 3955
tri 10073 3946 10082 3955 nw
tri 10153 3946 10162 3955 se
rect 10162 3946 10239 3955
tri 9851 3942 9855 3946 se
rect 9855 3942 9897 3946
tri 9897 3942 9901 3946 nw
tri 9937 3942 9941 3946 se
rect 9941 3942 9983 3946
tri 9983 3942 9987 3946 nw
tri 10023 3942 10027 3946 se
rect 10027 3942 10069 3946
tri 10069 3942 10073 3946 nw
tri 10149 3942 10153 3946 se
rect 10153 3942 10239 3946
tri 10239 3942 10253 3956 nw
tri 10492 3942 10506 3956 se
rect 10506 3942 10566 3956
tri 10566 3942 10585 3961 nw
tri 11590 3942 11609 3961 ne
rect 11609 3942 11638 3961
rect 11690 3942 11702 3994
rect 11754 3942 11760 3994
tri 12110 3975 12133 3998 se
rect 12133 3975 12184 3998
tri 12184 3975 12207 3998 nw
tri 12081 3946 12110 3975 se
rect 12110 3946 12155 3975
tri 12155 3946 12184 3975 nw
rect 8348 3938 8423 3942
tri 8423 3938 8427 3942 nw
tri 9847 3938 9851 3942 se
rect 9851 3938 9893 3942
tri 9893 3938 9897 3942 nw
tri 9933 3938 9937 3942 se
rect 9937 3938 9979 3942
tri 9979 3938 9983 3942 nw
tri 10019 3938 10023 3942 se
rect 10023 3938 10065 3942
tri 10065 3938 10069 3942 nw
tri 10145 3938 10149 3942 se
rect 10149 3938 10235 3942
tri 10235 3938 10239 3942 nw
tri 10489 3939 10492 3942 se
rect 10492 3939 10563 3942
tri 10563 3939 10566 3942 nw
tri 11609 3939 11612 3942 ne
rect 11612 3939 11760 3942
tri 10488 3938 10489 3939 se
rect 10489 3938 10562 3939
tri 10562 3938 10563 3939 nw
tri 11612 3938 11613 3939 ne
rect 11613 3938 11760 3939
tri 12073 3938 12081 3946 se
rect 12081 3938 12147 3946
tri 12147 3938 12155 3946 nw
rect 8348 3937 8400 3938
tri 8400 3915 8423 3938 nw
rect 8649 3886 8655 3938
rect 8707 3886 8719 3938
rect 8771 3886 8978 3938
rect 9030 3886 9042 3938
rect 9094 3886 9296 3938
rect 9348 3886 9360 3938
rect 9412 3886 9418 3938
tri 9841 3932 9847 3938 se
rect 9847 3936 9891 3938
tri 9891 3936 9893 3938 nw
tri 9931 3936 9933 3938 se
rect 9933 3936 9973 3938
rect 9847 3932 9887 3936
tri 9887 3932 9891 3936 nw
tri 9927 3932 9931 3936 se
rect 9931 3932 9973 3936
tri 9973 3932 9979 3938 nw
tri 10013 3932 10019 3938 se
rect 10019 3932 10059 3938
tri 10059 3932 10065 3938 nw
tri 10139 3932 10145 3938 se
rect 10145 3932 10229 3938
tri 10229 3932 10235 3938 nw
tri 10482 3932 10488 3938 se
rect 10488 3932 10556 3938
tri 10556 3932 10562 3938 nw
tri 12067 3932 12073 3938 se
rect 12073 3932 12141 3938
tri 12141 3932 12147 3938 nw
tri 9839 3930 9841 3932 se
rect 9841 3930 9885 3932
tri 9885 3930 9887 3932 nw
tri 9925 3930 9927 3932 se
rect 9927 3930 9968 3932
tri 9836 3927 9839 3930 se
rect 9839 3927 9882 3930
tri 9882 3927 9885 3930 nw
tri 9922 3927 9925 3930 se
rect 9925 3927 9968 3930
tri 9968 3927 9973 3932 nw
tri 10008 3927 10013 3932 se
rect 10013 3927 10054 3932
tri 10054 3927 10059 3932 nw
tri 10134 3927 10139 3932 se
rect 10139 3927 10224 3932
tri 10224 3927 10229 3932 nw
tri 10477 3927 10482 3932 se
rect 10482 3927 10551 3932
tri 10551 3927 10556 3932 nw
tri 12062 3927 12067 3932 se
rect 12067 3927 12136 3932
tri 12136 3927 12141 3932 nw
tri 9830 3921 9836 3927 se
rect 9836 3921 9876 3927
tri 9876 3921 9882 3927 nw
tri 9916 3921 9922 3927 se
rect 9922 3921 9962 3927
tri 9962 3921 9968 3927 nw
tri 10002 3921 10008 3927 se
rect 10008 3921 10048 3927
tri 10048 3921 10054 3927 nw
tri 10128 3921 10134 3927 se
rect 10134 3921 10218 3927
tri 10218 3921 10224 3927 nw
tri 10471 3921 10477 3927 se
rect 10477 3921 10545 3927
tri 10545 3921 10551 3927 nw
rect 10596 3921 11155 3927
tri 9824 3915 9830 3921 se
rect 9830 3915 9870 3921
tri 9870 3915 9876 3921 nw
tri 9910 3915 9916 3921 se
rect 9916 3915 9956 3921
tri 9956 3915 9962 3921 nw
tri 9996 3915 10002 3921 se
rect 10002 3915 10027 3921
tri 9809 3900 9824 3915 se
rect 9824 3900 9855 3915
tri 9855 3900 9870 3915 nw
tri 9895 3900 9910 3915 se
rect 9910 3900 9941 3915
tri 9941 3900 9956 3915 nw
tri 9981 3900 9996 3915 se
rect 9996 3900 10027 3915
tri 10027 3900 10048 3921 nw
tri 10107 3900 10128 3921 se
rect 10128 3900 10166 3921
tri 9795 3886 9809 3900 se
rect 9809 3890 9845 3900
tri 9845 3890 9855 3900 nw
tri 9885 3890 9895 3900 se
rect 9895 3890 9927 3900
rect 9809 3886 9841 3890
tri 9841 3886 9845 3890 nw
tri 9881 3886 9885 3890 se
rect 9885 3886 9927 3890
tri 9927 3886 9941 3900 nw
tri 9967 3886 9981 3900 se
rect 9981 3886 10013 3900
tri 10013 3886 10027 3900 nw
tri 10093 3886 10107 3900 se
rect 10107 3886 10166 3900
rect 8348 3879 8400 3885
tri 9793 3884 9795 3886 se
rect 9795 3884 9839 3886
tri 9839 3884 9841 3886 nw
tri 9879 3884 9881 3886 se
rect 9881 3884 9920 3886
tri 9788 3879 9793 3884 se
rect 9793 3879 9834 3884
tri 9834 3879 9839 3884 nw
tri 9874 3879 9879 3884 se
rect 9879 3879 9920 3884
tri 9920 3879 9927 3886 nw
tri 9960 3879 9967 3886 se
rect 9967 3879 10006 3886
tri 10006 3879 10013 3886 nw
tri 10086 3879 10093 3886 se
rect 10093 3879 10166 3886
tri 9778 3869 9788 3879 se
rect 9788 3869 9824 3879
tri 9824 3869 9834 3879 nw
tri 9864 3869 9874 3879 se
rect 9874 3875 9916 3879
tri 9916 3875 9920 3879 nw
tri 9956 3875 9960 3879 se
rect 9960 3875 9996 3879
rect 9874 3869 9910 3875
tri 9910 3869 9916 3875 nw
tri 9950 3869 9956 3875 se
rect 9956 3869 9996 3875
tri 9996 3869 10006 3879 nw
tri 10076 3869 10086 3879 se
rect 10086 3869 10166 3879
tri 10166 3869 10218 3921 nw
tri 10419 3869 10471 3921 se
rect 10471 3869 10493 3921
tri 10493 3869 10545 3921 nw
rect 10596 3869 11103 3921
tri 12039 3904 12062 3927 se
rect 12062 3904 12113 3927
tri 12113 3904 12136 3927 nw
tri 9775 3866 9778 3869 se
rect 9778 3866 9821 3869
tri 9821 3866 9824 3869 nw
tri 9861 3866 9864 3869 se
rect 9864 3866 9907 3869
tri 9907 3866 9910 3869 nw
tri 9947 3866 9950 3869 se
rect 9950 3866 9993 3869
tri 9993 3866 9996 3869 nw
tri 10073 3866 10076 3869 se
rect 10076 3866 10163 3869
tri 10163 3866 10166 3869 nw
tri 10416 3866 10419 3869 se
rect 10419 3866 10489 3869
tri 9774 3865 9775 3866 se
rect 9775 3865 9811 3866
tri 7672 3856 7681 3865 sw
tri 9765 3856 9774 3865 se
rect 9774 3856 9811 3865
tri 9811 3856 9821 3866 nw
tri 9851 3856 9861 3866 se
rect 9861 3856 9896 3866
rect 7624 3855 7681 3856
tri 7681 3855 7682 3856 sw
tri 8442 3855 8443 3856 se
rect 8443 3855 9810 3856
tri 9810 3855 9811 3856 nw
tri 9850 3855 9851 3856 se
rect 9851 3855 9896 3856
tri 9896 3855 9907 3866 nw
tri 9936 3855 9947 3866 se
rect 9947 3855 9982 3866
tri 9982 3855 9993 3866 nw
tri 10062 3855 10073 3866 se
rect 10073 3855 10152 3866
tri 10152 3855 10163 3866 nw
tri 10415 3865 10416 3866 se
rect 10416 3865 10489 3866
tri 10489 3865 10493 3869 nw
tri 10405 3855 10415 3865 se
rect 10415 3855 10479 3865
tri 10479 3855 10489 3865 nw
rect 10596 3855 11155 3869
rect 7624 3854 7682 3855
tri 7682 3854 7683 3855 sw
tri 8441 3854 8442 3855 se
rect 8442 3854 9809 3855
tri 9809 3854 9810 3855 nw
tri 9849 3854 9850 3855 se
rect 9850 3854 9895 3855
tri 9895 3854 9896 3855 nw
tri 9935 3854 9936 3855 se
rect 9936 3854 9981 3855
tri 9981 3854 9982 3855 nw
tri 10061 3854 10062 3855 se
rect 10062 3854 10100 3855
rect 7624 3853 7683 3854
tri 7683 3853 7684 3854 sw
tri 8440 3853 8441 3854 se
rect 8441 3853 9808 3854
tri 9808 3853 9809 3854 nw
tri 9848 3853 9849 3854 se
rect 9849 3853 9894 3854
tri 9894 3853 9895 3854 nw
tri 9934 3853 9935 3854 se
rect 9935 3853 9980 3854
tri 9980 3853 9981 3854 nw
tri 10060 3853 10061 3854 se
rect 10061 3853 10100 3854
rect 7624 3851 7684 3853
tri 7684 3851 7686 3853 sw
tri 8438 3851 8440 3853 se
rect 8440 3851 9806 3853
tri 9806 3851 9808 3853 nw
tri 9846 3851 9848 3853 se
rect 9848 3851 9892 3853
tri 9892 3851 9894 3853 nw
tri 9932 3851 9934 3853 se
rect 9934 3851 9978 3853
tri 9978 3851 9980 3853 nw
tri 10058 3851 10060 3853 se
rect 10060 3851 10100 3853
rect 7624 3823 7686 3851
tri 7686 3823 7714 3851 sw
tri 8410 3823 8438 3851 se
rect 8438 3823 9778 3851
tri 9778 3823 9806 3851 nw
tri 9818 3823 9846 3851 se
rect 9846 3829 9870 3851
tri 9870 3829 9892 3851 nw
tri 9910 3829 9932 3851 se
rect 9932 3829 9942 3851
rect 9846 3823 9864 3829
tri 9864 3823 9870 3829 nw
tri 9904 3823 9910 3829 se
rect 9910 3823 9942 3829
rect 7624 3822 7714 3823
tri 7714 3822 7715 3823 sw
tri 8409 3822 8410 3823 se
rect 8410 3822 9777 3823
tri 9777 3822 9778 3823 nw
tri 9817 3822 9818 3823 se
rect 9818 3822 9856 3823
rect 7624 3815 8457 3822
tri 8457 3815 8464 3822 nw
tri 9810 3815 9817 3822 se
rect 9817 3815 9856 3822
tri 9856 3815 9864 3823 nw
tri 9896 3815 9904 3823 se
rect 9904 3815 9942 3823
tri 9942 3815 9978 3851 nw
tri 10022 3815 10058 3851 se
rect 10058 3815 10100 3851
rect 7624 3808 8450 3815
tri 8450 3808 8457 3815 nw
tri 9803 3808 9810 3815 se
rect 9810 3808 9849 3815
tri 9849 3808 9856 3815 nw
tri 9889 3808 9896 3815 se
rect 9896 3808 9935 3815
tri 9935 3808 9942 3815 nw
tri 10015 3808 10022 3815 se
rect 10022 3808 10100 3815
rect 7624 3803 8445 3808
tri 8445 3803 8450 3808 nw
tri 9798 3803 9803 3808 se
rect 9803 3803 9844 3808
tri 9844 3803 9849 3808 nw
tri 9884 3803 9889 3808 se
rect 9889 3803 9930 3808
tri 9930 3803 9935 3808 nw
tri 10010 3803 10015 3808 se
rect 10015 3803 10100 3808
tri 10100 3803 10152 3855 nw
tri 10353 3803 10405 3855 se
rect 10405 3803 10427 3855
tri 10427 3803 10479 3855 nw
rect 10596 3803 11103 3855
tri 11712 3853 11763 3904 se
rect 11763 3853 11783 3904
tri 11711 3852 11712 3853 se
rect 11712 3852 11783 3853
rect 11835 3852 11847 3904
rect 11899 3852 11905 3904
tri 12036 3901 12039 3904 se
rect 12039 3901 12110 3904
tri 12110 3901 12113 3904 nw
tri 12015 3880 12036 3901 se
rect 12036 3880 12089 3901
tri 12089 3880 12110 3901 nw
tri 12001 3866 12015 3880 se
rect 12015 3866 12075 3880
tri 12075 3866 12089 3880 nw
tri 11987 3852 12001 3866 se
rect 12001 3852 12061 3866
tri 12061 3852 12075 3866 nw
tri 11710 3851 11711 3852 se
rect 11711 3851 11763 3852
tri 11689 3830 11710 3851 se
rect 11710 3830 11763 3851
tri 11763 3830 11785 3852 nw
tri 11965 3830 11987 3852 se
rect 11987 3830 12039 3852
tri 12039 3830 12061 3852 nw
tri 11674 3815 11689 3830 se
rect 11689 3815 11747 3830
tri 11673 3814 11674 3815 se
rect 11674 3814 11747 3815
tri 11747 3814 11763 3830 nw
tri 11962 3827 11965 3830 se
rect 11965 3827 12036 3830
tri 12036 3827 12039 3830 nw
tri 11949 3814 11962 3827 se
rect 11962 3814 12023 3827
tri 12023 3814 12036 3827 nw
rect 7624 3794 8436 3803
tri 8436 3794 8445 3803 nw
tri 9789 3794 9798 3803 se
rect 9798 3794 9835 3803
tri 9835 3794 9844 3803 nw
tri 9875 3794 9884 3803 se
rect 9884 3794 9911 3803
rect 7624 3786 8428 3794
tri 8428 3786 8436 3794 nw
tri 8489 3786 8497 3794 se
rect 8497 3786 9825 3794
tri 8488 3785 8489 3786 se
rect 8489 3785 9825 3786
tri 7552 3784 7553 3785 sw
tri 8487 3784 8488 3785 se
rect 8488 3784 9825 3785
tri 9825 3784 9835 3794 nw
tri 9865 3784 9875 3794 se
rect 9875 3784 9911 3794
tri 9911 3784 9930 3803 nw
tri 9991 3784 10010 3803 se
rect 10010 3784 10081 3803
tri 10081 3784 10100 3803 nw
tri 10341 3791 10353 3803 se
rect 10353 3791 10415 3803
tri 10415 3791 10427 3803 nw
rect 10596 3797 11155 3803
tri 11656 3797 11673 3814 se
rect 11673 3797 11717 3814
tri 10334 3784 10341 3791 se
rect 10341 3784 10408 3791
tri 10408 3784 10415 3791 nw
rect 10596 3784 10827 3797
tri 10827 3784 10840 3797 nw
tri 11643 3784 11656 3797 se
rect 11656 3784 11717 3797
tri 11717 3784 11747 3814 nw
tri 11919 3784 11949 3814 se
rect 11949 3784 11993 3814
tri 11993 3784 12023 3814 nw
rect 7500 3776 7553 3784
tri 7553 3776 7561 3784 sw
tri 8479 3776 8487 3784 se
rect 8487 3776 9817 3784
tri 9817 3776 9825 3784 nw
tri 9857 3776 9865 3784 se
rect 9865 3776 9903 3784
tri 9903 3776 9911 3784 nw
tri 9983 3776 9991 3784 se
rect 9991 3776 10073 3784
tri 10073 3776 10081 3784 nw
tri 10326 3776 10334 3784 se
rect 10334 3776 10395 3784
rect 7500 3771 7561 3776
tri 7561 3771 7566 3776 sw
tri 8474 3771 8479 3776 se
rect 8479 3771 9812 3776
tri 9812 3771 9817 3776 nw
tri 9852 3771 9857 3776 se
rect 9857 3771 9898 3776
tri 9898 3771 9903 3776 nw
tri 9978 3771 9983 3776 se
rect 9983 3771 10068 3776
tri 10068 3771 10073 3776 nw
tri 10321 3771 10326 3776 se
rect 10326 3771 10395 3776
tri 10395 3771 10408 3784 nw
rect 10596 3771 10814 3784
tri 10814 3771 10827 3784 nw
tri 11630 3771 11643 3784 se
rect 11643 3771 11704 3784
tri 11704 3771 11717 3784 nw
tri 11906 3771 11919 3784 se
rect 11919 3771 11980 3784
tri 11980 3771 11993 3784 nw
rect 7500 3762 7566 3771
tri 7566 3762 7575 3771 sw
tri 8465 3762 8474 3771 se
rect 8474 3762 9803 3771
tri 9803 3762 9812 3771 nw
tri 9843 3762 9852 3771 se
rect 9852 3762 9889 3771
tri 9889 3762 9898 3771 nw
tri 9969 3762 9978 3771 se
rect 9978 3762 10016 3771
rect 7500 3755 7575 3762
tri 7575 3755 7582 3762 sw
tri 8458 3755 8465 3762 se
rect 8465 3755 8523 3762
tri 8523 3755 8530 3762 nw
tri 9836 3755 9843 3762 se
rect 9843 3755 9861 3762
rect 7500 3734 8502 3755
tri 8502 3734 8523 3755 nw
tri 9815 3734 9836 3755 se
rect 9836 3734 9861 3755
tri 9861 3734 9889 3762 nw
tri 9941 3734 9969 3762 se
rect 9969 3734 10016 3762
rect 7500 3719 8487 3734
tri 8487 3719 8502 3734 nw
tri 8574 3719 8589 3734 se
rect 8589 3719 9846 3734
tri 9846 3719 9861 3734 nw
tri 9926 3719 9941 3734 se
rect 9941 3719 10016 3734
tri 10016 3719 10068 3771 nw
tri 10269 3719 10321 3771 se
rect 10321 3719 10343 3771
tri 10343 3719 10395 3771 nw
rect 10596 3756 10799 3771
tri 10799 3756 10814 3771 nw
tri 11615 3756 11630 3771 se
rect 11630 3756 11689 3771
tri 11689 3756 11704 3771 nw
tri 11891 3756 11906 3771 se
rect 11906 3756 11965 3771
tri 11965 3756 11980 3771 nw
rect 10596 3719 10762 3756
tri 10762 3719 10799 3756 nw
tri 11578 3719 11615 3756 se
rect 11615 3719 11652 3756
tri 11652 3719 11689 3756 nw
tri 11888 3753 11891 3756 se
rect 11891 3753 11962 3756
tri 11962 3753 11965 3756 nw
tri 11854 3719 11888 3753 se
rect 11888 3719 11928 3753
tri 11928 3719 11962 3753 nw
rect 7500 3718 8486 3719
tri 8486 3718 8487 3719 nw
tri 8573 3718 8574 3719 se
rect 8574 3718 9845 3719
tri 9845 3718 9846 3719 nw
tri 9925 3718 9926 3719 se
rect 9926 3718 10015 3719
tri 10015 3718 10016 3719 nw
tri 10268 3718 10269 3719 se
rect 10269 3718 10342 3719
tri 10342 3718 10343 3719 nw
rect 10596 3718 10761 3719
tri 10761 3718 10762 3719 nw
tri 11577 3718 11578 3719 se
rect 11578 3718 11651 3719
tri 11651 3718 11652 3719 nw
tri 11853 3718 11854 3719 se
rect 11854 3718 11927 3719
tri 11927 3718 11928 3719 nw
rect 7500 3710 8478 3718
tri 8478 3710 8486 3718 nw
tri 8565 3710 8573 3718 se
rect 8573 3710 9831 3718
tri 8559 3704 8565 3710 se
rect 8565 3704 9831 3710
tri 9831 3704 9845 3718 nw
tri 9911 3704 9925 3718 se
rect 9925 3704 10001 3718
tri 10001 3704 10015 3718 nw
tri 10267 3717 10268 3718 se
rect 10268 3717 10341 3718
tri 10341 3717 10342 3718 nw
tri 10254 3704 10267 3717 se
rect 10267 3704 10328 3717
tri 10328 3704 10341 3717 nw
rect 10596 3704 10747 3718
tri 10747 3704 10761 3718 nw
tri 11563 3704 11577 3718 se
rect 11577 3704 11637 3718
tri 11637 3704 11651 3718 nw
tri 11839 3704 11853 3718 se
rect 11853 3704 11913 3718
tri 11913 3704 11927 3718 nw
tri 8556 3701 8559 3704 se
rect 8559 3702 9829 3704
tri 9829 3702 9831 3704 nw
tri 9909 3702 9911 3704 se
rect 9911 3702 9998 3704
rect 8559 3701 8614 3702
tri 8614 3701 8615 3702 nw
tri 9908 3701 9909 3702 se
rect 9909 3701 9998 3702
tri 9998 3701 10001 3704 nw
tri 10251 3701 10254 3704 se
rect 10254 3701 10325 3704
tri 10325 3701 10328 3704 nw
rect 10596 3701 10744 3704
tri 10744 3701 10747 3704 nw
tri 11560 3701 11563 3704 se
rect 11563 3701 11634 3704
tri 11634 3701 11637 3704 nw
tri 11836 3701 11839 3704 se
rect 11839 3701 11910 3704
tri 11910 3701 11913 3704 nw
tri 8542 3687 8556 3701 se
rect 8556 3687 8600 3701
tri 8600 3687 8614 3701 nw
tri 9894 3687 9908 3701 se
rect 9908 3687 9983 3701
tri 8541 3686 8542 3687 se
rect 8542 3686 8599 3687
tri 8599 3686 8600 3687 nw
tri 9893 3686 9894 3687 se
rect 9894 3686 9983 3687
tri 9983 3686 9998 3701 nw
tri 10236 3686 10251 3701 se
rect 10251 3686 10288 3701
tri 8533 3678 8541 3686 se
rect 8541 3678 8589 3686
tri 1527 3676 1529 3678 sw
tri 8531 3676 8533 3678 se
rect 8533 3676 8589 3678
tri 8589 3676 8599 3686 nw
tri 9883 3676 9893 3686 se
rect 9893 3676 9961 3686
rect 1475 3673 1529 3676
tri 1529 3673 1532 3676 sw
tri 8528 3673 8531 3676 se
rect 8531 3673 8586 3676
tri 8586 3673 8589 3676 nw
tri 9880 3673 9883 3676 se
rect 9883 3673 9961 3676
rect 1475 3669 1532 3673
tri 1532 3669 1536 3673 sw
tri 8524 3669 8528 3673 se
rect 8528 3669 8582 3673
tri 8582 3669 8586 3673 nw
rect 1475 3667 1536 3669
tri 1536 3667 1538 3669 sw
tri 8522 3667 8524 3669 se
rect 8524 3667 8580 3669
tri 8580 3667 8582 3669 nw
rect 8646 3667 8698 3673
tri 9876 3669 9880 3673 se
rect 9880 3669 9961 3673
rect 1475 3653 1538 3667
tri 1538 3653 1552 3667 sw
tri 8508 3653 8522 3667 se
rect 8522 3653 8531 3667
rect 1475 3601 2553 3653
rect 2605 3601 2618 3653
rect 2670 3601 2682 3653
rect 2734 3601 2746 3653
rect 2798 3601 2810 3653
rect 2862 3601 2874 3653
rect 2926 3601 2938 3653
rect 2990 3601 3002 3653
rect 3054 3601 3066 3653
rect 3118 3601 3130 3653
rect 3182 3601 3194 3653
rect 3246 3601 3258 3653
rect 3310 3601 3322 3653
rect 3374 3601 3386 3653
rect 3438 3601 3450 3653
rect 3502 3601 3514 3653
rect 3566 3601 3578 3653
rect 3630 3601 3642 3653
rect 3694 3601 3706 3653
rect 3758 3601 3770 3653
rect 3822 3601 3834 3653
rect 3886 3601 3898 3653
rect 3950 3601 3962 3653
rect 4014 3601 4338 3653
rect 4390 3601 4433 3653
rect 4485 3601 4850 3653
rect 4902 3601 4921 3653
rect 4973 3601 4992 3653
rect 5044 3601 5062 3653
rect 5114 3601 5132 3653
rect 5184 3601 5202 3653
rect 5254 3601 5272 3653
rect 5324 3601 5342 3653
rect 5394 3601 5412 3653
rect 5464 3601 5482 3653
rect 5534 3601 5552 3653
rect 5604 3601 5649 3653
rect 5701 3601 5715 3653
rect 5767 3601 5780 3653
rect 5832 3601 5845 3653
rect 5897 3601 5910 3653
rect 5962 3601 5975 3653
rect 6027 3601 6040 3653
rect 6092 3601 6105 3653
rect 6157 3601 6170 3653
rect 6222 3601 6235 3653
rect 6287 3601 6410 3653
rect 6462 3601 6523 3653
rect 6575 3601 6674 3653
rect 6726 3601 6743 3653
rect 6795 3601 6801 3653
tri 8473 3618 8508 3653 se
rect 8508 3618 8531 3653
tri 8531 3618 8580 3667 nw
tri 8470 3615 8473 3618 se
rect 8473 3615 8528 3618
tri 8528 3615 8531 3618 nw
tri 8467 3612 8470 3615 se
rect 8470 3612 8525 3615
tri 8525 3612 8528 3615 nw
tri 8458 3603 8467 3612 se
rect 8467 3603 8516 3612
tri 8516 3603 8525 3612 nw
rect 8646 3603 8698 3615
rect 9013 3617 9019 3669
rect 9071 3617 9083 3669
rect 9135 3617 9141 3669
tri 9013 3614 9016 3617 ne
rect 9016 3616 9141 3617
rect 9016 3614 9139 3616
tri 9139 3614 9141 3616 nw
rect 9186 3617 9192 3669
rect 9244 3617 9256 3669
rect 9308 3617 9314 3669
tri 9374 3617 9426 3669 se
rect 9426 3617 9648 3669
rect 9700 3617 9712 3669
rect 9764 3617 9770 3669
tri 9871 3664 9876 3669 se
rect 9876 3664 9961 3669
tri 9961 3664 9983 3686 nw
tri 10214 3664 10236 3686 se
rect 10236 3664 10288 3686
tri 10288 3664 10325 3701 nw
rect 10596 3687 10730 3701
tri 10730 3687 10744 3701 nw
tri 11546 3687 11560 3701 se
rect 11560 3687 11615 3701
rect 10596 3682 10725 3687
tri 10725 3682 10730 3687 nw
tri 11541 3682 11546 3687 se
rect 11546 3682 11615 3687
tri 11615 3682 11634 3701 nw
rect 11836 3682 11891 3701
tri 11891 3682 11910 3701 nw
rect 10596 3664 10707 3682
tri 10707 3664 10725 3682 nw
tri 11523 3664 11541 3682 se
rect 11541 3664 11582 3682
tri 9824 3617 9871 3664 se
rect 9871 3617 9909 3664
tri 9186 3614 9189 3617 ne
tri 9016 3612 9018 3614 ne
rect 9018 3612 9137 3614
tri 9137 3612 9139 3614 nw
rect 9189 3612 9270 3617
tri 9270 3612 9275 3617 nw
tri 9369 3612 9374 3617 se
rect 9374 3612 9497 3617
tri 9497 3612 9502 3617 nw
tri 9819 3612 9824 3617 se
rect 9824 3612 9909 3617
tri 9909 3612 9961 3664 nw
tri 10018 3612 10070 3664 se
rect 10070 3612 10077 3664
rect 10129 3612 10141 3664
rect 10193 3649 10273 3664
tri 10273 3649 10288 3664 nw
rect 10596 3653 10696 3664
tri 10696 3653 10707 3664 nw
tri 11512 3653 11523 3664 se
rect 11523 3653 11582 3664
rect 10596 3649 10692 3653
tri 10692 3649 10696 3653 nw
tri 11508 3649 11512 3653 se
rect 11512 3649 11582 3653
tri 11582 3649 11615 3682 nw
rect 10193 3638 10262 3649
tri 10262 3638 10273 3649 nw
rect 10193 3631 10255 3638
tri 10255 3631 10262 3638 nw
rect 10193 3612 10236 3631
tri 10236 3612 10255 3631 nw
tri 8457 3602 8458 3603 se
rect 8458 3602 8515 3603
tri 8515 3602 8516 3603 nw
rect 8457 3601 8514 3602
tri 8514 3601 8515 3602 nw
rect 1475 3485 1527 3601
tri 1527 3576 1552 3601 nw
tri 1527 3485 1552 3510 sw
rect 1475 3433 1778 3485
rect 1830 3433 1844 3485
rect 1896 3433 1910 3485
rect 1962 3433 1976 3485
rect 2028 3433 2042 3485
rect 2094 3433 2108 3485
rect 2160 3433 2174 3485
rect 2226 3433 2240 3485
rect 2292 3433 2306 3485
rect 2358 3433 2372 3485
rect 2424 3433 2437 3485
rect 2489 3433 2502 3485
rect 2554 3433 2567 3485
rect 2619 3433 2632 3485
rect 2684 3433 2697 3485
rect 2749 3433 2762 3485
rect 2814 3433 2827 3485
rect 2879 3433 2892 3485
rect 2944 3433 2957 3485
rect 3009 3433 3022 3485
rect 3074 3433 3087 3485
rect 3139 3433 3152 3485
rect 3204 3433 3217 3485
rect 3269 3433 3282 3485
rect 3334 3433 3347 3485
rect 3399 3433 3412 3485
rect 3464 3433 3477 3485
rect 3529 3433 3542 3485
rect 3594 3433 3607 3485
rect 3659 3433 3672 3485
rect 3724 3433 3855 3485
rect 3907 3433 3922 3485
rect 3974 3433 3989 3485
rect 4041 3433 4056 3485
rect 4108 3433 4123 3485
rect 4175 3433 4189 3485
rect 4241 3433 4367 3485
rect 4419 3433 4434 3485
rect 4486 3433 4501 3485
rect 4553 3433 4568 3485
rect 4620 3433 4635 3485
rect 4687 3433 4701 3485
rect 4753 3433 4879 3485
rect 4931 3433 4986 3485
rect 5038 3433 5618 3485
rect 5670 3433 5684 3485
rect 5736 3433 5750 3485
rect 5802 3433 5816 3485
rect 5868 3433 5882 3485
rect 5934 3433 5948 3485
rect 6000 3433 6014 3485
rect 6066 3433 6079 3485
rect 6131 3433 6144 3485
rect 6196 3433 6209 3485
rect 6261 3433 6274 3485
rect 6326 3433 6339 3485
rect 6391 3433 6404 3485
rect 6456 3433 6469 3485
rect 6521 3433 6534 3485
rect 6586 3433 6674 3485
rect 6726 3433 6743 3485
rect 6795 3433 6801 3485
rect 1102 1773 1232 2436
tri 1232 2427 1241 2436 nw
rect 1334 2372 1386 2384
rect 1475 2376 1527 3433
tri 1527 3408 1552 3433 nw
rect 1575 3351 1581 3403
rect 1633 3397 6986 3403
rect 1633 3351 1974 3397
rect 1575 3345 1974 3351
rect 2026 3345 2486 3397
rect 2538 3369 2998 3397
rect 3050 3369 3510 3397
rect 2538 3345 2689 3369
rect 1575 3333 2689 3345
rect 1575 3327 1974 3333
rect 1575 3275 1581 3327
rect 1633 3281 1974 3327
rect 2026 3281 2486 3333
rect 2538 3313 2689 3333
rect 2745 3313 2771 3369
rect 2827 3313 2853 3369
rect 2909 3313 2935 3369
rect 2991 3345 2998 3369
rect 2991 3333 3017 3345
rect 2991 3313 2998 3333
rect 3073 3313 3099 3369
rect 3155 3313 3180 3369
rect 3236 3313 3261 3369
rect 3317 3313 3342 3369
rect 3398 3313 3423 3369
rect 3479 3313 3504 3369
rect 3562 3345 4022 3397
rect 4074 3345 4534 3397
rect 4586 3345 5046 3397
rect 5098 3345 5302 3397
rect 5354 3345 5558 3397
rect 5610 3345 6070 3397
rect 6122 3345 6582 3397
rect 6634 3351 6986 3397
rect 7038 3351 7085 3403
rect 7137 3351 7184 3403
rect 7236 3351 7283 3403
rect 7335 3351 7382 3403
rect 7434 3351 7712 3403
rect 7764 3351 7820 3403
rect 7872 3351 7878 3403
rect 6634 3345 7878 3351
rect 3560 3333 7878 3345
rect 2538 3281 2998 3313
rect 3050 3281 3510 3313
rect 3562 3281 4022 3333
rect 4074 3281 4534 3333
rect 4586 3281 5046 3333
rect 5098 3281 5302 3333
rect 5354 3281 5558 3333
rect 5610 3281 6070 3333
rect 6122 3281 6582 3333
rect 6634 3327 7878 3333
rect 6634 3281 6986 3327
rect 1633 3275 6986 3281
rect 7038 3275 7085 3327
rect 7137 3275 7184 3327
rect 7236 3275 7283 3327
rect 7335 3275 7382 3327
rect 7434 3275 7712 3327
rect 7764 3275 7820 3327
rect 7872 3275 7878 3327
tri 1575 3274 1576 3275 ne
rect 1576 3272 1799 3275
tri 1799 3272 1802 3275 nw
rect 1576 3248 1775 3272
tri 1775 3248 1799 3272 nw
tri 8433 3248 8457 3272 se
rect 8457 3248 8499 3601
tri 8499 3586 8514 3601 nw
rect 1576 3242 1769 3248
tri 1769 3242 1775 3248 nw
tri 8427 3242 8433 3248 se
rect 8433 3244 8499 3248
rect 8433 3242 8490 3244
rect 1576 3235 1762 3242
tri 1762 3235 1769 3242 nw
rect 1576 3117 1739 3235
tri 1739 3212 1762 3235 nw
rect 3657 3233 3713 3242
tri 8420 3235 8427 3242 se
rect 8427 3235 8490 3242
tri 8490 3235 8499 3244 nw
tri 9018 3601 9029 3612 ne
rect 9029 3601 9115 3612
tri 9029 3590 9040 3601 ne
rect 9040 3590 9115 3601
tri 9115 3590 9137 3612 nw
rect 9189 3608 9266 3612
tri 9266 3608 9270 3612 nw
tri 9365 3608 9369 3612 se
rect 9369 3608 9472 3612
rect 9189 3601 9259 3608
tri 9259 3601 9266 3608 nw
tri 9358 3601 9365 3608 se
rect 9365 3601 9472 3608
rect 2210 3177 3657 3181
tri 4360 3183 4409 3232 se
rect 4409 3184 5791 3232
rect 4409 3183 4438 3184
tri 4438 3183 4439 3184 nw
tri 5765 3183 5766 3184 ne
rect 5766 3183 5791 3184
tri 5791 3183 5840 3232 sw
rect 6283 3183 6289 3235
rect 6341 3183 6353 3235
rect 6405 3222 8477 3235
tri 8477 3222 8490 3235 nw
rect 6405 3220 8475 3222
tri 8475 3220 8477 3222 nw
rect 6405 3209 8464 3220
tri 8464 3209 8475 3220 nw
rect 6405 3183 8438 3209
tri 8438 3183 8464 3209 nw
rect 2210 3155 3713 3177
tri 4339 3162 4360 3183 se
rect 4360 3162 4417 3183
tri 4417 3162 4438 3183 nw
tri 5766 3162 5787 3183 ne
rect 5787 3167 5840 3183
tri 5840 3167 5856 3183 sw
rect 5787 3162 5856 3167
tri 5856 3162 5861 3167 sw
tri 4334 3157 4339 3162 se
rect 4339 3157 4412 3162
tri 4412 3157 4417 3162 nw
tri 5787 3158 5791 3162 ne
rect 5791 3158 5861 3162
tri 5791 3157 5792 3158 ne
rect 5792 3157 5861 3158
tri 8636 3157 8646 3167 se
rect 8646 3157 8698 3551
rect 9040 3579 9104 3590
tri 9104 3579 9115 3590 nw
rect 9040 3572 9097 3579
tri 9097 3572 9104 3579 nw
tri 8698 3157 8708 3167 sw
tri 4332 3155 4334 3157 se
rect 4334 3155 4410 3157
tri 4410 3155 4412 3157 nw
tri 5792 3155 5794 3157 ne
rect 5794 3155 5861 3157
tri 8634 3155 8636 3157 se
rect 8636 3155 8708 3157
tri 8708 3155 8710 3157 sw
rect 1576 3065 1582 3117
rect 1634 3065 1646 3117
rect 1698 3088 1739 3117
rect 1698 3065 1716 3088
tri 1716 3065 1739 3088 nw
rect 1958 3065 1964 3117
rect 2016 3065 2028 3117
rect 2080 3065 2086 3117
rect 2210 3099 2219 3155
rect 2275 3099 2299 3155
rect 2355 3153 3713 3155
tri 4331 3154 4332 3155 se
rect 4332 3154 4409 3155
tri 4409 3154 4410 3155 nw
tri 5794 3154 5795 3155 ne
rect 5795 3154 5861 3155
tri 8633 3154 8634 3155 se
rect 8634 3154 8710 3155
tri 8710 3154 8711 3155 sw
rect 2355 3099 3657 3153
rect 2210 3097 3657 3099
tri 4313 3136 4331 3154 se
rect 4331 3136 4391 3154
tri 4391 3136 4409 3154 nw
tri 5795 3144 5805 3154 ne
tri 4311 3134 4313 3136 se
rect 4313 3134 4389 3136
tri 4389 3134 4391 3136 nw
rect 5029 3134 5131 3136
rect 5187 3134 5260 3136
rect 5316 3134 5429 3136
rect 2210 3087 3713 3097
tri 4307 3130 4311 3134 se
rect 4311 3130 4385 3134
tri 4385 3130 4389 3134 nw
rect 1576 2789 1707 3065
tri 1707 3056 1716 3065 nw
rect 1958 3055 2031 3065
tri 2031 3055 2041 3065 nw
rect 1958 3054 2030 3055
tri 2030 3054 2031 3055 nw
rect 1958 3041 2017 3054
tri 2017 3041 2030 3054 nw
rect 1745 2989 1751 3041
rect 1803 2989 1815 3041
rect 1867 2989 1873 3041
tri 1790 2958 1821 2989 ne
tri 1707 2789 1717 2799 sw
rect 1576 2780 1717 2789
tri 1717 2780 1726 2789 sw
rect 1576 2729 1726 2780
tri 1726 2729 1777 2780 sw
rect 1576 2720 1777 2729
tri 1777 2720 1786 2729 sw
rect 1576 2646 1786 2720
rect 1576 2594 1734 2646
rect 1576 2582 1786 2594
rect 1576 2580 1734 2582
tri 1576 2530 1626 2580 ne
rect 1626 2530 1734 2580
tri 1626 2524 1632 2530 ne
rect 1632 2524 1786 2530
rect 1821 2646 1873 2989
tri 1911 2729 1958 2776 se
rect 1958 2756 2010 3041
tri 2010 3034 2017 3041 nw
rect 1958 2729 1983 2756
tri 1983 2729 2010 2756 nw
rect 1821 2582 1873 2594
rect 1821 2524 1873 2530
tri 1901 2719 1911 2729 se
rect 1911 2719 1973 2729
tri 1973 2719 1983 2729 nw
rect 1901 2646 1953 2719
tri 1953 2699 1973 2719 nw
rect 1901 2582 1953 2594
rect 1901 2524 1953 2530
tri 1632 2508 1648 2524 ne
rect 1648 2508 1786 2524
tri 1648 2456 1700 2508 ne
rect 1700 2456 1786 2508
tri 1786 2456 1838 2508 sw
tri 1700 2450 1706 2456 ne
rect 1706 2450 1838 2456
tri 1838 2450 1844 2456 sw
tri 1706 2415 1741 2450 ne
rect 1741 2415 2757 2450
tri 2757 2415 2792 2450 sw
tri 1527 2376 1566 2415 sw
tri 1741 2403 1753 2415 ne
rect 1753 2403 2792 2415
tri 2792 2403 2804 2415 sw
tri 1753 2396 1760 2403 ne
rect 1760 2396 2804 2403
tri 2721 2376 2741 2396 ne
rect 2741 2376 2804 2396
tri 1475 2364 1487 2376 ne
rect 1487 2364 1566 2376
tri 1566 2364 1578 2376 sw
tri 2741 2364 2753 2376 ne
rect 2753 2364 2804 2376
rect 1334 2314 1386 2320
rect 1487 2358 2692 2364
rect 1539 2312 2692 2358
tri 2753 2355 2762 2364 ne
rect 1539 2308 1582 2312
tri 1582 2308 1586 2312 nw
tri 2270 2308 2274 2312 ne
rect 2274 2308 2692 2312
rect 1539 2306 1554 2308
rect 1487 2294 1554 2306
rect 1539 2242 1554 2294
tri 1554 2280 1582 2308 nw
tri 2274 2280 2302 2308 ne
rect 2302 2280 2692 2308
rect 1487 2236 1554 2242
rect 1616 2274 1668 2280
rect 1821 2274 1873 2280
tri 1820 2226 1821 2227 se
tri 1668 2222 1672 2226 sw
tri 1816 2222 1820 2226 se
rect 1820 2222 1821 2226
tri 2302 2256 2326 2280 ne
rect 2326 2256 2692 2280
tri 2326 2246 2336 2256 ne
rect 2336 2246 2692 2256
tri 2336 2241 2341 2246 ne
rect 2341 2241 2692 2246
tri 2341 2236 2346 2241 ne
rect 2346 2236 2692 2241
rect 1616 2210 1672 2222
tri 1672 2210 1684 2222 sw
tri 1804 2210 1816 2222 se
rect 1816 2210 1873 2222
rect 1668 2192 1684 2210
tri 1684 2192 1702 2210 sw
tri 1786 2192 1804 2210 se
rect 1804 2192 1821 2210
rect 1668 2158 1821 2192
tri 2346 2189 2393 2236 ne
rect 2393 2189 2692 2236
tri 2393 2188 2394 2189 ne
rect 2394 2188 2692 2189
tri 2394 2166 2416 2188 ne
rect 1616 2152 1873 2158
rect 1658 2070 1664 2122
rect 1716 2070 1728 2122
rect 1780 2093 2280 2122
tri 2280 2093 2309 2122 sw
rect 1780 2088 2309 2093
tri 2309 2088 2314 2093 sw
rect 1780 2078 2314 2088
rect 1780 2070 1786 2078
tri 1786 2070 1794 2078 nw
tri 2247 2070 2255 2078 ne
rect 2255 2070 2314 2078
tri 2255 2045 2280 2070 ne
rect 2280 2045 2314 2070
tri 2314 2045 2357 2088 sw
tri 2280 2036 2289 2045 ne
rect 2289 2036 2357 2045
tri 2289 2022 2303 2036 ne
rect 2303 2022 2357 2036
tri 2303 2016 2309 2022 ne
rect 1102 1721 1108 1773
rect 1160 1721 1174 1773
rect 1226 1721 1232 1773
rect 1102 1615 1232 1721
rect 1102 1563 1108 1615
rect 1160 1563 1174 1615
rect 1226 1563 1232 1615
rect 1276 1798 1283 1850
rect 1335 1798 1347 1850
rect 1399 1798 1405 1850
rect 1276 1538 1405 1798
tri 1722 1735 1728 1741 se
rect 1728 1735 1784 1741
rect 1610 1732 1784 1735
rect 1610 1729 1728 1732
rect 1662 1677 1728 1729
rect 1610 1676 1728 1677
rect 1610 1665 1784 1676
rect 1662 1652 1784 1665
rect 1662 1613 1728 1652
rect 1610 1607 1728 1613
tri 1701 1591 1717 1607 ne
rect 1717 1596 1728 1607
rect 1717 1591 1784 1596
tri 1717 1587 1721 1591 ne
rect 1721 1587 1784 1591
rect 1820 1729 1953 1735
rect 1820 1677 1901 1729
rect 1820 1660 1953 1677
rect 1820 1608 1901 1660
rect 1820 1591 1953 1608
tri 1809 1539 1820 1550 se
rect 1820 1539 1901 1591
tri 1808 1538 1809 1539 se
rect 1809 1538 1953 1539
rect 1117 1487 1173 1496
rect 1276 1486 1283 1538
rect 1335 1486 1347 1538
rect 1399 1486 1405 1538
tri 1792 1522 1808 1538 se
rect 1808 1522 1953 1538
tri 1767 1497 1792 1522 se
rect 1792 1497 1901 1522
tri 1405 1486 1416 1497 sw
tri 1756 1486 1767 1497 se
rect 1767 1486 1901 1497
rect 1276 1470 1416 1486
tri 1416 1470 1432 1486 sw
tri 1740 1470 1756 1486 se
rect 1756 1470 1901 1486
rect 1276 1462 1432 1470
tri 1432 1462 1440 1470 sw
tri 1734 1464 1740 1470 se
rect 1740 1464 1953 1470
rect 1276 1460 1440 1462
tri 1276 1456 1280 1460 ne
rect 1280 1456 1440 1460
tri 1440 1456 1446 1462 sw
rect 1734 1456 1953 1464
rect 1117 1407 1173 1431
tri 1280 1404 1332 1456 ne
rect 1332 1404 1446 1456
tri 1446 1404 1498 1456 sw
rect 1786 1452 1953 1456
rect 1786 1404 1901 1452
tri 1332 1400 1336 1404 ne
rect 1336 1400 1498 1404
tri 1498 1400 1502 1404 sw
rect 1734 1400 1901 1404
tri 1336 1387 1349 1400 ne
rect 1349 1387 1502 1400
tri 1502 1387 1515 1400 sw
rect 1734 1391 1953 1400
rect 1734 1387 1949 1391
tri 1949 1387 1953 1391 nw
tri 1349 1381 1355 1387 ne
rect 1355 1381 1515 1387
tri 1515 1381 1521 1387 sw
rect 1734 1381 1943 1387
tri 1943 1381 1949 1387 nw
tri 1355 1377 1359 1381 ne
rect 1359 1377 1521 1381
tri 1521 1377 1525 1381 sw
rect 1734 1377 1929 1381
tri 1359 1357 1379 1377 ne
rect 1379 1357 1525 1377
tri 1525 1357 1545 1377 sw
tri 1100 1325 1117 1342 se
rect 1117 1325 1173 1351
tri 1379 1331 1405 1357 ne
rect 1405 1331 1545 1357
tri 1405 1325 1411 1331 ne
rect 1411 1325 1545 1331
tri 1098 1323 1100 1325 se
rect 1100 1323 1173 1325
rect 1098 1320 1173 1323
tri 1411 1320 1416 1325 ne
rect 1098 1303 1156 1320
tri 1156 1303 1173 1320 nw
rect 1098 1297 1150 1303
tri 1150 1297 1156 1303 nw
rect 1098 -587 1144 1297
tri 1144 1291 1150 1297 nw
rect 1256 1239 1262 1291
rect 1314 1239 1326 1291
rect 1378 1239 1384 1291
rect 1256 976 1384 1239
rect 1256 924 1262 976
rect 1314 924 1326 976
rect 1378 924 1384 976
rect 1174 811 1226 817
rect 1174 747 1226 759
rect 1174 581 1226 695
rect 1174 517 1226 529
rect 1174 -548 1226 465
tri 1174 -550 1176 -548 ne
rect 1176 -550 1226 -548
tri 1176 -554 1180 -550 ne
tri 1144 -587 1150 -581 sw
rect 1098 -593 1150 -587
rect 1098 -657 1150 -645
rect 1098 -715 1150 -709
tri 984 -1103 1011 -1076 se
rect 1011 -1103 1069 -1076
tri 983 -1104 984 -1103 se
rect 984 -1104 1069 -1103
rect 941 -1156 947 -1104
rect 999 -1156 1011 -1104
rect 1063 -1156 1069 -1104
tri 1174 -761 1180 -755 se
rect 1180 -761 1226 -550
rect 950 -1416 959 -1414
rect 1015 -1416 1039 -1414
rect 950 -1468 956 -1416
rect 1015 -1468 1035 -1416
rect 950 -1470 959 -1468
rect 1015 -1470 1039 -1468
rect 1095 -1470 1104 -1414
tri 1172 -1453 1174 -1451 se
rect 1174 -1453 1226 -761
rect 1256 47 1384 924
rect 1416 994 1545 1325
rect 1786 1367 1929 1377
tri 1929 1367 1943 1381 nw
rect 2309 1367 2357 2022
rect 2416 1910 2692 2188
rect 2416 1858 2422 1910
rect 2474 1858 2493 1910
rect 2545 1858 2564 1910
rect 2616 1858 2634 1910
rect 2686 1858 2692 1910
rect 2416 1439 2692 1858
rect 2416 1387 2422 1439
rect 2474 1387 2493 1439
rect 2545 1387 2564 1439
rect 2616 1387 2634 1439
rect 2686 1387 2692 1439
tri 2747 1387 2762 1402 se
rect 2762 1387 2804 2364
tri 4301 2308 4307 2314 se
rect 4307 2308 4363 3130
tri 4363 3108 4385 3130 nw
rect 5029 3082 5035 3134
rect 5087 3082 5102 3134
rect 5221 3082 5236 3134
rect 5355 3082 5371 3134
rect 5423 3082 5429 3134
tri 5029 3075 5036 3082 ne
rect 5036 3080 5131 3082
rect 5187 3080 5260 3082
rect 5316 3080 5422 3082
rect 5036 3075 5135 3080
tri 5135 3075 5140 3080 nw
tri 5312 3075 5317 3080 ne
rect 5317 3075 5422 3080
tri 5422 3075 5429 3082 nw
tri 5036 3065 5046 3075 ne
rect 5046 3065 5125 3075
tri 5125 3065 5135 3075 nw
tri 5317 3065 5327 3075 ne
rect 5327 3065 5412 3075
tri 5412 3065 5422 3075 nw
tri 5046 3055 5056 3065 ne
rect 5056 3055 5115 3065
tri 5115 3055 5125 3065 nw
tri 5327 3055 5337 3065 ne
rect 5337 3055 5402 3065
tri 5402 3055 5412 3065 nw
tri 5056 3054 5057 3055 ne
rect 5057 3054 5114 3055
tri 5114 3054 5115 3055 nw
tri 5337 3054 5338 3055 ne
rect 5338 3054 5401 3055
tri 5401 3054 5402 3055 nw
tri 5057 3053 5058 3054 ne
rect 5058 3053 5113 3054
tri 5113 3053 5114 3054 nw
tri 5338 3053 5339 3054 ne
rect 5339 3053 5400 3054
tri 5400 3053 5401 3054 nw
tri 5058 3052 5059 3053 ne
rect 5059 3052 5112 3053
tri 5112 3052 5113 3053 nw
tri 5339 3052 5340 3053 ne
rect 5340 3052 5396 3053
tri 4249 2256 4301 2308 se
rect 4301 2290 4363 2308
rect 4301 2256 4329 2290
tri 4329 2256 4363 2290 nw
rect 5059 3049 5109 3052
tri 5109 3049 5112 3052 nw
tri 5340 3049 5343 3052 ne
rect 5343 3049 5396 3052
tri 5396 3049 5400 3053 nw
rect 5059 3048 5108 3049
tri 5108 3048 5109 3049 nw
tri 5343 3048 5344 3049 ne
rect 5344 3048 5395 3049
tri 5395 3048 5396 3049 nw
tri 4248 2255 4249 2256 se
rect 4249 2255 4328 2256
tri 4328 2255 4329 2256 nw
rect 4248 2246 4319 2255
tri 4319 2246 4328 2255 nw
rect 4248 2241 4314 2246
tri 4314 2241 4319 2246 nw
tri 2741 1381 2747 1387 se
rect 2747 1381 2804 1387
tri 2732 1372 2741 1381 se
rect 2741 1372 2804 1381
tri 2357 1367 2362 1372 sw
tri 2727 1367 2732 1372 se
rect 2732 1367 2804 1372
rect 1786 1364 1926 1367
tri 1926 1364 1929 1367 nw
rect 2309 1364 2362 1367
tri 2362 1364 2365 1367 sw
tri 2724 1364 2727 1367 se
rect 2727 1364 2804 1367
rect 1786 1355 1917 1364
tri 1917 1355 1926 1364 nw
rect 2309 1355 2365 1364
tri 2365 1355 2374 1364 sw
tri 2715 1355 2724 1364 se
rect 2724 1358 2804 1364
rect 2724 1355 2801 1358
tri 2801 1355 2804 1358 nw
rect 3038 2093 3044 2145
rect 3096 2093 3115 2145
rect 3167 2093 3186 2145
rect 3238 2093 3256 2145
rect 3308 2093 3314 2145
rect 3038 1674 3314 2093
rect 3038 1622 3044 1674
rect 3096 1622 3115 1674
rect 3167 1622 3186 1674
rect 3238 1622 3256 1674
rect 3308 1622 3314 1674
rect 1786 1325 1914 1355
tri 1914 1352 1917 1355 nw
tri 1698 1239 1734 1275 se
rect 1734 1239 1914 1325
rect 2309 1347 2374 1355
tri 2374 1347 2382 1355 sw
tri 2707 1347 2715 1355 se
rect 2715 1347 2793 1355
tri 2793 1347 2801 1355 nw
rect 2309 1336 2782 1347
tri 2782 1336 2793 1347 nw
tri 2309 1303 2342 1336 ne
rect 2342 1303 2749 1336
tri 2749 1303 2782 1336 nw
tri 2342 1300 2345 1303 ne
rect 2345 1300 2746 1303
tri 2746 1300 2749 1303 nw
tri 1692 1233 1698 1239 se
rect 1698 1233 1914 1239
tri 1689 1230 1692 1233 se
rect 1692 1230 1914 1233
tri 1545 994 1546 995 sw
rect 1612 994 1914 1230
rect 3038 1202 3314 1622
rect 3863 1858 3869 1910
rect 3921 1858 3940 1910
rect 3992 1858 4011 1910
rect 4063 1858 4081 1910
rect 4133 1858 4139 1910
rect 3863 1439 4139 1858
rect 3863 1387 3869 1439
rect 3921 1387 3940 1439
rect 3992 1387 4011 1439
rect 4063 1387 4081 1439
rect 4133 1387 4139 1439
tri 4222 1207 4248 1233 se
rect 4248 1207 4304 2241
tri 4304 2231 4314 2241 nw
tri 4220 1205 4222 1207 se
rect 4222 1205 4304 1207
rect 3038 1150 3044 1202
rect 3096 1150 3115 1202
rect 3167 1150 3186 1202
rect 3238 1150 3256 1202
rect 3308 1150 3314 1202
tri 4190 1175 4220 1205 se
rect 4220 1175 4304 1205
rect 3660 1152 3716 1161
rect 1416 993 1546 994
tri 1546 993 1547 994 sw
tri 1612 993 1613 994 ne
rect 1613 993 1914 994
rect 1416 977 1547 993
tri 1547 977 1563 993 sw
tri 1739 977 1755 993 ne
rect 1755 977 1914 993
rect 1416 971 1563 977
tri 1563 971 1569 977 sw
tri 1755 971 1761 977 ne
rect 1761 971 1914 977
rect 1416 948 1569 971
tri 1569 948 1592 971 sw
tri 1761 948 1784 971 ne
rect 1416 946 1592 948
tri 1592 946 1594 948 sw
rect 1416 937 1667 946
rect 1416 881 1609 937
rect 1665 881 1667 937
rect 1416 857 1667 881
rect 1416 801 1609 857
rect 1665 801 1667 857
tri 1778 820 1784 826 se
rect 1784 820 1914 971
rect 3660 1072 3716 1096
rect 3851 1117 4304 1175
tri 3716 1065 3725 1074 sw
rect 3851 1065 3867 1117
rect 3919 1065 3931 1117
rect 3983 1107 4304 1117
rect 3983 1069 4266 1107
tri 4266 1069 4304 1107 nw
rect 4386 2189 4392 2241
rect 4444 2189 4476 2241
rect 4528 2189 4560 2241
rect 4612 2189 4644 2241
rect 4696 2189 4702 2241
rect 4386 2188 4447 2189
tri 4447 2188 4448 2189 nw
tri 4640 2188 4641 2189 ne
rect 4641 2188 4702 2189
rect 4386 2156 4415 2188
tri 4415 2156 4447 2188 nw
tri 4641 2156 4673 2188 ne
rect 4673 2156 4702 2188
rect 3983 1066 4263 1069
tri 4263 1066 4266 1069 nw
tri 4383 1066 4386 1069 se
rect 4386 1066 4414 2156
tri 4414 2155 4415 2156 nw
tri 4673 2155 4674 2156 ne
rect 4463 2088 4620 2094
rect 4515 2036 4568 2088
rect 4463 2022 4620 2036
rect 4515 2018 4620 2022
rect 4515 1970 4568 2018
rect 4463 1966 4568 1970
rect 4463 1955 4620 1966
rect 4515 1947 4620 1955
rect 4515 1903 4568 1947
rect 4463 1895 4568 1903
rect 4463 1888 4620 1895
rect 4515 1876 4620 1888
rect 4515 1836 4568 1876
rect 4463 1824 4568 1836
rect 4463 1821 4620 1824
rect 4515 1805 4620 1821
rect 4515 1769 4568 1805
rect 4463 1754 4568 1769
rect 4515 1753 4568 1754
rect 4515 1734 4620 1753
rect 4515 1702 4568 1734
rect 4463 1687 4568 1702
rect 4515 1682 4568 1687
rect 4515 1645 4620 1682
rect 4515 1635 4597 1645
rect 4463 1622 4597 1635
tri 4597 1622 4620 1645 nw
rect 4463 1620 4568 1622
rect 4515 1593 4568 1620
tri 4568 1593 4597 1622 nw
rect 4515 1568 4567 1593
tri 4567 1592 4568 1593 nw
rect 4463 1553 4567 1568
rect 4515 1501 4567 1553
rect 4463 1495 4567 1501
tri 4463 1491 4467 1495 ne
rect 3983 1065 4262 1066
tri 4262 1065 4263 1066 nw
tri 4382 1065 4383 1066 se
rect 4383 1065 4414 1066
rect 3716 1058 3725 1065
tri 3725 1058 3732 1065 sw
tri 4375 1058 4382 1065 se
rect 4382 1058 4414 1065
rect 3716 1056 3732 1058
tri 3732 1056 3734 1058 sw
tri 4373 1056 4375 1058 se
rect 4375 1056 4414 1058
rect 3716 1046 3734 1056
tri 3734 1046 3744 1056 sw
tri 4363 1046 4373 1056 se
rect 4373 1046 4414 1056
rect 3716 1035 3744 1046
tri 3744 1035 3755 1046 sw
tri 4352 1035 4363 1046 se
rect 4363 1035 4414 1046
rect 3716 1016 4414 1035
rect 3660 1007 4414 1016
rect 4467 1355 4567 1495
rect 4519 1303 4567 1355
rect 4467 1291 4567 1303
rect 4519 1239 4567 1291
tri 4463 1007 4467 1011 se
rect 4467 1007 4567 1239
rect 4674 1066 4702 2156
rect 5059 1110 5106 3048
tri 5106 3046 5108 3048 nw
tri 5344 3046 5346 3048 ne
rect 5160 2989 5166 3041
rect 5218 2989 5230 3041
rect 5282 2989 5288 3041
rect 5160 1153 5288 2989
rect 5346 1192 5393 3048
tri 5393 3046 5395 3048 nw
tri 5778 1155 5805 1182 se
rect 5805 1155 5861 3154
tri 8615 3136 8633 3154 se
rect 8633 3136 8711 3154
tri 8711 3136 8729 3154 sw
tri 8606 3127 8615 3136 se
rect 8615 3127 8729 3136
tri 8729 3127 8738 3136 sw
tri 8266 3099 8294 3127 se
rect 8294 3099 8881 3127
tri 8242 3075 8266 3099 se
rect 8266 3075 8881 3099
rect 8933 3075 8945 3127
rect 8997 3075 9003 3127
tri 8232 3065 8242 3075 se
rect 8242 3065 8296 3075
tri 8222 3055 8232 3065 se
rect 8232 3055 8296 3065
tri 8296 3055 8316 3075 nw
tri 8221 3054 8222 3055 se
rect 8222 3054 8295 3055
tri 8295 3054 8296 3055 nw
tri 8220 3053 8221 3054 se
rect 8221 3053 8294 3054
tri 8294 3053 8295 3054 nw
tri 8216 3049 8220 3053 se
rect 8220 3049 8289 3053
tri 8004 3048 8005 3049 se
rect 8005 3048 8109 3049
tri 8109 3048 8110 3049 sw
tri 8215 3048 8216 3049 se
rect 8216 3048 8289 3049
tri 8289 3048 8294 3053 nw
tri 7645 3041 7652 3048 se
rect 7652 3041 8255 3048
tri 7618 3014 7645 3041 se
rect 7645 3014 8255 3041
tri 8255 3014 8289 3048 nw
tri 7612 3008 7618 3014 se
rect 7618 3008 8249 3014
tri 8249 3008 8255 3014 nw
rect 8470 3008 8851 3014
tri 7578 2974 7612 3008 se
rect 7612 2996 8237 3008
tri 8237 2996 8249 3008 nw
rect 7612 2974 7652 2996
tri 7652 2974 7674 2996 nw
tri 7560 2956 7578 2974 se
rect 7578 2956 7634 2974
tri 7634 2956 7652 2974 nw
rect 8522 2962 8851 3008
rect 8903 2962 8915 3014
rect 8967 2962 8973 3014
tri 7548 2944 7560 2956 se
rect 7560 2944 7622 2956
tri 7622 2944 7634 2956 nw
rect 8470 2944 8522 2956
tri 7535 2931 7548 2944 se
rect 7548 2931 7609 2944
tri 7609 2931 7622 2944 nw
rect 6263 2533 6269 2585
rect 6321 2533 6349 2585
rect 6401 2533 6407 2585
tri 6263 2511 6285 2533 ne
tri 5288 1153 5290 1155 sw
tri 5776 1153 5778 1155 se
rect 5778 1153 5861 1155
rect 5160 1125 5290 1153
tri 5290 1125 5318 1153 sw
tri 5748 1125 5776 1153 se
rect 5776 1125 5861 1153
rect 5160 1118 5318 1125
tri 5318 1118 5325 1125 sw
rect 5160 1106 5518 1118
tri 5160 1069 5197 1106 ne
rect 5197 1069 5518 1106
tri 4702 1066 4705 1069 sw
tri 5197 1066 5200 1069 ne
rect 5200 1066 5518 1069
rect 5570 1066 5582 1118
rect 5634 1066 5640 1118
rect 5733 1073 5739 1125
rect 5791 1073 5803 1125
rect 5855 1073 5861 1125
rect 6048 2094 6054 2146
rect 6106 2094 6118 2146
rect 6170 2094 6176 2146
rect 6048 1674 6176 2094
rect 6048 1622 6054 1674
rect 6106 1622 6118 1674
rect 6170 1622 6176 1674
rect 6048 1123 6176 1622
rect 6048 1071 6054 1123
rect 6106 1071 6118 1123
rect 6170 1071 6176 1123
rect 6204 1349 6256 1355
rect 6204 1285 6256 1297
rect 6204 1110 6256 1233
rect 4674 1058 4705 1066
tri 4705 1058 4713 1066 sw
rect 4674 1056 4713 1058
tri 4713 1056 4715 1058 sw
rect 4674 1046 4715 1056
tri 4715 1046 4725 1056 sw
rect 6204 1046 6256 1058
rect 4674 1035 4725 1046
tri 4725 1035 4736 1046 sw
rect 3660 994 3709 1007
tri 3709 994 3722 1007 nw
tri 4450 994 4463 1007 se
rect 4463 994 4567 1007
tri 4567 994 4584 1011 sw
rect 4674 1007 6090 1035
tri 6090 1007 6118 1035 sw
tri 6078 995 6090 1007 ne
rect 6090 995 6118 1007
tri 6118 995 6130 1007 sw
tri 6090 994 6091 995 ne
rect 6091 994 6130 995
tri 6130 994 6131 995 sw
rect 3660 977 3692 994
tri 3692 977 3709 994 nw
tri 4433 977 4450 994 se
rect 4450 988 4584 994
tri 4584 988 4590 994 sw
tri 6091 988 6097 994 ne
rect 6097 988 6131 994
tri 6131 988 6137 994 sw
rect 6204 988 6256 994
rect 6285 1016 6407 2533
rect 6449 2533 6455 2585
rect 6507 2533 6519 2585
rect 6571 2533 6577 2585
rect 6449 1108 6577 2533
rect 7297 2533 7303 2585
rect 7355 2533 7367 2585
rect 7419 2533 7425 2585
rect 7141 2188 7147 2240
rect 7199 2188 7211 2240
rect 7263 2188 7269 2240
rect 6653 1858 6659 1910
rect 6711 1858 6723 1910
rect 6775 1858 6781 1910
tri 6653 1850 6661 1858 ne
rect 6661 1850 6765 1858
tri 6765 1850 6773 1858 nw
tri 6661 1835 6676 1850 ne
rect 6676 1835 6750 1850
tri 6750 1835 6765 1850 nw
tri 6676 1824 6687 1835 ne
rect 6687 1329 6739 1835
tri 6739 1824 6750 1835 nw
tri 7109 1741 7141 1773 se
rect 7141 1741 7260 2188
tri 7260 2179 7269 2188 nw
rect 7297 1971 7425 2533
tri 7498 2308 7535 2345 se
rect 7535 2308 7587 2931
tri 7587 2909 7609 2931 nw
tri 8522 2928 8556 2962 nw
rect 8470 2886 8522 2892
tri 9027 2866 9040 2879 se
rect 9040 2866 9094 3572
tri 9094 3569 9097 3572 nw
tri 9006 2845 9027 2866 se
rect 9027 2845 9094 2866
rect 7890 2788 9094 2845
rect 9189 2918 9241 3601
tri 9241 3583 9259 3601 nw
tri 9344 3587 9358 3601 se
rect 9358 3587 9472 3601
tri 9472 3587 9497 3612 nw
tri 9803 3596 9819 3612 se
rect 9819 3596 9893 3612
tri 9893 3596 9909 3612 nw
tri 10002 3596 10018 3612 se
rect 10018 3596 10082 3612
tri 9794 3587 9803 3596 se
rect 9803 3587 9876 3596
rect 9344 3441 9472 3587
tri 9786 3579 9794 3587 se
rect 9794 3579 9876 3587
tri 9876 3579 9893 3596 nw
tri 9985 3579 10002 3596 se
rect 10002 3579 10082 3596
tri 10082 3579 10115 3612 nw
tri 9779 3572 9786 3579 se
rect 9786 3572 9869 3579
tri 9869 3572 9876 3579 nw
tri 9978 3572 9985 3579 se
rect 9985 3572 10075 3579
tri 10075 3572 10082 3579 nw
tri 9763 3556 9779 3572 se
rect 9779 3556 9857 3572
tri 9857 3560 9869 3572 nw
tri 9973 3567 9978 3572 se
rect 9978 3567 10070 3572
tri 10070 3567 10075 3572 nw
tri 9966 3560 9973 3567 se
rect 9973 3560 10059 3567
tri 9962 3556 9966 3560 se
rect 9966 3556 10059 3560
tri 10059 3556 10070 3567 nw
tri 9725 3518 9763 3556 se
rect 9763 3518 9857 3556
tri 9713 3506 9725 3518 se
rect 9725 3506 9731 3518
tri 9673 3466 9713 3506 se
rect 9713 3466 9731 3506
rect 9783 3466 9799 3518
rect 9851 3466 9857 3518
tri 9955 3549 9962 3556 se
rect 9962 3549 10052 3556
tri 10052 3549 10059 3556 nw
tri 9671 3464 9673 3466 se
rect 9673 3464 9761 3466
tri 9761 3464 9763 3466 nw
rect 9344 3389 9350 3441
rect 9402 3389 9414 3441
rect 9466 3389 9472 3441
tri 9623 3416 9671 3464 se
rect 9671 3416 9713 3464
tri 9713 3416 9761 3464 nw
tri 9619 3412 9623 3416 se
rect 9623 3412 9709 3416
tri 9709 3412 9713 3416 nw
tri 9596 3389 9619 3412 se
rect 9619 3389 9698 3412
tri 9698 3401 9709 3412 nw
tri 9595 3388 9596 3389 se
rect 9596 3388 9698 3389
tri 9589 3382 9595 3388 se
rect 9595 3382 9698 3388
tri 9566 3359 9589 3382 se
rect 9589 3359 9698 3382
rect 9566 3209 9698 3359
rect 9566 3157 9572 3209
rect 9624 3157 9640 3209
rect 9692 3157 9698 3209
tri 9951 3157 9955 3161 se
rect 9955 3157 10015 3549
tri 10015 3512 10052 3549 nw
tri 9241 2918 9275 2952 sw
rect 9189 2866 9195 2918
rect 9247 2866 9259 2918
rect 9311 2866 9317 2918
rect 7890 2780 8065 2788
tri 8065 2780 8073 2788 nw
rect 7459 2256 7465 2308
rect 7517 2256 7529 2308
rect 7581 2256 7587 2308
tri 7496 2246 7506 2256 ne
rect 7506 2246 7587 2256
tri 7506 2217 7535 2246 ne
rect 7297 1919 7303 1971
rect 7355 1919 7367 1971
rect 7419 1919 7425 1971
tri 7107 1739 7109 1741 se
rect 7109 1739 7260 1741
rect 7001 1715 7260 1739
rect 7001 1663 7007 1715
rect 7059 1663 7105 1715
rect 7157 1663 7202 1715
rect 7254 1663 7260 1715
rect 7001 1639 7260 1663
rect 7535 1722 7587 2246
rect 7658 2533 7664 2585
rect 7716 2533 7728 2585
rect 7780 2533 7786 2585
rect 7658 2246 7786 2533
rect 7658 2194 7664 2246
rect 7716 2194 7728 2246
rect 7780 2194 7786 2246
rect 7890 1835 8035 2780
tri 8035 2750 8065 2780 nw
rect 8348 2729 8400 2735
tri 8400 2728 8407 2735 sw
rect 8400 2716 8407 2728
tri 8407 2716 8419 2728 sw
rect 8400 2710 8419 2716
tri 8419 2710 8425 2716 sw
rect 8400 2677 8868 2710
rect 8348 2665 8868 2677
rect 8087 2613 8093 2665
rect 8145 2613 8157 2665
rect 8209 2630 8248 2665
tri 8248 2630 8283 2665 sw
rect 8209 2613 8283 2630
tri 8283 2613 8300 2630 sw
rect 8400 2658 8868 2665
rect 8920 2658 8932 2710
rect 8984 2658 8990 2710
rect 8400 2640 8416 2658
tri 8416 2640 8434 2658 nw
rect 8400 2630 8406 2640
tri 8406 2630 8416 2640 nw
tri 8400 2624 8406 2630 nw
tri 8627 2624 8633 2630 se
rect 8633 2624 8865 2630
tri 8616 2613 8627 2624 se
rect 8627 2613 8865 2624
tri 8226 2578 8261 2613 ne
rect 8261 2578 8300 2613
tri 8300 2578 8335 2613 sw
rect 8348 2607 8400 2613
tri 8610 2607 8616 2613 se
rect 8616 2607 8865 2613
tri 8581 2578 8610 2607 se
rect 8610 2578 8865 2607
rect 8917 2578 8929 2630
rect 8981 2578 8987 2630
tri 8261 2560 8279 2578 ne
rect 8279 2566 8335 2578
tri 8335 2566 8347 2578 sw
tri 8569 2566 8581 2578 se
rect 8581 2566 8637 2578
rect 8279 2560 8637 2566
tri 8637 2560 8655 2578 nw
tri 8279 2539 8300 2560 ne
rect 8300 2539 8616 2560
tri 8616 2539 8637 2560 nw
tri 8300 2524 8315 2539 ne
rect 8315 2524 8591 2539
tri 8315 2514 8325 2524 ne
rect 8325 2514 8591 2524
tri 8591 2514 8616 2539 nw
rect 8090 2456 8096 2508
rect 8148 2456 8160 2508
rect 8212 2456 8218 2508
rect 8090 2220 8218 2456
tri 9167 2278 9189 2300 se
rect 9189 2278 9241 2866
tri 9241 2832 9275 2866 nw
rect 8601 2272 8653 2278
tri 8218 2220 8248 2250 sw
tri 8653 2266 8665 2278 sw
tri 9155 2266 9167 2278 se
rect 9167 2266 9241 2278
rect 8653 2220 9241 2266
rect 8090 2208 8248 2220
tri 8248 2208 8260 2220 sw
rect 8601 2214 9241 2220
rect 8601 2208 8653 2214
rect 8090 2196 8260 2208
tri 8090 2156 8130 2196 ne
rect 8130 2156 8260 2196
tri 8260 2156 8312 2208 sw
tri 8653 2180 8687 2214 nw
tri 8130 2138 8148 2156 ne
rect 8148 2150 8312 2156
tri 8312 2150 8318 2156 sw
rect 8601 2150 8653 2156
rect 8148 2138 8318 2150
tri 8318 2138 8330 2150 sw
tri 8148 2121 8165 2138 ne
rect 8165 2121 8330 2138
tri 8330 2121 8347 2138 sw
tri 8165 2086 8200 2121 ne
rect 8200 2086 9369 2121
tri 9369 2086 9404 2121 sw
tri 8200 2075 8211 2086 ne
rect 8211 2075 9404 2086
tri 9404 2075 9415 2086 sw
tri 8211 2068 8218 2075 ne
rect 8218 2068 9415 2075
tri 8218 2052 8234 2068 ne
rect 8234 2052 9415 2068
tri 9415 2052 9438 2075 sw
tri 8234 2033 8253 2052 ne
rect 8253 2033 9438 2052
tri 9299 2026 9306 2033 ne
rect 9306 2026 9438 2033
tri 9438 2026 9464 2052 sw
tri 9306 2013 9319 2026 ne
rect 9319 2013 9464 2026
tri 9319 1990 9342 2013 ne
rect 9342 1990 9401 2013
tri 9195 1984 9201 1990 se
rect 9201 1984 9253 1990
tri 9182 1971 9195 1984 se
rect 9195 1971 9201 1984
rect 8137 1919 8143 1971
rect 8195 1919 8207 1971
rect 8259 1932 9201 1971
tri 9342 1963 9369 1990 ne
rect 9369 1963 9401 1990
tri 9369 1961 9371 1963 ne
rect 9371 1961 9401 1963
rect 9453 1961 9464 2013
tri 9371 1956 9376 1961 ne
rect 8259 1920 9253 1932
rect 8259 1919 9201 1920
tri 9167 1885 9201 1919 ne
rect 9201 1862 9253 1868
rect 9376 1932 9464 1961
rect 9376 1880 9401 1932
rect 9453 1880 9464 1932
rect 7890 1783 7896 1835
rect 7948 1783 7977 1835
rect 8029 1783 8035 1835
rect 9376 1850 9464 1880
rect 9376 1798 9401 1850
rect 9453 1798 9464 1850
rect 9376 1784 9464 1798
rect 8598 1774 9255 1780
tri 7587 1722 7596 1731 sw
rect 8650 1722 9203 1774
rect 7535 1710 7596 1722
tri 7596 1710 7608 1722 sw
rect 8598 1710 9255 1722
rect 7535 1709 7608 1710
tri 7608 1709 7609 1710 sw
tri 7535 1658 7586 1709 ne
rect 7586 1658 7609 1709
tri 7609 1658 7660 1709 sw
rect 8650 1658 9203 1710
tri 7586 1652 7592 1658 ne
rect 7592 1652 7660 1658
tri 7660 1652 7666 1658 sw
rect 8598 1652 9255 1658
tri 7592 1645 7599 1652 ne
rect 7599 1645 7666 1652
tri 7666 1645 7673 1652 sw
tri 7107 1605 7141 1639 ne
rect 7141 1433 7260 1639
tri 7599 1635 7609 1645 ne
rect 7609 1635 7673 1645
tri 7673 1635 7683 1645 sw
tri 7609 1593 7651 1635 ne
rect 7651 1593 7683 1635
tri 7683 1593 7725 1635 sw
tri 7651 1561 7683 1593 ne
rect 7683 1561 7725 1593
tri 7725 1561 7757 1593 sw
tri 7683 1550 7694 1561 ne
rect 7694 1550 7757 1561
tri 7757 1550 7768 1561 sw
tri 7694 1544 7700 1550 ne
rect 7700 1544 7768 1550
tri 7768 1544 7774 1550 sw
tri 7700 1537 7707 1544 ne
rect 7707 1537 7774 1544
tri 7774 1537 7781 1544 sw
tri 7707 1514 7730 1537 ne
rect 7730 1514 7781 1537
tri 7781 1514 7804 1537 sw
tri 7730 1487 7757 1514 ne
rect 7757 1487 7804 1514
tri 7804 1487 7831 1514 sw
tri 7757 1462 7782 1487 ne
rect 7782 1462 7831 1487
tri 7831 1462 7856 1487 sw
tri 7782 1443 7801 1462 ne
rect 7801 1443 7856 1462
tri 7856 1443 7875 1462 sw
rect 7141 1381 7142 1433
rect 7194 1381 7208 1433
tri 7801 1413 7831 1443 ne
rect 7831 1413 7875 1443
tri 7875 1413 7905 1443 sw
tri 7831 1391 7853 1413 ne
rect 7853 1391 7905 1413
tri 7905 1391 7927 1413 sw
rect 7141 1364 7260 1381
tri 7853 1367 7877 1391 ne
rect 7877 1367 7927 1391
tri 7927 1367 7951 1391 sw
tri 6739 1329 6774 1364 sw
rect 6687 1323 7048 1329
rect 6687 1271 6996 1323
rect 6687 1263 7048 1271
tri 6934 1259 6938 1263 ne
rect 6938 1259 7048 1263
tri 6938 1207 6990 1259 ne
rect 6990 1207 6996 1259
tri 6990 1205 6992 1207 ne
rect 6992 1205 7048 1207
rect 6449 1056 6455 1108
rect 6507 1056 6519 1108
rect 6571 1056 6577 1108
rect 6802 1153 6808 1205
rect 6860 1153 6872 1205
rect 6924 1172 6930 1205
tri 6992 1201 6996 1205 ne
rect 6996 1201 7048 1205
rect 7141 1312 7142 1364
rect 7194 1312 7208 1364
tri 7877 1339 7905 1367 ne
rect 7905 1339 7951 1367
tri 7951 1339 7979 1367 sw
tri 7905 1315 7929 1339 ne
rect 7929 1315 7979 1339
tri 7979 1315 8003 1339 sw
rect 7141 1294 7260 1312
tri 7929 1299 7945 1315 ne
rect 7945 1299 8003 1315
rect 7141 1242 7142 1294
rect 7194 1242 7208 1294
rect 7141 1224 7260 1242
tri 6930 1172 6937 1179 sw
rect 7141 1172 7142 1224
rect 7194 1172 7208 1224
rect 7419 1293 7897 1299
rect 7419 1241 7501 1293
rect 7553 1241 7673 1293
rect 7725 1241 7845 1293
tri 7945 1282 7962 1299 ne
rect 7962 1282 8003 1299
tri 8003 1282 8036 1315 sw
tri 7962 1275 7969 1282 ne
rect 7969 1275 8036 1282
tri 8036 1275 8043 1282 sw
tri 7969 1265 7979 1275 ne
rect 7979 1265 8043 1275
tri 8043 1265 8053 1275 sw
rect 7419 1229 7897 1241
tri 7397 1177 7419 1199 se
rect 7419 1177 7501 1229
rect 7553 1177 7673 1229
rect 7725 1177 7845 1229
tri 7979 1223 8021 1265 ne
rect 8021 1223 8053 1265
tri 8053 1223 8095 1265 sw
tri 8021 1216 8028 1223 ne
rect 8028 1216 8095 1223
tri 8095 1216 8102 1223 sw
tri 8028 1191 8053 1216 ne
rect 8053 1191 8431 1216
rect 6924 1166 6937 1172
tri 6937 1166 6943 1172 sw
rect 7141 1166 7260 1172
tri 7386 1166 7397 1177 se
rect 7397 1171 7897 1177
tri 8053 1171 8073 1191 ne
rect 8073 1171 8431 1191
rect 7397 1166 7546 1171
rect 6924 1164 6943 1166
tri 6943 1164 6945 1166 sw
tri 7384 1164 7386 1166 se
rect 7386 1164 7546 1166
tri 7546 1164 7553 1171 nw
tri 8073 1164 8080 1171 ne
rect 8080 1164 8431 1171
rect 8483 1164 8509 1216
rect 8561 1164 8587 1216
rect 8639 1164 8665 1216
rect 8717 1164 8743 1216
rect 8795 1164 8801 1216
rect 6924 1153 6945 1164
rect 6802 1138 6945 1153
tri 6945 1138 6971 1164 sw
tri 7358 1138 7384 1164 se
rect 7384 1138 7520 1164
tri 7520 1138 7546 1164 nw
rect 6802 1125 7507 1138
tri 7507 1125 7520 1138 nw
tri 9556 1125 9566 1135 se
rect 9566 1125 9698 3157
tri 9948 3154 9951 3157 se
rect 9951 3154 10015 3157
tri 9930 3136 9948 3154 se
rect 9948 3136 10015 3154
tri 9921 3127 9930 3136 se
rect 9930 3127 10015 3136
rect 9887 3075 9893 3127
rect 9945 3075 9957 3127
rect 10009 3075 10015 3127
rect 10064 3055 10070 3107
rect 10122 3055 10134 3107
rect 10186 3055 10192 3107
rect 10064 3054 10131 3055
tri 10131 3054 10132 3055 nw
tri 10043 2918 10064 2939 se
rect 10064 2918 10104 3054
tri 10104 3027 10131 3054 nw
tri 10036 2911 10043 2918 se
rect 10043 2911 10104 2918
rect 9968 2871 10104 2911
rect 9968 2868 10033 2871
tri 10033 2868 10036 2871 nw
tri 9966 2170 9968 2172 se
rect 9968 2170 10008 2868
tri 10008 2843 10033 2868 nw
rect 10596 2664 10686 3649
tri 10686 3643 10692 3649 nw
tri 11502 3643 11508 3649 se
rect 11508 3643 11571 3649
tri 11497 3638 11502 3643 se
rect 11502 3638 11571 3643
tri 11571 3638 11582 3649 nw
tri 11490 3631 11497 3638 se
rect 11497 3631 11564 3638
tri 11564 3631 11571 3638 nw
tri 11467 3608 11490 3631 se
rect 11490 3608 11541 3631
tri 11541 3608 11564 3631 nw
tri 11460 3601 11467 3608 se
rect 11467 3601 11512 3608
tri 11438 3579 11460 3601 se
rect 11460 3579 11512 3601
tri 11512 3579 11541 3608 nw
tri 11431 3572 11438 3579 se
rect 11438 3572 11505 3579
tri 11505 3572 11512 3579 nw
tri 11415 3556 11431 3572 se
rect 11431 3556 11489 3572
tri 11489 3556 11505 3572 nw
rect 10717 3504 10723 3556
rect 10775 3504 10787 3556
rect 10839 3520 11453 3556
tri 11453 3520 11489 3556 nw
rect 10839 3506 11439 3520
tri 11439 3506 11453 3520 nw
rect 10839 3504 11437 3506
tri 11437 3504 11439 3506 nw
tri 11814 3465 11836 3487 se
rect 11836 3465 11888 3682
tri 11888 3679 11891 3682 nw
tri 11813 3464 11814 3465 se
rect 11814 3464 11887 3465
tri 11887 3464 11888 3465 nw
rect 11091 3412 11097 3464
rect 11149 3412 11161 3464
rect 11213 3412 11580 3464
rect 11632 3412 11644 3464
rect 11696 3412 11702 3464
tri 11761 3412 11813 3464 se
rect 11813 3412 11835 3464
tri 11835 3412 11887 3464 nw
tri 11751 3402 11761 3412 se
rect 11761 3402 11825 3412
tri 11825 3402 11835 3412 nw
tri 11737 3388 11751 3402 se
rect 11751 3388 11811 3402
tri 11811 3388 11825 3402 nw
tri 11731 3382 11737 3388 se
rect 11737 3382 11805 3388
tri 11805 3382 11811 3388 nw
tri 11679 3330 11731 3382 se
rect 11731 3330 11753 3382
tri 11753 3330 11805 3382 nw
tri 11677 3328 11679 3330 se
rect 11679 3328 11751 3330
tri 11751 3328 11753 3330 nw
tri 11649 3300 11677 3328 se
rect 11677 3300 11723 3328
tri 11723 3300 11751 3328 nw
tri 11603 3254 11649 3300 se
rect 11649 3254 11677 3300
tri 11677 3254 11723 3300 nw
tri 11597 3248 11603 3254 se
rect 11603 3248 11671 3254
tri 11671 3248 11677 3254 nw
tri 11571 3222 11597 3248 se
rect 11597 3222 11645 3248
tri 11645 3222 11671 3248 nw
tri 11569 3220 11571 3222 se
rect 11571 3220 11643 3222
tri 11643 3220 11645 3222 nw
rect 10791 3168 10797 3220
rect 10849 3168 10869 3220
rect 10921 3168 10941 3220
rect 10993 3168 11012 3220
rect 11064 3168 11083 3220
rect 11135 3168 11141 3220
tri 11567 3218 11569 3220 se
rect 11569 3218 11641 3220
tri 11641 3218 11643 3220 nw
tri 11529 3180 11567 3218 se
rect 11567 3180 11603 3218
tri 11603 3180 11641 3218 nw
tri 10879 3166 10881 3168 ne
rect 10881 3166 11141 3168
tri 11515 3166 11529 3180 se
rect 11529 3166 11589 3180
tri 11589 3166 11603 3180 nw
tri 10881 3154 10893 3166 ne
rect 10893 3154 11141 3166
tri 11503 3154 11515 3166 se
rect 11515 3154 11577 3166
tri 11577 3154 11589 3166 nw
tri 10893 3136 10911 3154 ne
rect 10911 3136 11141 3154
tri 11485 3136 11503 3154 se
rect 11503 3136 11559 3154
tri 11559 3136 11577 3154 nw
tri 10911 3116 10931 3136 ne
rect 10769 2816 10775 2868
rect 10827 2816 10839 2868
rect 10891 2816 10897 2868
tri 10686 2664 10697 2675 sw
rect 10596 2640 10697 2664
tri 10697 2640 10721 2664 sw
rect 10596 2630 10721 2640
tri 10721 2630 10731 2640 sw
rect 10092 2578 10098 2630
rect 10150 2578 10206 2630
rect 10258 2578 10314 2630
rect 10366 2578 10372 2630
rect 10596 2578 10602 2630
rect 10654 2578 10673 2630
rect 10725 2578 10731 2630
tri 10008 2170 10010 2172 sw
tri 9946 2150 9966 2170 se
rect 9966 2150 10010 2170
tri 9934 2138 9946 2150 se
rect 9946 2138 10010 2150
tri 10010 2138 10042 2170 sw
rect 9923 2086 9929 2138
rect 9981 2086 9993 2138
rect 10045 2086 10051 2138
rect 6802 1081 7463 1125
tri 7463 1081 7507 1125 nw
tri 9532 1101 9556 1125 se
rect 9556 1101 9698 1125
tri 7580 1081 7600 1101 se
rect 7600 1081 9698 1101
rect 6802 1079 7461 1081
tri 7461 1079 7463 1081 nw
tri 7578 1079 7580 1081 se
rect 7580 1079 9698 1081
rect 6802 1071 7453 1079
tri 7453 1071 7461 1079 nw
tri 7570 1071 7578 1079 se
rect 7578 1071 9698 1079
rect 6802 1027 7409 1071
tri 7409 1027 7453 1071 nw
tri 7526 1027 7570 1071 se
rect 7570 1049 9698 1071
rect 10092 1462 10372 2578
rect 10601 2170 10607 2222
rect 10659 2170 10671 2222
rect 10723 2170 10729 2222
rect 10769 2180 10897 2816
rect 10931 2395 11141 3136
tri 11477 3128 11485 3136 se
rect 11485 3128 11529 3136
rect 11477 2780 11529 3128
tri 11529 3106 11559 3136 nw
rect 12856 2962 12984 4067
rect 13077 4068 13083 4120
rect 13135 4068 13147 4120
rect 13199 4068 13205 4120
rect 13077 3464 13205 4068
rect 13077 3412 13083 3464
rect 13135 3412 13147 3464
rect 13199 3412 13205 3464
rect 13241 3464 13369 4211
rect 13241 3412 13247 3464
rect 13299 3412 13311 3464
rect 13363 3412 13369 3464
rect 12856 2910 12862 2962
rect 12914 2910 12926 2962
rect 12978 2910 12984 2962
rect 11477 2716 11529 2728
rect 11477 2658 11529 2664
tri 11141 2395 11205 2459 sw
rect 10931 2334 14187 2395
tri 10931 2235 11030 2334 ne
rect 11030 2235 14187 2334
tri 13744 2193 13786 2235 ne
rect 13786 2193 14187 2235
tri 10897 2180 10910 2193 sw
tri 13786 2180 13799 2193 ne
rect 10769 2170 10910 2180
tri 10910 2170 10920 2180 sw
rect 10769 2075 10920 2170
tri 10920 2075 11015 2170 sw
tri 10756 2052 10769 2065 se
rect 10769 2052 11015 2075
tri 11015 2052 11038 2075 sw
rect 10756 2000 10775 2052
rect 10827 2000 10839 2052
rect 10891 2000 10927 2052
rect 10979 2000 10992 2052
rect 11044 2000 11057 2052
rect 11109 2000 11122 2052
rect 11174 2000 11187 2052
rect 11239 2000 11252 2052
rect 11304 2000 11317 2052
rect 11369 2000 11382 2052
rect 11434 2000 11447 2052
rect 11499 2000 11512 2052
rect 11564 2000 11577 2052
rect 11629 2000 11642 2052
rect 11694 2000 11707 2052
rect 11759 2000 11772 2052
rect 11824 2000 11837 2052
rect 11889 2000 11901 2052
rect 11953 2000 11965 2052
rect 12017 2000 12029 2052
rect 12081 2000 12093 2052
rect 12145 2000 12157 2052
rect 12209 2000 12221 2052
rect 12273 2000 12285 2052
rect 12337 2000 12349 2052
rect 12401 2000 12413 2052
rect 12465 2000 12477 2052
rect 12529 2000 12541 2052
rect 12593 2000 12605 2052
rect 12657 2000 12669 2052
rect 12721 2000 12733 2052
rect 12785 2000 12797 2052
rect 12849 2000 12861 2052
rect 12913 2000 12925 2052
rect 12977 2000 12989 2052
rect 13041 2000 13053 2052
rect 13105 2000 13117 2052
rect 13169 2000 13181 2052
rect 13233 2000 13245 2052
rect 13297 2000 13309 2052
rect 13361 2000 13373 2052
rect 13425 2000 13437 2052
rect 13489 2000 13495 2052
rect 10756 1885 12417 2000
tri 12417 1885 12532 2000 nw
rect 10756 1833 10762 1885
rect 10814 1833 10829 1885
rect 10881 1833 10896 1885
rect 10948 1833 10963 1885
rect 11015 1833 11030 1885
rect 11082 1833 11097 1885
rect 11149 1833 11164 1885
rect 11216 1833 11231 1885
rect 11283 1833 11298 1885
rect 11350 1833 11365 1885
rect 11417 1833 11432 1885
rect 11484 1833 11499 1885
rect 11551 1833 11566 1885
rect 11618 1833 11633 1885
rect 11685 1833 11699 1885
rect 11751 1833 11765 1885
rect 11817 1833 11831 1885
rect 11883 1833 11897 1885
rect 11949 1833 11963 1885
rect 12015 1833 12029 1885
rect 12081 1833 12095 1885
rect 12147 1833 12161 1885
rect 12213 1833 12227 1885
rect 12279 1833 12293 1885
rect 12345 1833 12359 1885
rect 12411 1833 12417 1885
rect 10756 1805 12417 1833
rect 10756 1753 10762 1805
rect 10814 1753 10829 1805
rect 10881 1753 10896 1805
rect 10948 1753 10963 1805
rect 11015 1753 11030 1805
rect 11082 1753 11097 1805
rect 11149 1753 11164 1805
rect 11216 1753 11231 1805
rect 11283 1753 11298 1805
rect 11350 1753 11365 1805
rect 11417 1753 11432 1805
rect 11484 1753 11499 1805
rect 11551 1753 11566 1805
rect 11618 1753 11633 1805
rect 11685 1753 11699 1805
rect 11751 1753 11765 1805
rect 11817 1753 11831 1805
rect 11883 1753 11897 1805
rect 11949 1753 11963 1805
rect 12015 1753 12029 1805
rect 12081 1753 12095 1805
rect 12147 1753 12161 1805
rect 12213 1753 12227 1805
rect 12279 1753 12293 1805
rect 12345 1753 12359 1805
rect 12411 1753 12417 1805
rect 10756 1725 12417 1753
rect 10756 1673 10762 1725
rect 10814 1673 10829 1725
rect 10881 1673 10896 1725
rect 10948 1673 10963 1725
rect 11015 1673 11030 1725
rect 11082 1673 11097 1725
rect 11149 1673 11164 1725
rect 11216 1673 11231 1725
rect 11283 1673 11298 1725
rect 11350 1673 11365 1725
rect 11417 1673 11432 1725
rect 11484 1673 11499 1725
rect 11551 1673 11566 1725
rect 11618 1673 11633 1725
rect 11685 1673 11699 1725
rect 11751 1673 11765 1725
rect 11817 1673 11831 1725
rect 11883 1673 11897 1725
rect 11949 1673 11963 1725
rect 12015 1673 12029 1725
rect 12081 1673 12095 1725
rect 12147 1673 12161 1725
rect 12213 1673 12227 1725
rect 12279 1673 12293 1725
rect 12345 1673 12359 1725
rect 12411 1673 12417 1725
rect 10756 1645 12417 1673
rect 10756 1593 10762 1645
rect 10814 1593 10829 1645
rect 10881 1593 10896 1645
rect 10948 1593 10963 1645
rect 11015 1593 11030 1645
rect 11082 1593 11097 1645
rect 11149 1593 11164 1645
rect 11216 1593 11231 1645
rect 11283 1593 11298 1645
rect 11350 1593 11365 1645
rect 11417 1593 11432 1645
rect 11484 1593 11499 1645
rect 11551 1593 11566 1645
rect 11618 1593 11633 1645
rect 11685 1593 11699 1645
rect 11751 1593 11765 1645
rect 11817 1593 11831 1645
rect 11883 1593 11897 1645
rect 11949 1593 11963 1645
rect 12015 1593 12029 1645
rect 12081 1593 12095 1645
rect 12147 1593 12161 1645
rect 12213 1593 12227 1645
rect 12279 1593 12293 1645
rect 12345 1593 12359 1645
rect 12411 1593 12417 1645
tri 10372 1462 10377 1467 sw
rect 10092 1443 10377 1462
tri 10377 1443 10396 1462 sw
rect 10092 1391 10396 1443
tri 10396 1391 10448 1443 sw
rect 10092 1367 10448 1391
tri 10448 1367 10472 1391 sw
rect 10092 1315 10472 1367
tri 10472 1315 10524 1367 sw
rect 12258 1315 12264 1367
rect 12316 1315 12328 1367
rect 12380 1315 13501 1367
rect 13553 1315 13565 1367
rect 13617 1315 13623 1367
rect 13799 1315 14187 2193
rect 14437 1514 14565 4516
rect 16310 4075 16316 4127
rect 16368 4075 16380 4127
rect 16432 4075 16438 4127
rect 14697 3763 15253 3764
rect 14697 3707 14706 3763
rect 14762 3707 14827 3763
rect 14883 3707 14948 3763
rect 15004 3707 15068 3763
rect 15124 3707 15188 3763
rect 15244 3707 15253 3763
rect 14697 3663 15253 3707
rect 14697 3607 14706 3663
rect 14762 3607 14827 3663
rect 14883 3607 14948 3663
rect 15004 3607 15068 3663
rect 15124 3607 15188 3663
rect 15244 3607 15253 3663
rect 14697 3563 15253 3607
rect 14697 3507 14706 3563
rect 14762 3507 14827 3563
rect 14883 3507 14948 3563
rect 15004 3507 15068 3563
rect 15124 3507 15188 3563
rect 15244 3507 15253 3563
rect 14697 3506 15253 3507
rect 16310 3136 16438 4075
rect 14437 1462 14443 1514
rect 14495 1462 14507 1514
rect 14559 1462 14565 1514
rect 15825 3084 15831 3136
rect 15883 3084 15895 3136
rect 15947 3084 15953 3136
rect 16310 3084 16316 3136
rect 16368 3084 16380 3136
rect 16432 3084 16438 3136
rect 15825 1443 15953 3084
rect 16295 2909 16301 2961
rect 16353 2909 16365 2961
rect 16417 2909 16423 2961
tri 16327 2895 16341 2909 ne
rect 16341 2895 16409 2909
tri 16409 2895 16423 2909 nw
tri 16341 2883 16353 2895 ne
rect 16353 2883 16397 2895
tri 16397 2883 16409 2895 nw
tri 16353 2881 16355 2883 ne
rect 15825 1391 15831 1443
rect 15883 1391 15895 1443
rect 15947 1391 15953 1443
tri 14187 1315 14202 1330 sw
rect 10092 1282 10524 1315
tri 10524 1282 10557 1315 sw
rect 13799 1282 14202 1315
tri 14202 1282 14235 1315 sw
rect 10092 1275 10557 1282
tri 10557 1275 10564 1282 sw
rect 13799 1275 14235 1282
tri 14235 1275 14242 1282 sw
rect 10092 1259 10564 1275
tri 10564 1259 10580 1275 sw
rect 13799 1259 14242 1275
tri 14242 1259 14258 1275 sw
rect 10092 1223 13606 1259
tri 13606 1223 13642 1259 sw
rect 13799 1244 14258 1259
tri 14258 1244 14273 1259 sw
rect 13799 1223 15444 1244
tri 15444 1223 15465 1244 sw
rect 10092 1216 13642 1223
tri 13642 1216 13649 1223 sw
rect 13799 1216 15465 1223
tri 15465 1216 15472 1223 sw
rect 10092 1177 13649 1216
tri 13649 1177 13688 1216 sw
rect 13799 1177 15472 1216
tri 15472 1177 15511 1216 sw
rect 10092 1164 13688 1177
tri 13688 1164 13701 1177 sw
rect 13799 1164 15511 1177
tri 15511 1164 15524 1177 sw
rect 10092 1138 13701 1164
tri 13701 1138 13727 1164 sw
rect 13799 1138 15524 1164
tri 15524 1138 15550 1164 sw
rect 10092 1129 13727 1138
tri 13727 1129 13736 1138 sw
rect 7570 1027 7600 1049
tri 7600 1027 7622 1049 nw
rect 6802 1024 7406 1027
tri 7406 1024 7409 1027 nw
tri 7523 1024 7526 1027 se
rect 7526 1024 7588 1027
tri 7522 1023 7523 1024 se
rect 7523 1023 7588 1024
rect 4450 977 4590 988
tri 4590 977 4601 988 sw
tri 6097 977 6108 988 ne
rect 6108 977 6137 988
tri 6137 977 6148 988 sw
rect 2006 881 2015 937
rect 2071 881 2095 937
rect 2151 881 2194 937
tri 2090 855 2116 881 ne
rect 2116 855 2194 881
tri 2116 850 2121 855 ne
tri 1766 808 1778 820 se
rect 1778 808 1914 820
rect 1416 792 1667 801
tri 1753 795 1766 808 se
rect 1766 795 1914 808
tri 1750 792 1753 795 se
rect 1753 792 1914 795
rect 1416 763 1565 792
tri 1565 763 1594 792 nw
tri 1721 763 1750 792 se
rect 1750 763 1914 792
rect 1416 756 1558 763
tri 1558 756 1565 763 nw
tri 1714 756 1721 763 se
rect 1721 756 1914 763
rect 1416 754 1556 756
tri 1556 754 1558 756 nw
tri 1712 754 1714 756 se
rect 1714 754 1914 756
rect 1256 24 1320 47
tri 1320 24 1343 47 nw
rect 1256 -1190 1308 24
tri 1308 12 1320 24 nw
tri 1414 -53 1416 -51 se
rect 1416 -53 1545 754
tri 1545 743 1556 754 nw
tri 1701 743 1712 754 se
rect 1712 743 1914 754
tri 1660 702 1701 743 se
rect 1701 702 1914 743
rect 2121 795 2194 855
rect 3660 850 3688 977
tri 3688 973 3692 977 nw
rect 3778 971 6053 977
rect 3778 945 4237 971
rect 3778 889 3787 945
rect 3843 889 3867 945
rect 3923 919 4237 945
rect 4289 919 5173 971
rect 5225 919 5483 971
rect 5535 964 6053 971
tri 6053 964 6066 977 sw
tri 6108 964 6121 977 ne
rect 6121 964 6148 977
tri 6148 964 6161 977 sw
rect 6337 964 6407 1016
rect 5535 955 6066 964
tri 6066 955 6075 964 sw
tri 6121 955 6130 964 ne
rect 6130 955 6161 964
tri 6161 955 6170 964 sw
rect 5535 953 6075 955
tri 6075 953 6077 955 sw
tri 6130 953 6132 955 ne
rect 6132 953 6170 955
tri 6170 953 6172 955 sw
rect 5535 952 6077 953
tri 6077 952 6078 953 sw
tri 6132 952 6133 953 ne
rect 6133 952 6172 953
tri 6172 952 6173 953 sw
rect 6285 952 6407 964
rect 5535 919 6078 952
rect 3923 915 6078 919
tri 6078 915 6115 952 sw
tri 6133 915 6170 952 ne
rect 6170 915 6173 952
tri 6173 915 6210 952 sw
rect 3923 907 6115 915
rect 3923 889 4237 907
rect 3778 855 4237 889
rect 4289 855 5173 907
rect 5225 855 5483 907
rect 5535 900 6115 907
tri 6115 900 6130 915 sw
tri 6170 900 6185 915 ne
rect 6185 900 6210 915
tri 6210 900 6225 915 sw
rect 6337 901 6407 952
rect 6687 1017 6739 1023
tri 7514 1015 7522 1023 se
rect 7522 1015 7588 1023
tri 7588 1015 7600 1027 nw
rect 10092 1015 13736 1129
tri 7509 1010 7514 1015 se
rect 7514 1010 7582 1015
tri 6739 1009 6740 1010 sw
tri 7508 1009 7509 1010 se
rect 7509 1009 7582 1010
tri 7582 1009 7588 1015 nw
tri 13231 1009 13237 1015 ne
rect 13237 1009 13736 1015
rect 6739 996 6740 1009
tri 6740 996 6753 1009 sw
tri 7495 996 7508 1009 se
rect 7508 996 7569 1009
tri 7569 996 7582 1009 nw
tri 13237 996 13250 1009 ne
rect 13250 996 13736 1009
rect 6739 979 6753 996
tri 6753 979 6770 996 sw
tri 7478 979 7495 996 se
rect 7495 979 7552 996
tri 7552 979 7569 996 nw
tri 13250 979 13267 996 ne
rect 13267 979 13736 996
rect 6739 977 7550 979
tri 7550 977 7552 979 nw
tri 13267 977 13269 979 ne
rect 13269 977 13736 979
rect 6739 973 7546 977
tri 7546 973 7550 977 nw
tri 13269 973 13273 977 ne
rect 13273 973 13736 977
rect 6739 965 7517 973
rect 6687 953 7517 965
tri 6407 901 6430 924 sw
rect 6739 944 7517 953
tri 7517 944 7546 973 nw
tri 7569 944 7598 973 se
rect 7598 963 13154 973
tri 13154 963 13164 973 sw
tri 13273 963 13283 973 ne
rect 7598 944 13164 963
tri 13164 944 13183 963 sw
rect 6739 931 7504 944
tri 7504 931 7517 944 nw
tri 7556 931 7569 944 se
rect 7569 931 13183 944
tri 13183 931 13196 944 sw
rect 6739 927 7500 931
tri 7500 927 7504 931 nw
tri 7552 927 7556 931 se
rect 7556 927 13196 931
rect 6739 908 6751 927
tri 6751 908 6770 927 nw
tri 7533 908 7552 927 se
rect 7552 908 13196 927
tri 13196 908 13219 931 sw
rect 6337 900 6430 901
rect 5535 894 6130 900
tri 6130 894 6136 900 sw
tri 6185 894 6191 900 ne
rect 6191 894 6225 900
tri 6225 894 6231 900 sw
rect 6285 895 6430 900
tri 6430 895 6436 901 sw
rect 6687 895 6739 901
tri 6739 896 6751 908 nw
tri 7521 896 7533 908 se
rect 7533 896 13219 908
tri 7520 895 7521 896 se
rect 7521 895 13219 896
rect 6285 894 6436 895
tri 6436 894 6437 895 sw
tri 7519 894 7520 895 se
rect 7520 894 13219 895
rect 5535 879 6136 894
tri 6136 879 6151 894 sw
tri 6191 879 6206 894 ne
rect 6206 879 6231 894
tri 6231 879 6246 894 sw
rect 6285 893 6437 894
tri 6285 879 6299 893 ne
rect 6299 879 6437 893
tri 6437 879 6452 894 sw
tri 7504 879 7519 894 se
rect 7519 879 13219 894
rect 5535 875 6151 879
tri 6151 875 6155 879 sw
tri 6206 875 6210 879 ne
rect 6210 875 6246 879
tri 6246 875 6250 879 sw
tri 6299 875 6303 879 ne
rect 6303 875 6452 879
rect 5535 866 6155 875
tri 6155 866 6164 875 sw
tri 6210 866 6219 875 ne
rect 6219 866 6250 875
tri 6250 866 6259 875 sw
tri 6303 866 6312 875 ne
rect 6312 866 6452 875
tri 6452 866 6465 879 sw
tri 7491 866 7504 879 se
rect 7504 866 13219 879
rect 5535 855 6164 866
tri 3688 850 3692 854 sw
rect 3660 849 3692 850
tri 3692 849 3693 850 sw
rect 3778 849 6164 855
tri 6164 849 6181 866 sw
tri 6219 849 6236 866 ne
rect 6236 849 6259 866
tri 6259 849 6276 866 sw
tri 6312 849 6329 866 ne
rect 6329 849 6465 866
tri 6465 849 6482 866 sw
tri 7474 849 7491 866 se
rect 7491 849 13219 866
rect 3660 842 3693 849
tri 3693 842 3700 849 sw
tri 5999 842 6006 849 ne
rect 6006 842 6181 849
tri 6181 842 6188 849 sw
tri 6236 842 6243 849 ne
rect 6243 842 6276 849
tri 6276 842 6283 849 sw
tri 6329 842 6336 849 ne
rect 6336 842 6482 849
tri 6482 842 6489 849 sw
tri 7467 842 7474 849 se
rect 7474 847 13219 849
rect 7474 842 7641 847
tri 7641 842 7646 847 nw
tri 13014 842 13019 847 ne
rect 13019 842 13219 847
rect 3660 835 3700 842
tri 3700 835 3707 842 sw
tri 6006 835 6013 842 ne
rect 6013 835 6188 842
tri 6188 835 6195 842 sw
tri 6243 835 6250 842 ne
rect 6250 837 6283 842
tri 6283 837 6288 842 sw
tri 6336 837 6341 842 ne
rect 6341 837 6489 842
tri 6489 837 6494 842 sw
tri 7462 837 7467 842 se
rect 7467 837 7636 842
tri 7636 837 7641 842 nw
tri 13019 837 13024 842 ne
rect 13024 837 13219 842
rect 6250 835 6288 837
tri 6288 835 6290 837 sw
tri 6341 835 6343 837 ne
rect 6343 835 7613 837
rect 3660 820 3707 835
tri 3707 820 3722 835 sw
tri 6013 820 6028 835 ne
rect 6028 820 6195 835
rect 3660 808 5961 820
tri 5961 808 5973 820 sw
tri 6028 808 6040 820 ne
rect 6040 814 6195 820
tri 6195 814 6216 835 sw
tri 6250 814 6271 835 ne
rect 6271 814 6290 835
tri 6290 814 6311 835 sw
tri 6343 814 6364 835 ne
rect 6364 814 7613 835
tri 7613 814 7636 837 nw
tri 13024 814 13047 837 ne
rect 13047 814 13219 837
rect 6040 808 6216 814
tri 6216 808 6222 814 sw
tri 6271 808 6277 814 ne
rect 6277 808 6311 814
tri 6311 808 6317 814 sw
tri 6364 808 6370 814 ne
rect 6370 808 7607 814
tri 7607 808 7613 814 nw
rect 8431 808 12945 814
tri 2194 795 2196 797 sw
rect 3660 795 5973 808
tri 5973 795 5986 808 sw
tri 6040 795 6053 808 ne
rect 6053 795 6222 808
tri 6222 795 6235 808 sw
tri 6277 795 6290 808 ne
rect 6290 795 6317 808
tri 6317 795 6330 808 sw
tri 6370 795 6383 808 ne
rect 6383 795 7572 808
rect 2121 763 2196 795
tri 2196 763 2228 795 sw
rect 3660 792 5986 795
tri 5986 792 5989 795 sw
tri 6053 792 6056 795 ne
rect 6056 792 6235 795
tri 5949 780 5961 792 ne
rect 5961 780 5989 792
tri 5989 780 6001 792 sw
tri 6056 780 6068 792 ne
rect 6068 780 6235 792
tri 5961 763 5978 780 ne
rect 5978 763 6001 780
tri 6001 763 6018 780 sw
tri 6068 763 6085 780 ne
rect 6085 773 6235 780
tri 6235 773 6257 795 sw
tri 6290 773 6312 795 ne
rect 6312 773 6330 795
tri 6330 773 6352 795 sw
tri 6383 773 6405 795 ne
rect 6405 773 7572 795
tri 7572 773 7607 808 nw
rect 6085 763 6257 773
rect 2121 756 5792 763
tri 5792 756 5799 763 sw
tri 5978 756 5985 763 ne
rect 5985 756 6018 763
tri 6018 756 6025 763 sw
tri 6085 756 6092 763 ne
rect 6092 756 6257 763
tri 6257 756 6274 773 sw
tri 6312 756 6329 773 ne
rect 6329 771 6352 773
tri 6352 771 6354 773 sw
tri 6405 771 6407 773 ne
rect 6407 771 7570 773
tri 7570 771 7572 773 nw
tri 7807 771 7809 773 se
rect 7809 771 8239 773
rect 6329 769 6354 771
tri 6354 769 6356 771 sw
tri 6407 769 6409 771 ne
rect 6409 769 7568 771
tri 7568 769 7570 771 nw
tri 7805 769 7807 771 se
rect 7807 769 8239 771
rect 6329 756 6356 769
tri 6356 756 6369 769 sw
tri 7792 756 7805 769 se
rect 7805 756 8239 769
tri 8239 756 8256 773 sw
rect 8483 764 8743 808
rect 8483 756 8509 764
tri 8509 756 8517 764 nw
tri 8709 756 8717 764 ne
rect 8717 756 8743 764
rect 8795 790 12945 808
tri 12945 790 12969 814 sw
tri 13047 801 13060 814 ne
rect 8795 782 12969 790
tri 12969 782 12977 790 sw
rect 8795 764 12977 782
rect 8795 756 8813 764
rect 2121 754 5799 756
tri 5799 754 5801 756 sw
tri 5985 754 5987 756 ne
rect 5987 754 6025 756
tri 6025 754 6027 756 sw
tri 6092 754 6094 756 ne
rect 6094 754 6274 756
tri 6274 754 6276 756 sw
tri 6329 755 6330 756 ne
rect 6330 755 6369 756
tri 6369 755 6370 756 sw
tri 7791 755 7792 756 se
rect 7792 755 8256 756
tri 6330 754 6331 755 ne
rect 6331 754 6370 755
tri 6370 754 6371 755 sw
tri 7790 754 7791 755 se
rect 7791 754 8256 755
tri 8256 754 8258 756 sw
rect 2121 741 5662 754
tri 2121 702 2160 741 ne
rect 2160 702 5662 741
rect 5714 702 5729 754
rect 5781 753 5801 754
tri 5801 753 5802 754 sw
tri 5987 753 5988 754 ne
rect 5988 753 6027 754
tri 6027 753 6028 754 sw
tri 6094 753 6095 754 ne
rect 6095 753 6276 754
rect 5781 748 5802 753
tri 5802 748 5807 753 sw
tri 5988 748 5993 753 ne
rect 5993 748 6028 753
tri 6028 748 6033 753 sw
tri 6095 748 6100 753 ne
rect 6100 748 6276 753
tri 6276 748 6282 754 sw
tri 6331 748 6337 754 ne
rect 6337 748 6371 754
tri 6371 748 6377 754 sw
tri 7784 748 7790 754 se
rect 7790 748 8258 754
tri 8258 748 8264 754 sw
rect 8431 748 8501 756
tri 8501 748 8509 756 nw
tri 8717 748 8725 756 ne
rect 8725 748 8813 756
tri 8813 748 8829 764 nw
tri 12893 748 12909 764 ne
rect 12909 748 12977 764
rect 5781 744 5807 748
tri 5807 744 5811 748 sw
tri 5993 744 5997 748 ne
rect 5997 744 6033 748
tri 6033 744 6037 748 sw
tri 6100 744 6104 748 ne
rect 6104 744 6282 748
tri 6282 744 6286 748 sw
tri 6337 744 6341 748 ne
rect 6341 744 6377 748
tri 6377 744 6381 748 sw
tri 7780 744 7784 748 se
rect 7784 744 8264 748
tri 8264 744 8268 748 sw
rect 8431 744 8497 748
tri 8497 744 8501 748 nw
tri 8725 744 8729 748 ne
rect 8729 744 8801 748
rect 5781 714 5811 744
tri 5811 714 5841 744 sw
tri 5997 740 6001 744 ne
rect 6001 740 6037 744
tri 6037 740 6041 744 sw
tri 6104 740 6108 744 ne
rect 6108 740 6286 744
tri 6001 714 6027 740 ne
rect 6027 714 6041 740
tri 6041 714 6067 740 sw
tri 6108 714 6134 740 ne
rect 6134 714 6286 740
tri 6286 714 6316 744 sw
tri 6341 715 6370 744 ne
rect 6370 720 6381 744
tri 6381 720 6405 744 sw
tri 7756 720 7780 744 se
rect 7780 720 8268 744
rect 6370 715 6405 720
tri 6405 715 6410 720 sw
tri 7751 715 7756 720 se
rect 7756 715 8268 720
tri 6370 714 6371 715 ne
rect 6371 714 6410 715
tri 6410 714 6411 715 sw
tri 7750 714 7751 715 se
rect 7751 714 8268 715
rect 5781 702 5841 714
tri 5841 702 5853 714 sw
tri 6027 702 6039 714 ne
rect 6039 702 6067 714
tri 6067 702 6079 714 sw
tri 6134 702 6146 714 ne
rect 6146 702 6316 714
tri 6316 702 6328 714 sw
tri 6371 703 6382 714 ne
rect 6382 711 6411 714
tri 6411 711 6414 714 sw
tri 7747 711 7750 714 se
rect 7750 711 7758 714
rect 6382 703 7377 711
tri 6382 702 6383 703 ne
rect 6383 702 7377 703
tri 7738 702 7747 711 se
rect 7747 702 7758 711
tri 1632 674 1660 702 se
rect 1660 674 1914 702
tri 5755 674 5783 702 ne
rect 5783 674 5853 702
tri 5853 674 5881 702 sw
tri 6039 700 6041 702 ne
rect 6041 700 6079 702
tri 6079 700 6081 702 sw
tri 6146 700 6148 702 ne
rect 6148 700 6328 702
tri 6041 674 6067 700 ne
rect 6067 674 6081 700
tri 6081 674 6107 700 sw
tri 6148 674 6174 700 ne
rect 6174 674 6328 700
tri 6328 674 6356 702 sw
tri 6383 683 6402 702 ne
rect 6402 683 7377 702
tri 7719 683 7738 702 se
rect 7738 683 7758 702
tri 7710 674 7719 683 se
rect 7719 674 7758 683
tri 1626 668 1632 674 se
rect 1632 668 1914 674
tri 1407 -60 1414 -53 se
rect 1414 -60 1545 -53
tri 1355 -112 1407 -60 se
rect 1407 -112 1545 -60
tri 1350 -117 1355 -112 se
rect 1355 -117 1545 -112
tri 1339 -128 1350 -117 se
rect 1350 -128 1545 -117
rect 1256 -1254 1308 -1242
rect 1256 -1312 1308 -1306
tri 1337 -130 1339 -128 se
rect 1339 -130 1545 -128
rect 1337 -1024 1545 -130
tri 1612 654 1626 668 se
rect 1626 654 1914 668
rect 1612 623 1914 654
rect 1612 616 1907 623
tri 1907 616 1914 623 nw
rect 2004 669 5721 674
rect 1612 604 1895 616
tri 1895 604 1907 616 nw
rect 1612 260 1849 604
tri 1849 558 1895 604 nw
rect 2004 533 2013 669
rect 2149 668 5721 669
rect 2149 616 3177 668
rect 3229 616 3489 668
rect 3541 616 3925 668
rect 3977 662 5721 668
tri 5721 662 5733 674 sw
tri 5783 662 5795 674 ne
rect 5795 662 5881 674
tri 5881 662 5893 674 sw
tri 6067 662 6079 674 ne
rect 6079 662 6107 674
tri 6107 662 6119 674 sw
tri 6174 662 6186 674 ne
rect 6186 662 6356 674
tri 6356 662 6368 674 sw
tri 7698 662 7710 674 se
rect 7710 662 7758 674
rect 7810 702 8268 714
tri 8268 702 8310 744 sw
rect 7810 692 8310 702
tri 8310 692 8320 702 sw
tri 8483 730 8497 744 nw
tri 8729 730 8743 744 ne
rect 7810 686 8320 692
tri 8320 686 8326 692 sw
rect 8431 686 8483 692
rect 8795 736 8801 744
tri 8801 736 8813 748 nw
tri 12909 736 12921 748 ne
rect 12921 736 12977 748
tri 8795 730 8801 736 nw
tri 8902 730 8908 736 se
rect 8908 730 12857 736
tri 12857 730 12863 736 sw
tri 12921 730 12927 736 ne
tri 8870 698 8902 730 se
rect 8902 698 12863 730
tri 12863 698 12895 730 sw
rect 8743 686 8795 692
tri 8858 686 8870 698 se
rect 8870 686 12895 698
rect 7810 674 8326 686
tri 8326 674 8338 686 sw
tri 8846 674 8858 686 se
rect 8858 674 9025 686
rect 7810 671 8338 674
tri 8338 671 8341 674 sw
tri 8843 671 8846 674 se
rect 8846 671 9025 674
tri 9025 671 9040 686 nw
tri 12811 671 12826 686 ne
rect 12826 671 12895 686
rect 7810 662 8341 671
rect 3977 655 5733 662
tri 5733 655 5740 662 sw
tri 5795 655 5802 662 ne
rect 5802 655 5893 662
tri 5893 655 5900 662 sw
tri 6079 660 6081 662 ne
rect 6081 660 6119 662
tri 6119 660 6121 662 sw
tri 6186 660 6188 662 ne
rect 6188 660 6368 662
tri 6081 655 6086 660 ne
rect 6086 655 6121 660
tri 6121 655 6126 660 sw
tri 6188 655 6193 660 ne
rect 6193 655 6368 660
tri 6368 655 6375 662 sw
tri 7691 655 7698 662 se
rect 7698 655 8341 662
tri 8341 655 8357 671 sw
tri 8827 655 8843 671 se
rect 8843 655 8973 671
rect 3977 616 5740 655
rect 2149 604 5740 616
rect 2149 552 3177 604
rect 3229 552 3489 604
rect 3541 552 3925 604
rect 3977 603 5740 604
tri 5740 603 5792 655 sw
tri 5802 603 5854 655 ne
rect 5854 603 5902 655
rect 5954 603 5969 655
rect 6021 603 6027 655
tri 6086 650 6091 655 ne
rect 6091 653 6126 655
tri 6126 653 6128 655 sw
tri 6193 653 6195 655 ne
rect 6195 653 6375 655
tri 6375 653 6377 655 sw
tri 7689 653 7691 655 se
rect 7691 653 8357 655
tri 8357 653 8359 655 sw
tri 8825 653 8827 655 se
rect 8827 653 8973 655
rect 6091 650 6128 653
tri 6128 650 6131 653 sw
tri 6195 650 6198 653 ne
rect 6198 650 7377 653
tri 7686 650 7689 653 se
rect 7689 650 8359 653
tri 6091 647 6094 650 ne
rect 6094 647 6131 650
tri 6131 647 6134 650 sw
tri 6198 647 6201 650 ne
rect 6201 647 7377 650
tri 6094 620 6121 647 ne
rect 6121 620 6134 647
tri 6134 620 6161 647 sw
tri 6201 620 6228 647 ne
rect 6228 620 6563 647
tri 6121 603 6138 620 ne
rect 6138 603 6161 620
tri 6161 603 6178 620 sw
tri 6228 603 6245 620 ne
rect 6245 603 6563 620
rect 3977 595 5792 603
tri 5792 595 5800 603 sw
tri 6138 595 6146 603 ne
rect 6146 595 6178 603
tri 6178 595 6186 603 sw
tri 6245 595 6253 603 ne
rect 6253 595 6563 603
rect 6615 595 7325 647
tri 7646 610 7686 650 se
rect 7686 610 7758 650
rect 3977 583 5525 595
tri 5525 583 5537 595 nw
tri 5636 583 5648 595 ne
rect 5648 583 5800 595
tri 5800 583 5812 595 sw
tri 6146 583 6158 595 ne
rect 6158 583 6186 595
tri 6186 583 6198 595 sw
tri 6253 583 6265 595 ne
rect 6265 583 7377 595
rect 3977 566 5508 583
tri 5508 566 5525 583 nw
tri 5648 566 5665 583 ne
rect 5665 566 5812 583
tri 5812 566 5829 583 sw
tri 6158 580 6161 583 ne
rect 6161 580 6198 583
tri 6198 580 6201 583 sw
tri 6265 580 6268 583 ne
rect 6268 580 6563 583
tri 6161 566 6175 580 ne
rect 6175 566 6201 580
tri 6201 566 6215 580 sw
tri 6268 566 6282 580 ne
rect 6282 566 6563 580
rect 3977 558 5500 566
tri 5500 558 5508 566 nw
tri 5665 564 5667 566 ne
rect 5667 564 6131 566
rect 5567 558 5619 564
rect 3977 552 5488 558
rect 2149 546 5488 552
tri 5488 546 5500 558 nw
rect 2149 533 2158 546
tri 2158 533 2171 546 nw
tri 5554 533 5567 546 se
tri 5536 515 5554 533 se
rect 5554 515 5567 533
rect 2371 463 2377 515
rect 2429 463 2441 515
rect 2493 463 2718 515
rect 2770 463 2782 515
rect 2834 463 2994 515
rect 3046 463 3058 515
rect 3110 463 3342 515
rect 3394 463 3406 515
rect 3458 463 3618 515
rect 3670 463 3682 515
rect 3734 463 3740 515
tri 5531 510 5536 515 se
rect 5536 510 5567 515
tri 5528 507 5531 510 se
rect 5531 507 5567 510
rect 3846 476 4056 482
rect 3898 424 4004 476
rect 4703 455 4709 507
rect 4761 455 4773 507
rect 4825 506 5567 507
tri 5667 546 5685 564 ne
rect 5685 546 6131 564
tri 6131 546 6151 566 sw
tri 6175 546 6195 566 ne
rect 6195 546 6215 566
tri 6215 546 6235 566 sw
tri 6282 546 6302 566 ne
rect 6302 546 6563 566
tri 5685 533 5698 546 ne
rect 5698 540 6151 546
tri 6151 540 6157 546 sw
tri 6195 540 6201 546 ne
rect 6201 540 6235 546
tri 6235 540 6241 546 sw
tri 6302 540 6308 546 ne
rect 6308 540 6563 546
rect 5698 533 6157 540
tri 5698 531 5700 533 ne
rect 5700 531 6157 533
tri 6157 531 6166 540 sw
tri 6201 531 6210 540 ne
rect 6210 531 6241 540
tri 6241 531 6250 540 sw
tri 6308 531 6317 540 ne
rect 6317 531 6563 540
rect 6615 531 7325 583
tri 5700 515 5716 531 ne
rect 5716 522 6166 531
tri 6166 522 6175 531 sw
tri 6210 522 6219 531 ne
rect 6219 525 6250 531
tri 6250 525 6256 531 sw
tri 6317 525 6323 531 ne
rect 6323 525 7377 531
rect 7414 604 7758 610
rect 7466 552 7586 604
rect 7638 598 7758 604
rect 7810 645 8359 650
rect 7810 619 7837 645
tri 7837 619 7863 645 nw
tri 8185 619 8211 645 ne
rect 8211 619 8359 645
tri 8359 619 8393 653 sw
tri 8791 619 8825 653 se
rect 8825 619 8973 653
tri 8973 619 9025 671 nw
tri 12826 652 12845 671 ne
rect 7810 618 7836 619
tri 7836 618 7837 619 nw
tri 8211 618 8212 619 ne
rect 8212 618 8393 619
tri 8393 618 8394 619 sw
tri 8790 618 8791 619 se
rect 8791 618 8972 619
tri 8972 618 8973 619 nw
rect 9055 618 10355 624
rect 7810 610 7828 618
tri 7828 610 7836 618 nw
tri 8212 610 8220 618 ne
rect 8220 610 8394 618
tri 8394 610 8402 618 sw
tri 8782 610 8790 618 se
rect 8790 610 8964 618
tri 8964 610 8972 618 nw
rect 7638 592 7810 598
tri 7810 592 7828 610 nw
tri 8220 592 8238 610 ne
rect 8238 592 8945 610
rect 7638 566 7784 592
tri 7784 566 7810 592 nw
tri 8238 591 8239 592 ne
rect 8239 591 8945 592
tri 8945 591 8964 610 nw
tri 8239 566 8264 591 ne
rect 8264 566 8920 591
tri 8920 566 8945 591 nw
rect 9107 566 9367 618
rect 9419 566 9679 618
rect 9731 566 9991 618
rect 10043 566 10303 618
rect 7638 554 7772 566
tri 7772 554 7784 566 nw
tri 8264 554 8276 566 ne
rect 8276 554 8908 566
tri 8908 554 8920 566 nw
rect 9055 554 10355 566
rect 7638 552 7748 554
rect 7414 540 7748 552
rect 6219 522 6256 525
tri 6256 522 6259 525 sw
rect 5716 515 6175 522
tri 6175 515 6182 522 sw
tri 6219 515 6226 522 ne
rect 6226 515 6259 522
tri 6259 515 6266 522 sw
tri 5716 510 5721 515 ne
rect 5721 510 6182 515
rect 4825 494 5619 506
rect 4825 455 5567 494
tri 5548 442 5561 455 ne
rect 5561 442 5567 455
tri 5721 490 5741 510 ne
rect 5741 500 6182 510
tri 6182 500 6197 515 sw
tri 6226 500 6241 515 ne
rect 6241 500 6266 515
tri 6266 500 6281 515 sw
rect 5741 490 6197 500
tri 6197 490 6207 500 sw
tri 5741 463 5768 490 ne
rect 5768 463 6085 490
tri 5768 459 5772 463 ne
rect 5772 459 6085 463
tri 5561 440 5563 442 ne
rect 5563 440 5619 442
tri 4056 438 4058 440 sw
tri 5563 438 5565 440 ne
rect 5565 438 5619 440
tri 5772 438 5793 459 ne
rect 5793 438 6085 459
rect 6137 438 6149 490
rect 6201 438 6207 490
tri 6241 488 6253 500 ne
rect 6253 495 6281 500
tri 6281 495 6286 500 sw
rect 6253 488 7377 495
tri 6253 487 6254 488 ne
rect 6254 487 7377 488
tri 6254 478 6263 487 ne
rect 6263 478 7377 487
rect 7466 488 7586 540
rect 7638 530 7748 540
tri 7748 530 7772 554 nw
tri 8276 536 8294 554 ne
rect 8294 536 8876 554
rect 7929 530 7981 536
rect 7638 525 7743 530
tri 7743 525 7748 530 nw
rect 7638 522 7740 525
tri 7740 522 7743 525 nw
rect 7638 515 7733 522
tri 7733 515 7740 522 nw
rect 7638 488 7700 515
rect 7414 482 7700 488
tri 7700 482 7733 515 nw
tri 6263 467 6274 478 ne
rect 6274 467 7377 478
tri 8294 525 8305 536 ne
rect 8305 525 8876 536
tri 8305 522 8308 525 ne
rect 8308 522 8876 525
tri 8876 522 8908 554 nw
tri 8308 515 8315 522 ne
rect 8315 515 8869 522
tri 8869 515 8876 522 nw
tri 8315 502 8328 515 ne
rect 8328 502 8856 515
tri 8856 502 8869 515 nw
rect 9107 502 9367 554
rect 9419 502 9679 554
rect 9731 502 9991 554
rect 10043 502 10303 554
tri 12752 516 12758 522 se
rect 12758 516 12810 522
tri 12751 515 12752 516 se
rect 12752 515 12758 516
tri 8328 482 8348 502 ne
rect 8348 482 8836 502
tri 8836 482 8856 502 nw
rect 9055 496 10355 502
tri 12732 496 12751 515 se
rect 12751 496 12758 515
tri 12718 482 12732 496 se
rect 12732 482 12758 496
rect 7929 466 7981 478
tri 7927 438 7929 440 se
rect 4056 436 4058 438
tri 4058 436 4060 438 sw
tri 5565 436 5567 438 ne
rect 5567 436 5619 438
tri 7925 436 7927 438 se
rect 7927 436 7929 438
rect 4056 424 4060 436
rect 3846 414 4060 424
tri 4060 414 4082 436 sw
tri 7903 414 7925 436 se
rect 7925 414 7929 436
tri 12700 464 12718 482 se
rect 12718 464 12758 482
tri 12699 463 12700 464 se
rect 12700 463 12810 464
tri 12695 459 12699 463 se
rect 12699 459 12810 463
tri 12688 452 12695 459 se
rect 12695 452 12810 459
rect 3846 412 4082 414
rect 3254 394 3306 400
rect 3898 360 4004 412
rect 4056 408 4082 412
tri 4082 408 4088 414 sw
tri 7897 408 7903 414 se
rect 7903 408 7981 414
rect 4056 406 4088 408
tri 4088 406 4090 408 sw
tri 7895 406 7897 408 se
rect 7897 406 7979 408
tri 7979 406 7981 408 nw
rect 8010 446 8062 452
tri 12684 448 12688 452 se
rect 12688 448 12810 452
rect 4056 394 7967 406
tri 7967 394 7979 406 nw
tri 12669 433 12684 448 se
rect 12684 433 12810 448
tri 12662 426 12669 433 se
rect 12669 426 12758 433
rect 4056 382 7955 394
tri 7955 382 7967 394 nw
rect 8010 382 8062 394
rect 4056 360 7927 382
tri 3306 354 3310 358 sw
rect 3846 354 7927 360
tri 7927 354 7955 382 nw
rect 3306 349 3310 354
tri 3310 349 3315 354 sw
rect 3306 342 3315 349
rect 3254 330 3315 342
tri 3315 330 3334 349 sw
tri 7991 330 8010 349 se
rect 2630 312 2682 318
tri 1849 260 1889 300 sw
rect 3306 324 3334 330
tri 3334 324 3340 330 sw
tri 7985 324 7991 330 se
rect 7991 324 8062 330
rect 3306 318 8062 324
rect 9834 420 9886 426
rect 9834 350 9886 368
rect 3306 312 8056 318
tri 8056 312 8062 318 nw
rect 8090 312 8142 318
rect 3306 292 8036 312
tri 8036 292 8056 312 nw
rect 3306 278 8016 292
tri 2682 272 2686 276 sw
rect 3254 272 8016 278
tri 8016 272 8036 292 nw
tri 8086 272 8090 276 se
rect 2682 260 2686 272
tri 2686 260 2698 272 sw
tri 8074 260 8086 272 se
rect 8086 260 8090 272
rect 9834 292 9886 298
rect 9920 420 12758 426
rect 9920 368 10146 420
rect 10198 368 10458 420
rect 10510 381 12758 420
rect 10510 368 12810 381
rect 9920 350 12810 368
rect 9920 298 10146 350
rect 10198 298 10458 350
rect 10510 298 12758 350
rect 9920 292 12810 298
rect 1612 248 1889 260
tri 1889 248 1901 260 sw
rect 1612 231 1901 248
tri 1901 231 1918 248 sw
rect 1612 212 1918 231
rect 1612 160 1866 212
rect 1612 144 1918 160
rect 1612 92 1866 144
rect 2063 240 2119 249
rect 2630 248 2698 260
tri 2698 248 2710 260 sw
tri 8062 248 8074 260 se
rect 8074 248 8142 260
rect 2682 242 2710 248
tri 2710 242 2716 248 sw
tri 8056 242 8062 248 se
rect 8062 242 8090 248
rect 2682 196 8090 242
rect 2630 190 8142 196
rect 2063 169 2065 184
rect 2117 169 2119 184
rect 2063 160 2119 169
rect 2063 95 2119 104
rect 2421 154 12737 160
rect 2421 102 2553 154
rect 2605 102 2865 154
rect 2917 102 3769 154
rect 3821 102 4081 154
rect 4133 102 4393 154
rect 4445 102 4549 154
rect 4601 102 4861 154
rect 4913 102 5017 154
rect 5069 102 5329 154
rect 5381 102 5814 154
rect 5866 102 6407 154
rect 6459 102 6843 154
rect 6895 102 7142 154
rect 7194 102 7208 154
rect 7260 102 8171 154
rect 8223 102 8275 154
rect 8327 102 8587 154
rect 8639 102 8899 154
rect 8951 102 9211 154
rect 9263 102 9523 154
rect 9575 151 12737 154
rect 9575 102 10595 151
rect 2421 99 10595 102
rect 10647 99 10728 151
rect 10780 99 11184 151
rect 11236 99 11640 151
rect 11692 99 12097 151
rect 12149 99 12438 151
rect 12490 99 12520 151
rect 12572 99 12602 151
rect 12654 99 12684 151
rect 12736 99 12737 151
rect 1612 76 1918 92
rect 1612 24 1866 76
rect 1612 8 1918 24
rect 1612 -44 1866 8
rect 1612 -60 1918 -44
rect 2421 89 12737 99
rect 12845 129 12895 671
rect 12927 155 12977 736
rect 13060 228 13219 814
rect 13283 842 13736 973
rect 13283 790 13289 842
rect 13341 790 13354 842
rect 13406 790 13419 842
rect 13471 790 13484 842
rect 13536 790 13549 842
rect 13601 790 13614 842
rect 13666 790 13678 842
rect 13730 790 13736 842
rect 13283 369 13736 790
rect 13283 317 13289 369
rect 13341 317 13354 369
rect 13406 317 13419 369
rect 13471 317 13484 369
rect 13536 317 13549 369
rect 13601 317 13614 369
rect 13666 317 13678 369
rect 13730 317 13736 369
rect 13799 1125 15550 1138
tri 15550 1125 15563 1138 sw
rect 13799 1081 15563 1125
tri 15563 1081 15607 1125 sw
rect 13799 1079 15607 1081
rect 13799 1027 13805 1079
rect 13857 1027 13873 1079
rect 13925 1027 13941 1079
rect 13993 1027 14008 1079
rect 14060 1027 14075 1079
rect 14127 1027 14142 1079
rect 14194 1027 14209 1079
rect 14261 1027 14276 1079
rect 14328 1027 14343 1079
rect 14395 1027 14410 1079
rect 14462 1027 14477 1079
rect 14529 1027 14544 1079
rect 14596 1027 14611 1079
rect 14663 1027 14678 1079
rect 14730 1027 14745 1079
rect 14797 1027 14812 1079
rect 14864 1027 14879 1079
rect 14931 1027 14946 1079
rect 14998 1067 15607 1079
tri 15607 1067 15621 1081 sw
rect 14998 1061 15976 1067
rect 14998 1027 15452 1061
rect 13799 1009 15452 1027
rect 15504 1009 15924 1061
rect 13799 996 15976 1009
rect 13799 944 15452 996
rect 15504 944 15924 996
rect 13799 931 15976 944
rect 13799 920 15452 931
rect 13799 879 14412 920
tri 14412 879 14453 920 nw
tri 15198 879 15239 920 ne
rect 15239 879 15452 920
rect 15504 879 15924 931
rect 13799 866 14399 879
tri 14399 866 14412 879 nw
tri 15239 866 15252 879 ne
rect 15252 866 15976 879
rect 13799 845 14378 866
tri 14378 845 14399 866 nw
tri 15252 845 15273 866 ne
rect 15273 845 15452 866
rect 13799 842 14375 845
tri 14375 842 14378 845 nw
rect 14478 842 15028 845
rect 13799 606 14357 842
tri 14357 824 14375 842 nw
rect 13799 554 13805 606
rect 13857 554 13876 606
rect 13928 554 13947 606
rect 13999 554 14018 606
rect 14070 554 14089 606
rect 14141 554 14159 606
rect 14211 554 14229 606
rect 14281 554 14299 606
rect 14351 554 14357 606
tri 13219 228 13247 256 sw
rect 13799 228 14357 554
rect 14478 790 14484 842
rect 14536 790 14555 842
rect 14607 790 14626 842
rect 14678 790 14697 842
rect 14749 790 14768 842
rect 14820 790 14838 842
rect 14890 790 14908 842
rect 14960 814 15028 842
tri 15028 814 15059 845 sw
tri 15273 814 15304 845 ne
rect 15304 814 15452 845
rect 15504 814 15924 866
rect 14960 800 15059 814
tri 15059 800 15073 814 sw
tri 15304 800 15318 814 ne
rect 15318 800 15976 814
rect 14960 790 15073 800
rect 14478 748 15073 790
tri 15073 748 15125 800 sw
tri 15318 748 15370 800 ne
rect 15370 748 15452 800
rect 15504 748 15924 800
rect 14478 742 15125 748
tri 15125 742 15131 748 sw
tri 15370 742 15376 748 ne
rect 15376 742 15976 748
rect 14478 687 15131 742
tri 15131 687 15186 742 sw
rect 14478 671 16215 687
rect 14478 619 15214 671
rect 15266 619 15687 671
rect 15739 619 16159 671
rect 16211 619 16215 671
rect 14478 597 16215 619
rect 14478 545 15214 597
rect 15266 545 15687 597
rect 15739 545 16159 597
rect 16211 545 16215 597
rect 14478 523 16215 545
rect 14478 471 15214 523
rect 15266 471 15687 523
rect 15739 471 16159 523
rect 16211 471 16215 523
rect 14478 448 16215 471
rect 14478 396 15214 448
rect 15266 396 15687 448
rect 15739 396 16159 448
rect 16211 396 16215 448
rect 14478 373 16215 396
rect 14478 369 15214 373
rect 14478 317 14484 369
rect 14536 317 14555 369
rect 14607 317 14626 369
rect 14678 317 14697 369
rect 14749 317 14768 369
rect 14820 317 14838 369
rect 14890 317 14908 369
rect 14960 321 15214 369
rect 15266 321 15687 373
rect 15739 321 16159 373
rect 16211 321 16215 373
tri 16335 326 16355 346 se
rect 16355 328 16395 2883
tri 16395 2881 16397 2883 nw
rect 16630 2692 16666 4553
rect 16698 2895 16734 4568
rect 16766 2982 16802 4605
rect 17051 4590 17057 4642
rect 17109 4590 17121 4642
rect 17173 4590 17254 4642
rect 17523 4620 17529 4672
rect 17581 4620 17593 4672
rect 17645 4620 17651 4672
rect 18720 4653 18848 4827
tri 18848 4826 18849 4827 nw
rect 19753 4788 20024 4827
rect 19753 4736 19755 4788
rect 19807 4736 19819 4788
rect 19871 4736 19883 4788
rect 19935 4736 19947 4788
rect 19999 4736 20024 4788
rect 19753 4735 20024 4736
rect 19753 4730 20085 4735
tri 20085 4730 20090 4735 nw
rect 19753 4693 20048 4730
tri 20048 4693 20085 4730 nw
rect 19753 4692 20047 4693
tri 20047 4692 20048 4693 nw
rect 19753 4686 20024 4692
tri 17523 4611 17532 4620 ne
rect 17532 4611 17603 4620
tri 17603 4611 17612 4620 nw
tri 17160 4573 17177 4590 ne
rect 17177 4573 17254 4590
tri 17177 4569 17181 4573 ne
rect 17181 4569 17254 4573
tri 17181 4568 17182 4569 ne
rect 17182 4568 17254 4569
tri 17182 4556 17194 4568 ne
rect 17194 4556 17254 4568
tri 17194 4548 17202 4556 ne
rect 16837 4222 16925 4278
rect 16837 4121 16889 4222
tri 16889 4186 16925 4222 nw
rect 16990 4077 16996 4129
rect 17048 4077 17062 4129
rect 17114 4077 17120 4129
rect 16837 4055 16889 4069
rect 16837 3997 16889 4003
tri 16996 3248 17000 3252 se
rect 17000 3248 17052 4077
tri 16983 3235 16996 3248 se
rect 16996 3235 17052 3248
tri 16970 3222 16983 3235 se
rect 16983 3222 17052 3235
tri 16966 3218 16970 3222 se
rect 16970 3218 17052 3222
rect 16924 3166 16930 3218
rect 16982 3166 16994 3218
rect 17046 3166 17052 3218
tri 16924 3157 16933 3166 ne
rect 16933 3154 17040 3166
tri 17040 3154 17052 3166 nw
rect 17107 3932 17159 3938
rect 17107 3866 17159 3880
rect 16933 3128 17014 3154
tri 17014 3128 17040 3154 nw
rect 16933 3123 17009 3128
tri 17009 3123 17014 3128 nw
tri 16802 2982 16819 2999 sw
rect 16766 2972 16819 2982
tri 16819 2972 16829 2982 sw
rect 16766 2920 16772 2972
rect 16824 2920 16836 2972
rect 16888 2920 16894 2972
tri 16734 2895 16748 2909 sw
rect 16698 2883 16748 2895
tri 16748 2883 16760 2895 sw
rect 16698 2875 16764 2883
tri 16698 2831 16742 2875 ne
rect 16742 2831 16764 2875
rect 16816 2831 16828 2883
rect 16880 2831 16886 2883
rect 16933 2737 16985 3123
tri 16985 3099 17009 3123 nw
tri 17103 3084 17107 3088 se
rect 17107 3084 17159 3814
tri 17090 3071 17103 3084 se
rect 17103 3071 17159 3084
tri 17083 3064 17090 3071 se
rect 17090 3064 17159 3071
tri 17078 3059 17083 3064 se
rect 17083 3059 17159 3064
tri 17073 3054 17078 3059 se
rect 17078 3054 17159 3059
rect 17031 3002 17037 3054
rect 17089 3002 17101 3054
rect 17153 3002 17159 3054
tri 17167 2789 17202 2824 se
rect 17202 2789 17254 4556
rect 17532 4601 17593 4611
tri 17593 4601 17603 4611 nw
rect 18720 4601 18726 4653
rect 18778 4601 18790 4653
rect 18842 4601 18848 4653
tri 16985 2737 16993 2745 sw
rect 17126 2737 17132 2789
rect 17184 2737 17196 2789
rect 17248 2737 17254 2789
rect 17292 3330 17298 3382
rect 17350 3330 17362 3382
rect 17414 3330 17420 3382
rect 17292 3222 17420 3330
rect 17292 3170 17298 3222
rect 17350 3170 17362 3222
rect 17414 3170 17420 3222
rect 16933 2730 16993 2737
tri 16993 2730 17000 2737 sw
rect 16933 2723 17000 2730
tri 16933 2717 16939 2723 ne
rect 16939 2717 17000 2723
tri 17000 2717 17013 2730 sw
tri 16666 2692 16691 2717 sw
tri 16939 2692 16964 2717 ne
rect 16964 2692 17013 2717
tri 17013 2692 17038 2717 sw
rect 16630 2687 16773 2692
tri 16630 2640 16677 2687 ne
rect 16677 2640 16773 2687
rect 16825 2640 16837 2692
rect 16889 2640 16895 2692
tri 16964 2656 17000 2692 ne
rect 17000 2656 17038 2692
tri 17038 2656 17074 2692 sw
tri 17000 2640 17016 2656 ne
rect 17016 2640 17074 2656
tri 17074 2640 17090 2656 sw
tri 17016 2612 17044 2640 ne
rect 17044 2612 17090 2640
tri 17090 2612 17118 2640 sw
rect 17292 2612 17420 3170
tri 17044 2582 17074 2612 ne
rect 17074 2582 17118 2612
tri 17118 2582 17148 2612 sw
tri 17074 2560 17096 2582 ne
rect 17096 2560 17148 2582
tri 17148 2560 17170 2582 sw
rect 17292 2560 17298 2612
rect 17350 2560 17362 2612
rect 17414 2560 17420 2612
rect 17451 3123 17503 3129
rect 17451 3059 17503 3071
tri 17096 2508 17148 2560 ne
rect 17148 2508 17170 2560
tri 17170 2508 17222 2560 sw
tri 17148 2486 17170 2508 ne
rect 17170 2497 17222 2508
tri 17136 2332 17170 2366 se
rect 16535 1760 16739 1766
rect 16587 1708 16611 1760
rect 16663 1708 16687 1760
rect 16535 1681 16739 1708
rect 16587 1629 16611 1681
rect 16663 1629 16687 1681
rect 16535 1602 16739 1629
rect 16587 1550 16611 1602
rect 16663 1550 16687 1602
rect 16535 1474 16739 1550
tri 17444 1474 17451 1481 se
rect 17451 1474 17503 3007
rect 17532 2185 17584 4601
tri 17584 4592 17593 4601 nw
rect 18947 4600 19004 4656
rect 19060 4600 19084 4656
rect 19140 4600 19149 4656
rect 19753 4634 19964 4686
rect 20016 4634 20024 4686
tri 20024 4669 20047 4692 nw
rect 19753 4621 20024 4634
rect 18405 4474 18414 4530
rect 18470 4474 18494 4530
rect 18550 4474 18559 4530
rect 18405 4473 18553 4474
tri 18553 4473 18554 4474 nw
tri 18405 4439 18439 4473 ne
rect 18439 4439 18519 4473
tri 18519 4439 18553 4473 nw
tri 18439 4432 18446 4439 ne
rect 17675 4062 17727 4069
rect 17675 3998 17727 4010
rect 17675 3222 17727 3946
rect 17759 4030 17765 4082
rect 17817 4030 17839 4082
rect 17891 4030 17912 4082
rect 17964 4030 17970 4082
rect 17759 3373 17970 4030
rect 17759 3300 17897 3373
tri 17897 3300 17970 3373 nw
rect 17759 3248 17765 3300
rect 17817 3248 17839 3300
rect 17891 3248 17897 3300
tri 17727 3222 17741 3236 sw
rect 17675 3221 17741 3222
tri 17675 3213 17683 3221 ne
rect 17683 3213 17741 3221
tri 17741 3213 17750 3222 sw
tri 17683 3173 17723 3213 ne
rect 17723 3173 17801 3213
tri 17801 3173 17841 3213 sw
tri 17723 3170 17726 3173 ne
rect 17726 3170 17841 3173
tri 17726 3169 17727 3170 ne
rect 17727 3169 17841 3170
tri 17727 3165 17731 3169 ne
rect 17731 3165 17841 3169
tri 17770 3154 17781 3165 ne
rect 17781 3154 17841 3165
tri 17781 3146 17789 3154 ne
rect 17613 3128 17665 3134
rect 17613 3064 17665 3076
rect 17613 1545 17665 3012
rect 17789 2982 17841 3154
rect 18104 3154 18156 3160
rect 18104 3088 18156 3102
tri 17841 2982 17883 3024 sw
rect 17789 2930 17795 2982
rect 17847 2930 17859 2982
rect 17911 2930 17917 2982
tri 18086 2895 18104 2913 se
rect 18104 2895 18156 3036
rect 18273 3154 18325 3160
rect 18273 3088 18325 3102
tri 18156 2895 18171 2910 sw
tri 18074 2883 18086 2895 se
rect 18086 2883 18171 2895
tri 18171 2883 18183 2895 sw
rect 18060 2831 18066 2883
rect 18118 2831 18132 2883
rect 18184 2831 18190 2883
tri 18270 2739 18273 2742 se
rect 18273 2739 18325 3036
rect 18446 2739 18512 4439
tri 18512 4432 18519 4439 nw
rect 18582 3961 18588 4013
rect 18640 3961 18652 4013
rect 18704 3961 18710 4013
tri 18564 3526 18582 3544 se
rect 18582 3526 18710 3961
rect 18760 3836 18766 3888
rect 18818 3836 18833 3888
rect 18885 3836 18891 3888
tri 18760 3835 18761 3836 ne
tri 18560 3522 18564 3526 se
rect 18564 3522 18710 3526
tri 18710 3522 18714 3526 sw
rect 18560 3466 18569 3522
rect 18625 3466 18649 3522
rect 18705 3466 18714 3522
rect 18560 3464 18714 3466
rect 18560 3460 18710 3464
tri 18710 3460 18714 3464 nw
rect 18761 3464 18891 3836
rect 18761 3412 18767 3464
rect 18819 3412 18833 3464
rect 18885 3412 18891 3464
rect 18583 3154 18635 3160
rect 18583 3088 18635 3102
rect 18583 3030 18635 3036
tri 18583 3025 18588 3030 ne
rect 18588 3025 18630 3030
tri 18630 3025 18635 3030 nw
rect 18733 3154 18785 3160
rect 18733 3088 18785 3102
rect 18733 3030 18785 3036
rect 18733 3027 18782 3030
tri 18782 3027 18785 3030 nw
rect 18821 3153 18873 3159
rect 18821 3087 18873 3101
rect 18821 3029 18873 3035
rect 18821 3027 18871 3029
tri 18871 3027 18873 3029 nw
tri 18733 3025 18735 3027 ne
rect 18735 3025 18779 3027
tri 18238 2707 18270 2739 se
rect 18270 2707 18325 2739
tri 18223 2692 18238 2707 se
rect 18238 2692 18325 2707
tri 18325 2692 18340 2707 sw
rect 18212 2640 18218 2692
rect 18270 2640 18282 2692
rect 18334 2640 18340 2692
rect 18395 2687 18401 2739
rect 18453 2687 18492 2739
rect 18544 2687 18550 2739
tri 18585 2640 18588 2643 se
rect 18588 2640 18627 3025
tri 18627 3022 18630 3025 nw
tri 18735 3024 18736 3025 ne
rect 18736 3024 18779 3025
tri 18779 3024 18782 3027 nw
rect 18821 3024 18868 3027
tri 18868 3024 18871 3027 nw
rect 18736 3022 18777 3024
tri 18777 3022 18779 3024 nw
rect 18821 3022 18866 3024
tri 18866 3022 18868 3024 nw
tri 18556 2611 18585 2640 se
rect 18585 2611 18627 2640
tri 18110 2587 18134 2611 se
rect 18134 2590 18627 2611
rect 18134 2587 18624 2590
tri 18624 2587 18627 2590 nw
rect 18110 2560 18597 2587
tri 18597 2560 18624 2587 nw
tri 18735 2560 18736 2561 se
rect 18736 2560 18775 3022
tri 18775 3020 18777 3022 nw
rect 18821 3020 18864 3022
tri 18864 3020 18866 3022 nw
tri 18053 2116 18110 2173 se
rect 18110 2155 18149 2560
tri 18149 2529 18180 2560 nw
tri 18704 2529 18735 2560 se
rect 18735 2529 18775 2560
rect 18110 2126 18120 2155
tri 18120 2126 18149 2155 nw
tri 18184 2505 18208 2529 se
rect 18208 2508 18775 2529
rect 18208 2505 18772 2508
tri 18772 2505 18775 2508 nw
rect 18184 2478 18745 2505
tri 18745 2478 18772 2505 nw
tri 18110 2116 18120 2126 nw
tri 18174 2116 18184 2126 se
rect 18184 2116 18223 2478
tri 18223 2451 18250 2478 nw
tri 18797 2451 18821 2475 se
rect 18821 2451 18860 3020
tri 18860 3016 18864 3020 nw
tri 18789 2443 18797 2451 se
rect 18797 2443 18860 2451
tri 18022 2085 18053 2116 se
rect 18053 2085 18079 2116
tri 18079 2085 18110 2116 nw
tri 18143 2085 18174 2116 se
rect 18174 2108 18223 2116
rect 18174 2085 18190 2108
rect 18022 2075 18069 2085
tri 18069 2075 18079 2085 nw
tri 18133 2075 18143 2085 se
rect 18143 2075 18190 2085
tri 18190 2075 18223 2108 nw
tri 18261 2411 18293 2443 se
rect 18293 2422 18860 2443
rect 18293 2411 18849 2422
tri 18849 2411 18860 2422 nw
rect 18947 2895 19011 4600
rect 19753 4569 19964 4621
rect 20016 4569 20024 4621
rect 19753 4556 20024 4569
rect 19753 4504 19964 4556
rect 20016 4504 20024 4556
rect 19753 4491 20024 4504
rect 19753 4439 19964 4491
rect 20016 4439 20024 4491
rect 19753 4426 20024 4439
rect 19753 4374 19964 4426
rect 20016 4374 20024 4426
rect 19753 4361 20024 4374
rect 19753 4309 19964 4361
rect 20016 4309 20024 4361
rect 19753 4296 20024 4309
rect 19753 4244 19964 4296
rect 20016 4244 20024 4296
rect 19753 4231 20024 4244
rect 19753 4179 19964 4231
rect 20016 4179 20024 4231
rect 19753 4166 20024 4179
rect 19753 4114 19964 4166
rect 20016 4114 20024 4166
rect 19259 4098 19311 4104
rect 19259 4034 19311 4046
rect 19259 3976 19311 3982
rect 19753 4100 20024 4114
rect 19753 4048 19964 4100
rect 20016 4048 20024 4100
rect 19753 4034 20024 4048
rect 19753 3982 19964 4034
rect 20016 3982 20024 4034
rect 19753 3968 20024 3982
rect 19753 3916 19964 3968
rect 20016 3916 20024 3968
rect 19753 3902 20024 3916
rect 19753 3850 19964 3902
rect 20016 3850 20024 3902
rect 19753 3836 20024 3850
rect 19753 3784 19964 3836
rect 20016 3784 20024 3836
rect 19082 3719 19088 3771
rect 19140 3719 19165 3771
rect 19217 3719 19242 3771
rect 19294 3719 19300 3771
rect 19082 3701 19300 3719
rect 19082 3649 19088 3701
rect 19140 3649 19165 3701
rect 19217 3649 19242 3701
rect 19294 3649 19300 3701
rect 19082 3631 19300 3649
rect 19082 3579 19088 3631
rect 19140 3579 19165 3631
rect 19217 3579 19242 3631
rect 19294 3579 19300 3631
rect 19753 3770 20024 3784
rect 19753 3718 19964 3770
rect 20016 3718 20024 3770
rect 19753 3704 20024 3718
rect 19753 3652 19964 3704
rect 20016 3652 20024 3704
rect 19753 3638 20024 3652
rect 19753 3586 19964 3638
rect 20016 3586 20024 3638
rect 19753 3572 20024 3586
rect 19753 3520 19964 3572
rect 20016 3520 20024 3572
rect 19753 3506 20024 3520
tri 19729 3454 19753 3478 se
rect 19753 3454 19964 3506
rect 20016 3454 20024 3506
tri 19715 3440 19729 3454 se
rect 19729 3440 20024 3454
tri 19663 3388 19715 3440 se
rect 19715 3388 19964 3440
rect 20016 3388 20024 3440
tri 19657 3382 19663 3388 se
rect 19663 3382 20024 3388
tri 19655 3380 19657 3382 se
rect 19657 3380 20024 3382
rect 19378 3227 20024 3380
tri 19011 2895 19059 2943 sw
rect 18947 2843 18953 2895
rect 19005 2843 19044 2895
rect 19096 2843 19102 2895
rect 18261 2392 18830 2411
tri 18830 2392 18849 2411 nw
tri 17665 1545 17695 1575 sw
rect 17613 1544 17695 1545
tri 17695 1544 17696 1545 sw
rect 17613 1537 17696 1544
tri 17696 1537 17703 1544 sw
rect 17613 1485 17619 1537
rect 17671 1485 17683 1537
rect 17735 1485 17741 1537
tri 17413 1443 17444 1474 se
rect 17444 1443 17503 1474
rect 17375 1391 17381 1443
rect 17433 1391 17445 1443
rect 17497 1391 17503 1443
tri 17985 1282 18022 1319 se
rect 18022 1282 18061 2075
tri 18061 2067 18069 2075 nw
tri 18127 2069 18133 2075 se
rect 18133 2069 18184 2075
tri 18184 2069 18190 2075 nw
tri 18125 2067 18127 2069 se
rect 18127 2067 18153 2069
tri 17984 1281 17985 1282 se
rect 17985 1281 18061 1282
tri 17978 1275 17984 1281 se
rect 17984 1275 18061 1281
rect 17933 1223 17939 1275
rect 17991 1223 18003 1275
rect 18055 1223 18061 1275
tri 18096 2038 18125 2067 se
rect 18125 2038 18153 2067
tri 18153 2038 18184 2069 nw
tri 18259 2038 18261 2040 se
rect 18261 2038 18300 2392
tri 18300 2359 18333 2392 nw
tri 18693 2246 18727 2280 ne
tri 18609 2154 18643 2188 ne
tri 18521 2075 18543 2097 ne
rect 18543 2075 18555 2097
tri 18543 2069 18549 2075 ne
rect 18549 2069 18555 2075
tri 18549 2063 18555 2069 ne
rect 18096 2023 18138 2038
tri 18138 2023 18153 2038 nw
tri 18244 2023 18259 2038 se
rect 18259 2023 18300 2038
tri 18065 1177 18096 1208 se
rect 18096 1177 18135 2023
tri 18135 2020 18138 2023 nw
tri 18241 2020 18244 2023 se
rect 18244 2022 18300 2023
rect 18244 2020 18261 2022
tri 18204 1983 18241 2020 se
rect 18241 1983 18261 2020
tri 18261 1983 18300 2022 nw
rect 18007 1125 18013 1177
rect 18065 1125 18077 1177
rect 18129 1125 18135 1177
tri 18173 1952 18204 1983 se
rect 18204 1952 18230 1983
tri 18230 1952 18261 1983 nw
tri 18145 1081 18173 1109 se
rect 18173 1081 18212 1952
tri 18212 1934 18230 1952 nw
tri 18894 1860 18947 1913 se
rect 18947 1860 19018 2843
tri 19018 2801 19060 2843 nw
rect 25328 2075 25337 2077
rect 25393 2075 25417 2077
rect 25328 2023 25334 2075
rect 25393 2023 25398 2075
rect 25328 2021 25337 2023
rect 25393 2021 25417 2023
rect 25473 2021 25482 2077
rect 18864 1804 18873 1860
rect 18929 1804 18953 1860
rect 19009 1804 19018 1860
rect 18869 1703 18875 1755
rect 18927 1703 18941 1755
rect 18993 1703 19007 1755
rect 19059 1703 19073 1755
rect 19125 1703 19139 1755
rect 19191 1703 20436 1755
rect 18869 1655 20436 1703
rect 18869 1603 18875 1655
rect 18927 1603 18941 1655
rect 18993 1603 19007 1655
rect 19059 1603 19073 1655
rect 19125 1603 19139 1655
rect 19191 1603 20436 1655
tri 20166 1575 20194 1603 ne
rect 20194 1575 20436 1603
tri 20436 1575 20616 1755 sw
rect 23947 1575 24004 1577
tri 24004 1575 24006 1577 sw
tri 20194 1549 20220 1575 ne
rect 20220 1549 20616 1575
tri 20616 1549 20642 1575 sw
rect 23947 1568 24006 1575
tri 20220 1545 20224 1549 ne
rect 20224 1545 20884 1549
tri 20224 1544 20225 1545 ne
rect 20225 1544 20884 1545
tri 20225 1537 20232 1544 ne
rect 20232 1537 20519 1544
tri 20232 1492 20277 1537 ne
rect 20277 1492 20519 1537
rect 20571 1492 20592 1544
rect 20644 1492 20665 1544
rect 20717 1492 20738 1544
rect 20790 1492 20810 1544
rect 20862 1492 20884 1544
tri 20277 1490 20279 1492 ne
rect 20279 1490 20884 1492
tri 20279 1485 20284 1490 ne
rect 20284 1485 20884 1490
tri 20284 1474 20295 1485 ne
rect 20295 1474 20884 1485
tri 20295 1422 20347 1474 ne
rect 20347 1422 20519 1474
rect 20571 1422 20592 1474
rect 20644 1422 20665 1474
rect 20717 1422 20738 1474
rect 20790 1422 20810 1474
rect 20862 1422 20884 1474
rect 24003 1549 24006 1568
tri 24006 1549 24032 1575 sw
rect 24003 1542 24032 1549
tri 24032 1542 24039 1549 sw
rect 24003 1512 25239 1542
rect 23947 1490 25239 1512
rect 25291 1490 25303 1542
rect 25355 1490 25361 1542
rect 23947 1488 24003 1490
tri 24003 1454 24039 1490 nw
rect 23947 1423 24003 1432
tri 20347 1404 20365 1422 ne
rect 20365 1404 20884 1422
tri 20365 1352 20417 1404 ne
rect 20417 1352 20519 1404
rect 20571 1352 20592 1404
rect 20644 1352 20665 1404
rect 20717 1352 20738 1404
rect 20790 1352 20810 1404
rect 20862 1352 20884 1404
tri 20417 1334 20435 1352 ne
rect 20435 1334 20884 1352
tri 20435 1333 20436 1334 ne
rect 20436 1333 20519 1334
tri 20436 1282 20487 1333 ne
rect 20487 1282 20519 1333
rect 20571 1282 20592 1334
rect 20644 1282 20665 1334
rect 20717 1282 20738 1334
rect 20790 1282 20810 1334
rect 20862 1282 20884 1334
tri 24218 1324 24260 1366 se
rect 24260 1324 25239 1366
tri 20487 1281 20488 1282 ne
rect 20488 1281 20884 1282
tri 20488 1274 20495 1281 ne
rect 20495 1274 20884 1281
rect 23942 1268 23951 1324
rect 24007 1268 24031 1324
rect 24087 1314 25239 1324
rect 25291 1314 25303 1366
rect 25355 1314 25361 1366
rect 24087 1268 24246 1314
tri 24246 1268 24292 1314 nw
tri 18212 1081 18239 1108 sw
rect 18122 1029 18128 1081
rect 18180 1029 18192 1081
rect 18244 1029 18250 1081
rect 18531 346 18537 398
rect 18589 346 18601 398
rect 18653 346 18659 398
rect 16355 326 16393 328
tri 16393 326 16395 328 nw
rect 14960 317 16215 321
rect 14478 315 16215 317
tri 16324 315 16335 326 se
rect 16335 315 16355 326
tri 16301 292 16324 315 se
rect 16324 292 16355 315
tri 16291 282 16301 292 se
rect 16301 288 16355 292
tri 16355 288 16393 326 nw
rect 16301 282 16349 288
tri 16349 282 16355 288 nw
tri 16277 268 16291 282 se
rect 16291 268 16335 282
tri 16335 268 16349 282 nw
tri 19029 268 19043 282 se
rect 19043 268 19161 282
rect 13060 193 13247 228
tri 13060 176 13077 193 ne
rect 13077 176 13247 193
tri 13247 176 13299 228 sw
rect 13799 176 13805 228
rect 13857 176 13876 228
rect 13928 176 13947 228
rect 13999 176 14018 228
rect 14070 176 14089 228
rect 14141 176 14159 228
rect 14211 176 14229 228
rect 14281 176 14299 228
rect 14351 176 14357 228
rect 15895 216 15901 268
rect 15953 216 15971 268
rect 16023 230 16297 268
tri 16297 230 16335 268 nw
tri 18991 230 19029 268 se
rect 19029 230 19161 268
rect 19213 230 19227 282
rect 19279 230 19354 282
rect 16023 227 16294 230
tri 16294 227 16297 230 nw
tri 18988 227 18991 230 se
rect 18991 227 19354 230
rect 16023 216 16029 227
tri 16029 216 16040 227 nw
tri 18977 216 18988 227 se
rect 18988 216 19354 227
tri 18967 206 18977 216 se
rect 18977 206 19354 216
tri 18937 176 18967 206 se
rect 18967 176 19161 206
tri 13077 175 13078 176 ne
rect 13078 175 13299 176
tri 13299 175 13300 176 sw
tri 18936 175 18937 176 se
rect 18937 175 19161 176
tri 12927 154 12928 155 ne
rect 12928 154 12977 155
tri 12977 154 12998 175 sw
tri 13078 154 13099 175 ne
rect 13099 154 13300 175
tri 13300 154 13321 175 sw
tri 18915 154 18936 175 se
rect 18936 154 19161 175
rect 19213 154 19227 206
rect 19279 154 19354 206
tri 12928 131 12951 154 ne
rect 12951 135 12998 154
tri 12998 135 13017 154 sw
tri 13099 135 13118 154 ne
rect 13118 135 13321 154
tri 13321 135 13340 154 sw
tri 18896 135 18915 154 se
rect 18915 135 19071 154
rect 12951 131 13017 135
tri 13017 131 13021 135 sw
tri 13118 131 13122 135 ne
rect 13122 131 13340 135
tri 13340 131 13344 135 sw
tri 16183 131 16187 135 se
rect 16187 131 16240 135
tri 12895 129 12897 131 sw
tri 12951 129 12953 131 ne
rect 12953 129 13021 131
tri 13021 129 13023 131 sw
tri 13122 129 13124 131 ne
rect 13124 129 13344 131
tri 13344 129 13346 131 sw
tri 16181 129 16183 131 se
rect 16183 129 16240 131
rect 12845 111 12897 129
tri 12845 97 12859 111 ne
rect 12859 105 12897 111
tri 12897 105 12921 129 sw
tri 12953 105 12977 129 ne
rect 12977 105 13023 129
tri 13023 105 13047 129 sw
tri 13124 124 13129 129 ne
rect 13129 124 13346 129
tri 13346 124 13351 129 sw
tri 16176 124 16181 129 se
rect 16181 124 16187 129
tri 13129 105 13148 124 ne
rect 13148 105 16187 124
rect 12859 97 12921 105
tri 12921 97 12929 105 sw
tri 12977 97 12985 105 ne
rect 12985 97 13047 105
tri 13047 97 13055 105 sw
tri 13148 97 13156 105 ne
rect 13156 97 16187 105
rect 2421 37 2553 89
rect 2605 37 2865 89
rect 2917 37 3769 89
rect 3821 37 4081 89
rect 4133 37 4393 89
rect 4445 37 4549 89
rect 4601 37 4861 89
rect 4913 37 5017 89
rect 5069 37 5329 89
rect 5381 37 5814 89
rect 5866 37 6407 89
rect 6459 37 6843 89
rect 6895 84 12737 89
rect 6895 37 7142 84
rect 2421 32 7142 37
rect 7194 32 7208 84
rect 7260 72 12737 84
tri 12859 77 12879 97 ne
rect 12879 77 12929 97
tri 12929 77 12949 97 sw
tri 12985 77 13005 97 ne
rect 13005 92 13055 97
tri 13055 92 13060 97 sw
tri 13156 92 13161 97 ne
rect 13161 92 16187 97
rect 13005 77 13060 92
tri 13060 77 13075 92 sw
tri 13161 77 13176 92 ne
rect 13176 77 16187 92
rect 16239 128 16240 129
tri 16240 128 16247 135 sw
tri 18889 128 18896 135 se
rect 18896 128 19071 135
tri 19071 128 19097 154 nw
rect 16239 124 16247 128
tri 16247 124 16251 128 sw
tri 18885 124 18889 128 se
rect 18889 124 19067 128
tri 19067 124 19071 128 nw
tri 22731 124 22735 128 se
rect 22735 124 22861 859
rect 16239 123 16251 124
tri 16251 123 16252 124 sw
tri 18302 123 18303 124 se
rect 18303 123 19066 124
tri 19066 123 19067 124 nw
tri 22730 123 22731 124 se
rect 22731 123 22861 124
rect 16239 94 19037 123
tri 19037 94 19066 123 nw
tri 22701 94 22730 123 se
rect 22730 94 22861 123
rect 16239 77 18983 94
rect 7260 32 8171 72
rect 2421 24 8171 32
rect 2421 -28 2553 24
rect 2605 -28 2865 24
rect 2917 -28 3769 24
rect 3821 -28 4081 24
rect 4133 -28 4393 24
rect 4445 -28 4549 24
rect 4601 -28 4861 24
rect 4913 -28 5017 24
rect 5069 -28 5329 24
rect 5381 -28 5814 24
rect 5866 -28 6407 24
rect 6459 -28 6843 24
rect 6895 20 8171 24
rect 8223 20 8275 72
rect 8327 20 8587 72
rect 8639 20 8899 72
rect 8951 20 9211 72
rect 9263 20 9523 72
rect 9575 57 12737 72
tri 12879 61 12895 77 ne
rect 12895 61 12949 77
rect 9575 20 10595 57
rect 6895 13 10595 20
rect 6895 -28 7142 13
rect 2421 -39 7142 -28
rect 7194 -39 7208 13
rect 7260 5 10595 13
rect 10647 5 10728 57
rect 10780 5 11184 57
rect 11236 5 11640 57
rect 11692 5 12097 57
rect 12149 5 12438 57
rect 12490 5 12520 57
rect 12572 5 12602 57
rect 12654 5 12684 57
rect 12736 5 12737 57
tri 12895 56 12900 61 ne
rect 12900 56 12949 61
tri 12949 56 12970 77 sw
tri 13005 56 13026 77 ne
rect 13026 56 13075 77
tri 13075 56 13096 77 sw
tri 13176 56 13197 77 ne
rect 13197 56 18983 77
tri 12900 27 12929 56 ne
rect 12929 49 12970 56
tri 12970 49 12977 56 sw
tri 13026 49 13033 56 ne
rect 13033 49 13096 56
rect 12929 35 12977 49
tri 12977 35 12991 49 sw
tri 13033 35 13047 49 ne
rect 13047 35 13096 49
tri 13096 35 13117 56 sw
tri 13197 35 13218 56 ne
rect 13218 35 16187 56
rect 12929 27 12991 35
tri 12991 27 12999 35 sw
tri 13047 27 13055 35 ne
rect 13055 34 13117 35
tri 13117 34 13118 35 sw
tri 13218 34 13219 35 ne
rect 13219 34 16187 35
rect 13055 27 13118 34
tri 13118 27 13125 34 sw
tri 13219 27 13226 34 ne
rect 13226 27 16187 34
rect 7260 -11 12737 5
tri 12929 4 12952 27 ne
rect 12952 4 12999 27
tri 12999 4 13022 27 sw
tri 13055 4 13078 27 ne
rect 13078 4 13125 27
tri 13125 4 13148 27 sw
tri 13226 4 13249 27 ne
rect 13249 4 16187 27
rect 16239 40 18983 56
tri 18983 40 19037 94 nw
rect 19106 40 19289 94
rect 22655 40 22861 94
rect 16239 6 18949 40
tri 18949 6 18983 40 nw
rect 16239 4 18941 6
rect 7260 -39 8171 -11
rect 2421 -46 8171 -39
rect 1612 -112 1866 -60
rect 1612 -128 1918 -112
rect 1612 -180 1866 -128
rect 1948 -53 2273 -47
rect 2000 -105 2221 -53
rect 1948 -117 2273 -105
rect 2000 -169 2221 -117
rect 2421 -98 2748 -46
rect 2800 -98 2813 -46
rect 2865 -98 2878 -46
rect 2930 -98 2943 -46
rect 2995 -98 3008 -46
rect 3060 -98 3073 -46
rect 3125 -98 3138 -46
rect 3190 -98 3203 -46
rect 3255 -98 3268 -46
rect 3320 -98 3333 -46
rect 3385 -98 3398 -46
rect 3450 -98 3463 -46
rect 3515 -98 3528 -46
rect 3580 -98 3593 -46
rect 3645 -98 3658 -46
rect 3710 -98 3723 -46
rect 3775 -98 3788 -46
rect 3840 -98 3853 -46
rect 3905 -98 3918 -46
rect 3970 -98 3983 -46
rect 4035 -98 4048 -46
rect 4100 -98 4113 -46
rect 4165 -98 4178 -46
rect 4230 -98 4243 -46
rect 4295 -98 4308 -46
rect 4360 -98 4373 -46
rect 4425 -98 4438 -46
rect 4490 -98 4503 -46
rect 4555 -98 4568 -46
rect 4620 -98 4632 -46
rect 4684 -98 4696 -46
rect 4748 -98 4760 -46
rect 4812 -98 4824 -46
rect 4876 -98 4888 -46
rect 4940 -98 4952 -46
rect 5004 -98 5016 -46
rect 5068 -98 5080 -46
rect 5132 -98 5144 -46
rect 5196 -98 5208 -46
rect 5260 -98 5272 -46
rect 5324 -98 5336 -46
rect 5388 -98 5400 -46
rect 5452 -98 5464 -46
rect 5516 -98 5528 -46
rect 5580 -98 5592 -46
rect 5644 -98 5680 -46
rect 5732 -98 5745 -46
rect 5797 -98 5810 -46
rect 5862 -98 5875 -46
rect 5927 -98 5940 -46
rect 5992 -98 6005 -46
rect 6057 -98 6070 -46
rect 6122 -98 6135 -46
rect 6187 -98 6200 -46
rect 6252 -98 6265 -46
rect 6317 -98 6330 -46
rect 6382 -98 6395 -46
rect 6447 -98 6460 -46
rect 6512 -98 6525 -46
rect 6577 -98 6590 -46
rect 6642 -98 6655 -46
rect 6707 -98 6720 -46
rect 6772 -98 6785 -46
rect 6837 -98 6850 -46
rect 6902 -58 8171 -46
rect 6902 -98 7142 -58
rect 2421 -110 7142 -98
rect 7194 -110 7208 -58
rect 7260 -63 8171 -58
rect 8223 -63 8275 -11
rect 8327 -63 8587 -11
rect 8639 -63 8899 -11
rect 8951 -63 9211 -11
rect 9263 -63 9523 -11
rect 9575 -38 12737 -11
rect 9575 -63 10595 -38
rect 7260 -90 10595 -63
rect 10647 -90 10728 -38
rect 10780 -90 11184 -38
rect 11236 -90 11640 -38
rect 11692 -90 12097 -38
rect 12149 -90 12438 -38
rect 12490 -90 12520 -38
rect 12572 -90 12602 -38
rect 12654 -90 12684 -38
rect 12736 -90 12737 -38
tri 12952 -42 12998 4 ne
rect 12998 -2 13022 4
tri 13022 -2 13028 4 sw
tri 13078 -2 13084 4 ne
rect 13084 -2 13148 4
tri 13148 -2 13154 4 sw
tri 13249 -2 13255 4 ne
rect 13255 -2 18941 4
tri 18941 -2 18949 6 nw
rect 12998 -21 13028 -2
tri 13028 -21 13047 -2 sw
tri 13084 -21 13103 -2 ne
rect 13103 -21 13154 -2
rect 12998 -35 13047 -21
tri 13047 -35 13061 -21 sw
tri 13103 -35 13117 -21 ne
rect 13117 -35 13154 -21
tri 13154 -35 13187 -2 sw
tri 16587 -4 16589 -2 ne
rect 16589 -4 18939 -2
tri 18939 -4 18941 -2 nw
rect 12998 -36 13061 -35
tri 13061 -36 13062 -35 sw
tri 13117 -36 13118 -35 ne
rect 13118 -36 16557 -35
tri 16557 -36 16558 -35 sw
rect 12998 -42 13062 -36
tri 13062 -42 13068 -36 sw
tri 13118 -42 13124 -36 ne
rect 13124 -42 18914 -36
tri 12998 -43 12999 -42 ne
rect 12999 -43 13068 -42
tri 13068 -43 13069 -42 sw
tri 13124 -43 13125 -42 ne
rect 13125 -43 18862 -42
tri 12999 -69 13025 -43 ne
rect 13025 -69 13069 -43
tri 13069 -69 13095 -43 sw
tri 13125 -69 13151 -43 ne
rect 13151 -69 18862 -43
rect 7260 -110 12737 -90
tri 13025 -94 13050 -69 ne
rect 13050 -85 13095 -69
tri 13095 -85 13111 -69 sw
tri 13151 -85 13167 -69 ne
rect 13167 -85 18862 -69
rect 13050 -94 13111 -85
tri 13111 -94 13120 -85 sw
tri 18828 -94 18837 -85 ne
rect 18837 -94 18862 -85
tri 13050 -106 13062 -94 ne
rect 13062 -106 13120 -94
tri 13120 -106 13132 -94 sw
tri 18837 -106 18849 -94 ne
rect 18849 -106 18914 -94
rect 2421 -137 12737 -110
tri 13062 -113 13069 -106 ne
rect 13069 -113 13132 -106
tri 13132 -113 13139 -106 sw
tri 18849 -113 18856 -106 ne
rect 18856 -113 18862 -106
tri 13069 -114 13070 -113 ne
rect 13070 -114 16508 -113
tri 16508 -114 16509 -113 sw
tri 18856 -114 18857 -113 ne
rect 18857 -114 18862 -113
tri 13070 -116 13072 -114 ne
rect 13072 -116 18803 -114
tri 13072 -120 13076 -116 ne
rect 13076 -120 18803 -116
tri 18857 -119 18862 -114 ne
tri 13076 -137 13093 -120 ne
rect 13093 -137 18751 -120
tri 13093 -163 13119 -137 ne
rect 13119 -163 18751 -137
tri 18672 -164 18673 -163 ne
rect 18673 -164 18751 -163
rect 1948 -175 2273 -169
tri 18673 -172 18681 -164 ne
rect 18681 -172 18751 -164
rect 18862 -164 18914 -158
tri 18681 -175 18684 -172 ne
rect 18684 -175 18803 -172
rect 1612 -196 1918 -180
tri 18684 -184 18693 -175 ne
rect 18693 -184 18803 -175
tri 18693 -191 18700 -184 ne
rect 18700 -191 18751 -184
rect 1612 -248 1866 -196
tri 13008 -227 13044 -191 se
rect 13044 -227 18362 -191
rect 1612 -265 1918 -248
rect 1612 -317 1866 -265
rect 1612 -334 1918 -317
rect 1612 -386 1866 -334
rect 1612 -420 1918 -386
rect 2221 -279 2227 -227
rect 2279 -279 2291 -227
rect 2343 -279 2349 -227
tri 12993 -242 13008 -227 se
rect 13008 -228 18362 -227
rect 13008 -242 13050 -228
tri 13050 -242 13064 -228 nw
tri 18341 -242 18355 -228 ne
rect 18355 -242 18362 -228
tri 12992 -243 12993 -242 se
rect 12993 -243 13049 -242
tri 13049 -243 13050 -242 nw
tri 18355 -243 18356 -242 ne
rect 18356 -243 18362 -242
rect 18414 -243 18426 -191
rect 18478 -243 18484 -191
rect 18522 -197 18574 -191
tri 12987 -248 12992 -243 se
rect 12992 -248 13044 -243
tri 13044 -248 13049 -243 nw
tri 12986 -249 12987 -248 se
rect 12987 -249 13043 -248
tri 13043 -249 13044 -248 nw
tri 18521 -249 18522 -248 se
tri 18700 -236 18745 -191 ne
rect 18745 -236 18751 -191
tri 18745 -242 18751 -236 ne
rect 18751 -242 18803 -236
tri 12974 -261 12986 -249 se
rect 12986 -261 13031 -249
tri 13031 -261 13043 -249 nw
tri 18509 -261 18521 -249 se
rect 18521 -261 18574 -249
tri 12956 -279 12974 -261 se
rect 12974 -279 12987 -261
tri 2191 -420 2221 -390 se
rect 2221 -420 2273 -279
tri 2273 -313 2307 -279 nw
tri 12930 -305 12956 -279 se
rect 12956 -305 12987 -279
tri 12987 -305 13031 -261 nw
tri 18488 -282 18509 -261 se
rect 18509 -282 18522 -261
tri 12924 -311 12930 -305 se
rect 12930 -311 12981 -305
tri 12981 -311 12987 -305 nw
tri 7443 -313 7445 -311 se
rect 7445 -313 12979 -311
tri 12979 -313 12981 -311 nw
tri 2189 -422 2191 -420 se
rect 2191 -422 2273 -420
rect 2132 -428 2273 -422
rect 2184 -465 2273 -428
tri 7408 -348 7443 -313 se
rect 7443 -348 12944 -313
tri 12944 -348 12979 -313 nw
rect 18354 -338 18382 -282
rect 18438 -338 18462 -282
rect 18518 -313 18522 -282
rect 18518 -319 18574 -313
rect 18518 -338 18555 -319
tri 18555 -338 18574 -319 nw
rect 2132 -492 2184 -480
tri 2184 -503 2222 -465 nw
rect 2132 -550 2184 -544
rect 3660 -703 3716 -694
rect 1610 -766 1662 -760
tri 3628 -793 3660 -761 se
rect 3660 -783 3716 -759
tri 7380 -767 7408 -739 se
rect 7408 -760 7463 -348
tri 7463 -392 7507 -348 nw
rect 7408 -767 7456 -760
tri 7456 -767 7463 -760 nw
tri 1662 -801 1670 -793 sw
tri 3626 -795 3628 -793 se
rect 3628 -795 3660 -793
rect 1779 -801 3660 -795
rect 1662 -818 1670 -801
rect 1610 -830 1670 -818
rect 1662 -853 1670 -830
tri 1670 -853 1722 -801 sw
rect 1831 -839 3660 -801
rect 1831 -848 3716 -839
tri 4165 -830 4228 -767 se
rect 4228 -813 7410 -767
tri 7410 -813 7456 -767 nw
tri 19074 -813 19106 -781 se
rect 19106 -813 19232 40
tri 22701 6 22735 40 ne
rect 4228 -830 4257 -813
tri 4257 -830 4274 -813 nw
tri 19057 -830 19074 -813 se
rect 19074 -830 19232 -813
rect 4165 -848 4239 -830
tri 4239 -848 4257 -830 nw
tri 19054 -833 19057 -830 se
rect 19057 -833 19232 -830
tri 19039 -848 19054 -833 se
rect 19054 -848 19217 -833
tri 19217 -848 19232 -833 nw
rect 1662 -865 1722 -853
tri 1722 -865 1734 -853 sw
rect 1779 -865 1831 -853
rect 1662 -882 1734 -865
tri 1734 -882 1751 -865 sw
rect 1610 -888 1751 -882
tri 1687 -916 1715 -888 ne
rect 1337 -1076 1343 -1024
rect 1395 -1076 1415 -1024
rect 1467 -1076 1487 -1024
rect 1539 -1076 1545 -1024
rect 1337 -1337 1545 -1076
rect 1628 -941 1680 -935
rect 1628 -1005 1680 -993
rect 1628 -1156 1680 -1057
rect 1715 -1135 1751 -888
tri 1831 -877 1860 -848 nw
tri 1912 -890 1914 -888 se
rect 1914 -890 3787 -888
rect 1779 -923 1831 -917
rect 1860 -896 3787 -890
rect 1912 -944 3787 -896
rect 3843 -944 3867 -888
rect 3923 -944 3932 -888
rect 3995 -889 4051 -880
rect 1912 -947 1941 -944
tri 1941 -947 1944 -944 nw
rect 1860 -960 1912 -948
tri 1912 -976 1941 -947 nw
tri 3966 -976 3995 -947 se
rect 3995 -969 4051 -945
tri 3961 -981 3966 -976 se
rect 3966 -981 3995 -976
rect 1860 -1018 1912 -1012
rect 1949 -987 3995 -981
rect 2001 -1025 3995 -987
rect 2001 -1034 4051 -1025
tri 4160 -1034 4165 -1029 se
rect 4165 -1034 4236 -848
tri 4236 -851 4239 -848 nw
tri 19036 -851 19039 -848 se
rect 19039 -851 19214 -848
tri 19214 -851 19217 -848 nw
rect 2001 -1038 2030 -1034
tri 2030 -1038 2034 -1034 nw
tri 4156 -1038 4160 -1034 se
rect 4160 -1038 4236 -1034
tri 18955 -932 19036 -851 se
rect 19036 -932 19081 -851
rect 2001 -1039 2016 -1038
rect 1949 -1051 2016 -1039
rect 2001 -1052 2016 -1051
tri 2016 -1052 2030 -1038 nw
tri 4142 -1052 4156 -1038 se
rect 4156 -1052 4236 -1038
tri 16891 -1052 16905 -1038 se
rect 16905 -1052 16911 -1038
rect 2001 -1066 2002 -1052
tri 2002 -1066 2016 -1052 nw
tri 4128 -1066 4142 -1052 se
rect 4142 -1066 4236 -1052
tri 2001 -1067 2002 -1066 nw
rect 1949 -1109 2001 -1103
rect 2225 -1118 2231 -1066
rect 2283 -1118 2295 -1066
rect 2347 -1082 4236 -1066
tri 7058 -1076 7082 -1052 se
rect 7082 -1076 16911 -1052
rect 2347 -1090 4228 -1082
tri 4228 -1090 4236 -1082 nw
tri 7044 -1090 7058 -1076 se
rect 7058 -1088 16911 -1076
rect 7058 -1090 7096 -1088
tri 7096 -1090 7098 -1088 nw
tri 16903 -1090 16905 -1088 ne
rect 16905 -1090 16911 -1088
rect 16963 -1090 16975 -1038
rect 17027 -1090 17033 -1038
rect 17096 -1090 17102 -1038
rect 17154 -1090 17166 -1038
rect 17218 -1090 17224 -1038
rect 2347 -1104 4214 -1090
tri 4214 -1104 4228 -1090 nw
tri 7030 -1104 7044 -1090 se
rect 7044 -1104 7082 -1090
tri 7082 -1104 7096 -1090 nw
tri 17082 -1104 17096 -1090 se
rect 17096 -1104 17224 -1090
rect 2347 -1118 4200 -1104
tri 4200 -1118 4214 -1104 nw
tri 7016 -1118 7030 -1104 se
rect 7030 -1118 7066 -1104
tri 7015 -1119 7016 -1118 se
rect 7016 -1119 7066 -1118
tri 1751 -1135 1767 -1119 sw
tri 6999 -1135 7015 -1119 se
rect 7015 -1120 7066 -1119
tri 7066 -1120 7082 -1104 nw
tri 17066 -1120 17082 -1104 se
rect 17082 -1120 17224 -1104
rect 7015 -1126 7060 -1120
tri 7060 -1126 7066 -1120 nw
tri 7106 -1126 7112 -1120 se
rect 7112 -1126 17224 -1120
rect 7015 -1135 7030 -1126
tri 1715 -1146 1726 -1135 ne
rect 1726 -1146 1767 -1135
tri 1680 -1156 1690 -1146 sw
tri 1726 -1156 1736 -1146 ne
rect 1736 -1156 1767 -1146
tri 1767 -1156 1788 -1135 sw
tri 6978 -1156 6999 -1135 se
rect 6999 -1156 7030 -1135
tri 7030 -1156 7060 -1126 nw
tri 7076 -1156 7106 -1126 se
rect 7106 -1133 17224 -1126
rect 7106 -1153 17204 -1133
tri 17204 -1153 17224 -1133 nw
rect 17258 -1090 17264 -1038
rect 17316 -1090 17328 -1038
rect 17380 -1090 17386 -1038
rect 7106 -1156 17201 -1153
tri 17201 -1156 17204 -1153 nw
tri 17255 -1156 17258 -1153 se
rect 17258 -1156 17386 -1090
rect 1628 -1158 1690 -1156
tri 1628 -1191 1661 -1158 ne
rect 1661 -1184 1690 -1158
tri 1690 -1184 1718 -1156 sw
tri 1736 -1184 1764 -1156 ne
rect 1764 -1184 1788 -1156
tri 1788 -1184 1816 -1156 sw
tri 6950 -1184 6978 -1156 se
rect 6978 -1172 7014 -1156
tri 7014 -1172 7030 -1156 nw
tri 7060 -1172 7076 -1156 se
rect 7076 -1172 7112 -1156
tri 7112 -1172 7128 -1156 nw
tri 17239 -1172 17255 -1156 se
rect 17255 -1172 17386 -1156
rect 6978 -1178 7008 -1172
tri 7008 -1178 7014 -1172 nw
tri 7054 -1178 7060 -1172 se
rect 7060 -1178 7096 -1172
rect 6978 -1184 6999 -1178
rect 1661 -1187 1718 -1184
tri 1718 -1187 1721 -1184 sw
tri 1764 -1187 1767 -1184 ne
rect 1767 -1187 1816 -1184
tri 1816 -1187 1819 -1184 sw
tri 6947 -1187 6950 -1184 se
rect 6950 -1187 6999 -1184
tri 6999 -1187 7008 -1178 nw
tri 7045 -1187 7054 -1178 se
rect 7054 -1187 7096 -1178
rect 1661 -1191 1721 -1187
tri 1721 -1191 1725 -1187 sw
tri 1767 -1191 1771 -1187 ne
rect 1771 -1191 6963 -1187
tri 1661 -1210 1680 -1191 ne
rect 1680 -1209 1725 -1191
tri 1725 -1209 1743 -1191 sw
tri 1771 -1209 1789 -1191 ne
rect 1789 -1209 6963 -1191
rect 1680 -1210 1743 -1209
tri 1680 -1255 1725 -1210 ne
rect 1725 -1223 1743 -1210
tri 1743 -1223 1757 -1209 sw
tri 1789 -1223 1803 -1209 ne
rect 1803 -1223 6963 -1209
tri 6963 -1223 6999 -1187 nw
tri 7009 -1223 7045 -1187 se
rect 7045 -1188 7096 -1187
tri 7096 -1188 7112 -1172 nw
tri 17223 -1188 17239 -1172 se
rect 17239 -1188 17386 -1172
rect 7045 -1194 7090 -1188
tri 7090 -1194 7096 -1188 nw
tri 7136 -1194 7142 -1188 se
rect 7142 -1194 17386 -1188
rect 7045 -1223 7060 -1194
rect 1725 -1224 1757 -1223
tri 1757 -1224 1758 -1223 sw
tri 7008 -1224 7009 -1223 se
rect 7009 -1224 7060 -1223
tri 7060 -1224 7090 -1194 nw
tri 7106 -1224 7136 -1194 se
rect 7136 -1224 17386 -1194
rect 1725 -1255 1758 -1224
tri 1758 -1255 1789 -1224 sw
tri 6977 -1255 7008 -1224 se
rect 7008 -1240 7044 -1224
tri 7044 -1240 7060 -1224 nw
tri 7090 -1240 7106 -1224 se
rect 7106 -1240 7142 -1224
tri 7142 -1240 7158 -1224 nw
rect 7008 -1246 7038 -1240
tri 7038 -1246 7044 -1240 nw
tri 7084 -1246 7090 -1240 se
rect 7008 -1255 7029 -1246
tri 7029 -1255 7038 -1246 nw
tri 7075 -1255 7084 -1246 se
rect 7084 -1255 7090 -1246
tri 1725 -1291 1761 -1255 ne
rect 1761 -1291 6993 -1255
tri 6993 -1291 7029 -1255 nw
tri 7039 -1291 7075 -1255 se
rect 7075 -1291 7090 -1255
tri 7038 -1292 7039 -1291 se
rect 7039 -1292 7090 -1291
tri 7090 -1292 7142 -1240 nw
tri 7018 -1312 7038 -1292 se
rect 7038 -1312 7059 -1292
tri 7017 -1313 7018 -1312 se
rect 7018 -1313 7059 -1312
rect 1337 -1389 1343 -1337
rect 1395 -1389 1415 -1337
rect 1467 -1389 1487 -1337
rect 1539 -1389 1545 -1337
tri 1155 -1470 1172 -1453 se
rect 1172 -1462 1226 -1453
tri 1226 -1462 1235 -1453 sw
rect 1172 -1470 1235 -1462
tri 1135 -1490 1155 -1470 se
rect 1155 -1490 1235 -1470
tri 1235 -1490 1263 -1462 sw
rect 1135 -1542 1141 -1490
rect 1193 -1542 1205 -1490
rect 1257 -1542 1263 -1490
tri 1298 -1632 1337 -1593 se
rect 1337 -1632 1545 -1389
rect 1609 -1319 1661 -1313
tri 1661 -1323 1671 -1313 sw
tri 7007 -1323 7017 -1313 se
rect 7017 -1323 7059 -1313
tri 7059 -1323 7090 -1292 nw
rect 1661 -1359 7023 -1323
tri 7023 -1359 7059 -1323 nw
rect 1661 -1371 1683 -1359
rect 1609 -1374 1683 -1371
tri 1683 -1374 1698 -1359 nw
rect 1609 -1398 1661 -1374
tri 1661 -1396 1683 -1374 nw
rect 1609 -1456 1661 -1450
rect 18955 -1408 19081 -932
tri 19081 -984 19214 -851 nw
tri 19081 -1408 19115 -1374 sw
tri 22701 -1408 22735 -1374 se
rect 22735 -1408 22861 40
rect 18955 -1462 19289 -1408
rect 22655 -1462 22861 -1408
rect 18955 -1490 19087 -1462
tri 19087 -1490 19115 -1462 nw
tri 22701 -1490 22729 -1462 ne
rect 22729 -1490 22861 -1462
tri 1284 -1646 1298 -1632 se
rect 1298 -1646 1545 -1632
rect 1613 -1501 2184 -1495
rect 1665 -1553 2132 -1501
rect 1613 -1580 2184 -1553
rect 1665 -1632 2132 -1580
rect 1613 -1638 2184 -1632
tri 1232 -1698 1284 -1646 se
rect 1284 -1698 1343 -1646
rect 1395 -1698 1415 -1646
rect 1467 -1698 1487 -1646
rect 1539 -1698 1545 -1646
tri 1190 -1740 1232 -1698 se
rect 1232 -1708 1545 -1698
rect 1232 -1740 1513 -1708
tri 1513 -1740 1545 -1708 nw
rect 2227 -1740 2279 -1734
tri 1138 -1792 1190 -1740 se
rect 1190 -1792 1461 -1740
tri 1461 -1792 1513 -1740 nw
tri 2202 -1792 2227 -1767 se
tri 1126 -1804 1138 -1792 se
rect 1138 -1804 1449 -1792
tri 1449 -1804 1461 -1792 nw
tri 2190 -1804 2202 -1792 se
rect 2202 -1804 2279 -1792
tri 1116 -1814 1126 -1804 se
rect 1126 -1808 1445 -1804
tri 1445 -1808 1449 -1804 nw
tri 2186 -1808 2190 -1804 se
rect 2190 -1808 2227 -1804
rect 1126 -1814 1439 -1808
tri 1439 -1814 1445 -1808 nw
rect 1501 -1814 2227 -1808
tri 1089 -1841 1116 -1814 se
rect 1116 -1841 1412 -1814
tri 1412 -1841 1439 -1814 nw
rect 1036 -1850 1387 -1841
rect 1092 -1866 1387 -1850
tri 1387 -1866 1412 -1841 nw
rect 1553 -1856 2227 -1814
rect 1553 -1862 2279 -1856
rect 1092 -1878 1375 -1866
tri 1375 -1878 1387 -1866 nw
rect 1501 -1878 1553 -1866
rect 1092 -1906 1323 -1878
rect 1036 -1930 1323 -1906
tri 1323 -1930 1375 -1878 nw
tri 1553 -1892 1583 -1862 nw
rect 1036 -1945 1319 -1930
tri 1319 -1934 1323 -1930 nw
rect 1501 -1936 1553 -1930
rect 1092 -1958 1319 -1945
rect 1092 -2001 1117 -1958
tri 907 -2010 911 -2006 sw
rect 1036 -2010 1117 -2001
rect 1169 -2010 1189 -1958
rect 1241 -2010 1261 -1958
rect 1313 -2010 1319 -1958
rect 859 -2040 911 -2010
tri 911 -2040 941 -2010 sw
rect 859 -2092 865 -2040
rect 917 -2092 929 -2040
rect 981 -2092 987 -2040
rect 1036 -2041 1319 -2010
rect 693 -2149 745 -2137
rect 693 -2207 745 -2201
rect 1092 -2097 1319 -2041
rect 1036 -2137 1319 -2097
rect 1092 -2150 1319 -2137
rect 1092 -2193 1110 -2150
rect 1036 -2202 1110 -2193
rect 1162 -2202 1185 -2150
rect 1237 -2202 1260 -2150
rect 1312 -2202 1319 -2150
rect 18955 -2910 19081 -1490
tri 19081 -1496 19087 -1490 nw
tri 22729 -1496 22735 -1490 ne
tri 19081 -2910 19115 -2876 sw
tri 22701 -2910 22735 -2876 se
rect 22735 -2910 22861 -1490
rect 18955 -2964 19289 -2910
rect 22655 -2964 22861 -2910
rect 395 -3432 744 -3426
rect 447 -3484 692 -3432
rect 395 -3496 744 -3484
rect 447 -3548 692 -3496
rect 395 -3554 744 -3548
rect 395 -4229 1918 -4227
rect 395 -4233 1697 -4229
rect 395 -4285 398 -4233
rect 450 -4285 1030 -4233
rect 1082 -4281 1697 -4233
rect 1749 -4234 1778 -4229
rect 1830 -4234 1859 -4229
rect 1830 -4281 1844 -4234
rect 1911 -4281 1918 -4229
rect 1082 -4285 1729 -4281
rect 395 -4290 1729 -4285
rect 1785 -4290 1844 -4281
rect 1900 -4290 1918 -4281
rect 395 -4299 1918 -4290
rect 395 -4351 398 -4299
rect 450 -4351 1030 -4299
rect 1082 -4351 1697 -4299
rect 1749 -4351 1778 -4299
rect 1830 -4351 1859 -4299
rect 1911 -4351 1918 -4299
rect 395 -4356 1918 -4351
rect 395 -4365 1729 -4356
rect 395 -4417 398 -4365
rect 450 -4417 1030 -4365
rect 1082 -4369 1729 -4365
rect 1785 -4369 1844 -4356
rect 1900 -4369 1918 -4356
rect 1082 -4417 1697 -4369
rect 1830 -4412 1844 -4369
rect 395 -4421 1697 -4417
rect 1749 -4421 1778 -4412
rect 1830 -4421 1859 -4412
rect 1911 -4421 1918 -4369
rect 395 -4423 1918 -4421
rect 18955 -4412 19081 -2964
tri 19081 -2998 19115 -2964 nw
tri 22701 -2998 22735 -2964 ne
tri 19081 -4412 19115 -4378 sw
tri 22701 -4412 22735 -4378 se
rect 22735 -4412 22861 -2964
rect 18955 -4466 19289 -4412
rect 22655 -4466 22861 -4412
rect 1036 -5455 1092 -5446
rect 1036 -5535 1092 -5511
rect 1036 -5635 1092 -5591
tri 996 -5677 1036 -5637 se
rect 1036 -5677 1050 -5635
tri 1050 -5677 1092 -5635 nw
tri 958 -5715 996 -5677 se
tri 942 -6463 958 -6447 se
rect 958 -6463 996 -5715
tri 996 -5731 1050 -5677 nw
rect 18955 -5914 19081 -4466
tri 19081 -4500 19115 -4466 nw
tri 22701 -4500 22735 -4466 ne
tri 19081 -5914 19115 -5880 sw
tri 22701 -5914 22735 -5880 se
rect 22735 -5914 22861 -4466
tri 889 -6516 942 -6463 se
rect 942 -6498 961 -6463
tri 961 -6498 996 -6463 nw
rect 1040 -5941 1096 -5932
rect 1040 -6021 1096 -5997
rect 1040 -6496 1096 -6077
rect 942 -6514 945 -6498
tri 945 -6514 961 -6498 nw
tri 1024 -6514 1040 -6498 se
rect 1040 -6514 1078 -6496
tri 1078 -6514 1096 -6496 nw
rect 18955 -5968 19289 -5914
rect 22655 -5968 22861 -5914
rect 942 -6516 943 -6514
tri 943 -6516 945 -6514 nw
tri 1022 -6516 1024 -6514 se
tri 835 -6570 889 -6516 se
rect 889 -6568 891 -6516
tri 891 -6568 943 -6516 nw
tri 970 -6568 1022 -6516 se
rect 1022 -6568 1024 -6516
tri 1024 -6568 1078 -6514 nw
tri 889 -6570 891 -6568 nw
tri 968 -6570 970 -6568 se
tri 781 -6624 835 -6570 se
rect 835 -6622 837 -6570
tri 837 -6622 889 -6570 nw
tri 916 -6622 968 -6570 se
rect 968 -6622 970 -6570
tri 970 -6622 1024 -6568 nw
tri 835 -6624 837 -6622 nw
tri 914 -6624 916 -6622 se
tri 743 -6662 781 -6624 se
rect 781 -6662 783 -6624
rect 743 -6676 783 -6662
tri 783 -6676 835 -6624 nw
tri 862 -6676 914 -6624 se
rect 914 -6676 916 -6624
tri 916 -6676 970 -6622 nw
tri 727 -11345 743 -11329 se
rect 743 -11345 781 -6676
tri 781 -6678 783 -6676 nw
tri 860 -6678 862 -6676 se
tri 674 -11398 727 -11345 se
rect 727 -11395 731 -11345
tri 731 -11395 781 -11345 nw
tri 824 -6714 860 -6678 se
rect 860 -6714 862 -6678
rect 727 -11398 728 -11395
tri 728 -11398 731 -11395 nw
tri 821 -11398 824 -11395 se
rect 824 -11398 862 -6714
tri 862 -6730 916 -6676 nw
rect 18955 -7416 19081 -5968
tri 19081 -6002 19115 -5968 nw
tri 22701 -6002 22735 -5968 ne
tri 19081 -7416 19115 -7382 sw
tri 22701 -7416 22735 -7382 se
rect 22735 -7416 22861 -5968
rect 18955 -7470 19289 -7416
rect 22655 -7470 22861 -7416
rect 18955 -8918 19081 -7470
tri 19081 -7504 19115 -7470 nw
tri 22701 -7504 22735 -7470 ne
tri 19081 -8918 19115 -8884 sw
tri 22701 -8918 22735 -8884 se
rect 22735 -8918 22861 -7470
rect 18955 -8972 19289 -8918
rect 22655 -8972 22861 -8918
rect 2610 -9602 2666 -9593
tri 2608 -9677 2610 -9675 se
rect 2610 -9677 2612 -9658
rect 2664 -9677 2666 -9658
tri 2596 -9689 2608 -9677 se
rect 2608 -9682 2666 -9677
rect 2608 -9689 2610 -9682
tri 2590 -9695 2596 -9689 se
rect 2596 -9695 2610 -9689
tri 2422 -9741 2468 -9695 se
rect 2468 -9738 2610 -9695
rect 2468 -9741 2612 -9738
rect 2664 -9741 2666 -9738
tri 2416 -9747 2422 -9741 se
rect 2422 -9747 2666 -9741
tri 2414 -9749 2416 -9747 se
rect 2416 -9749 2488 -9747
tri 2488 -9749 2490 -9747 nw
rect 2771 -9749 2823 -9743
tri 2394 -9769 2414 -9749 se
rect 2414 -9769 2468 -9749
tri 2468 -9769 2488 -9749 nw
tri 2389 -9774 2394 -9769 se
rect 2394 -9774 2463 -9769
tri 2463 -9774 2468 -9769 nw
rect 2389 -9778 2459 -9774
tri 2459 -9778 2463 -9774 nw
rect 2389 -10868 2441 -9778
tri 2441 -9796 2459 -9778 nw
tri 2753 -9796 2771 -9778 se
tri 2748 -9801 2753 -9796 se
rect 2753 -9801 2771 -9796
tri 2736 -9813 2748 -9801 se
rect 2748 -9813 2823 -9801
tri 2730 -9819 2736 -9813 se
rect 2736 -9819 2771 -9813
tri 2504 -9865 2550 -9819 se
rect 2550 -9865 2771 -9819
tri 2498 -9871 2504 -9865 se
rect 2504 -9871 2823 -9865
tri 2476 -9893 2498 -9871 se
rect 2498 -9893 2550 -9871
tri 2550 -9893 2572 -9871 nw
rect 2389 -10932 2441 -10920
rect 2389 -10990 2441 -10984
tri 2473 -9896 2476 -9893 se
rect 2476 -9896 2547 -9893
tri 2547 -9896 2550 -9893 nw
rect 2473 -10951 2525 -9896
tri 2525 -9918 2547 -9896 nw
rect 2641 -10223 2650 -10221
rect 2706 -10223 2730 -10221
rect 2641 -10275 2647 -10223
rect 2706 -10275 2711 -10223
rect 2641 -10277 2650 -10275
rect 2706 -10277 2730 -10275
rect 2786 -10277 2795 -10221
rect 2473 -11015 2525 -11003
rect 18955 -10420 19081 -8972
tri 19081 -9006 19115 -8972 nw
tri 22701 -9006 22735 -8972 ne
tri 19081 -10420 19115 -10386 sw
tri 22701 -10420 22735 -10386 se
rect 22735 -10420 22861 -8972
rect 18955 -10474 19289 -10420
rect 22655 -10474 22861 -10420
rect 2473 -11073 2525 -11067
tri 18925 -11073 18955 -11043 se
rect 18955 -11073 19081 -10474
tri 19081 -10508 19115 -10474 nw
tri 22701 -10508 22735 -10474 ne
tri 620 -11452 674 -11398 se
rect 674 -11411 715 -11398
tri 715 -11411 728 -11398 nw
tri 808 -11411 821 -11398 se
rect 821 -11411 862 -11398
rect 674 -11412 714 -11411
tri 714 -11412 715 -11411 nw
tri 807 -11412 808 -11411 se
rect 808 -11412 861 -11411
tri 861 -11412 862 -11411 nw
tri 18791 -11207 18925 -11073 se
rect 18925 -11207 19081 -11073
tri 674 -11452 714 -11412 nw
tri 767 -11452 807 -11412 se
tri 566 -11506 620 -11452 se
rect 620 -11466 660 -11452
tri 660 -11466 674 -11452 nw
tri 753 -11466 767 -11452 se
rect 767 -11466 807 -11452
tri 807 -11466 861 -11412 nw
tri 620 -11506 660 -11466 nw
tri 713 -11506 753 -11466 se
tri 512 -11560 566 -11506 se
rect 566 -11520 606 -11506
tri 606 -11520 620 -11506 nw
tri 699 -11520 713 -11506 se
rect 713 -11520 753 -11506
tri 753 -11520 807 -11466 nw
tri 566 -11560 606 -11520 nw
tri 659 -11560 699 -11520 se
tri 458 -11614 512 -11560 se
rect 512 -11574 552 -11560
tri 552 -11574 566 -11560 nw
tri 645 -11574 659 -11560 se
rect 659 -11574 699 -11560
tri 699 -11574 753 -11520 nw
tri 512 -11614 552 -11574 nw
tri 605 -11614 645 -11574 se
tri 404 -11668 458 -11614 se
rect 458 -11628 498 -11614
tri 498 -11628 512 -11614 nw
tri 591 -11628 605 -11614 se
rect 605 -11628 645 -11614
tri 645 -11628 699 -11574 nw
tri 458 -11668 498 -11628 nw
tri 551 -11668 591 -11628 se
tri 366 -11706 404 -11668 se
rect 404 -11682 444 -11668
tri 444 -11682 458 -11668 nw
tri 537 -11682 551 -11668 se
rect 551 -11682 591 -11668
tri 591 -11682 645 -11628 nw
tri 350 -13373 366 -13357 se
rect 366 -13373 404 -11706
tri 404 -11722 444 -11682 nw
tri 497 -11722 537 -11682 se
tri 483 -11736 497 -11722 se
rect 497 -11736 537 -11722
tri 537 -11736 591 -11682 nw
tri 336 -13387 350 -13373 se
rect 350 -13387 390 -13373
tri 390 -13387 404 -13373 nw
tri 445 -11774 483 -11736 se
tri 298 -13425 336 -13387 se
rect 298 -14040 336 -13425
tri 336 -13441 390 -13387 nw
tri 429 -13473 445 -13457 se
rect 445 -13473 483 -11774
tri 483 -11790 537 -11736 nw
rect 18791 -11922 19081 -11207
tri 19081 -11922 19115 -11888 sw
tri 22701 -11922 22735 -11888 se
rect 22735 -11922 22861 -10474
rect 3649 -11936 3701 -11930
rect 3649 -12000 3701 -11988
rect 3558 -12019 3610 -12013
rect 3558 -12083 3610 -12071
tri 3531 -12305 3558 -12278 se
rect 3558 -12300 3610 -12135
rect 3558 -12305 3605 -12300
tri 3605 -12305 3610 -12300 nw
tri 3484 -12352 3531 -12305 se
rect 3531 -12344 3566 -12305
tri 3566 -12344 3605 -12305 nw
tri 3610 -12344 3649 -12305 se
rect 3649 -12327 3701 -12052
rect 18791 -11976 19289 -11922
rect 22655 -11976 22861 -11922
rect 18791 -12156 19069 -11976
tri 19069 -12073 19166 -11976 nw
rect 3531 -12352 3558 -12344
tri 3558 -12352 3566 -12344 nw
tri 3602 -12352 3610 -12344 se
rect 3610 -12352 3649 -12344
tri 3457 -12379 3484 -12352 se
rect 3484 -12379 3531 -12352
tri 3531 -12379 3558 -12352 nw
tri 3575 -12379 3602 -12352 se
rect 3602 -12379 3649 -12352
tri 3649 -12379 3701 -12327 nw
tri 3410 -12426 3457 -12379 se
rect 3457 -12396 3514 -12379
tri 3514 -12396 3531 -12379 nw
tri 3558 -12396 3575 -12379 se
rect 3457 -12426 3484 -12396
tri 3484 -12426 3514 -12396 nw
tri 3528 -12426 3558 -12396 se
rect 3558 -12426 3575 -12396
tri 3383 -12453 3410 -12426 se
rect 3410 -12453 3457 -12426
tri 3457 -12453 3484 -12426 nw
tri 3501 -12453 3528 -12426 se
rect 3528 -12453 3575 -12426
tri 3575 -12453 3649 -12379 nw
tri 3336 -12500 3383 -12453 se
rect 3383 -12470 3440 -12453
tri 3440 -12470 3457 -12453 nw
tri 3484 -12470 3501 -12453 se
rect 3383 -12500 3410 -12470
tri 3410 -12500 3440 -12470 nw
tri 3454 -12500 3484 -12470 se
rect 3484 -12500 3501 -12470
tri 423 -13479 429 -13473 se
rect 429 -13479 477 -13473
tri 477 -13479 483 -13473 nw
tri 3323 -12513 3336 -12500 se
rect 3336 -12513 3397 -12500
tri 3397 -12513 3410 -12500 nw
tri 3441 -12513 3454 -12500 se
rect 3454 -12513 3501 -12500
rect 3323 -12527 3383 -12513
tri 3383 -12527 3397 -12513 nw
tri 3427 -12527 3441 -12513 se
rect 3441 -12527 3501 -12513
tri 3501 -12527 3575 -12453 nw
tri 385 -13517 423 -13479 se
rect 385 -13936 423 -13517
tri 423 -13533 477 -13479 nw
tri 423 -13936 429 -13930 sw
rect 385 -13946 429 -13936
tri 385 -13990 429 -13946 ne
tri 429 -13990 483 -13936 sw
tri 429 -14006 445 -13990 ne
tri 336 -14040 344 -14032 sw
rect 298 -14048 344 -14040
tri 298 -14094 344 -14048 ne
tri 344 -14094 398 -14040 sw
tri 344 -14110 360 -14094 ne
tri 344 -16955 360 -16939 se
rect 360 -16955 398 -14094
tri 293 -17006 344 -16955 se
rect 344 -17006 347 -16955
tri 347 -17006 398 -16955 nw
tri 255 -17044 293 -17006 se
rect 293 -17024 329 -17006
tri 329 -17024 347 -17006 nw
rect 293 -17040 313 -17024
tri 313 -17040 329 -17024 nw
tri 429 -17040 445 -17024 se
rect 445 -17040 483 -13990
tri 3298 -14298 3323 -14273 se
rect 3323 -14283 3375 -12527
tri 3375 -12535 3383 -12527 nw
tri 3419 -12535 3427 -12527 se
rect 3427 -12535 3485 -12527
rect 3323 -14298 3360 -14283
tri 3360 -14298 3375 -14283 nw
tri 3411 -12543 3419 -12535 se
rect 3419 -12543 3485 -12535
tri 3485 -12543 3501 -12527 nw
tri 3261 -14335 3298 -14298 se
rect 3298 -14334 3324 -14298
tri 3324 -14334 3360 -14298 nw
tri 3375 -14334 3411 -14298 se
rect 3411 -14304 3463 -12543
tri 3463 -12565 3485 -12543 nw
rect 3298 -14335 3323 -14334
tri 3323 -14335 3324 -14334 nw
tri 3374 -14335 3375 -14334 se
rect 3375 -14335 3411 -14334
tri 3240 -14356 3261 -14335 se
rect 3261 -14356 3302 -14335
tri 3302 -14356 3323 -14335 nw
tri 3353 -14356 3374 -14335 se
rect 3374 -14356 3411 -14335
tri 3411 -14356 3463 -14304 nw
tri 3219 -14377 3240 -14356 se
rect 3240 -14377 3281 -14356
tri 3281 -14377 3302 -14356 nw
tri 3332 -14377 3353 -14356 se
tri 3202 -14680 3219 -14663 se
rect 3219 -14680 3252 -14377
tri 3252 -14406 3281 -14377 nw
tri 3303 -14406 3332 -14377 se
rect 3332 -14406 3353 -14377
tri 3295 -14414 3303 -14406 se
rect 3303 -14414 3353 -14406
tri 3353 -14414 3411 -14356 nw
tri 3282 -14427 3295 -14414 se
rect 3295 -14427 3340 -14414
tri 3340 -14427 3353 -14414 nw
tri 3252 -14680 3254 -14678 sw
rect 3202 -14686 3254 -14680
rect 3202 -14750 3254 -14738
rect 3202 -14808 3254 -14802
tri 3202 -14825 3219 -14808 ne
rect 255 -17659 293 -17044
tri 293 -17060 313 -17040 nw
tri 409 -17060 429 -17040 se
rect 429 -17060 436 -17040
tri 382 -17087 409 -17060 se
rect 409 -17087 436 -17060
tri 436 -17087 483 -17040 nw
tri 344 -17125 382 -17087 se
rect 382 -17090 433 -17087
tri 433 -17090 436 -17087 nw
rect 382 -17125 387 -17090
rect 344 -17136 387 -17125
tri 387 -17136 433 -17090 nw
tri 3173 -17136 3219 -17090 se
rect 3219 -17103 3252 -14808
tri 3252 -14810 3254 -14808 nw
tri 3219 -17136 3252 -17103 nw
rect 344 -17596 382 -17136
tri 382 -17141 387 -17136 nw
tri 3168 -17141 3173 -17136 se
rect 3173 -17141 3184 -17136
tri 3138 -17171 3168 -17141 se
rect 3168 -17171 3184 -17141
tri 3184 -17171 3219 -17136 nw
tri 3127 -17182 3138 -17171 se
rect 3138 -17182 3173 -17171
tri 3173 -17182 3184 -17171 nw
tri 3271 -17182 3282 -17171 se
rect 3282 -17182 3316 -14427
tri 3316 -14451 3340 -14427 nw
tri 3090 -17219 3127 -17182 se
rect 3127 -17219 3140 -17182
tri 3140 -17215 3173 -17182 nw
tri 3238 -17215 3271 -17182 se
rect 3271 -17185 3316 -17182
rect 3271 -17215 3282 -17185
tri 3234 -17219 3238 -17215 se
rect 3238 -17219 3282 -17215
tri 3282 -17219 3316 -17185 nw
tri 3088 -17221 3090 -17219 se
rect 3090 -17221 3140 -17219
rect 3088 -17422 3140 -17221
tri 3186 -17267 3234 -17219 se
tri 3234 -17267 3282 -17219 nw
rect 3088 -17488 3140 -17474
rect 3088 -17546 3140 -17540
tri 3173 -17280 3186 -17267 se
rect 3186 -17280 3225 -17267
tri 3225 -17276 3234 -17267 nw
rect 3173 -17425 3225 -17280
rect 3173 -17489 3225 -17477
rect 3173 -17547 3225 -17541
tri 344 -17627 375 -17596 ne
rect 375 -17627 382 -17596
tri 382 -17627 429 -17580 sw
tri 375 -17634 382 -17627 ne
rect 382 -17634 429 -17627
tri 382 -17643 391 -17634 ne
rect 391 -17643 429 -17634
tri 255 -17695 291 -17659 ne
rect 291 -17681 293 -17659
tri 293 -17681 331 -17643 sw
tri 391 -17681 429 -17643 ne
tri 429 -17681 483 -17627 sw
rect 291 -17695 331 -17681
tri 331 -17695 345 -17681 sw
tri 429 -17695 443 -17681 ne
rect 443 -17695 483 -17681
tri 291 -17697 293 -17695 ne
rect 293 -17697 345 -17695
tri 345 -17697 347 -17695 sw
tri 443 -17697 445 -17695 ne
tri 293 -17749 345 -17697 ne
rect 345 -17749 347 -17697
tri 347 -17749 399 -17697 sw
tri 345 -17765 361 -17749 ne
rect 361 -19428 399 -17749
rect 445 -19402 483 -17695
tri 2468 -18696 2492 -18672 se
rect 2492 -18696 2498 -18672
rect 2468 -18724 2498 -18696
rect 2550 -18724 2562 -18672
rect 2614 -18724 2620 -18672
tri 483 -19402 493 -19392 sw
rect 445 -19408 493 -19402
tri 445 -19419 456 -19408 ne
rect 456 -19419 493 -19408
tri 399 -19428 408 -19419 sw
tri 456 -19428 465 -19419 ne
rect 465 -19422 493 -19419
tri 493 -19422 513 -19402 sw
tri 2448 -19422 2468 -19402 se
rect 2468 -19418 2506 -18724
tri 2506 -18761 2543 -18724 nw
rect 2468 -19422 2502 -19418
tri 2502 -19422 2506 -19418 nw
rect 2561 -18794 2613 -18788
rect 2561 -18858 2613 -18846
rect 465 -19424 513 -19422
tri 513 -19424 515 -19422 sw
tri 2446 -19424 2448 -19422 se
rect 2448 -19424 2500 -19422
tri 2500 -19424 2502 -19422 nw
tri 2559 -19424 2561 -19422 se
rect 2561 -19424 2613 -18910
rect 465 -19428 515 -19424
tri 515 -19428 519 -19424 sw
tri 2442 -19428 2446 -19424 se
rect 2446 -19428 2468 -19424
rect 361 -19435 408 -19428
tri 361 -19451 377 -19435 ne
rect 377 -19446 408 -19435
tri 408 -19446 426 -19428 sw
tri 465 -19446 483 -19428 ne
rect 483 -19446 780 -19428
rect 377 -19451 426 -19446
tri 426 -19451 431 -19446 sw
tri 483 -19451 488 -19446 ne
rect 488 -19451 780 -19446
tri 377 -19473 399 -19451 ne
rect 399 -19466 431 -19451
tri 431 -19466 446 -19451 sw
tri 488 -19466 503 -19451 ne
rect 503 -19456 780 -19451
tri 780 -19456 808 -19428 sw
tri 2414 -19456 2442 -19428 se
rect 2442 -19456 2468 -19428
tri 2468 -19456 2500 -19424 nw
tri 2527 -19456 2559 -19424 se
rect 2559 -19456 2570 -19424
rect 503 -19466 808 -19456
tri 808 -19466 818 -19456 sw
tri 2404 -19466 2414 -19456 se
rect 2414 -19466 2457 -19456
rect 399 -19473 446 -19466
tri 399 -19505 431 -19473 ne
rect 431 -19505 446 -19473
tri 446 -19505 485 -19466 sw
tri 764 -19505 803 -19466 ne
rect 803 -19467 818 -19466
tri 818 -19467 819 -19466 sw
tri 2403 -19467 2404 -19466 se
rect 2404 -19467 2457 -19466
tri 2457 -19467 2468 -19456 nw
tri 2516 -19467 2527 -19456 se
rect 2527 -19467 2570 -19456
tri 2570 -19467 2613 -19424 nw
rect 803 -19505 819 -19467
tri 431 -19537 463 -19505 ne
rect 463 -19520 743 -19505
tri 743 -19520 758 -19505 sw
tri 803 -19520 818 -19505 ne
rect 818 -19510 819 -19505
tri 819 -19510 862 -19467 sw
tri 2360 -19510 2403 -19467 se
rect 2403 -19510 2414 -19467
tri 2414 -19510 2457 -19467 nw
tri 2473 -19510 2516 -19467 se
rect 818 -19520 862 -19510
tri 862 -19520 872 -19510 sw
tri 2350 -19520 2360 -19510 se
rect 2360 -19520 2404 -19510
tri 2404 -19520 2414 -19510 nw
tri 2463 -19520 2473 -19510 se
rect 2473 -19520 2516 -19510
rect 463 -19521 758 -19520
tri 758 -19521 759 -19520 sw
tri 818 -19521 819 -19520 ne
rect 819 -19521 2403 -19520
tri 2403 -19521 2404 -19520 nw
tri 2462 -19521 2463 -19520 se
rect 2463 -19521 2516 -19520
tri 2516 -19521 2570 -19467 nw
rect 463 -19537 759 -19521
tri 759 -19537 775 -19521 sw
tri 819 -19537 835 -19521 ne
rect 835 -19537 2366 -19521
tri 463 -19543 469 -19537 ne
rect 469 -19543 775 -19537
tri 727 -19591 775 -19543 ne
tri 775 -19558 796 -19537 sw
tri 835 -19558 856 -19537 ne
rect 856 -19558 2366 -19537
tri 2366 -19558 2403 -19521 nw
tri 2425 -19558 2462 -19521 se
rect 775 -19559 796 -19558
tri 796 -19559 797 -19558 sw
rect 1789 -19559 2365 -19558
tri 2365 -19559 2366 -19558 nw
tri 2424 -19559 2425 -19558 se
rect 2425 -19559 2462 -19558
rect 775 -19575 797 -19559
tri 797 -19575 813 -19559 sw
tri 2408 -19575 2424 -19559 se
rect 2424 -19575 2462 -19559
tri 2462 -19575 2516 -19521 nw
rect 775 -19591 813 -19575
tri 813 -19591 829 -19575 sw
tri 2392 -19591 2408 -19575 se
tri 775 -19629 813 -19591 ne
rect 813 -19629 2408 -19591
tri 2408 -19629 2462 -19575 nw
rect 1790 -19630 2348 -19629
<< via2 >>
rect 18729 4852 18785 4908
rect 18809 4852 18865 4908
rect 777 475 833 531
rect 777 395 833 451
rect 1111 2451 1167 2507
rect 1191 2451 1247 2507
rect 2689 4355 2742 4379
rect 2742 4355 2745 4379
rect 2771 4355 2794 4379
rect 2794 4355 2827 4379
rect 2689 4343 2745 4355
rect 2771 4343 2827 4355
rect 2689 4323 2742 4343
rect 2742 4323 2745 4343
rect 2771 4323 2794 4343
rect 2794 4323 2827 4343
rect 2853 4323 2909 4379
rect 2935 4323 2991 4379
rect 3017 4323 3073 4379
rect 3099 4323 3155 4379
rect 3180 4323 3236 4379
rect 3261 4355 3306 4379
rect 3306 4355 3317 4379
rect 3261 4343 3317 4355
rect 3261 4323 3306 4343
rect 3306 4323 3317 4343
rect 3342 4323 3398 4379
rect 3423 4323 3479 4379
rect 3504 4323 3560 4379
rect 2689 3757 2742 3777
rect 2742 3757 2745 3777
rect 2771 3757 2794 3777
rect 2794 3757 2827 3777
rect 2689 3745 2745 3757
rect 2771 3745 2827 3757
rect 2689 3721 2742 3745
rect 2742 3721 2745 3745
rect 2771 3721 2794 3745
rect 2794 3721 2827 3745
rect 2853 3721 2909 3777
rect 2935 3721 2991 3777
rect 3017 3721 3073 3777
rect 3099 3721 3155 3777
rect 3180 3721 3236 3777
rect 3261 3757 3306 3777
rect 3306 3757 3317 3777
rect 3261 3745 3317 3757
rect 3261 3721 3306 3745
rect 3306 3721 3317 3745
rect 3342 3721 3398 3777
rect 3423 3721 3479 3777
rect 3504 3721 3560 3777
rect 2689 3313 2745 3369
rect 2771 3313 2827 3369
rect 2853 3313 2909 3369
rect 2935 3313 2991 3369
rect 3017 3345 3050 3369
rect 3050 3345 3073 3369
rect 3017 3333 3073 3345
rect 3017 3313 3050 3333
rect 3050 3313 3073 3333
rect 3099 3313 3155 3369
rect 3180 3313 3236 3369
rect 3261 3313 3317 3369
rect 3342 3313 3398 3369
rect 3423 3313 3479 3369
rect 3504 3345 3510 3369
rect 3510 3345 3560 3369
rect 3504 3333 3560 3345
rect 3504 3313 3510 3333
rect 3510 3313 3560 3333
rect 3657 3177 3713 3233
rect 2219 3099 2275 3155
rect 2299 3099 2355 3155
rect 3657 3097 3713 3153
rect 5131 3134 5187 3136
rect 5260 3134 5316 3136
rect 1728 1676 1784 1732
rect 1728 1596 1784 1652
rect 1117 1431 1173 1487
rect 1117 1351 1173 1407
rect 959 -1416 1015 -1414
rect 1039 -1416 1095 -1414
rect 959 -1468 1008 -1416
rect 1008 -1468 1015 -1416
rect 1039 -1468 1087 -1416
rect 1087 -1468 1095 -1416
rect 959 -1470 1015 -1468
rect 1039 -1470 1095 -1468
rect 5131 3082 5154 3134
rect 5154 3082 5169 3134
rect 5169 3082 5187 3134
rect 5260 3082 5288 3134
rect 5288 3082 5303 3134
rect 5303 3082 5316 3134
rect 5131 3080 5187 3082
rect 5260 3080 5316 3082
rect 1609 881 1665 937
rect 1609 801 1665 857
rect 3660 1096 3716 1152
rect 3660 1016 3716 1072
rect 14706 3707 14762 3763
rect 14827 3707 14883 3763
rect 14948 3707 15004 3763
rect 15068 3707 15124 3763
rect 15188 3707 15244 3763
rect 14706 3607 14762 3663
rect 14827 3607 14883 3663
rect 14948 3607 15004 3663
rect 15068 3607 15124 3663
rect 15188 3607 15244 3663
rect 14706 3507 14762 3563
rect 14827 3507 14883 3563
rect 14948 3507 15004 3563
rect 15068 3507 15124 3563
rect 15188 3507 15244 3563
rect 2015 881 2071 937
rect 2095 881 2151 937
rect 3787 889 3843 945
rect 3867 889 3923 945
rect 2013 533 2149 669
rect 2063 221 2119 240
rect 2063 184 2065 221
rect 2065 184 2117 221
rect 2117 184 2119 221
rect 2063 157 2119 160
rect 2063 105 2065 157
rect 2065 105 2117 157
rect 2117 105 2119 157
rect 2063 104 2119 105
rect 19004 4600 19060 4656
rect 19084 4600 19140 4656
rect 18414 4474 18470 4530
rect 18494 4474 18550 4530
rect 18569 3466 18625 3522
rect 18649 3466 18705 3522
rect 25337 2075 25393 2077
rect 25417 2075 25473 2077
rect 25337 2023 25386 2075
rect 25386 2023 25393 2075
rect 25417 2023 25450 2075
rect 25450 2023 25473 2075
rect 25337 2021 25393 2023
rect 25417 2021 25473 2023
rect 18873 1804 18929 1860
rect 18953 1804 19009 1860
rect 23947 1512 24003 1568
rect 23947 1432 24003 1488
rect 23951 1268 24007 1324
rect 24031 1268 24087 1324
rect 18382 -338 18438 -282
rect 18462 -338 18518 -282
rect 3660 -759 3716 -703
rect 3660 -839 3716 -783
rect 3787 -944 3843 -888
rect 3867 -944 3923 -888
rect 3995 -945 4051 -889
rect 3995 -1025 4051 -969
rect 1036 -1906 1092 -1850
rect 1036 -2001 1092 -1945
rect 1036 -2097 1092 -2041
rect 1036 -2193 1092 -2137
rect 1729 -4281 1749 -4234
rect 1749 -4281 1778 -4234
rect 1778 -4281 1785 -4234
rect 1844 -4281 1859 -4234
rect 1859 -4281 1900 -4234
rect 1729 -4290 1785 -4281
rect 1844 -4290 1900 -4281
rect 1729 -4369 1785 -4356
rect 1844 -4369 1900 -4356
rect 1729 -4412 1749 -4369
rect 1749 -4412 1778 -4369
rect 1778 -4412 1785 -4369
rect 1844 -4412 1859 -4369
rect 1859 -4412 1900 -4369
rect 1036 -5511 1092 -5455
rect 1036 -5591 1092 -5535
rect 1040 -5997 1096 -5941
rect 1040 -6077 1096 -6021
rect 2610 -9625 2666 -9602
rect 2610 -9658 2612 -9625
rect 2612 -9658 2664 -9625
rect 2664 -9658 2666 -9625
rect 2610 -9689 2666 -9682
rect 2610 -9738 2612 -9689
rect 2612 -9738 2664 -9689
rect 2664 -9738 2666 -9689
rect 2650 -10223 2706 -10221
rect 2730 -10223 2786 -10221
rect 2650 -10275 2699 -10223
rect 2699 -10275 2706 -10223
rect 2730 -10275 2763 -10223
rect 2763 -10275 2786 -10223
rect 2650 -10277 2706 -10275
rect 2730 -10277 2786 -10275
<< metal3 >>
rect 18724 4908 23859 4913
rect 18724 4852 18729 4908
rect 18785 4852 18809 4908
rect 18865 4878 23859 4908
tri 23859 4878 23894 4913 sw
rect 18865 4852 23894 4878
rect 18724 4847 23894 4852
tri 23831 4808 23870 4847 ne
rect 23870 4808 23894 4847
tri 3960 4748 4020 4808 se
rect 4020 4784 16534 4808
tri 16534 4784 16558 4808 sw
tri 23870 4784 23894 4808 ne
tri 23894 4784 23988 4878 sw
rect 4020 4748 16558 4784
tri 16558 4748 16594 4784 sw
tri 23894 4748 23930 4784 ne
rect 23930 4748 23988 4784
tri 3926 4714 3960 4748 se
rect 3960 4742 16594 4748
rect 3960 4714 4020 4742
tri 4020 4714 4048 4742 nw
tri 16508 4714 16536 4742 ne
rect 16536 4714 16594 4742
tri 3868 4656 3926 4714 se
rect 3926 4656 3962 4714
tri 3962 4656 4020 4714 nw
tri 16536 4656 16594 4714 ne
tri 16594 4690 16652 4748 sw
tri 23930 4690 23988 4748 ne
tri 23988 4690 24082 4784 sw
rect 16594 4661 16652 4690
tri 16652 4661 16681 4690 sw
tri 23988 4661 24017 4690 ne
rect 24017 4661 24082 4690
rect 16594 4656 16681 4661
tri 16681 4656 16686 4661 sw
tri 18994 4656 18999 4661 se
rect 18999 4656 19145 4661
tri 3832 4620 3868 4656 se
rect 3868 4620 3926 4656
tri 3926 4620 3962 4656 nw
tri 16594 4620 16630 4656 ne
rect 16630 4620 19004 4656
tri 3812 4600 3832 4620 se
rect 3832 4600 3906 4620
tri 3906 4600 3926 4620 nw
tri 16630 4600 16650 4620 ne
rect 16650 4600 19004 4620
rect 19060 4600 19084 4656
rect 19140 4600 19145 4656
tri 3807 4595 3812 4600 se
rect 3812 4595 3901 4600
tri 3901 4595 3906 4600 nw
tri 16650 4595 16655 4600 ne
rect 16655 4595 19145 4600
tri 24017 4596 24082 4661 ne
tri 24082 4596 24176 4690 sw
tri 24082 4595 24083 4596 ne
rect 24083 4595 24176 4596
tri 3747 4535 3807 4595 se
rect 3807 4535 3841 4595
tri 3841 4535 3901 4595 nw
tri 24083 4535 24143 4595 ne
rect 24143 4535 24176 4595
tri 3742 4530 3747 4535 se
rect 3747 4530 3836 4535
tri 3836 4530 3841 4535 nw
rect 18409 4530 18555 4535
tri 3738 4526 3742 4530 se
rect 3742 4526 3832 4530
tri 3832 4526 3836 4530 nw
tri 3686 4474 3738 4526 se
rect 3738 4474 3780 4526
tri 3780 4474 3832 4526 nw
rect 18409 4474 18414 4530
rect 18470 4474 18494 4530
rect 18550 4474 18555 4530
tri 24143 4502 24176 4535 ne
tri 24176 4502 24270 4596 sw
tri 3681 4469 3686 4474 se
rect 3686 4469 3775 4474
tri 3775 4469 3780 4474 nw
rect 18409 4469 18555 4474
tri 24176 4469 24209 4502 ne
rect 24209 4469 24270 4502
tri 3652 4440 3681 4469 se
rect 3681 4440 3746 4469
tri 3746 4440 3775 4469 nw
tri 24209 4440 24238 4469 ne
rect 24238 4440 24270 4469
rect 3652 4418 3724 4440
tri 3724 4418 3746 4440 nw
tri 24238 4418 24260 4440 ne
rect 24260 4418 24270 4440
rect 2684 4379 3565 4418
rect 2684 4323 2689 4379
rect 2745 4323 2771 4379
rect 2827 4323 2853 4379
rect 2909 4323 2935 4379
rect 2991 4323 3017 4379
rect 3073 4323 3099 4379
rect 3155 4323 3180 4379
rect 3236 4323 3261 4379
rect 3317 4323 3342 4379
rect 3398 4323 3423 4379
rect 3479 4323 3504 4379
rect 3560 4323 3565 4379
rect 2684 4284 3565 4323
rect 2684 3777 3565 3816
rect 2684 3721 2689 3777
rect 2745 3721 2771 3777
rect 2827 3721 2853 3777
rect 2909 3721 2935 3777
rect 2991 3721 3017 3777
rect 3073 3721 3099 3777
rect 3155 3721 3180 3777
rect 3236 3721 3261 3777
rect 3317 3721 3342 3777
rect 3398 3721 3423 3777
rect 3479 3721 3504 3777
rect 3560 3721 3565 3777
rect 2684 3682 3565 3721
rect 2684 3369 3565 3408
rect 2684 3313 2689 3369
rect 2745 3313 2771 3369
rect 2827 3313 2853 3369
rect 2909 3313 2935 3369
rect 2991 3313 3017 3369
rect 3073 3313 3099 3369
rect 3155 3313 3180 3369
rect 3236 3313 3261 3369
rect 3317 3313 3342 3369
rect 3398 3313 3423 3369
rect 3479 3313 3504 3369
rect 3560 3313 3565 3369
rect 2684 3274 3565 3313
rect 3652 3233 3718 4418
tri 3718 4412 3724 4418 nw
tri 24260 4412 24266 4418 ne
rect 24266 4412 24270 4418
tri 24266 4408 24270 4412 ne
tri 24270 4408 24364 4502 sw
tri 24270 4314 24364 4408 ne
tri 24364 4314 24458 4408 sw
tri 24364 4220 24458 4314 ne
tri 24458 4220 24552 4314 sw
tri 24458 4126 24552 4220 ne
tri 24552 4126 24646 4220 sw
tri 24552 4032 24646 4126 ne
tri 24646 4032 24740 4126 sw
tri 24646 3938 24740 4032 ne
tri 24740 3938 24834 4032 sw
tri 24740 3844 24834 3938 ne
tri 24834 3844 24928 3938 sw
tri 24834 3822 24856 3844 ne
rect 24856 3822 24928 3844
rect 14578 3758 14584 3822
rect 14648 3763 14728 3822
rect 14792 3763 14871 3822
rect 14935 3763 15014 3822
rect 15078 3763 15157 3822
rect 15221 3763 15300 3822
rect 14648 3758 14706 3763
rect 14792 3758 14827 3763
rect 14935 3758 14948 3763
rect 14578 3707 14706 3758
rect 14762 3707 14827 3758
rect 14883 3707 14948 3758
rect 15004 3758 15014 3763
rect 15124 3758 15157 3763
rect 15244 3758 15300 3763
rect 15364 3758 15370 3822
rect 15004 3707 15068 3758
rect 15124 3707 15188 3758
rect 15244 3707 15370 3758
tri 24856 3750 24928 3822 ne
tri 24928 3750 25022 3844 sw
rect 14578 3686 15370 3707
rect 14578 3622 14584 3686
rect 14648 3663 14728 3686
rect 14792 3663 14871 3686
rect 14935 3663 15014 3686
rect 15078 3663 15157 3686
rect 15221 3663 15300 3686
rect 14648 3622 14706 3663
rect 14792 3622 14827 3663
rect 14935 3622 14948 3663
rect 14578 3607 14706 3622
rect 14762 3607 14827 3622
rect 14883 3607 14948 3622
rect 15004 3622 15014 3663
rect 15124 3622 15157 3663
rect 15244 3622 15300 3663
rect 15364 3622 15370 3686
tri 24928 3656 25022 3750 ne
tri 25022 3656 25116 3750 sw
tri 25022 3653 25025 3656 ne
rect 25025 3653 25116 3656
rect 15004 3607 15068 3622
rect 15124 3607 15188 3622
rect 15244 3607 15370 3622
rect 14578 3563 15370 3607
rect 18383 3619 23164 3653
tri 23164 3619 23198 3653 sw
tri 25025 3619 25059 3653 ne
rect 25059 3619 25116 3653
rect 18383 3587 23198 3619
rect 14578 3550 14706 3563
rect 14762 3550 14827 3563
rect 14883 3550 14948 3563
rect 14578 3486 14584 3550
rect 14648 3507 14706 3550
rect 14792 3507 14827 3550
rect 14935 3507 14948 3550
rect 15004 3550 15068 3563
rect 15124 3550 15188 3563
rect 15244 3550 15370 3563
rect 15004 3507 15014 3550
rect 15124 3507 15157 3550
rect 15244 3507 15300 3550
rect 14648 3486 14728 3507
rect 14792 3486 14871 3507
rect 14935 3486 15014 3507
rect 15078 3486 15157 3507
rect 15221 3486 15300 3507
rect 15364 3486 15370 3550
tri 23136 3527 23196 3587 ne
rect 23196 3562 23198 3587
tri 23198 3562 23255 3619 sw
tri 25059 3562 25116 3619 ne
tri 25116 3562 25210 3656 sw
rect 23196 3527 23255 3562
tri 23255 3527 23290 3562 sw
tri 25116 3527 25151 3562 ne
rect 25151 3527 25210 3562
rect 18383 3525 23107 3527
tri 23107 3525 23109 3527 sw
tri 23196 3525 23198 3527 ne
rect 23198 3525 23290 3527
tri 23290 3525 23292 3527 sw
tri 25151 3525 25153 3527 ne
rect 25153 3525 25210 3527
rect 18383 3522 23109 3525
rect 18383 3466 18569 3522
rect 18625 3466 18649 3522
rect 18705 3472 23109 3522
tri 23109 3472 23162 3525 sw
tri 23198 3472 23251 3525 ne
rect 23251 3472 23292 3525
tri 23292 3472 23345 3525 sw
tri 25153 3472 25206 3525 ne
rect 25206 3472 25210 3525
rect 18705 3468 23162 3472
tri 23162 3468 23166 3472 sw
tri 23251 3468 23255 3472 ne
rect 23255 3468 23345 3472
tri 23345 3468 23349 3472 sw
tri 25206 3468 25210 3472 ne
tri 25210 3468 25304 3562 sw
rect 18705 3466 23166 3468
rect 18383 3461 23166 3466
tri 23166 3461 23173 3468 sw
tri 23255 3461 23262 3468 ne
rect 23262 3461 23349 3468
tri 23349 3461 23356 3468 sw
tri 25210 3461 25217 3468 ne
rect 25217 3461 25304 3468
tri 23079 3378 23162 3461 ne
rect 23162 3436 23173 3461
tri 23173 3436 23198 3461 sw
tri 23262 3436 23287 3461 ne
rect 23287 3436 23356 3461
rect 23162 3431 23198 3436
tri 23198 3431 23203 3436 sw
tri 23287 3431 23292 3436 ne
rect 23292 3431 23356 3436
tri 23356 3431 23386 3461 sw
tri 25217 3431 25247 3461 ne
rect 25247 3431 25304 3461
rect 23162 3378 23203 3431
tri 23203 3378 23256 3431 sw
tri 23292 3378 23345 3431 ne
rect 23345 3378 23386 3431
tri 23386 3378 23439 3431 sw
tri 25247 3378 25300 3431 ne
rect 25300 3378 25304 3431
tri 23162 3284 23256 3378 ne
tri 23256 3374 23260 3378 sw
tri 23345 3374 23349 3378 ne
rect 23349 3374 23439 3378
tri 23439 3374 23443 3378 sw
tri 25300 3374 25304 3378 ne
tri 25304 3374 25398 3468 sw
rect 23256 3346 23260 3374
tri 23260 3346 23288 3374 sw
tri 23349 3346 23377 3374 ne
rect 23377 3346 23443 3374
tri 23443 3346 23471 3374 sw
tri 25304 3346 25332 3374 ne
rect 23256 3342 23288 3346
tri 23288 3342 23292 3346 sw
tri 23377 3342 23381 3346 ne
rect 23381 3342 23471 3346
rect 23256 3337 23292 3342
tri 23292 3337 23297 3342 sw
tri 23381 3337 23386 3342 ne
rect 23386 3337 23471 3342
tri 23471 3337 23480 3346 sw
rect 23256 3284 23297 3337
tri 23297 3284 23350 3337 sw
tri 23386 3284 23439 3337 ne
rect 23439 3284 23480 3337
tri 23480 3284 23533 3337 sw
rect 3652 3177 3657 3233
rect 3713 3177 3718 3233
tri 23256 3190 23350 3284 ne
tri 23350 3248 23386 3284 sw
tri 23439 3248 23475 3284 ne
rect 23475 3248 23533 3284
rect 23350 3243 23386 3248
tri 23386 3243 23391 3248 sw
tri 23475 3243 23480 3248 ne
rect 23480 3243 23533 3248
tri 23533 3243 23574 3284 sw
rect 23350 3190 23391 3243
tri 23391 3190 23444 3243 sw
tri 23480 3190 23533 3243 ne
rect 23533 3190 23574 3243
tri 23574 3190 23627 3243 sw
tri 1691 3155 1696 3160 se
rect 1696 3155 2360 3160
tri 1636 3100 1691 3155 se
rect 1691 3100 2219 3155
rect 1636 3099 2219 3100
rect 2275 3099 2299 3155
rect 2355 3099 2360 3155
rect 1636 3094 2360 3099
rect 3652 3153 3718 3177
rect 3652 3097 3657 3153
rect 3713 3097 3718 3153
tri 23350 3141 23399 3190 ne
rect 23399 3154 23444 3190
tri 23444 3154 23480 3190 sw
tri 23533 3154 23569 3190 ne
rect 23569 3154 23627 3190
rect 23399 3149 23480 3154
tri 23480 3149 23485 3154 sw
tri 23569 3149 23574 3154 ne
rect 23574 3149 23627 3154
tri 23627 3149 23668 3190 sw
rect 23399 3141 23485 3149
tri 23485 3141 23493 3149 sw
tri 23574 3141 23582 3149 ne
rect 23582 3141 23668 3149
tri 23668 3141 23676 3149 sw
rect 1636 3087 1766 3094
tri 1766 3087 1773 3094 nw
rect 3652 3087 3718 3097
rect 5126 3136 5321 3141
rect 1636 3080 1759 3087
tri 1759 3080 1766 3087 nw
rect 5126 3080 5131 3136
rect 5187 3080 5260 3136
rect 5316 3080 5321 3136
tri 23399 3096 23444 3141 ne
rect 23444 3096 23493 3141
tri 23493 3096 23538 3141 sw
tri 23582 3096 23627 3141 ne
rect 23627 3096 23676 3141
tri 23676 3096 23721 3141 sw
tri 1542 2564 1636 2658 se
rect 1636 2630 1702 3080
tri 1702 3023 1759 3080 nw
tri 1636 2564 1702 2630 nw
tri 1490 2512 1542 2564 se
tri 1042 2507 1047 2512 se
rect 1047 2507 1252 2512
tri 986 2451 1042 2507 se
rect 1042 2451 1111 2507
rect 1167 2451 1191 2507
rect 1247 2451 1252 2507
tri 1448 2470 1490 2512 se
rect 1490 2470 1542 2512
tri 1542 2470 1636 2564 nw
tri 968 2433 986 2451 se
rect 986 2446 1252 2451
tri 1424 2446 1448 2470 se
rect 986 2433 1062 2446
tri 1062 2433 1075 2446 nw
tri 1411 2433 1424 2446 se
rect 1424 2433 1448 2446
rect 772 531 838 536
rect 772 475 777 531
rect 833 475 838 531
rect 772 451 838 475
rect 772 395 777 451
rect 833 395 838 451
rect 772 -1409 838 395
rect 968 21 1034 2433
tri 1034 2405 1062 2433 nw
tri 1383 2405 1411 2433 se
rect 1411 2405 1448 2433
tri 1354 2376 1383 2405 se
rect 1383 2376 1448 2405
tri 1448 2376 1542 2470 nw
tri 1260 2282 1354 2376 se
tri 1354 2282 1448 2376 nw
tri 1166 2188 1260 2282 se
tri 1260 2188 1354 2282 nw
tri 1112 2134 1166 2188 se
rect 1166 2134 1206 2188
tri 1206 2134 1260 2188 nw
rect 1112 1487 1178 2134
tri 1178 2106 1206 2134 nw
rect 1723 1732 1914 1741
rect 1723 1676 1728 1732
rect 1784 1676 1914 1732
rect 1723 1652 1914 1676
rect 1723 1596 1728 1652
rect 1784 1596 1914 1652
rect 1723 1585 1914 1596
tri 1723 1568 1740 1585 ne
rect 1740 1568 1914 1585
tri 1740 1524 1784 1568 ne
rect 1112 1431 1117 1487
rect 1173 1431 1178 1487
rect 1112 1407 1178 1431
rect 1112 1351 1117 1407
rect 1173 1351 1178 1407
rect 1112 1341 1178 1351
rect 1784 1152 1914 1568
tri 1914 1152 1926 1164 sw
rect 3655 1152 4056 1157
rect 1784 1096 1926 1152
tri 1926 1096 1982 1152 sw
rect 3655 1096 3660 1152
rect 3716 1096 4056 1152
rect 1784 1072 1982 1096
tri 1982 1072 2006 1096 sw
rect 3655 1072 4056 1096
rect 1784 1040 2006 1072
tri 1784 1016 1808 1040 ne
rect 1808 1016 2006 1040
tri 2006 1016 2062 1072 sw
rect 3655 1016 3660 1072
rect 3716 1032 4056 1072
rect 5126 1047 5321 3080
tri 23444 3002 23538 3096 ne
tri 23538 3060 23574 3096 sw
tri 23627 3060 23663 3096 ne
rect 23663 3060 23721 3096
rect 23538 3055 23574 3060
tri 23574 3055 23579 3060 sw
tri 23663 3055 23668 3060 ne
rect 23668 3055 23721 3060
tri 23721 3055 23762 3096 sw
rect 23538 3002 23579 3055
tri 23579 3002 23632 3055 sw
tri 23668 3002 23721 3055 ne
rect 23721 3002 23762 3055
tri 23762 3002 23815 3055 sw
tri 23538 2908 23632 3002 ne
tri 23632 2966 23668 3002 sw
tri 23721 2966 23757 3002 ne
rect 23757 2966 23815 3002
rect 23632 2961 23668 2966
tri 23668 2961 23673 2966 sw
tri 23757 2961 23762 2966 ne
rect 23762 2961 23815 2966
tri 23815 2961 23856 3002 sw
rect 23632 2908 23673 2961
tri 23673 2908 23726 2961 sw
tri 23762 2908 23815 2961 ne
rect 23815 2908 23856 2961
tri 23856 2908 23909 2961 sw
tri 23632 2814 23726 2908 ne
tri 23726 2872 23762 2908 sw
tri 23815 2872 23851 2908 ne
rect 23851 2872 23909 2908
rect 23726 2867 23762 2872
tri 23762 2867 23767 2872 sw
tri 23851 2867 23856 2872 ne
rect 23856 2867 23909 2872
tri 23909 2867 23950 2908 sw
rect 23726 2814 23767 2867
tri 23767 2814 23820 2867 sw
tri 23856 2814 23909 2867 ne
rect 23909 2814 23950 2867
tri 23950 2814 24003 2867 sw
tri 23726 2720 23820 2814 ne
tri 23820 2778 23856 2814 sw
tri 23909 2778 23945 2814 ne
rect 23945 2778 24003 2814
rect 23820 2773 23856 2778
tri 23856 2773 23861 2778 sw
tri 23945 2773 23950 2778 ne
rect 23950 2773 24003 2778
tri 24003 2773 24044 2814 sw
rect 23820 2720 23861 2773
tri 23861 2720 23914 2773 sw
tri 23950 2720 24003 2773 ne
rect 24003 2720 24044 2773
tri 24044 2720 24097 2773 sw
tri 23820 2626 23914 2720 ne
tri 23914 2684 23950 2720 sw
tri 24003 2684 24039 2720 ne
rect 24039 2684 24097 2720
rect 23914 2679 23950 2684
tri 23950 2679 23955 2684 sw
tri 24039 2679 24044 2684 ne
rect 24044 2679 24097 2684
tri 24097 2679 24138 2720 sw
rect 23914 2626 23955 2679
tri 23955 2626 24008 2679 sw
tri 24044 2651 24072 2679 ne
tri 23914 2598 23942 2626 ne
tri 18605 1865 18607 1867 se
rect 18607 1865 19026 1867
tri 18600 1860 18605 1865 se
rect 18605 1860 19026 1865
tri 18544 1804 18600 1860 se
rect 18600 1804 18873 1860
rect 18929 1804 18953 1860
rect 19009 1804 19026 1860
tri 18539 1799 18544 1804 se
rect 18544 1799 19026 1804
tri 18489 1749 18539 1799 se
rect 18539 1794 19026 1799
rect 18539 1749 18607 1794
tri 18607 1749 18652 1794 nw
tri 18444 1704 18489 1749 se
rect 18489 1704 18562 1749
tri 18562 1704 18607 1749 nw
rect 3716 1016 3733 1032
tri 1808 945 1879 1016 ne
rect 1879 961 2062 1016
tri 2062 961 2117 1016 sw
rect 3655 1011 3733 1016
tri 3733 1011 3754 1032 nw
tri 3955 1011 3976 1032 ne
rect 3976 1011 4056 1032
rect 1879 945 2117 961
tri 2117 945 2133 961 sw
tri 1879 942 1882 945 ne
rect 1882 942 2133 945
tri 2133 942 2136 945 sw
rect 1604 937 1670 942
tri 1882 937 1887 942 ne
rect 1887 937 2156 942
rect 1604 881 1609 937
rect 1665 881 1670 937
tri 1887 910 1914 937 ne
rect 1914 910 2015 937
tri 1914 881 1943 910 ne
rect 1943 881 2015 910
rect 2071 881 2095 937
rect 2151 881 2156 937
rect 1604 857 1670 881
tri 1943 876 1948 881 ne
rect 1948 876 2156 881
rect 1604 801 1609 857
rect 1665 801 1670 857
rect 1604 796 1670 801
tri 1670 796 1712 838 sw
rect 1604 718 1712 796
tri 1604 674 1648 718 ne
rect 1648 674 1712 718
tri 1712 674 1834 796 sw
tri 1648 669 1653 674 ne
rect 1653 669 2154 674
tri 1653 652 1670 669 ne
rect 1670 652 2013 669
tri 1670 546 1776 652 ne
rect 1776 546 2013 652
tri 1990 533 2003 546 ne
rect 2003 533 2013 546
rect 2149 533 2154 669
tri 2003 528 2008 533 ne
rect 2008 528 2154 533
rect 968 -43 969 21
rect 1033 -43 1034 21
rect 968 -59 1034 -43
rect 968 -123 969 -59
rect 1033 -123 1034 -59
rect 968 -129 1034 -123
rect 2058 240 2124 245
rect 2058 184 2063 240
rect 2119 184 2124 240
rect 2058 160 2124 184
rect 2058 104 2063 160
rect 2119 104 2124 160
tri 838 -1409 877 -1370 sw
rect 772 -1414 1100 -1409
rect 772 -1425 959 -1414
tri 772 -1470 817 -1425 ne
rect 817 -1470 959 -1425
rect 1015 -1470 1039 -1414
rect 1095 -1470 1100 -1414
tri 817 -1475 822 -1470 ne
rect 822 -1475 1100 -1470
rect 1031 -1850 1097 -1817
rect 1031 -1906 1036 -1850
rect 1092 -1906 1097 -1850
rect 1031 -1945 1097 -1906
rect 1031 -2001 1036 -1945
rect 1092 -2001 1097 -1945
rect 1031 -2041 1097 -2001
rect 1031 -2097 1036 -2041
rect 1092 -2097 1097 -2041
rect 2058 -1912 2124 104
rect 3655 -703 3721 1011
tri 3721 999 3733 1011 nw
tri 3976 999 3988 1011 ne
rect 3988 999 4056 1011
tri 3988 997 3990 999 ne
rect 3655 -759 3660 -703
rect 3716 -759 3721 -703
rect 3655 -783 3721 -759
rect 3655 -839 3660 -783
rect 3716 -839 3721 -783
rect 3655 -848 3721 -839
rect 3782 945 3928 950
rect 3782 889 3787 945
rect 3843 889 3867 945
rect 3923 889 3928 945
rect 3782 -888 3928 889
rect 3782 -944 3787 -888
rect 3843 -944 3867 -888
rect 3923 -944 3928 -888
rect 3782 -949 3928 -944
rect 3990 -889 4056 999
tri 18401 -277 18444 -234 se
rect 18444 -277 18523 1704
tri 18523 1665 18562 1704 nw
rect 23942 1568 24008 2626
rect 23942 1512 23947 1568
rect 24003 1512 24008 1568
rect 23942 1488 24008 1512
rect 23942 1432 23947 1488
rect 24003 1432 24008 1488
rect 23942 1427 24008 1432
tri 24022 1329 24072 1379 se
rect 24072 1329 24138 2679
rect 25332 2082 25398 3374
tri 25398 2082 25464 2148 sw
rect 25332 2077 25478 2082
rect 25332 2021 25337 2077
rect 25393 2021 25417 2077
rect 25473 2021 25478 2077
rect 25332 2016 25478 2021
rect 23946 1324 24138 1329
rect 23946 1268 23951 1324
rect 24007 1268 24031 1324
rect 24087 1268 24138 1324
rect 23946 1263 24138 1268
rect 19300 600 19306 664
rect 19370 600 19388 664
rect 19452 600 19470 664
rect 19534 600 19552 664
rect 19616 600 19634 664
rect 19698 600 19716 664
rect 19780 600 19798 664
rect 19862 600 19880 664
rect 19944 600 19962 664
rect 20026 600 20044 664
rect 20108 600 20126 664
rect 20190 600 20208 664
rect 20272 600 20290 664
rect 20354 600 20372 664
rect 20436 600 20454 664
rect 20518 600 20536 664
rect 20600 600 20618 664
rect 20682 600 20700 664
rect 20764 600 20782 664
rect 20846 600 20864 664
rect 20928 600 20946 664
rect 21010 600 21028 664
rect 21092 600 21110 664
rect 21174 600 21192 664
rect 21256 600 21274 664
rect 21338 600 21356 664
rect 21420 600 21438 664
rect 21502 600 21520 664
rect 21584 600 21601 664
rect 21665 600 21682 664
rect 21746 600 21763 664
rect 21827 600 21844 664
rect 21908 600 21925 664
rect 21989 600 22006 664
rect 22070 600 22087 664
rect 22151 600 22168 664
rect 22232 600 22249 664
rect 22313 600 22330 664
rect 22394 600 22411 664
rect 22475 600 22492 664
rect 22556 600 22573 664
rect 22637 600 22643 664
rect 19300 584 22643 600
rect 19300 520 19306 584
rect 19370 520 19388 584
rect 19452 520 19470 584
rect 19534 520 19552 584
rect 19616 520 19634 584
rect 19698 520 19716 584
rect 19780 520 19798 584
rect 19862 520 19880 584
rect 19944 520 19962 584
rect 20026 520 20044 584
rect 20108 520 20126 584
rect 20190 520 20208 584
rect 20272 520 20290 584
rect 20354 520 20372 584
rect 20436 520 20454 584
rect 20518 520 20536 584
rect 20600 520 20618 584
rect 20682 520 20700 584
rect 20764 520 20782 584
rect 20846 520 20864 584
rect 20928 520 20946 584
rect 21010 520 21028 584
rect 21092 520 21110 584
rect 21174 520 21192 584
rect 21256 520 21274 584
rect 21338 520 21356 584
rect 21420 520 21438 584
rect 21502 520 21520 584
rect 21584 520 21601 584
rect 21665 520 21682 584
rect 21746 520 21763 584
rect 21827 520 21844 584
rect 21908 520 21925 584
rect 21989 520 22006 584
rect 22070 520 22087 584
rect 22151 520 22168 584
rect 22232 520 22249 584
rect 22313 520 22330 584
rect 22394 520 22411 584
rect 22475 520 22492 584
rect 22556 520 22573 584
rect 22637 520 22643 584
rect 19300 504 22643 520
rect 19300 440 19306 504
rect 19370 440 19388 504
rect 19452 440 19470 504
rect 19534 440 19552 504
rect 19616 440 19634 504
rect 19698 440 19716 504
rect 19780 440 19798 504
rect 19862 440 19880 504
rect 19944 440 19962 504
rect 20026 440 20044 504
rect 20108 440 20126 504
rect 20190 440 20208 504
rect 20272 440 20290 504
rect 20354 440 20372 504
rect 20436 440 20454 504
rect 20518 440 20536 504
rect 20600 440 20618 504
rect 20682 440 20700 504
rect 20764 440 20782 504
rect 20846 440 20864 504
rect 20928 440 20946 504
rect 21010 440 21028 504
rect 21092 440 21110 504
rect 21174 440 21192 504
rect 21256 440 21274 504
rect 21338 440 21356 504
rect 21420 440 21438 504
rect 21502 440 21520 504
rect 21584 440 21601 504
rect 21665 440 21682 504
rect 21746 440 21763 504
rect 21827 440 21844 504
rect 21908 440 21925 504
rect 21989 440 22006 504
rect 22070 440 22087 504
rect 22151 440 22168 504
rect 22232 440 22249 504
rect 22313 440 22330 504
rect 22394 440 22411 504
rect 22475 440 22492 504
rect 22556 440 22573 504
rect 22637 440 22643 504
rect 19300 424 22643 440
rect 19300 360 19306 424
rect 19370 360 19388 424
rect 19452 360 19470 424
rect 19534 360 19552 424
rect 19616 360 19634 424
rect 19698 360 19716 424
rect 19780 360 19798 424
rect 19862 360 19880 424
rect 19944 360 19962 424
rect 20026 360 20044 424
rect 20108 360 20126 424
rect 20190 360 20208 424
rect 20272 360 20290 424
rect 20354 360 20372 424
rect 20436 360 20454 424
rect 20518 360 20536 424
rect 20600 360 20618 424
rect 20682 360 20700 424
rect 20764 360 20782 424
rect 20846 360 20864 424
rect 20928 360 20946 424
rect 21010 360 21028 424
rect 21092 360 21110 424
rect 21174 360 21192 424
rect 21256 360 21274 424
rect 21338 360 21356 424
rect 21420 360 21438 424
rect 21502 360 21520 424
rect 21584 360 21601 424
rect 21665 360 21682 424
rect 21746 360 21763 424
rect 21827 360 21844 424
rect 21908 360 21925 424
rect 21989 360 22006 424
rect 22070 360 22087 424
rect 22151 360 22168 424
rect 22232 360 22249 424
rect 22313 360 22330 424
rect 22394 360 22411 424
rect 22475 360 22492 424
rect 22556 360 22573 424
rect 22637 360 22643 424
rect 19300 344 22643 360
rect 19300 280 19306 344
rect 19370 280 19388 344
rect 19452 280 19470 344
rect 19534 280 19552 344
rect 19616 280 19634 344
rect 19698 280 19716 344
rect 19780 280 19798 344
rect 19862 280 19880 344
rect 19944 280 19962 344
rect 20026 280 20044 344
rect 20108 280 20126 344
rect 20190 280 20208 344
rect 20272 280 20290 344
rect 20354 280 20372 344
rect 20436 280 20454 344
rect 20518 280 20536 344
rect 20600 280 20618 344
rect 20682 280 20700 344
rect 20764 280 20782 344
rect 20846 280 20864 344
rect 20928 280 20946 344
rect 21010 280 21028 344
rect 21092 280 21110 344
rect 21174 280 21192 344
rect 21256 280 21274 344
rect 21338 280 21356 344
rect 21420 280 21438 344
rect 21502 280 21520 344
rect 21584 280 21601 344
rect 21665 280 21682 344
rect 21746 280 21763 344
rect 21827 280 21844 344
rect 21908 280 21925 344
rect 21989 280 22006 344
rect 22070 280 22087 344
rect 22151 280 22168 344
rect 22232 280 22249 344
rect 22313 280 22330 344
rect 22394 280 22411 344
rect 22475 280 22492 344
rect 22556 280 22573 344
rect 22637 280 22643 344
rect 19300 264 22643 280
rect 19300 200 19306 264
rect 19370 200 19388 264
rect 19452 200 19470 264
rect 19534 200 19552 264
rect 19616 200 19634 264
rect 19698 200 19716 264
rect 19780 200 19798 264
rect 19862 200 19880 264
rect 19944 200 19962 264
rect 20026 200 20044 264
rect 20108 200 20126 264
rect 20190 200 20208 264
rect 20272 200 20290 264
rect 20354 200 20372 264
rect 20436 200 20454 264
rect 20518 200 20536 264
rect 20600 200 20618 264
rect 20682 200 20700 264
rect 20764 200 20782 264
rect 20846 200 20864 264
rect 20928 200 20946 264
rect 21010 200 21028 264
rect 21092 200 21110 264
rect 21174 200 21192 264
rect 21256 200 21274 264
rect 21338 200 21356 264
rect 21420 200 21438 264
rect 21502 200 21520 264
rect 21584 200 21601 264
rect 21665 200 21682 264
rect 21746 200 21763 264
rect 21827 200 21844 264
rect 21908 200 21925 264
rect 21989 200 22006 264
rect 22070 200 22087 264
rect 22151 200 22168 264
rect 22232 200 22249 264
rect 22313 200 22330 264
rect 22394 200 22411 264
rect 22475 200 22492 264
rect 22556 200 22573 264
rect 22637 200 22643 264
rect 18377 -282 18523 -277
rect 18377 -338 18382 -282
rect 18438 -338 18462 -282
rect 18518 -338 18523 -282
rect 18377 -343 18523 -338
rect 3990 -945 3995 -889
rect 4051 -945 4056 -889
rect 3990 -969 4056 -945
rect 3990 -1025 3995 -969
rect 4051 -1025 4056 -969
rect 3990 -1030 4056 -1025
rect 21348 -1242 21941 -797
rect 2058 -1976 2059 -1912
rect 2123 -1976 2124 -1912
rect 2058 -1992 2124 -1976
rect 2058 -2056 2059 -1992
rect 2123 -2056 2124 -1992
rect 2058 -2062 2124 -2056
rect 1031 -2137 1097 -2097
rect 1031 -2193 1036 -2137
rect 1092 -2193 1097 -2137
rect 1031 -5455 1097 -2193
rect 1724 -4234 1905 -4229
rect 1724 -4290 1729 -4234
rect 1785 -4290 1844 -4234
rect 1900 -4290 1905 -4234
rect 1724 -4356 1905 -4290
rect 1724 -4412 1729 -4356
rect 1785 -4412 1844 -4356
rect 1900 -4412 1905 -4356
rect 1724 -4417 1905 -4412
rect 1031 -5511 1036 -5455
rect 1092 -5511 1097 -5455
rect 1031 -5535 1097 -5511
rect 1031 -5591 1036 -5535
rect 1092 -5591 1097 -5535
rect 1031 -5596 1097 -5591
rect 1036 -5932 1100 -5926
rect 1035 -5996 1036 -5936
rect 1100 -5996 1101 -5936
rect 1035 -5997 1040 -5996
rect 1096 -5997 1101 -5996
rect 1035 -6012 1101 -5997
rect 1035 -6076 1036 -6012
rect 1100 -6076 1101 -6012
rect 1035 -6077 1040 -6076
rect 1096 -6077 1101 -6076
rect 1035 -6082 1101 -6077
rect 2605 -9593 2669 -9587
rect 2669 -9657 2671 -9597
rect 2605 -9658 2610 -9657
rect 2666 -9658 2671 -9657
rect 2605 -9673 2671 -9658
rect 2669 -9737 2671 -9673
rect 2605 -9738 2610 -9737
rect 2666 -9738 2671 -9737
rect 2605 -9743 2671 -9738
rect 2645 -10221 2791 -10216
rect 2645 -10277 2650 -10221
rect 2706 -10277 2730 -10221
rect 2786 -10277 2791 -10221
rect 2645 -10282 2791 -10277
<< via3 >>
rect 14584 3758 14648 3822
rect 14728 3763 14792 3822
rect 14871 3763 14935 3822
rect 15014 3763 15078 3822
rect 15157 3763 15221 3822
rect 14728 3758 14762 3763
rect 14762 3758 14792 3763
rect 14871 3758 14883 3763
rect 14883 3758 14935 3763
rect 15014 3758 15068 3763
rect 15068 3758 15078 3763
rect 15157 3758 15188 3763
rect 15188 3758 15221 3763
rect 15300 3758 15364 3822
rect 14584 3622 14648 3686
rect 14728 3663 14792 3686
rect 14871 3663 14935 3686
rect 15014 3663 15078 3686
rect 15157 3663 15221 3686
rect 14728 3622 14762 3663
rect 14762 3622 14792 3663
rect 14871 3622 14883 3663
rect 14883 3622 14935 3663
rect 15014 3622 15068 3663
rect 15068 3622 15078 3663
rect 15157 3622 15188 3663
rect 15188 3622 15221 3663
rect 15300 3622 15364 3686
rect 14584 3486 14648 3550
rect 14728 3507 14762 3550
rect 14762 3507 14792 3550
rect 14871 3507 14883 3550
rect 14883 3507 14935 3550
rect 15014 3507 15068 3550
rect 15068 3507 15078 3550
rect 15157 3507 15188 3550
rect 15188 3507 15221 3550
rect 14728 3486 14792 3507
rect 14871 3486 14935 3507
rect 15014 3486 15078 3507
rect 15157 3486 15221 3507
rect 15300 3486 15364 3550
rect 969 -43 1033 21
rect 969 -123 1033 -59
rect 19306 600 19370 664
rect 19388 600 19452 664
rect 19470 600 19534 664
rect 19552 600 19616 664
rect 19634 600 19698 664
rect 19716 600 19780 664
rect 19798 600 19862 664
rect 19880 600 19944 664
rect 19962 600 20026 664
rect 20044 600 20108 664
rect 20126 600 20190 664
rect 20208 600 20272 664
rect 20290 600 20354 664
rect 20372 600 20436 664
rect 20454 600 20518 664
rect 20536 600 20600 664
rect 20618 600 20682 664
rect 20700 600 20764 664
rect 20782 600 20846 664
rect 20864 600 20928 664
rect 20946 600 21010 664
rect 21028 600 21092 664
rect 21110 600 21174 664
rect 21192 600 21256 664
rect 21274 600 21338 664
rect 21356 600 21420 664
rect 21438 600 21502 664
rect 21520 600 21584 664
rect 21601 600 21665 664
rect 21682 600 21746 664
rect 21763 600 21827 664
rect 21844 600 21908 664
rect 21925 600 21989 664
rect 22006 600 22070 664
rect 22087 600 22151 664
rect 22168 600 22232 664
rect 22249 600 22313 664
rect 22330 600 22394 664
rect 22411 600 22475 664
rect 22492 600 22556 664
rect 22573 600 22637 664
rect 19306 520 19370 584
rect 19388 520 19452 584
rect 19470 520 19534 584
rect 19552 520 19616 584
rect 19634 520 19698 584
rect 19716 520 19780 584
rect 19798 520 19862 584
rect 19880 520 19944 584
rect 19962 520 20026 584
rect 20044 520 20108 584
rect 20126 520 20190 584
rect 20208 520 20272 584
rect 20290 520 20354 584
rect 20372 520 20436 584
rect 20454 520 20518 584
rect 20536 520 20600 584
rect 20618 520 20682 584
rect 20700 520 20764 584
rect 20782 520 20846 584
rect 20864 520 20928 584
rect 20946 520 21010 584
rect 21028 520 21092 584
rect 21110 520 21174 584
rect 21192 520 21256 584
rect 21274 520 21338 584
rect 21356 520 21420 584
rect 21438 520 21502 584
rect 21520 520 21584 584
rect 21601 520 21665 584
rect 21682 520 21746 584
rect 21763 520 21827 584
rect 21844 520 21908 584
rect 21925 520 21989 584
rect 22006 520 22070 584
rect 22087 520 22151 584
rect 22168 520 22232 584
rect 22249 520 22313 584
rect 22330 520 22394 584
rect 22411 520 22475 584
rect 22492 520 22556 584
rect 22573 520 22637 584
rect 19306 440 19370 504
rect 19388 440 19452 504
rect 19470 440 19534 504
rect 19552 440 19616 504
rect 19634 440 19698 504
rect 19716 440 19780 504
rect 19798 440 19862 504
rect 19880 440 19944 504
rect 19962 440 20026 504
rect 20044 440 20108 504
rect 20126 440 20190 504
rect 20208 440 20272 504
rect 20290 440 20354 504
rect 20372 440 20436 504
rect 20454 440 20518 504
rect 20536 440 20600 504
rect 20618 440 20682 504
rect 20700 440 20764 504
rect 20782 440 20846 504
rect 20864 440 20928 504
rect 20946 440 21010 504
rect 21028 440 21092 504
rect 21110 440 21174 504
rect 21192 440 21256 504
rect 21274 440 21338 504
rect 21356 440 21420 504
rect 21438 440 21502 504
rect 21520 440 21584 504
rect 21601 440 21665 504
rect 21682 440 21746 504
rect 21763 440 21827 504
rect 21844 440 21908 504
rect 21925 440 21989 504
rect 22006 440 22070 504
rect 22087 440 22151 504
rect 22168 440 22232 504
rect 22249 440 22313 504
rect 22330 440 22394 504
rect 22411 440 22475 504
rect 22492 440 22556 504
rect 22573 440 22637 504
rect 19306 360 19370 424
rect 19388 360 19452 424
rect 19470 360 19534 424
rect 19552 360 19616 424
rect 19634 360 19698 424
rect 19716 360 19780 424
rect 19798 360 19862 424
rect 19880 360 19944 424
rect 19962 360 20026 424
rect 20044 360 20108 424
rect 20126 360 20190 424
rect 20208 360 20272 424
rect 20290 360 20354 424
rect 20372 360 20436 424
rect 20454 360 20518 424
rect 20536 360 20600 424
rect 20618 360 20682 424
rect 20700 360 20764 424
rect 20782 360 20846 424
rect 20864 360 20928 424
rect 20946 360 21010 424
rect 21028 360 21092 424
rect 21110 360 21174 424
rect 21192 360 21256 424
rect 21274 360 21338 424
rect 21356 360 21420 424
rect 21438 360 21502 424
rect 21520 360 21584 424
rect 21601 360 21665 424
rect 21682 360 21746 424
rect 21763 360 21827 424
rect 21844 360 21908 424
rect 21925 360 21989 424
rect 22006 360 22070 424
rect 22087 360 22151 424
rect 22168 360 22232 424
rect 22249 360 22313 424
rect 22330 360 22394 424
rect 22411 360 22475 424
rect 22492 360 22556 424
rect 22573 360 22637 424
rect 19306 280 19370 344
rect 19388 280 19452 344
rect 19470 280 19534 344
rect 19552 280 19616 344
rect 19634 280 19698 344
rect 19716 280 19780 344
rect 19798 280 19862 344
rect 19880 280 19944 344
rect 19962 280 20026 344
rect 20044 280 20108 344
rect 20126 280 20190 344
rect 20208 280 20272 344
rect 20290 280 20354 344
rect 20372 280 20436 344
rect 20454 280 20518 344
rect 20536 280 20600 344
rect 20618 280 20682 344
rect 20700 280 20764 344
rect 20782 280 20846 344
rect 20864 280 20928 344
rect 20946 280 21010 344
rect 21028 280 21092 344
rect 21110 280 21174 344
rect 21192 280 21256 344
rect 21274 280 21338 344
rect 21356 280 21420 344
rect 21438 280 21502 344
rect 21520 280 21584 344
rect 21601 280 21665 344
rect 21682 280 21746 344
rect 21763 280 21827 344
rect 21844 280 21908 344
rect 21925 280 21989 344
rect 22006 280 22070 344
rect 22087 280 22151 344
rect 22168 280 22232 344
rect 22249 280 22313 344
rect 22330 280 22394 344
rect 22411 280 22475 344
rect 22492 280 22556 344
rect 22573 280 22637 344
rect 19306 200 19370 264
rect 19388 200 19452 264
rect 19470 200 19534 264
rect 19552 200 19616 264
rect 19634 200 19698 264
rect 19716 200 19780 264
rect 19798 200 19862 264
rect 19880 200 19944 264
rect 19962 200 20026 264
rect 20044 200 20108 264
rect 20126 200 20190 264
rect 20208 200 20272 264
rect 20290 200 20354 264
rect 20372 200 20436 264
rect 20454 200 20518 264
rect 20536 200 20600 264
rect 20618 200 20682 264
rect 20700 200 20764 264
rect 20782 200 20846 264
rect 20864 200 20928 264
rect 20946 200 21010 264
rect 21028 200 21092 264
rect 21110 200 21174 264
rect 21192 200 21256 264
rect 21274 200 21338 264
rect 21356 200 21420 264
rect 21438 200 21502 264
rect 21520 200 21584 264
rect 21601 200 21665 264
rect 21682 200 21746 264
rect 21763 200 21827 264
rect 21844 200 21908 264
rect 21925 200 21989 264
rect 22006 200 22070 264
rect 22087 200 22151 264
rect 22168 200 22232 264
rect 22249 200 22313 264
rect 22330 200 22394 264
rect 22411 200 22475 264
rect 22492 200 22556 264
rect 22573 200 22637 264
rect 2059 -1976 2123 -1912
rect 2059 -2056 2123 -1992
rect 1036 -5941 1100 -5932
rect 1036 -5996 1040 -5941
rect 1040 -5996 1096 -5941
rect 1096 -5996 1100 -5941
rect 1036 -6021 1100 -6012
rect 1036 -6076 1040 -6021
rect 1040 -6076 1096 -6021
rect 1096 -6076 1100 -6021
rect 2605 -9602 2669 -9593
rect 2605 -9657 2610 -9602
rect 2610 -9657 2666 -9602
rect 2666 -9657 2669 -9602
rect 2605 -9682 2669 -9673
rect 2605 -9737 2610 -9682
rect 2610 -9737 2666 -9682
rect 2666 -9737 2669 -9682
<< metal4 >>
rect 14583 3822 15365 3823
rect 14583 3758 14584 3822
rect 14648 3758 14728 3822
rect 14792 3758 14871 3822
rect 14935 3758 15014 3822
rect 15078 3758 15157 3822
rect 15221 3758 15300 3822
rect 15364 3758 15365 3822
rect 14583 3686 15365 3758
rect 14583 3622 14584 3686
rect 14648 3622 14728 3686
rect 14792 3622 14871 3686
rect 14935 3622 15014 3686
rect 15078 3622 15157 3686
rect 15221 3622 15300 3686
rect 15364 3622 15365 3686
rect 14583 3550 15365 3622
rect 14583 3486 14584 3550
rect 14648 3486 14728 3550
rect 14792 3486 14871 3550
rect 14935 3486 15014 3550
rect 15078 3486 15157 3550
rect 15221 3486 15300 3550
rect 15364 3486 15365 3550
rect 14583 3485 15365 3486
rect 19305 664 22638 665
rect 19305 600 19306 664
rect 19370 600 19388 664
rect 19452 600 19470 664
rect 19534 600 19552 664
rect 19616 600 19634 664
rect 19698 600 19716 664
rect 19780 600 19798 664
rect 19862 600 19880 664
rect 19944 600 19962 664
rect 20026 600 20044 664
rect 20108 600 20126 664
rect 20190 600 20208 664
rect 20272 600 20290 664
rect 20354 600 20372 664
rect 20436 600 20454 664
rect 20518 600 20536 664
rect 20600 600 20618 664
rect 20682 600 20700 664
rect 20764 600 20782 664
rect 20846 600 20864 664
rect 20928 600 20946 664
rect 21010 600 21028 664
rect 21092 600 21110 664
rect 21174 600 21192 664
rect 21256 600 21274 664
rect 21338 600 21356 664
rect 21420 600 21438 664
rect 21502 600 21520 664
rect 21584 600 21601 664
rect 21665 600 21682 664
rect 21746 600 21763 664
rect 21827 600 21844 664
rect 21908 600 21925 664
rect 21989 600 22006 664
rect 22070 600 22087 664
rect 22151 600 22168 664
rect 22232 600 22249 664
rect 22313 600 22330 664
rect 22394 600 22411 664
rect 22475 600 22492 664
rect 22556 600 22573 664
rect 22637 600 22638 664
rect 19305 584 22638 600
rect 19305 520 19306 584
rect 19370 520 19388 584
rect 19452 520 19470 584
rect 19534 520 19552 584
rect 19616 520 19634 584
rect 19698 520 19716 584
rect 19780 520 19798 584
rect 19862 520 19880 584
rect 19944 520 19962 584
rect 20026 520 20044 584
rect 20108 520 20126 584
rect 20190 520 20208 584
rect 20272 520 20290 584
rect 20354 520 20372 584
rect 20436 520 20454 584
rect 20518 520 20536 584
rect 20600 520 20618 584
rect 20682 520 20700 584
rect 20764 520 20782 584
rect 20846 520 20864 584
rect 20928 520 20946 584
rect 21010 520 21028 584
rect 21092 520 21110 584
rect 21174 520 21192 584
rect 21256 520 21274 584
rect 21338 520 21356 584
rect 21420 520 21438 584
rect 21502 520 21520 584
rect 21584 520 21601 584
rect 21665 520 21682 584
rect 21746 520 21763 584
rect 21827 520 21844 584
rect 21908 520 21925 584
rect 21989 520 22006 584
rect 22070 520 22087 584
rect 22151 520 22168 584
rect 22232 520 22249 584
rect 22313 520 22330 584
rect 22394 520 22411 584
rect 22475 520 22492 584
rect 22556 520 22573 584
rect 22637 520 22638 584
rect 19305 504 22638 520
rect 19305 440 19306 504
rect 19370 440 19388 504
rect 19452 440 19470 504
rect 19534 440 19552 504
rect 19616 440 19634 504
rect 19698 440 19716 504
rect 19780 440 19798 504
rect 19862 440 19880 504
rect 19944 440 19962 504
rect 20026 440 20044 504
rect 20108 440 20126 504
rect 20190 440 20208 504
rect 20272 440 20290 504
rect 20354 440 20372 504
rect 20436 440 20454 504
rect 20518 440 20536 504
rect 20600 440 20618 504
rect 20682 440 20700 504
rect 20764 440 20782 504
rect 20846 440 20864 504
rect 20928 440 20946 504
rect 21010 440 21028 504
rect 21092 440 21110 504
rect 21174 440 21192 504
rect 21256 440 21274 504
rect 21338 440 21356 504
rect 21420 440 21438 504
rect 21502 440 21520 504
rect 21584 440 21601 504
rect 21665 440 21682 504
rect 21746 440 21763 504
rect 21827 440 21844 504
rect 21908 440 21925 504
rect 21989 440 22006 504
rect 22070 440 22087 504
rect 22151 440 22168 504
rect 22232 440 22249 504
rect 22313 440 22330 504
rect 22394 440 22411 504
rect 22475 440 22492 504
rect 22556 440 22573 504
rect 22637 440 22638 504
rect 19305 424 22638 440
rect 19305 360 19306 424
rect 19370 360 19388 424
rect 19452 360 19470 424
rect 19534 360 19552 424
rect 19616 360 19634 424
rect 19698 360 19716 424
rect 19780 360 19798 424
rect 19862 360 19880 424
rect 19944 360 19962 424
rect 20026 360 20044 424
rect 20108 360 20126 424
rect 20190 360 20208 424
rect 20272 360 20290 424
rect 20354 360 20372 424
rect 20436 360 20454 424
rect 20518 360 20536 424
rect 20600 360 20618 424
rect 20682 360 20700 424
rect 20764 360 20782 424
rect 20846 360 20864 424
rect 20928 360 20946 424
rect 21010 360 21028 424
rect 21092 360 21110 424
rect 21174 360 21192 424
rect 21256 360 21274 424
rect 21338 360 21356 424
rect 21420 360 21438 424
rect 21502 360 21520 424
rect 21584 360 21601 424
rect 21665 360 21682 424
rect 21746 360 21763 424
rect 21827 360 21844 424
rect 21908 360 21925 424
rect 21989 360 22006 424
rect 22070 360 22087 424
rect 22151 360 22168 424
rect 22232 360 22249 424
rect 22313 360 22330 424
rect 22394 360 22411 424
rect 22475 360 22492 424
rect 22556 360 22573 424
rect 22637 360 22638 424
rect 19305 344 22638 360
rect 19305 280 19306 344
rect 19370 280 19388 344
rect 19452 280 19470 344
rect 19534 280 19552 344
rect 19616 280 19634 344
rect 19698 280 19716 344
rect 19780 280 19798 344
rect 19862 280 19880 344
rect 19944 280 19962 344
rect 20026 280 20044 344
rect 20108 280 20126 344
rect 20190 280 20208 344
rect 20272 280 20290 344
rect 20354 280 20372 344
rect 20436 280 20454 344
rect 20518 280 20536 344
rect 20600 280 20618 344
rect 20682 280 20700 344
rect 20764 280 20782 344
rect 20846 280 20864 344
rect 20928 280 20946 344
rect 21010 280 21028 344
rect 21092 280 21110 344
rect 21174 280 21192 344
rect 21256 280 21274 344
rect 21338 280 21356 344
rect 21420 280 21438 344
rect 21502 280 21520 344
rect 21584 280 21601 344
rect 21665 280 21682 344
rect 21746 280 21763 344
rect 21827 280 21844 344
rect 21908 280 21925 344
rect 21989 280 22006 344
rect 22070 280 22087 344
rect 22151 280 22168 344
rect 22232 280 22249 344
rect 22313 280 22330 344
rect 22394 280 22411 344
rect 22475 280 22492 344
rect 22556 280 22573 344
rect 22637 280 22638 344
rect 19305 264 22638 280
rect 19305 200 19306 264
rect 19370 200 19388 264
rect 19452 200 19470 264
rect 19534 200 19552 264
rect 19616 200 19634 264
rect 19698 200 19716 264
rect 19780 200 19798 264
rect 19862 200 19880 264
rect 19944 200 19962 264
rect 20026 200 20044 264
rect 20108 200 20126 264
rect 20190 200 20208 264
rect 20272 200 20290 264
rect 20354 200 20372 264
rect 20436 200 20454 264
rect 20518 200 20536 264
rect 20600 200 20618 264
rect 20682 200 20700 264
rect 20764 200 20782 264
rect 20846 200 20864 264
rect 20928 200 20946 264
rect 21010 200 21028 264
rect 21092 200 21110 264
rect 21174 200 21192 264
rect 21256 200 21274 264
rect 21338 200 21356 264
rect 21420 200 21438 264
rect 21502 200 21520 264
rect 21584 200 21601 264
rect 21665 200 21682 264
rect 21746 200 21763 264
rect 21827 200 21844 264
rect 21908 200 21925 264
rect 21989 200 22006 264
rect 22070 200 22087 264
rect 22151 200 22168 264
rect 22232 200 22249 264
rect 22313 200 22330 264
rect 22394 200 22411 264
rect 22475 200 22492 264
rect 22556 200 22573 264
rect 22637 200 22638 264
rect 19305 199 22638 200
rect 968 21 1034 22
rect 968 -43 969 21
rect 1033 -43 1034 21
rect 968 -44 1034 -43
tri 1034 -44 1100 22 sw
rect 968 -55 2377 -44
tri 2377 -55 2388 -44 sw
rect 968 -59 2388 -55
rect 968 -123 969 -59
rect 1033 -123 2388 -59
rect 968 -124 2388 -123
tri 2388 -124 2457 -55 sw
tri 2343 -169 2388 -124 ne
rect 2388 -169 2457 -124
tri 2457 -169 2502 -124 sw
tri 2388 -283 2502 -169 ne
tri 2502 -283 2616 -169 sw
tri 2502 -317 2536 -283 ne
rect 2058 -1912 2124 -1911
rect 2058 -1976 2059 -1912
rect 2123 -1976 2124 -1912
rect 2058 -1992 2124 -1976
rect 2058 -2056 2059 -1992
rect 2123 -2056 2124 -1992
tri 1994 -5931 2058 -5867 se
rect 2058 -5895 2124 -2056
rect 2058 -5931 2088 -5895
tri 2088 -5931 2124 -5895 nw
rect 1035 -5932 2022 -5931
rect 1035 -5996 1036 -5932
rect 1100 -5996 2022 -5932
rect 1035 -5997 2022 -5996
tri 2022 -5997 2088 -5931 nw
rect 1035 -6012 1101 -5997
rect 1035 -6076 1036 -6012
rect 1100 -6076 1101 -6012
rect 1035 -6077 1101 -6076
rect 2536 -9592 2616 -283
tri 2616 -9592 2670 -9538 sw
rect 2536 -9593 2670 -9592
rect 2536 -9657 2605 -9593
rect 2669 -9657 2670 -9593
rect 2536 -9673 2670 -9657
rect 2536 -9737 2605 -9673
rect 2669 -9737 2670 -9673
rect 2536 -9747 2670 -9737
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_0
timestamp 1694700623
transform 0 -1 25729 1 0 1574
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_1
timestamp 1694700623
transform 1 0 18855 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2_1  sky130_fd_io__com_inv_x1_dnwv2_1_0
timestamp 1694700623
transform 1 0 17503 0 1 1972
box 825 -1510 2624 1229
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_2
timestamp 1694700623
transform -1 0 13096 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_3
timestamp 1694700623
transform -1 0 16993 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_4
timestamp 1694700623
transform 1 0 16895 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_5
timestamp 1694700623
transform 1 0 19509 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_6
timestamp 1694700623
transform -1 0 13777 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_7
timestamp 1694700623
transform -1 0 15385 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_8
timestamp 1694700623
transform -1 0 17945 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_9
timestamp 1694700623
transform -1 0 16189 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_10
timestamp 1694700623
transform -1 0 14581 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_inv_x1_dnwv2  sky130_fd_io__com_inv_x1_dnwv2_11
timestamp 1694700623
transform 1 0 12522 0 1 3686
box -47 -115 316 1292
use sky130_fd_io__com_nand2_dnwv2  sky130_fd_io__com_nand2_dnwv2_0
timestamp 1694700623
transform 1 0 19166 0 1 3783
box -57 -212 483 1195
use sky130_fd_io__com_nand2_dnwv2  sky130_fd_io__com_nand2_dnwv2_1
timestamp 1694700623
transform -1 0 17636 0 1 3783
box -57 -212 483 1195
use sky130_fd_io__com_nand2_dnwv2  sky130_fd_io__com_nand2_dnwv2_2
timestamp 1694700623
transform 1 0 12179 0 1 3783
box -57 -212 483 1195
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_0
timestamp 1694700623
transform 0 -1 25713 -1 0 1943
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2_1  sky130_fd_io__com_nor2_dnwv2_1_0
timestamp 1694700623
transform 1 0 16626 0 1 2029
box 468 -1391 3211 1172
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_1
timestamp 1694700623
transform 1 0 12727 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_2
timestamp 1694700623
transform -1 0 16964 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_3
timestamp 1694700623
transform -1 0 16160 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_4
timestamp 1694700623
transform -1 0 18720 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_5
timestamp 1694700623
transform -1 0 14552 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_6
timestamp 1694700623
transform -1 0 15356 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__com_nor2_dnwv2  sky130_fd_io__com_nor2_dnwv2_7
timestamp 1694700623
transform 1 0 18080 0 1 3702
box 229 -131 791 1276
use sky130_fd_io__nor3_dnw  sky130_fd_io__nor3_dnw_0
timestamp 1694700623
transform 1 0 11395 0 1 3702
box 25 -131 791 1276
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_0
timestamp 1694700623
transform -1 0 22655 0 1 -717
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_1
timestamp 1694700623
transform 1 0 19289 0 1 -717
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_2
timestamp 1694700623
transform -1 0 22655 0 1 -6725
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_3
timestamp 1694700623
transform 1 0 19289 0 1 -6725
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_4
timestamp 1694700623
transform -1 0 22655 0 -1 -3655
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_5
timestamp 1694700623
transform 1 0 19289 0 -1 -3655
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_6
timestamp 1694700623
transform -1 0 22655 0 1 -3721
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_7
timestamp 1694700623
transform 1 0 19289 0 1 -3721
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_8
timestamp 1694700623
transform 1 0 19289 0 -1 -651
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_9
timestamp 1694700623
transform -1 0 22655 0 -1 -651
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_10
timestamp 1694700623
transform -1 0 22655 0 1 -9729
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_11
timestamp 1694700623
transform 1 0 19289 0 1 -9729
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_12
timestamp 1694700623
transform 1 0 19289 0 -1 -6659
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_13
timestamp 1694700623
transform -1 0 22655 0 1 -12733
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_14
timestamp 1694700623
transform -1 0 22655 0 -1 -6659
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_15
timestamp 1694700623
transform 1 0 19289 0 -1 -9663
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_16
timestamp 1694700623
transform 1 0 19289 0 1 -12733
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3_17
timestamp 1694700623
transform -1 0 22655 0 -1 -9663
box 0 0 1716 1568
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_0
timestamp 1694700623
transform 1 0 6874 0 -1 1954
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808230  sky130_fd_pr__nfet_01v8__example_55959141808230_0
timestamp 1694700623
transform 1 0 2669 0 1 -10184
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808231  sky130_fd_pr__nfet_01v8__example_55959141808231_0
timestamp 1694700623
transform 1 0 12828 0 1 748
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808232  sky130_fd_pr__nfet_01v8__example_55959141808232_0
timestamp 1694700623
transform 0 1 7503 1 0 2092
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808234  sky130_fd_pr__nfet_01v8__example_55959141808234_0
timestamp 1694700623
transform 0 -1 18596 1 0 37
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808235  sky130_fd_pr__nfet_01v8__example_55959141808235_0
timestamp 1694700623
transform 1 0 5071 0 1 16
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808235  sky130_fd_pr__nfet_01v8__example_55959141808235_1
timestamp 1694700623
transform 1 0 4603 0 1 16
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808236  sky130_fd_pr__nfet_01v8__example_55959141808236_0
timestamp 1694700623
transform 0 -1 6662 1 0 1204
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808238  sky130_fd_pr__nfet_01v8__example_55959141808238_0
timestamp 1694700623
transform 0 -1 6662 -1 0 2092
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808239  sky130_fd_pr__nfet_01v8__example_55959141808239_0
timestamp 1694700623
transform -1 0 8897 0 1 -52
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808241  sky130_fd_pr__nfet_01v8__example_55959141808241_0
timestamp 1694700623
transform 1 0 15268 0 -1 294
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808244  sky130_fd_pr__nfet_01v8__example_55959141808244_0
timestamp 1694700623
transform 1 0 15268 0 1 479
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808244  sky130_fd_pr__nfet_01v8__example_55959141808244_1
timestamp 1694700623
transform 1 0 15268 0 -1 1034
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808245  sky130_fd_pr__nfet_01v8__example_55959141808245_0
timestamp 1694700623
transform -1 0 12550 0 1 -52
box -1 0 1769 1
use sky130_fd_pr__nfet_01v8__example_55959141808246  sky130_fd_pr__nfet_01v8__example_55959141808246_0
timestamp 1694700623
transform -1 0 9677 0 1 -52
box -1 0 725 1
use sky130_fd_pr__nfet_01v8__example_55959141808246  sky130_fd_pr__nfet_01v8__example_55959141808246_1
timestamp 1694700623
transform -1 0 10457 0 1 -52
box -1 0 725 1
use sky130_fd_pr__nfet_01v8__example_55959141808247  sky130_fd_pr__nfet_01v8__example_55959141808247_0
timestamp 1694700623
transform 0 1 13076 -1 0 1024
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808247  sky130_fd_pr__nfet_01v8__example_55959141808247_1
timestamp 1694700623
transform 0 1 2424 1 0 1204
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1694700623
transform 1 0 4447 0 1 16
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808249  sky130_fd_pr__nfet_01v8__example_55959141808249_0
timestamp 1694700623
transform 1 0 7469 0 1 -9
box -1 0 375 1
use sky130_fd_pr__nfet_01v8__example_55959141808252  sky130_fd_pr__nfet_01v8__example_55959141808252_0
timestamp 1694700623
transform 1 0 6741 0 1 16
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808252  sky130_fd_pr__nfet_01v8__example_55959141808252_1
timestamp 1694700623
transform 1 0 15929 0 1 -823
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808252  sky130_fd_pr__nfet_01v8__example_55959141808252_2
timestamp 1694700623
transform 1 0 3823 0 1 16
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808252  sky130_fd_pr__nfet_01v8__example_55959141808252_3
timestamp 1694700623
transform 1 0 4135 0 1 16
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808253  sky130_fd_pr__nfet_01v8__example_55959141808253_0
timestamp 1694700623
transform 1 0 3075 0 1 16
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808254  sky130_fd_pr__nfet_01v8__example_55959141808254_0
timestamp 1694700623
transform 1 0 2451 0 1 16
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808255  sky130_fd_pr__nfet_01v8__example_55959141808255_0
timestamp 1694700623
transform 1 0 5713 0 1 16
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808256  sky130_fd_pr__nfet_01v8__example_55959141808256_0
timestamp 1694700623
transform -1 0 6125 0 1 16
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808256  sky130_fd_pr__nfet_01v8__example_55959141808256_1
timestamp 1694700623
transform 1 0 6461 0 1 16
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808256  sky130_fd_pr__nfet_01v8__example_55959141808256_2
timestamp 1694700623
transform -1 0 6281 0 1 16
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808257  sky130_fd_pr__nfet_01v8__example_55959141808257_0
timestamp 1694700623
transform -1 0 8474 0 1 1656
box -1 0 1601 1
use sky130_fd_pr__pfet_01v8__example_5595914180813  sky130_fd_pr__pfet_01v8__example_5595914180813_0
timestamp 1694700623
transform 0 -1 17571 1 0 3064
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1694700623
transform 1 0 3068 0 -1 -17100
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_0
timestamp 1694700623
transform 1 0 2625 0 1 -18915
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808192  sky130_fd_pr__pfet_01v8__example_55959141808192_0
timestamp 1694700623
transform 1 0 10624 0 1 3477
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808193  sky130_fd_pr__pfet_01v8__example_55959141808193_0
timestamp 1694700623
transform 0 -1 19086 1 0 2738
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808195  sky130_fd_pr__pfet_01v8__example_55959141808195_0
timestamp 1694700623
transform -1 0 18889 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808195  sky130_fd_pr__pfet_01v8__example_55959141808195_1
timestamp 1694700623
transform -1 0 17943 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808195  sky130_fd_pr__pfet_01v8__example_55959141808195_2
timestamp 1694700623
transform 1 0 17999 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808195  sky130_fd_pr__pfet_01v8__example_55959141808195_3
timestamp 1694700623
transform 1 0 18945 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808196  sky130_fd_pr__pfet_01v8__example_55959141808196_0
timestamp 1694700623
transform 0 1 574 1 0 -1959
box -1 0 881 1
use sky130_fd_pr__pfet_01v8__example_55959141808198  sky130_fd_pr__pfet_01v8__example_55959141808198_0
timestamp 1694700623
transform 0 1 574 1 0 -738
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808199  sky130_fd_pr__pfet_01v8__example_55959141808199_0
timestamp 1694700623
transform -1 0 18427 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808199  sky130_fd_pr__pfet_01v8__example_55959141808199_1
timestamp 1694700623
transform 1 0 18483 0 1 3034
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808201  sky130_fd_pr__pfet_01v8__example_55959141808201_0
timestamp 1694700623
transform 0 1 574 1 0 -2271
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808203  sky130_fd_pr__pfet_01v8__example_55959141808203_0
timestamp 1694700623
transform 0 1 574 1 0 822
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808203  sky130_fd_pr__pfet_01v8__example_55959141808203_1
timestamp 1694700623
transform 0 1 574 1 0 -114
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808203  sky130_fd_pr__pfet_01v8__example_55959141808203_2
timestamp 1694700623
transform 0 1 574 1 0 -582
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808203  sky130_fd_pr__pfet_01v8__example_55959141808203_3
timestamp 1694700623
transform 0 1 574 1 0 354
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808204  sky130_fd_pr__pfet_01v8__example_55959141808204_0
timestamp 1694700623
transform 0 1 574 1 0 42
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808204  sky130_fd_pr__pfet_01v8__example_55959141808204_1
timestamp 1694700623
transform 0 1 574 1 0 978
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808204  sky130_fd_pr__pfet_01v8__example_55959141808204_2
timestamp 1694700623
transform 0 1 574 1 0 510
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808204  sky130_fd_pr__pfet_01v8__example_55959141808204_3
timestamp 1694700623
transform 0 1 574 1 0 -426
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808205  sky130_fd_pr__pfet_01v8__example_55959141808205_0
timestamp 1694700623
transform 0 -1 11152 1 0 3225
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_0
timestamp 1694700623
transform 1 0 6892 0 -1 3809
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_1
timestamp 1694700623
transform 1 0 6892 0 1 3281
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_2
timestamp 1694700623
transform 1 0 6892 0 1 4291
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_3
timestamp 1694700623
transform 1 0 6892 0 -1 4819
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_4
timestamp 1694700623
transform -1 0 1716 0 -1 4819
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_5
timestamp 1694700623
transform -1 0 1716 0 -1 3809
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_6
timestamp 1694700623
transform -1 0 1716 0 1 3281
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808206  sky130_fd_pr__pfet_01v8__example_55959141808206_7
timestamp 1694700623
transform -1 0 1716 0 1 4291
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_0
timestamp 1694700623
transform 1 0 6636 0 -1 3809
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_1
timestamp 1694700623
transform 1 0 6636 0 1 3281
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_2
timestamp 1694700623
transform 1 0 6636 0 1 4291
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_3
timestamp 1694700623
transform 1 0 6636 0 -1 4819
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_4
timestamp 1694700623
transform -1 0 1972 0 -1 4819
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_5
timestamp 1694700623
transform -1 0 1972 0 -1 3809
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_6
timestamp 1694700623
transform -1 0 1972 0 1 3281
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_7
timestamp 1694700623
transform -1 0 2228 0 -1 4819
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_8
timestamp 1694700623
transform -1 0 2228 0 1 4291
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_9
timestamp 1694700623
transform -1 0 1972 0 1 4291
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_10
timestamp 1694700623
transform -1 0 2228 0 -1 3809
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808208  sky130_fd_pr__pfet_01v8__example_55959141808208_11
timestamp 1694700623
transform -1 0 2228 0 1 3281
box -1 0 201 1
use sky130_fd_pr__pfet_01v8__example_55959141808209  sky130_fd_pr__pfet_01v8__example_55959141808209_0
timestamp 1694700623
transform -1 0 6580 0 -1 3809
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808209  sky130_fd_pr__pfet_01v8__example_55959141808209_1
timestamp 1694700623
transform -1 0 6580 0 1 3281
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808209  sky130_fd_pr__pfet_01v8__example_55959141808209_2
timestamp 1694700623
transform -1 0 6580 0 1 4291
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808209  sky130_fd_pr__pfet_01v8__example_55959141808209_3
timestamp 1694700623
transform -1 0 6580 0 -1 4819
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808211  sky130_fd_pr__pfet_01v8__example_55959141808211_0
timestamp 1694700623
transform 1 0 10376 0 -1 4804
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808213  sky130_fd_pr__pfet_01v8__example_55959141808213_0
timestamp 1694700623
transform 0 1 8893 -1 0 3464
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808214  sky130_fd_pr__pfet_01v8__example_55959141808214_0
timestamp 1694700623
transform 0 1 574 -1 0 2388
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808215  sky130_fd_pr__pfet_01v8__example_55959141808215_0
timestamp 1694700623
transform 1 0 8759 0 -1 4804
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808215  sky130_fd_pr__pfet_01v8__example_55959141808215_1
timestamp 1694700623
transform 0 1 574 1 0 1540
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808216  sky130_fd_pr__pfet_01v8__example_55959141808216_0
timestamp 1694700623
transform -1 0 11100 0 -1 4804
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808216  sky130_fd_pr__pfet_01v8__example_55959141808216_1
timestamp 1694700623
transform -1 0 9887 0 -1 4804
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808216  sky130_fd_pr__pfet_01v8__example_55959141808216_2
timestamp 1694700623
transform 1 0 9943 0 -1 4804
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808216  sky130_fd_pr__pfet_01v8__example_55959141808216_3
timestamp 1694700623
transform 1 0 9507 0 -1 4804
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808217  sky130_fd_pr__pfet_01v8__example_55959141808217_0
timestamp 1694700623
transform 1 0 9071 0 -1 4804
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808218  sky130_fd_pr__pfet_01v8__example_55959141808218_0
timestamp 1694700623
transform -1 0 3764 0 1 3281
box -1 0 1481 1
use sky130_fd_pr__pfet_01v8__example_55959141808220  sky130_fd_pr__pfet_01v8__example_55959141808220_0
timestamp 1694700623
transform -1 0 6068 0 1 3281
box -1 0 1225 1
use sky130_fd_pr__pfet_01v8__example_55959141808221  sky130_fd_pr__pfet_01v8__example_55959141808221_0
timestamp 1694700623
transform -1 0 2996 0 -1 3809
box -1 0 713 1
use sky130_fd_pr__pfet_01v8__example_55959141808222  sky130_fd_pr__pfet_01v8__example_55959141808222_0
timestamp 1694700623
transform -1 0 6068 0 -1 3809
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808223  sky130_fd_pr__pfet_01v8__example_55959141808223_0
timestamp 1694700623
transform -1 0 4788 0 1 4291
box -1 0 969 1
use sky130_fd_pr__pfet_01v8__example_55959141808223  sky130_fd_pr__pfet_01v8__example_55959141808223_1
timestamp 1694700623
transform -1 0 3252 0 1 4291
box -1 0 969 1
use sky130_fd_pr__pfet_01v8__example_55959141808223  sky130_fd_pr__pfet_01v8__example_55959141808223_2
timestamp 1694700623
transform -1 0 4788 0 1 3281
box -1 0 969 1
use sky130_fd_pr__pfet_01v8__example_55959141808224  sky130_fd_pr__pfet_01v8__example_55959141808224_0
timestamp 1694700623
transform -1 0 3764 0 1 4291
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808224  sky130_fd_pr__pfet_01v8__example_55959141808224_1
timestamp 1694700623
transform -1 0 5300 0 1 4291
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808224  sky130_fd_pr__pfet_01v8__example_55959141808224_2
timestamp 1694700623
transform -1 0 3508 0 -1 3809
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808224  sky130_fd_pr__pfet_01v8__example_55959141808224_3
timestamp 1694700623
transform -1 0 5556 0 -1 3809
box -1 0 457 1
use sky130_fd_pr__pfet_01v8__example_55959141808226  sky130_fd_pr__pfet_01v8__example_55959141808226_0
timestamp 1694700623
transform -1 0 6068 0 1 4291
box -1 0 713 1
use sky130_fd_pr__pfet_01v8__example_55959141808227  sky130_fd_pr__pfet_01v8__example_55959141808227_0
timestamp 1694700623
transform -1 0 3508 0 -1 4819
box -1 0 1225 1
use sky130_fd_pr__pfet_01v8__example_55959141808228  sky130_fd_pr__pfet_01v8__example_55959141808228_0
timestamp 1694700623
transform -1 0 5044 0 -1 3809
box -1 0 1481 1
use sky130_fd_pr__pfet_01v8__example_55959141808228  sky130_fd_pr__pfet_01v8__example_55959141808228_1
timestamp 1694700623
transform -1 0 5044 0 -1 4819
box -1 0 1481 1
use sky130_fd_pr__pfet_01v8__example_55959141808229  sky130_fd_pr__pfet_01v8__example_55959141808229_0
timestamp 1694700623
transform -1 0 6068 0 -1 4819
box -1 0 969 1
use sky130_fd_pr__res_bent_nd__example_55959141808186  sky130_fd_pr__res_bent_nd__example_55959141808186_0
timestamp 1694700623
transform 1 0 10668 0 -1 2221
box -42 -501 -38 22
use sky130_fd_pr__res_bent_nd__example_55959141808188  sky130_fd_pr__res_bent_nd__example_55959141808188_0
timestamp 1694700623
transform 0 -1 615 1 0 -10922
box -42 -327 7512 22
use sky130_fd_pr__res_bent_po__example_55959141808185  sky130_fd_pr__res_bent_po__example_55959141808185_0
timestamp 1694700623
transform -1 0 18874 0 -1 -12843
box -50 -1242 -45 9
<< labels >>
flabel metal2 s 4888 -129 5043 160 3 FreeSans 520 180 0 0 VGND_IO
port 2 nsew
flabel metal2 s 2077 555 2249 637 3 FreeSans 520 0 0 0 PD_H[3]
port 3 nsew
flabel metal2 s 22750 -1548 22858 -1180 3 FreeSans 520 0 0 0 PAD_CAP
port 4 nsew
flabel metal2 s 11333 4756 11702 4958 3 FreeSans 520 90 0 0 VCC_IO
port 5 nsew
flabel metal2 s 18968 -1544 19076 -1176 3 FreeSans 520 180 0 0 PAD_CAP
port 4 nsew
flabel metal2 s 3088 -17325 3140 -17284 3 FreeSans 520 0 0 0 PUG_H
port 6 nsew
flabel metal3 s 2695 -10265 2735 -10236 0 FreeSans 200 0 0 0 NGHS_H
port 8 nsew
flabel metal3 s 1951 885 2102 961 3 FreeSans 520 0 0 0 PD_H[2]
port 9 nsew
flabel metal3 s 21348 -1242 21941 -797 3 FreeSans 520 270 0 0 VGND_IO
port 2 nsew
flabel metal3 s 18456 3587 18497 3653 3 FreeSans 520 90 0 0 SLEW_CTL_H[0]
port 10 nsew
flabel locali s 18469 4070 18505 4106 3 FreeSans 520 90 0 0 SLEW_CTL_H[1]
port 12 nsew
flabel locali s 19260 4017 19316 4061 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[0]
port 13 nsew
flabel locali s 16848 4024 16880 4068 3 FreeSans 520 90 0 0 DRVLO_H_N
port 14 nsew
flabel locali s 18105 4088 18135 4117 3 FreeSans 520 90 0 0 I2C_MODE_H_N
port 15 nsew
flabel locali s 11972 4081 12003 4119 3 FreeSans 520 90 0 0 PD_DIS_H
port 16 nsew
flabel locali s 17014 4031 17045 4071 3 FreeSans 520 90 0 0 PDEN_H_N[1]
port 17 nsew
flabel locali s 18283 4076 18318 4111 3 FreeSans 520 90 0 0 SLOW_H_N
port 18 nsew
flabel metal1 s 18571 4744 19157 4946 3 FreeSans 520 90 0 0 VCC_IO
port 5 nsew
flabel metal1 s 18630 3590 19225 3745 3 FreeSans 520 90 0 0 VGND_IO
port 2 nsew
flabel metal1 s 17406 4571 17436 4637 3 FreeSans 520 90 0 0 EN_CMOS_B
port 20 nsew
flabel metal1 s 19916 2647 19948 2732 3 FreeSans 520 0 0 0 NSW_EN_INT
port 21 nsew
flabel metal1 s 20525 1380 20588 1458 3 FreeSans 520 0 0 0 VSSD
port 22 nsew
flabel metal1 s 11560 3636 11602 3678 3 FreeSans 520 90 0 0 OE_I_H_N
port 23 nsew
flabel metal1 s 19460 3457 19539 3489 3 FreeSans 520 180 0 0 SLEW_CTL_H_N[1]
port 24 nsew
flabel metal1 s 25673 1280 25828 1875 3 FreeSans 520 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 24462 1352 24664 1938 3 FreeSans 520 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 18656 136 18699 169 3 FreeSans 520 0 0 0 PGHS_H
port 25 nsew
flabel comment s 729 2798 729 2798 0 FreeSans 440 0 0 0 B
flabel comment s 4932 3754 4932 3754 0 FreeSans 800 0 0 0 A
flabel comment s 4687 3754 4687 3754 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 5465 3754 5465 3754 0 FreeSans 800 0 0 0 C
flabel comment s 642 2795 642 2795 0 FreeSans 440 0 0 0 C
flabel comment s 809 2801 809 2801 0 FreeSans 440 0 0 0 E
flabel comment s 561 2804 561 2804 0 FreeSans 440 0 0 0 D
flabel comment s 5195 3754 5195 3754 0 FreeSans 800 0 0 0 A
flabel comment s 3659 3758 3659 3758 0 FreeSans 800 0 0 0 A
flabel comment s 2123 3755 2123 3755 0 FreeSans 800 0 0 0 B
flabel comment s 6198 3754 6198 3754 0 FreeSans 800 0 0 0 B
flabel comment s 6468 3754 6468 3754 0 FreeSans 800 0 0 0 B
flabel comment s 11813 4088 11813 4088 0 FreeSans 200 270 0 0 NSW_ENB
flabel comment s 1360 3019 1360 3019 0 FreeSans 440 0 0 0 A
flabel comment s 12006 4084 12006 4084 0 FreeSans 200 270 0 0 PD_DIS_H
flabel comment s 723 4019 723 4019 0 FreeSans 440 180 0 0 B
flabel comment s 761 4255 761 4255 0 FreeSans 440 180 0 0 E
flabel comment s 2363 4148 2363 4148 0 FreeSans 440 180 0 0 NET367
flabel comment s 2337 3960 2337 3960 0 FreeSans 440 180 0 0 NC
flabel comment s 19463 4038 19463 4038 0 FreeSans 200 90 0 0 SLEW_CTL_H_N[1]
flabel comment s 19278 4042 19278 4042 0 FreeSans 200 90 0 0 SLEW_CTL_H_N[0]
flabel comment s 19742 4089 19742 4089 0 FreeSans 200 90 0 0 MODE0B
flabel comment s 18334 4034 18334 4034 0 FreeSans 200 90 0 0 SLEW_CTL_H[1]
flabel comment s 18516 4046 18516 4046 0 FreeSans 200 90 0 0 SLEW_CTL_H[0]
flabel comment s 18524 3860 18524 3860 0 FreeSans 200 0 0 0 MODE2B
flabel comment s 18421 4744 18421 4744 0 FreeSans 200 90 0 0 MODE2B
flabel comment s 18146 4108 18146 4108 0 FreeSans 200 90 0 0 SLOW_H_N
flabel comment s 17968 4107 17968 4107 0 FreeSans 200 90 0 0 I2C_MODE_H_N
flabel comment s 16709 4055 16709 4055 0 FreeSans 200 90 0 0 DRVLO_H_N
flabel comment s 16970 4683 16970 4683 0 FreeSans 200 90 0 0 PDEN_H<1>
flabel comment s 16622 4669 16622 4669 0 FreeSans 200 90 0 0 DRVLO_H
flabel comment s 17553 4699 17553 4699 0 FreeSans 200 90 0 0 NSW_ENB
flabel comment s 16879 4063 16879 4063 0 FreeSans 200 90 0 0 PDEN_H_N[1]
flabel comment s 17269 4701 17269 4701 0 FreeSans 200 90 0 0 EN_CMOS_B
flabel comment s 17866 4699 17866 4699 0 FreeSans 200 90 0 0 NSW_EN
flabel comment s 15791 4694 15791 4694 0 FreeSans 200 90 0 0 DRVLO_H_N_I2C
flabel comment s 14983 4613 14983 4613 0 FreeSans 200 90 0 0 DRVLO_H_N_I2C_0
flabel comment s 15589 4109 15589 4109 0 FreeSans 200 90 0 0 DRVLO_H_N_I2C
flabel comment s 15410 4092 15410 4092 0 FreeSans 200 90 0 0 MODE0B
flabel comment s 12333 4028 12333 4028 0 FreeSans 200 90 0 0 VDELAY
flabel comment s 1341 1696 1341 1696 0 FreeSans 200 270 0 0 PD_H[3]
flabel comment s 2713 1051 2713 1051 0 FreeSans 200 0 0 0 PDEN_H<1>
flabel comment s 3344 1053 3344 1053 0 FreeSans 200 0 0 0 DRVLO_H_N
flabel comment s 3955 1052 3955 1052 0 FreeSans 200 0 0 0 PDEN_H_N[1]
flabel comment s 2393 3755 2393 3755 0 FreeSans 800 0 0 0 B
flabel comment s 4173 3757 4173 3757 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 4443 3756 4443 3756 0 FreeSans 800 0 0 0 D
flabel comment s 3396 3758 3396 3758 0 FreeSans 800 0 0 0 A
flabel comment s 3929 3758 3929 3758 0 FreeSans 800 0 0 0 A
flabel comment s 5979 3754 5979 3754 0 FreeSans 800 0 0 0 B
flabel comment s 5709 3754 5709 3754 0 FreeSans 800 0 0 0 C
flabel comment s 4662 904 4662 904 0 FreeSans 200 0 0 0 RES1
flabel comment s 7734 552 7734 552 0 FreeSans 200 0 0 0 RES2
flabel comment s 1495 2995 1495 2995 0 FreeSans 400 90 0 0 BIASP
flabel comment s 1380 749 1380 749 0 FreeSans 200 90 0 0 PD_H[3]
flabel comment s 1086 1806 1086 1806 0 FreeSans 200 90 0 0 NSW_ENB
flabel comment s 5640 745 5640 745 0 FreeSans 200 90 0 0 PD_H[2]
flabel comment s 13385 4613 13385 4613 0 FreeSans 200 90 0 0 DRVLO_H_N_I2C_2
flabel comment s 14185 4613 14185 4613 0 FreeSans 200 90 0 0 DRVLO_H_N_I2C_1
flabel comment s 9146 1417 9146 1417 0 FreeSans 440 90 0 0 2VTN
flabel comment s 11377 3445 11377 3445 0 FreeSans 200 0 0 0 DRVLO_H_N_I2C
flabel comment s 725 -88 725 -88 0 FreeSans 200 90 0 0 B
flabel comment s 723 -1596 723 -1596 0 FreeSans 200 90 0 0 D
flabel comment s 1843 2592 1843 2592 0 FreeSans 400 90 0 0 BIASP1
flabel comment s 18825 3860 18825 3860 0 FreeSans 200 0 0 0 MODE4B
flabel comment s 3272 -174 3272 -174 0 FreeSans 200 0 0 0 CONDIODE
flabel comment s 10257 2539 10257 2539 0 FreeSans 440 0 0 0 D
flabel comment s 11946 3567 11946 3567 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 7816 630 7816 630 0 FreeSans 200 0 0 0 RES2
flabel comment s 1870 3338 1870 3338 0 FreeSans 800 0 0 0 E
flabel comment s 18986 2925 18986 2925 0 FreeSans 600 0 0 0 NE
flabel comment s 18761 2924 18761 2924 0 FreeSans 600 0 0 0 ND
flabel comment s 964 2801 964 2801 0 FreeSans 440 0 0 0 F
flabel comment s 6727 4763 6727 4763 0 FreeSans 800 0 0 0 E
flabel comment s 1875 4350 1875 4350 0 FreeSans 800 0 0 0 B
flabel comment s 18605 2652 18605 2652 0 FreeSans 600 0 0 0 NC
flabel comment s 2337 4064 2337 4064 0 FreeSans 440 180 0 0 NA
flabel comment s 8430 3109 8430 3109 0 FreeSans 600 0 0 0 ENB
flabel comment s 1329 1025 1329 1025 0 FreeSans 400 0 0 0 CAS5
flabel comment s 2123 4763 2123 4763 0 FreeSans 800 0 0 0 F
flabel comment s 2393 4763 2393 4763 0 FreeSans 800 0 0 0 F
flabel comment s 2907 4763 2907 4763 0 FreeSans 800 0 0 0 F
flabel comment s 2637 4763 2637 4763 0 FreeSans 800 0 0 0 F
flabel comment s 3396 4763 3396 4763 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 3126 4763 3126 4763 0 FreeSans 800 0 0 0 C
flabel comment s 4173 4763 4173 4763 0 FreeSans 800 0 0 0 D
flabel comment s 4443 4763 4443 4763 0 FreeSans 800 0 0 0 D
flabel comment s 4662 4763 4662 4763 0 FreeSans 800 0 0 0 D
flabel comment s 4932 4763 4932 4763 0 FreeSans 800 0 0 0 D
flabel comment s 3659 4763 3659 4763 0 FreeSans 800 0 0 0 D
flabel comment s 3929 4763 3929 4763 0 FreeSans 800 0 0 0 D
flabel comment s 5709 4763 5709 4763 0 FreeSans 800 0 0 0 E
flabel comment s 5979 4763 5979 4763 0 FreeSans 800 0 0 0 E
flabel comment s 6198 4763 6198 4763 0 FreeSans 800 0 0 0 E
flabel comment s 6468 4763 6468 4763 0 FreeSans 800 0 0 0 E
flabel comment s 5195 4763 5195 4763 0 FreeSans 800 0 0 0 E
flabel comment s 5465 4763 5465 4763 0 FreeSans 800 0 0 0 E
flabel comment s 2123 3338 2123 3338 0 FreeSans 800 0 0 0 E
flabel comment s 2393 3338 2393 3338 0 FreeSans 800 0 0 0 E
flabel comment s 2637 3338 2637 3338 0 FreeSans 800 0 0 0 E
flabel comment s 2907 3338 2907 3338 0 FreeSans 800 0 0 0 E
flabel comment s 3126 3338 3126 3338 0 FreeSans 800 0 0 0 E
flabel comment s 3396 3338 3396 3338 0 FreeSans 800 0 0 0 E
flabel comment s 3659 3338 3659 3338 0 FreeSans 800 0 0 0 D
flabel comment s 3929 3338 3929 3338 0 FreeSans 800 0 0 0 D
flabel comment s 4173 3338 4173 3338 0 FreeSans 800 0 0 0 D
flabel comment s 4443 3338 4443 3338 0 FreeSans 800 0 0 0 D
flabel comment s 4662 3338 4662 3338 0 FreeSans 800 0 0 0 D
flabel comment s 4932 3338 4932 3338 0 FreeSans 800 0 0 0 D
flabel comment s 5195 3338 5195 3338 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 5465 3338 5465 3338 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 5709 3338 5709 3338 0 FreeSans 800 0 0 0 F
flabel comment s 5979 3338 5979 3338 0 FreeSans 800 0 0 0 F
flabel comment s 6198 3338 6198 3338 0 FreeSans 800 0 0 0 F
flabel comment s 6468 3338 6468 3338 0 FreeSans 800 0 0 0 F
flabel comment s 2123 4350 2123 4350 0 FreeSans 800 0 0 0 B
flabel comment s 2393 4350 2393 4350 0 FreeSans 800 0 0 0 B
flabel comment s 2637 4350 2637 4350 0 FreeSans 800 0 0 0 B
flabel comment s 2907 4350 2907 4350 0 FreeSans 800 0 0 0 C
flabel comment s 3126 4350 3126 4350 0 FreeSans 800 0 0 0 C
flabel comment s 3396 4350 3396 4350 0 FreeSans 800 0 0 0 A
flabel comment s 3659 4350 3659 4350 0 FreeSans 800 0 0 0 A
flabel comment s 3929 4350 3929 4350 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 4173 4350 4173 4350 0 FreeSans 800 0 0 0 D
flabel comment s 4443 4350 4443 4350 0 FreeSans 200 0 0 0 DUMMY
flabel comment s 4662 4350 4662 4350 0 FreeSans 800 0 0 0 A
flabel comment s 4932 4350 4932 4350 0 FreeSans 800 0 0 0 A
flabel comment s 5195 4350 5195 4350 0 FreeSans 800 0 0 0 A
flabel comment s 5465 4350 5465 4350 0 FreeSans 800 0 0 0 B
flabel comment s 5709 4350 5709 4350 0 FreeSans 800 0 0 0 B
flabel comment s 5979 4350 5979 4350 0 FreeSans 800 0 0 0 B
flabel comment s 6198 4350 6198 4350 0 FreeSans 800 0 0 0 B
flabel comment s 6468 4350 6468 4350 0 FreeSans 800 0 0 0 B
flabel comment s 2637 3755 2637 3755 0 FreeSans 800 0 0 0 B
flabel comment s 2907 3755 2907 3755 0 FreeSans 800 0 0 0 B
flabel comment s 3126 3755 3126 3755 0 FreeSans 800 0 0 0 B
flabel comment s 25986 1800 25986 1800 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 760 212 760 212 0 FreeSans 400 0 0 0 CAS3
flabel comment s 1452 -764 1452 -764 0 FreeSans 400 0 0 0 PD_H[3]
<< properties >>
string GDS_END 38168744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37335308
<< end >>
