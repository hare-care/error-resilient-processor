magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1559 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 961 47 991 177
rect 1115 47 1145 177
rect 1199 47 1229 177
rect 1283 47 1313 177
rect 1367 47 1397 177
rect 1451 47 1481 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 483 297 513 497
rect 567 297 597 497
rect 651 297 681 497
rect 735 297 765 497
rect 927 297 957 497
rect 1011 297 1041 497
rect 1199 297 1229 497
rect 1283 297 1313 497
rect 1367 297 1397 497
rect 1451 297 1481 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 47 163 127
rect 193 89 247 177
rect 193 55 203 89
rect 237 55 247 89
rect 193 47 247 55
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 47 331 127
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 467 93 519 177
rect 467 59 475 93
rect 509 59 519 93
rect 467 47 519 59
rect 549 169 603 177
rect 549 135 559 169
rect 593 135 603 169
rect 549 47 603 135
rect 633 157 687 177
rect 633 123 643 157
rect 677 123 687 157
rect 633 89 687 123
rect 633 55 643 89
rect 677 55 687 89
rect 633 47 687 55
rect 717 169 771 177
rect 717 135 727 169
rect 761 135 771 169
rect 717 47 771 135
rect 801 93 853 177
rect 801 59 811 93
rect 845 59 853 93
rect 801 47 853 59
rect 909 161 961 177
rect 909 127 917 161
rect 951 127 961 161
rect 909 47 961 127
rect 991 89 1115 177
rect 991 55 1002 89
rect 1036 55 1070 89
rect 1104 55 1115 89
rect 991 47 1115 55
rect 1145 161 1199 177
rect 1145 127 1155 161
rect 1189 127 1199 161
rect 1145 47 1199 127
rect 1229 89 1283 177
rect 1229 55 1239 89
rect 1273 55 1283 89
rect 1229 47 1283 55
rect 1313 161 1367 177
rect 1313 127 1323 161
rect 1357 127 1367 161
rect 1313 47 1367 127
rect 1397 89 1451 177
rect 1397 55 1407 89
rect 1441 55 1451 89
rect 1397 47 1451 55
rect 1481 161 1533 177
rect 1481 127 1491 161
rect 1525 127 1533 161
rect 1481 47 1533 127
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 448 163 497
rect 109 414 119 448
rect 153 414 163 448
rect 109 380 163 414
rect 109 346 119 380
rect 153 346 163 380
rect 109 297 163 346
rect 193 489 247 497
rect 193 455 203 489
rect 237 455 247 489
rect 193 421 247 455
rect 193 387 203 421
rect 237 387 247 421
rect 193 297 247 387
rect 277 448 331 497
rect 277 414 287 448
rect 321 414 331 448
rect 277 380 331 414
rect 277 346 287 380
rect 321 346 331 380
rect 277 297 331 346
rect 361 489 483 497
rect 361 387 371 489
rect 473 387 483 489
rect 361 297 483 387
rect 513 448 567 497
rect 513 414 523 448
rect 557 414 567 448
rect 513 380 567 414
rect 513 346 523 380
rect 557 346 567 380
rect 513 297 567 346
rect 597 489 651 497
rect 597 455 607 489
rect 641 455 651 489
rect 597 421 651 455
rect 597 387 607 421
rect 641 387 651 421
rect 597 297 651 387
rect 681 448 735 497
rect 681 414 691 448
rect 725 414 735 448
rect 681 380 735 414
rect 681 346 691 380
rect 725 346 735 380
rect 681 297 735 346
rect 765 429 817 497
rect 765 395 775 429
rect 809 395 817 429
rect 765 297 817 395
rect 875 429 927 497
rect 875 395 883 429
rect 917 395 927 429
rect 875 297 927 395
rect 957 380 1011 497
rect 957 346 967 380
rect 1001 346 1011 380
rect 957 297 1011 346
rect 1041 378 1093 497
rect 1041 344 1051 378
rect 1085 344 1093 378
rect 1041 297 1093 344
rect 1147 380 1199 497
rect 1147 346 1155 380
rect 1189 346 1199 380
rect 1147 297 1199 346
rect 1229 489 1283 497
rect 1229 455 1239 489
rect 1273 455 1283 489
rect 1229 421 1283 455
rect 1229 387 1239 421
rect 1273 387 1283 421
rect 1229 297 1283 387
rect 1313 380 1367 497
rect 1313 346 1323 380
rect 1357 346 1367 380
rect 1313 297 1367 346
rect 1397 489 1451 497
rect 1397 455 1407 489
rect 1441 455 1451 489
rect 1397 421 1451 455
rect 1397 387 1407 421
rect 1441 387 1451 421
rect 1397 297 1451 387
rect 1481 448 1533 497
rect 1481 414 1491 448
rect 1525 414 1533 448
rect 1481 380 1533 414
rect 1481 346 1491 380
rect 1525 346 1533 380
rect 1481 297 1533 346
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 203 55 237 89
rect 287 127 321 161
rect 371 59 405 93
rect 475 59 509 93
rect 559 135 593 169
rect 643 123 677 157
rect 643 55 677 89
rect 727 135 761 169
rect 811 59 845 93
rect 917 127 951 161
rect 1002 55 1036 89
rect 1070 55 1104 89
rect 1155 127 1189 161
rect 1239 55 1273 89
rect 1323 127 1357 161
rect 1407 55 1441 89
rect 1491 127 1525 161
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 414 153 448
rect 119 346 153 380
rect 203 455 237 489
rect 203 387 237 421
rect 287 414 321 448
rect 287 346 321 380
rect 371 387 473 489
rect 523 414 557 448
rect 523 346 557 380
rect 607 455 641 489
rect 607 387 641 421
rect 691 414 725 448
rect 691 346 725 380
rect 775 395 809 429
rect 883 395 917 429
rect 967 346 1001 380
rect 1051 344 1085 378
rect 1155 346 1189 380
rect 1239 455 1273 489
rect 1239 387 1273 421
rect 1323 346 1357 380
rect 1407 455 1441 489
rect 1407 387 1441 421
rect 1491 414 1525 448
rect 1491 346 1525 380
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 483 497 513 523
rect 567 497 597 523
rect 651 497 681 523
rect 735 497 765 523
rect 927 497 957 523
rect 1011 497 1041 523
rect 1199 497 1229 523
rect 1283 497 1313 523
rect 1367 497 1397 523
rect 1451 497 1481 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 249 389 265
rect 483 259 513 297
rect 567 259 597 297
rect 651 282 681 297
rect 735 282 765 297
rect 651 265 777 282
rect 651 260 801 265
rect 653 259 801 260
rect 79 215 203 249
rect 237 215 271 249
rect 305 215 339 249
rect 373 215 389 249
rect 79 199 389 215
rect 464 249 597 259
rect 655 258 801 259
rect 657 257 801 258
rect 658 256 801 257
rect 659 255 801 256
rect 661 254 801 255
rect 662 253 801 254
rect 663 252 801 253
rect 464 215 547 249
rect 581 222 597 249
rect 687 249 801 252
rect 581 215 633 222
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 464 192 633 215
rect 519 177 549 192
rect 603 177 633 192
rect 687 215 723 249
rect 757 215 801 249
rect 687 199 801 215
rect 927 259 957 297
rect 1011 259 1041 297
rect 1199 259 1229 297
rect 1283 259 1313 297
rect 927 249 1145 259
rect 927 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1145 249
rect 927 205 1145 215
rect 687 177 717 199
rect 771 177 801 199
rect 961 177 991 205
rect 1115 177 1145 205
rect 1199 249 1313 259
rect 1199 215 1223 249
rect 1257 215 1313 249
rect 1199 205 1313 215
rect 1199 177 1229 205
rect 1283 177 1313 205
rect 1367 259 1397 297
rect 1451 261 1481 297
rect 1451 259 1524 261
rect 1367 249 1524 259
rect 1367 215 1406 249
rect 1440 215 1474 249
rect 1508 215 1524 249
rect 1367 205 1524 215
rect 1367 177 1397 205
rect 1451 203 1524 205
rect 1451 177 1481 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 961 21 991 47
rect 1115 21 1145 47
rect 1199 21 1229 47
rect 1283 21 1313 47
rect 1367 21 1397 47
rect 1451 21 1481 47
<< polycont >>
rect 203 215 237 249
rect 271 215 305 249
rect 339 215 373 249
rect 547 215 581 249
rect 723 215 757 249
rect 947 215 981 249
rect 1015 215 1049 249
rect 1083 215 1117 249
rect 1223 215 1257 249
rect 1406 215 1440 249
rect 1474 215 1508 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 485 85 527
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 297 85 315
rect 119 448 153 493
rect 119 380 153 414
rect 187 489 253 527
rect 187 455 203 489
rect 237 455 253 489
rect 187 421 253 455
rect 187 387 203 421
rect 237 387 253 421
rect 187 379 253 387
rect 287 448 321 493
rect 287 380 321 414
rect 119 345 153 346
rect 355 489 489 527
rect 355 387 371 489
rect 473 387 489 489
rect 355 379 489 387
rect 523 448 557 493
rect 523 380 557 414
rect 287 345 321 346
rect 591 489 657 527
rect 591 455 607 489
rect 641 455 657 489
rect 591 421 657 455
rect 591 387 607 421
rect 641 387 657 421
rect 591 379 657 387
rect 691 448 725 493
rect 691 380 725 414
rect 523 345 557 346
rect 771 429 809 527
rect 771 395 775 429
rect 771 379 809 395
rect 867 489 1289 493
rect 867 459 1239 489
rect 867 429 933 459
rect 867 395 883 429
rect 917 395 933 429
rect 867 379 933 395
rect 967 380 1001 425
rect 691 345 725 346
rect 967 345 1001 346
rect 119 297 321 345
rect 355 297 1001 345
rect 1051 378 1105 459
rect 1223 455 1239 459
rect 1273 455 1289 489
rect 1085 344 1105 378
rect 1051 297 1105 344
rect 1139 380 1189 425
rect 1139 346 1155 380
rect 1223 421 1289 455
rect 1391 489 1457 527
rect 1391 455 1407 489
rect 1441 455 1457 489
rect 1223 387 1239 421
rect 1273 387 1289 421
rect 1223 379 1289 387
rect 1323 380 1357 425
rect 1139 345 1189 346
rect 1391 421 1457 455
rect 1391 387 1407 421
rect 1441 387 1457 421
rect 1391 379 1457 387
rect 1491 448 1547 493
rect 1525 414 1547 448
rect 1491 380 1547 414
rect 1323 345 1357 346
rect 1525 346 1547 380
rect 1491 345 1547 346
rect 1139 297 1547 345
rect 119 263 153 297
rect 355 263 389 297
rect 17 211 153 263
rect 187 249 389 263
rect 187 215 203 249
rect 237 215 271 249
rect 305 215 339 249
rect 373 215 389 249
rect 187 211 389 215
rect 423 249 616 263
rect 423 215 547 249
rect 581 215 616 249
rect 423 211 616 215
rect 650 249 895 263
rect 650 215 723 249
rect 757 215 895 249
rect 650 211 895 215
rect 931 249 1170 263
rect 931 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1170 249
rect 931 211 1170 215
rect 1204 249 1354 263
rect 1204 215 1223 249
rect 1257 215 1354 249
rect 1204 211 1354 215
rect 1390 249 1547 263
rect 1390 215 1406 249
rect 1440 215 1474 249
rect 1508 215 1547 249
rect 1390 211 1547 215
rect 119 177 153 211
rect 355 177 389 211
rect 17 161 85 177
rect 17 127 35 161
rect 69 127 85 161
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 17 85 59
rect 119 161 321 177
rect 153 143 287 161
rect 119 51 153 127
rect 355 169 609 177
rect 355 143 559 169
rect 439 135 559 143
rect 593 135 609 169
rect 643 157 677 177
rect 187 89 253 109
rect 187 55 203 89
rect 237 55 253 89
rect 187 17 253 55
rect 287 51 321 127
rect 711 169 1547 177
rect 711 135 727 169
rect 761 161 1547 169
rect 761 135 917 161
rect 355 93 405 109
rect 643 101 677 123
rect 897 127 917 135
rect 951 135 1155 161
rect 355 59 371 93
rect 355 17 405 59
rect 439 93 861 101
rect 439 59 475 93
rect 509 89 811 93
rect 509 59 643 89
rect 439 55 643 59
rect 677 59 811 89
rect 845 59 861 93
rect 677 55 861 59
rect 439 51 861 55
rect 897 51 951 127
rect 1189 135 1323 161
rect 985 89 1121 101
rect 985 55 1002 89
rect 1036 55 1070 89
rect 1104 55 1121 89
rect 985 17 1121 55
rect 1155 51 1189 127
rect 1357 135 1491 161
rect 1223 89 1289 101
rect 1223 55 1239 89
rect 1273 55 1289 89
rect 1223 17 1289 55
rect 1323 51 1357 127
rect 1525 127 1547 161
rect 1391 89 1457 101
rect 1391 55 1407 89
rect 1441 55 1457 89
rect 1391 17 1457 55
rect 1491 51 1547 127
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1502 221 1536 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1410 221 1444 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1318 221 1352 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1134 221 1168 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 1226 221 1260 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o311a_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 904470
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 892178
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.820 0.000 
<< end >>
