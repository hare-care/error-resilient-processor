magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< pwell >>
rect 90 486 106 503
<< metal1 >>
rect -88 912 396 918
rect -88 860 -36 912
rect 16 860 28 912
rect 80 860 92 912
rect 144 860 156 912
rect 208 860 220 912
rect 272 860 284 912
rect 336 860 396 912
rect -88 854 396 860
rect -88 809 -34 854
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 92 -34 117
rect 0 64 28 826
rect 56 92 84 854
rect 112 64 140 826
rect 168 92 196 854
rect 224 64 252 826
rect 280 92 308 854
rect 342 809 396 854
rect 342 757 343 809
rect 395 757 396 809
rect 342 745 396 757
rect 342 693 343 745
rect 395 693 396 745
rect 342 681 396 693
rect 342 629 343 681
rect 395 629 396 681
rect 342 617 396 629
rect 342 565 343 617
rect 395 565 396 617
rect 342 553 396 565
rect 342 501 343 553
rect 395 501 396 553
rect 342 489 396 501
rect 342 437 343 489
rect 395 437 396 489
rect 342 425 396 437
rect 342 373 343 425
rect 395 373 396 425
rect 342 361 396 373
rect 342 309 343 361
rect 395 309 396 361
rect 342 297 396 309
rect 342 245 343 297
rect 395 245 396 297
rect 342 233 396 245
rect 342 181 343 233
rect 395 181 396 233
rect 342 169 396 181
rect 342 117 343 169
rect 395 117 396 169
rect 342 92 396 117
rect 0 58 308 64
rect 0 6 28 58
rect 80 6 92 58
rect 144 6 156 58
rect 208 6 220 58
rect 272 6 308 58
rect 0 0 308 6
<< via1 >>
rect -36 860 16 912
rect 28 860 80 912
rect 92 860 144 912
rect 156 860 208 912
rect 220 860 272 912
rect 284 860 336 912
rect -87 757 -35 809
rect -87 693 -35 745
rect -87 629 -35 681
rect -87 565 -35 617
rect -87 501 -35 553
rect -87 437 -35 489
rect -87 373 -35 425
rect -87 309 -35 361
rect -87 245 -35 297
rect -87 181 -35 233
rect -87 117 -35 169
rect 343 757 395 809
rect 343 693 395 745
rect 343 629 395 681
rect 343 565 395 617
rect 343 501 395 553
rect 343 437 395 489
rect 343 373 395 425
rect 343 309 395 361
rect 343 245 395 297
rect 343 181 395 233
rect 343 117 395 169
rect 28 6 80 58
rect 92 6 144 58
rect 156 6 208 58
rect 220 6 272 58
<< metal2 >>
rect -88 912 396 918
rect -88 860 -36 912
rect 16 860 28 912
rect 80 860 92 912
rect 144 860 156 912
rect 208 860 220 912
rect 272 860 284 912
rect 336 860 396 912
rect -88 854 396 860
rect -88 809 -34 854
rect -88 757 -87 809
rect -35 757 -34 809
rect -88 745 -34 757
rect -88 693 -87 745
rect -35 693 -34 745
rect -88 681 -34 693
rect -88 629 -87 681
rect -35 629 -34 681
rect -88 617 -34 629
rect -88 565 -87 617
rect -35 565 -34 617
rect -88 553 -34 565
rect -88 501 -87 553
rect -35 501 -34 553
rect -88 489 -34 501
rect -88 437 -87 489
rect -35 437 -34 489
rect -88 425 -34 437
rect -88 373 -87 425
rect -35 373 -34 425
rect -88 361 -34 373
rect -88 309 -87 361
rect -35 309 -34 361
rect -88 297 -34 309
rect -88 245 -87 297
rect -35 245 -34 297
rect -88 233 -34 245
rect -88 181 -87 233
rect -35 181 -34 233
rect -88 169 -34 181
rect -88 117 -87 169
rect -35 117 -34 169
rect -88 92 -34 117
rect 0 92 28 854
rect 56 64 84 826
rect 112 92 140 854
rect 168 64 196 826
rect 224 92 252 854
rect 280 64 308 826
rect 342 809 396 854
rect 342 757 343 809
rect 395 757 396 809
rect 342 745 396 757
rect 342 693 343 745
rect 395 693 396 745
rect 342 681 396 693
rect 342 629 343 681
rect 395 629 396 681
rect 342 617 396 629
rect 342 565 343 617
rect 395 565 396 617
rect 342 553 396 565
rect 342 501 343 553
rect 395 501 396 553
rect 342 489 396 501
rect 342 437 343 489
rect 395 437 396 489
rect 342 425 396 437
rect 342 373 343 425
rect 395 373 396 425
rect 342 361 396 373
rect 342 309 343 361
rect 395 309 396 361
rect 342 297 396 309
rect 342 245 343 297
rect 395 245 396 297
rect 342 233 396 245
rect 342 181 343 233
rect 395 181 396 233
rect 342 169 396 181
rect 342 117 343 169
rect 395 117 396 169
rect 342 92 396 117
rect 0 58 308 64
rect 0 6 28 58
rect 80 6 92 58
rect 144 6 156 58
rect 208 6 220 58
rect 272 6 308 58
rect 0 0 308 6
<< labels >>
flabel metal2 s 172 110 194 137 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 116 781 137 807 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 90 486 106 503 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 4180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 148
string device primitive
<< end >>
