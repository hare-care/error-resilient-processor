magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 704 157 886 201
rect 1193 157 1547 203
rect 1 21 1547 157
rect 29 -17 63 21
<< locali >>
rect 18 195 88 325
rect 274 143 330 333
rect 1377 315 1443 484
rect 1377 299 1455 315
rect 1412 289 1455 299
rect 1421 173 1455 289
rect 1410 165 1455 173
rect 1379 148 1455 165
rect 1379 61 1445 148
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 240 493
rect 288 435 341 527
rect 375 408 425 493
rect 467 438 688 472
rect 364 382 425 408
rect 364 161 398 382
rect 432 225 480 344
rect 514 331 620 404
rect 514 191 548 331
rect 654 315 688 438
rect 722 367 756 527
rect 790 427 840 493
rect 885 433 1062 467
rect 654 297 756 315
rect 364 135 409 161
rect 443 147 548 191
rect 582 263 756 297
rect 291 17 341 109
rect 375 107 409 135
rect 582 107 616 263
rect 722 249 756 263
rect 658 213 698 219
rect 790 213 824 427
rect 858 249 896 393
rect 658 153 824 213
rect 930 207 994 399
rect 375 73 442 107
rect 481 73 616 107
rect 680 17 754 117
rect 790 107 824 153
rect 901 141 994 207
rect 1028 265 1062 433
rect 1098 427 1161 527
rect 1207 381 1275 493
rect 1096 306 1275 381
rect 1309 325 1343 527
rect 1237 265 1275 306
rect 1477 344 1511 527
rect 1028 199 1203 265
rect 1237 199 1387 265
rect 1028 107 1062 199
rect 1237 165 1277 199
rect 790 73 871 107
rect 905 73 1062 107
rect 1117 17 1159 123
rect 1211 60 1277 165
rect 1311 17 1345 139
rect 1479 17 1513 120
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 114 388 172 397
rect 534 388 592 397
rect 848 388 906 397
rect 114 360 906 388
rect 114 351 172 360
rect 534 351 592 360
rect 848 351 906 360
rect 193 320 251 329
rect 431 320 489 329
rect 935 320 993 329
rect 193 292 993 320
rect 193 283 251 292
rect 431 283 489 292
rect 935 283 993 292
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 274 143 330 333 6 D
port 2 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1547 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1193 157 1547 203 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 704 157 886 201 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1379 61 1445 148 6 Q
port 7 nsew signal output
rlabel locali s 1379 148 1455 165 6 Q
port 7 nsew signal output
rlabel locali s 1410 165 1455 173 6 Q
port 7 nsew signal output
rlabel locali s 1421 173 1455 289 6 Q
port 7 nsew signal output
rlabel locali s 1412 289 1455 299 6 Q
port 7 nsew signal output
rlabel locali s 1377 299 1455 315 6 Q
port 7 nsew signal output
rlabel locali s 1377 315 1443 484 6 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2633870
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2621364
<< end >>
