magic
tech sky130B
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1694700623
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_0
timestamp 1694700623
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_1
timestamp 1694700623
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48406188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48404228
<< end >>
