magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 450 897
<< pwell >>
rect 16 43 378 295
rect -26 -43 410 43
<< mvnmos >>
rect 95 119 295 269
<< mvpmos >>
rect 95 541 295 741
<< mvndiff >>
rect 42 169 95 269
rect 42 135 50 169
rect 84 135 95 169
rect 42 119 95 135
rect 295 250 352 269
rect 295 216 306 250
rect 340 216 352 250
rect 295 179 352 216
rect 295 145 306 179
rect 340 145 352 179
rect 295 119 352 145
<< mvpdiff >>
rect 42 729 95 741
rect 42 695 50 729
rect 84 695 95 729
rect 42 658 95 695
rect 42 624 50 658
rect 84 624 95 658
rect 42 587 95 624
rect 42 553 50 587
rect 84 553 95 587
rect 42 541 95 553
rect 295 729 352 741
rect 295 695 306 729
rect 340 695 352 729
rect 295 658 352 695
rect 295 624 306 658
rect 340 624 352 658
rect 295 587 352 624
rect 295 553 306 587
rect 340 553 352 587
rect 295 541 352 553
<< mvndiffc >>
rect 50 135 84 169
rect 306 216 340 250
rect 306 145 340 179
<< mvpdiffc >>
rect 50 695 84 729
rect 50 624 84 658
rect 50 553 84 587
rect 306 695 340 729
rect 306 624 340 658
rect 306 553 340 587
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
<< poly >>
rect 95 741 295 767
rect 95 515 295 541
rect 95 390 161 515
rect 95 356 111 390
rect 145 356 161 390
rect 95 340 161 356
rect 203 390 295 406
rect 203 356 219 390
rect 253 356 295 390
rect 203 295 295 356
rect 95 269 295 295
rect 95 81 295 119
<< polycont >>
rect 111 356 145 390
rect 219 356 253 390
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 50 746 340 751
rect 50 729 99 746
rect 84 712 99 729
rect 133 712 172 746
rect 206 712 260 746
rect 294 729 340 746
rect 294 712 306 729
rect 84 695 306 712
rect 50 658 340 695
rect 84 624 306 658
rect 50 587 340 624
rect 84 553 306 587
rect 50 537 340 553
rect 95 390 161 406
rect 95 356 111 390
rect 145 356 161 390
rect 95 250 161 356
rect 203 390 269 537
rect 203 356 219 390
rect 253 356 269 390
rect 203 340 269 356
rect 95 216 306 250
rect 340 216 356 250
rect 95 179 356 216
rect 95 169 306 179
rect 34 135 50 169
rect 84 145 306 169
rect 340 145 356 179
rect 84 135 356 145
rect 34 113 356 135
rect 34 79 43 113
rect 77 79 131 113
rect 165 79 219 113
rect 253 79 302 113
rect 336 79 356 113
rect 34 73 356 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 99 712 133 746
rect 172 712 206 746
rect 260 712 294 746
rect 43 79 77 113
rect 131 79 165 113
rect 219 79 253 113
rect 302 79 336 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 831 384 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 0 791 384 797
rect 0 746 384 763
rect 0 712 99 746
rect 133 712 172 746
rect 206 712 260 746
rect 294 712 384 746
rect 0 689 384 712
rect 0 113 384 125
rect 0 79 43 113
rect 77 79 131 113
rect 165 79 219 113
rect 253 79 302 113
rect 336 79 384 113
rect 0 51 384 79
rect 0 17 384 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -23 384 -17
<< labels >>
rlabel comment s 0 0 0 0 4 decap_4
flabel metal1 s 0 0 384 23 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel metal1 s 0 51 384 125 0 FreeSans 340 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 s 192 11 192 11 0 FreeSans 340 0 0 0 VNB
flabel metal1 s 0 689 384 763 0 FreeSans 340 0 0 0 VPWR
port 4 nsew power bidirectional
flabel metal1 s 0 791 384 814 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel metal1 s 192 802 192 802 0 FreeSans 340 0 0 0 VPB
<< properties >>
string FIXED_BBOX 0 0 384 814
string GDS_END 959862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 955112
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
