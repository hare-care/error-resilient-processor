magic
tech sky130A
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_1
timestamp 1694700623
transform 1 0 180 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 37249434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37248444
<< end >>
