magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -179 2150 195 2250
rect -179 1403 -14 2150
rect 6101 2150 6352 2250
rect 4038 -369 4747 -10
rect 5762 -133 6121 568
<< pwell >>
rect 2477 1941 3819 2231
rect 5803 673 6081 865
rect 3741 -328 3933 -50
rect 6257 145 6401 891
<< mvnmos >>
rect 5882 699 6002 839
rect 3767 -249 3907 -129
<< mvpmos >>
rect 5882 301 6002 501
rect 5882 33 6002 233
rect 4105 -249 4305 -129
rect 4373 -249 4573 -129
<< mvndiff >>
rect 5829 813 5882 839
rect 5829 779 5837 813
rect 5871 779 5882 813
rect 5829 745 5882 779
rect 5829 711 5837 745
rect 5871 711 5882 745
rect 5829 699 5882 711
rect 6002 813 6055 839
rect 6002 779 6013 813
rect 6047 779 6055 813
rect 6002 745 6055 779
rect 6002 711 6013 745
rect 6047 711 6055 745
rect 6002 699 6055 711
rect 3767 -84 3907 -76
rect 3767 -118 3793 -84
rect 3827 -118 3861 -84
rect 3895 -118 3907 -84
rect 3767 -129 3907 -118
rect 3767 -260 3907 -249
rect 3767 -294 3793 -260
rect 3827 -294 3861 -260
rect 3895 -294 3907 -260
rect 3767 -302 3907 -294
<< mvpdiff >>
rect 5829 483 5882 501
rect 5829 449 5837 483
rect 5871 449 5882 483
rect 5829 415 5882 449
rect 5829 381 5837 415
rect 5871 381 5882 415
rect 5829 347 5882 381
rect 5829 313 5837 347
rect 5871 313 5882 347
rect 5829 301 5882 313
rect 6002 483 6055 501
rect 6002 449 6013 483
rect 6047 449 6055 483
rect 6002 415 6055 449
rect 6002 381 6013 415
rect 6047 381 6055 415
rect 6002 347 6055 381
rect 6002 313 6013 347
rect 6047 313 6055 347
rect 6002 301 6055 313
rect 5829 221 5882 233
rect 5829 187 5837 221
rect 5871 187 5882 221
rect 5829 153 5882 187
rect 5829 119 5837 153
rect 5871 119 5882 153
rect 5829 85 5882 119
rect 5829 51 5837 85
rect 5871 51 5882 85
rect 5829 33 5882 51
rect 6002 221 6055 233
rect 6002 187 6013 221
rect 6047 187 6055 221
rect 6002 153 6055 187
rect 6002 119 6013 153
rect 6047 119 6055 153
rect 6002 85 6055 119
rect 6002 51 6013 85
rect 6047 51 6055 85
rect 6002 33 6055 51
rect 4105 -84 4305 -76
rect 4105 -118 4123 -84
rect 4157 -118 4191 -84
rect 4225 -118 4259 -84
rect 4293 -118 4305 -84
rect 4105 -129 4305 -118
rect 4373 -84 4573 -76
rect 4373 -118 4385 -84
rect 4419 -118 4453 -84
rect 4487 -118 4521 -84
rect 4555 -118 4573 -84
rect 4373 -129 4573 -118
rect 4105 -260 4305 -249
rect 4105 -294 4123 -260
rect 4157 -294 4191 -260
rect 4225 -294 4259 -260
rect 4293 -294 4305 -260
rect 4105 -302 4305 -294
rect 4373 -260 4573 -249
rect 4373 -294 4385 -260
rect 4419 -294 4453 -260
rect 4487 -294 4521 -260
rect 4555 -294 4573 -260
rect 4373 -302 4573 -294
<< mvndiffc >>
rect 5837 779 5871 813
rect 5837 711 5871 745
rect 6013 779 6047 813
rect 6013 711 6047 745
rect 3793 -118 3827 -84
rect 3861 -118 3895 -84
rect 3793 -294 3827 -260
rect 3861 -294 3895 -260
<< mvpdiffc >>
rect 5837 449 5871 483
rect 5837 381 5871 415
rect 5837 313 5871 347
rect 6013 449 6047 483
rect 6013 381 6047 415
rect 6013 313 6047 347
rect 5837 187 5871 221
rect 5837 119 5871 153
rect 5837 51 5871 85
rect 6013 187 6047 221
rect 6013 119 6047 153
rect 6013 51 6047 85
rect 4123 -118 4157 -84
rect 4191 -118 4225 -84
rect 4259 -118 4293 -84
rect 4385 -118 4419 -84
rect 4453 -118 4487 -84
rect 4521 -118 4555 -84
rect 4123 -294 4157 -260
rect 4191 -294 4225 -260
rect 4259 -294 4293 -260
rect 4385 -294 4419 -260
rect 4453 -294 4487 -260
rect 4521 -294 4555 -260
<< psubdiff >>
rect 2503 2171 2596 2205
rect 2630 2171 2669 2205
rect 2703 2171 2741 2205
rect 2775 2171 2813 2205
rect 2847 2171 2885 2205
rect 2919 2171 2957 2205
rect 2991 2171 3029 2205
rect 3063 2171 3101 2205
rect 3135 2171 3173 2205
rect 3207 2171 3245 2205
rect 3279 2171 3317 2205
rect 3351 2171 3389 2205
rect 3423 2171 3461 2205
rect 3495 2171 3533 2205
rect 3567 2171 3605 2205
rect 3639 2171 3677 2205
rect 3711 2171 3793 2205
rect 2503 2137 3793 2171
rect 2503 2103 2596 2137
rect 2630 2103 2669 2137
rect 2703 2103 2741 2137
rect 2775 2103 2813 2137
rect 2847 2103 2885 2137
rect 2919 2103 2957 2137
rect 2991 2103 3029 2137
rect 3063 2103 3101 2137
rect 3135 2103 3173 2137
rect 3207 2103 3245 2137
rect 3279 2103 3317 2137
rect 3351 2103 3389 2137
rect 3423 2103 3461 2137
rect 3495 2103 3533 2137
rect 3567 2103 3605 2137
rect 3639 2103 3677 2137
rect 3711 2103 3793 2137
rect 2503 2069 3793 2103
rect 2503 2035 2596 2069
rect 2630 2035 2669 2069
rect 2703 2035 2741 2069
rect 2775 2035 2813 2069
rect 2847 2035 2885 2069
rect 2919 2035 2957 2069
rect 2991 2035 3029 2069
rect 3063 2035 3101 2069
rect 3135 2035 3173 2069
rect 3207 2035 3245 2069
rect 3279 2035 3317 2069
rect 3351 2035 3389 2069
rect 3423 2035 3461 2069
rect 3495 2035 3533 2069
rect 3567 2035 3605 2069
rect 3639 2035 3677 2069
rect 3711 2035 3793 2069
rect 2503 2001 3793 2035
rect 2503 1967 2596 2001
rect 2630 1967 2669 2001
rect 2703 1967 2741 2001
rect 2775 1967 2813 2001
rect 2847 1967 2885 2001
rect 2919 1967 2957 2001
rect 2991 1967 3029 2001
rect 3063 1967 3101 2001
rect 3135 1967 3173 2001
rect 3207 1967 3245 2001
rect 3279 1967 3317 2001
rect 3351 1967 3389 2001
rect 3423 1967 3461 2001
rect 3495 1967 3533 2001
rect 3567 1967 3605 2001
rect 3639 1967 3677 2001
rect 3711 1967 3793 2001
rect 6283 841 6375 865
rect 6283 807 6307 841
rect 6341 807 6375 841
rect 6283 773 6375 807
rect 6283 739 6307 773
rect 6341 739 6375 773
rect 6283 705 6375 739
rect 6283 671 6307 705
rect 6341 671 6375 705
rect 6283 637 6375 671
rect 6283 603 6307 637
rect 6341 603 6375 637
rect 6283 569 6375 603
rect 6283 535 6307 569
rect 6341 535 6375 569
rect 6283 501 6375 535
rect 6283 467 6307 501
rect 6341 467 6375 501
rect 6283 433 6375 467
rect 6283 399 6307 433
rect 6341 399 6375 433
rect 6283 365 6375 399
rect 6283 331 6307 365
rect 6341 331 6375 365
rect 6283 297 6375 331
rect 6283 263 6307 297
rect 6341 263 6375 297
rect 6283 229 6375 263
rect 6283 195 6307 229
rect 6341 195 6375 229
rect 6283 171 6375 195
<< mvnsubdiff >>
rect 4647 -100 4681 -76
rect 5798 -97 5822 -63
rect 5856 -97 5890 -63
rect 5924 -97 5958 -63
rect 5992 -97 6027 -63
rect 6061 -97 6085 -63
rect 4647 -170 4681 -134
rect 4647 -240 4681 -204
rect 4647 -298 4681 -274
<< psubdiffcont >>
rect 2596 2171 2630 2205
rect 2669 2171 2703 2205
rect 2741 2171 2775 2205
rect 2813 2171 2847 2205
rect 2885 2171 2919 2205
rect 2957 2171 2991 2205
rect 3029 2171 3063 2205
rect 3101 2171 3135 2205
rect 3173 2171 3207 2205
rect 3245 2171 3279 2205
rect 3317 2171 3351 2205
rect 3389 2171 3423 2205
rect 3461 2171 3495 2205
rect 3533 2171 3567 2205
rect 3605 2171 3639 2205
rect 3677 2171 3711 2205
rect 2596 2103 2630 2137
rect 2669 2103 2703 2137
rect 2741 2103 2775 2137
rect 2813 2103 2847 2137
rect 2885 2103 2919 2137
rect 2957 2103 2991 2137
rect 3029 2103 3063 2137
rect 3101 2103 3135 2137
rect 3173 2103 3207 2137
rect 3245 2103 3279 2137
rect 3317 2103 3351 2137
rect 3389 2103 3423 2137
rect 3461 2103 3495 2137
rect 3533 2103 3567 2137
rect 3605 2103 3639 2137
rect 3677 2103 3711 2137
rect 2596 2035 2630 2069
rect 2669 2035 2703 2069
rect 2741 2035 2775 2069
rect 2813 2035 2847 2069
rect 2885 2035 2919 2069
rect 2957 2035 2991 2069
rect 3029 2035 3063 2069
rect 3101 2035 3135 2069
rect 3173 2035 3207 2069
rect 3245 2035 3279 2069
rect 3317 2035 3351 2069
rect 3389 2035 3423 2069
rect 3461 2035 3495 2069
rect 3533 2035 3567 2069
rect 3605 2035 3639 2069
rect 3677 2035 3711 2069
rect 2596 1967 2630 2001
rect 2669 1967 2703 2001
rect 2741 1967 2775 2001
rect 2813 1967 2847 2001
rect 2885 1967 2919 2001
rect 2957 1967 2991 2001
rect 3029 1967 3063 2001
rect 3101 1967 3135 2001
rect 3173 1967 3207 2001
rect 3245 1967 3279 2001
rect 3317 1967 3351 2001
rect 3389 1967 3423 2001
rect 3461 1967 3495 2001
rect 3533 1967 3567 2001
rect 3605 1967 3639 2001
rect 3677 1967 3711 2001
rect 6307 807 6341 841
rect 6307 739 6341 773
rect 6307 671 6341 705
rect 6307 603 6341 637
rect 6307 535 6341 569
rect 6307 467 6341 501
rect 6307 399 6341 433
rect 6307 331 6341 365
rect 6307 263 6341 297
rect 6307 195 6341 229
<< mvnsubdiffcont >>
rect 5822 -97 5856 -63
rect 5890 -97 5924 -63
rect 5958 -97 5992 -63
rect 6027 -97 6061 -63
rect 4647 -134 4681 -100
rect 4647 -204 4681 -170
rect 4647 -274 4681 -240
<< poly >>
rect 5882 839 6002 865
rect 5882 651 6002 699
rect 5882 617 5926 651
rect 5960 617 6002 651
rect 5882 583 6002 617
rect 5882 549 5926 583
rect 5960 549 6002 583
rect 5882 501 6002 549
rect 5882 233 6002 301
rect 5882 7 6002 33
rect 3741 -249 3767 -129
rect 3907 -171 4105 -129
rect 3907 -205 3955 -171
rect 3989 -205 4023 -171
rect 4057 -205 4105 -171
rect 3907 -249 4105 -205
rect 4305 -249 4373 -129
rect 4573 -249 4599 -129
<< polycont >>
rect 5926 617 5960 651
rect 5926 549 5960 583
rect 3955 -205 3989 -171
rect 4023 -205 4057 -171
<< locali >>
rect 2537 2171 2596 2205
rect 2630 2171 2669 2205
rect 2703 2171 2741 2205
rect 2775 2171 2813 2205
rect 2847 2171 2885 2205
rect 2919 2171 2957 2205
rect 2991 2171 3029 2205
rect 3063 2171 3101 2205
rect 3135 2171 3173 2205
rect 3207 2171 3245 2205
rect 3279 2171 3317 2205
rect 3351 2171 3389 2205
rect 3423 2171 3461 2205
rect 3495 2171 3533 2205
rect 3567 2171 3605 2205
rect 3639 2171 3677 2205
rect 3711 2171 3759 2205
rect 2537 2137 3759 2171
rect 2537 2103 2596 2137
rect 2630 2103 2669 2137
rect 2703 2103 2741 2137
rect 2775 2103 2813 2137
rect 2847 2103 2885 2137
rect 2919 2103 2957 2137
rect 2991 2103 3029 2137
rect 3063 2103 3101 2137
rect 3135 2103 3173 2137
rect 3207 2103 3245 2137
rect 3279 2103 3317 2137
rect 3351 2103 3389 2137
rect 3423 2103 3461 2137
rect 3495 2103 3533 2137
rect 3567 2103 3605 2137
rect 3639 2103 3677 2137
rect 3711 2103 3759 2137
rect 2537 2069 3759 2103
rect 2537 2035 2596 2069
rect 2630 2035 2669 2069
rect 2703 2035 2741 2069
rect 2775 2035 2813 2069
rect 2847 2035 2885 2069
rect 2919 2035 2957 2069
rect 2991 2035 3029 2069
rect 3063 2035 3101 2069
rect 3135 2035 3173 2069
rect 3207 2035 3245 2069
rect 3279 2035 3317 2069
rect 3351 2035 3389 2069
rect 3423 2035 3461 2069
rect 3495 2035 3533 2069
rect 3567 2035 3605 2069
rect 3639 2035 3677 2069
rect 3711 2035 3759 2069
rect 2537 2001 3759 2035
rect 2537 1967 2596 2001
rect 2630 1967 2669 2001
rect 2703 1967 2741 2001
rect 2775 1999 2813 2001
rect 2780 1967 2813 1999
rect 2847 1967 2885 2001
rect 2919 1999 2957 2001
rect 2919 1967 2948 1999
rect 2991 1967 3029 2001
rect 3063 1967 3101 2001
rect 3135 1999 3173 2001
rect 3163 1967 3173 1999
rect 3207 1967 3245 2001
rect 3279 1999 3317 2001
rect 3279 1967 3314 1999
rect 3351 1967 3389 2001
rect 3423 1967 3461 2001
rect 3495 1999 3533 2001
rect 3495 1967 3513 1999
rect 3567 1967 3605 2001
rect 3639 1967 3677 2001
rect 3711 1967 3759 2001
rect 2780 1965 2802 1967
rect 2982 1965 3004 1967
rect 3163 1965 3185 1967
rect 3348 1965 3370 1967
rect 3547 1965 3569 1967
rect 413 1188 448 1234
rect 5831 1136 5869 1170
rect 5197 768 5271 1086
rect 5197 734 5217 768
rect 5251 734 5271 768
rect 5197 696 5271 734
rect 5197 662 5217 696
rect 5251 662 5271 696
rect 4599 622 4653 632
rect 1491 601 1541 621
rect 1491 567 1498 601
rect 1532 567 1541 601
rect 1491 529 1541 567
rect 1491 495 1498 529
rect 1532 495 1541 529
rect 822 -63 1153 141
rect 1491 95 1541 495
rect 1643 601 1697 621
rect 1643 567 1653 601
rect 1687 567 1697 601
rect 1643 529 1697 567
rect 1643 495 1653 529
rect 1687 495 1697 529
rect 1643 95 1697 495
rect 4599 588 4610 622
rect 4644 588 4653 622
rect 4599 550 4653 588
rect 4599 516 4610 550
rect 4644 516 4653 550
rect 4599 95 4653 516
rect 4755 622 4804 632
rect 4755 588 4763 622
rect 4797 588 4804 622
rect 4755 550 4804 588
rect 4755 516 4763 550
rect 4797 516 4804 550
rect 4755 95 4804 516
rect 5197 267 5271 662
rect 5373 1062 5447 1086
rect 5373 1028 5393 1062
rect 5427 1028 5447 1062
rect 5373 990 5447 1028
rect 5373 956 5393 990
rect 5427 956 5447 990
rect 7050 1002 7084 1040
rect 5373 267 5447 956
rect 6284 841 6375 862
rect 5837 813 5871 828
rect 5837 745 5871 756
rect 5837 695 5871 711
rect 6013 813 6047 829
rect 6013 745 6047 779
rect 5703 617 5926 651
rect 5960 617 5976 651
rect 5703 583 5976 617
rect 5703 549 5926 583
rect 5960 549 5976 583
rect 6013 620 6047 711
rect 5703 160 5769 549
rect 6013 548 6047 586
rect 5630 154 5769 160
rect 5630 120 5642 154
rect 5676 120 5723 154
rect 5757 120 5769 154
rect 5630 114 5769 120
rect 5837 483 5935 499
rect 5871 449 5935 483
rect 5837 415 5935 449
rect 5871 375 5935 415
rect 5837 347 5935 375
rect 5871 303 5935 347
rect 5837 265 5935 303
rect 5871 231 5935 265
rect 5837 221 5935 231
rect 5871 187 5935 221
rect 5837 153 5935 187
rect 5871 119 5935 153
rect 1719 61 1817 95
rect 5837 85 5935 119
rect 5871 51 5935 85
rect 822 -97 834 -63
rect 868 -97 925 -63
rect 959 -97 1016 -63
rect 1050 -97 1107 -63
rect 1141 -97 1153 -63
rect 822 -100 1153 -97
rect 3517 -26 4573 -23
rect 3551 -60 3589 -26
rect 3623 -60 4573 -26
rect 3517 -84 4573 -60
rect 5837 -63 5935 51
rect 6013 483 6047 514
rect 6013 415 6047 449
rect 6013 347 6047 381
rect 6013 221 6047 313
rect 6013 153 6047 187
rect 6284 807 6307 841
rect 6341 807 6375 841
rect 6284 773 6375 807
rect 6284 739 6307 773
rect 6341 739 6375 773
rect 6284 705 6375 739
rect 6284 671 6307 705
rect 6341 671 6375 705
rect 6284 637 6375 671
rect 6284 603 6307 637
rect 6341 603 6375 637
rect 6284 569 6375 603
rect 6284 535 6307 569
rect 6341 535 6375 569
rect 6284 501 6375 535
rect 6284 467 6307 501
rect 6341 467 6375 501
rect 6284 433 6375 467
rect 6284 399 6307 433
rect 6341 399 6375 433
rect 6284 365 6375 399
rect 6284 331 6307 365
rect 6341 331 6375 365
rect 6284 297 6375 331
rect 6284 263 6307 297
rect 6341 263 6375 297
rect 6284 229 6375 263
rect 6284 195 6307 229
rect 6341 223 6375 229
rect 6341 204 8068 223
rect 8102 204 8142 238
rect 8176 204 8216 238
rect 8250 204 8290 238
rect 8324 204 8364 238
rect 8398 204 8438 238
rect 8472 204 8512 238
rect 8546 204 8586 238
rect 8620 204 8660 238
rect 8694 204 8734 238
rect 8768 204 8808 238
rect 8842 204 8882 238
rect 8916 204 8956 238
rect 8990 204 9030 238
rect 9064 204 9104 238
rect 9138 204 9178 238
rect 9212 204 9252 238
rect 9286 204 9326 238
rect 9360 204 9400 238
rect 9434 204 9475 238
rect 9509 204 9550 238
rect 9584 204 9625 238
rect 9659 204 9700 238
rect 9734 204 9775 238
rect 9809 204 9850 238
rect 9884 204 9925 238
rect 9959 204 10000 238
rect 10034 204 10075 238
rect 10109 204 12098 223
rect 6341 195 12098 204
rect 6284 185 12098 195
rect 6284 133 10419 185
rect 11067 133 12098 185
rect 6013 85 6047 119
rect 10133 53 10419 133
rect 6013 33 6047 51
rect 3517 -116 3793 -84
rect 3777 -118 3793 -116
rect 3827 -118 3861 -84
rect 3895 -118 4123 -84
rect 4157 -118 4191 -84
rect 4225 -118 4259 -84
rect 4293 -118 4385 -84
rect 4419 -118 4453 -84
rect 4487 -118 4521 -84
rect 4555 -118 4573 -84
rect 4647 -100 4681 -76
rect 5798 -97 5822 -63
rect 5856 -97 5890 -63
rect 5924 -97 5958 -63
rect 5992 -97 6027 -63
rect 6061 -97 6085 -63
rect 3955 -158 4430 -152
rect 3955 -171 4303 -158
rect 3989 -205 4023 -171
rect 4057 -192 4303 -171
rect 4337 -192 4384 -158
rect 4418 -192 4430 -158
rect 4057 -205 4430 -192
rect 3955 -226 4430 -205
rect 4647 -170 4681 -134
rect 4647 -233 4681 -204
rect 3777 -294 3793 -260
rect 3827 -294 3861 -260
rect 3895 -294 3911 -260
rect 3777 -428 3911 -294
rect 4107 -294 4123 -260
rect 4157 -294 4191 -260
rect 4225 -294 4259 -260
rect 4293 -294 4385 -260
rect 4419 -294 4453 -260
rect 4487 -294 4521 -260
rect 4555 -274 4647 -260
rect 4681 -267 4719 -233
rect 4555 -294 4681 -274
rect 4107 -333 4681 -294
<< viali >>
rect 2746 1967 2775 1999
rect 2775 1967 2780 1999
rect 2948 1967 2957 1999
rect 2957 1967 2982 1999
rect 3129 1967 3135 1999
rect 3135 1967 3163 1999
rect 3314 1967 3317 1999
rect 3317 1967 3348 1999
rect 3513 1967 3533 1999
rect 3533 1967 3547 1999
rect 2746 1965 2780 1967
rect 2948 1965 2982 1967
rect 3129 1965 3163 1967
rect 3314 1965 3348 1967
rect 3513 1965 3547 1967
rect 5797 1136 5831 1170
rect 5869 1136 5903 1170
rect 11785 1107 12323 1213
rect 5217 734 5251 768
rect 5217 662 5251 696
rect 1498 567 1532 601
rect 1498 495 1532 529
rect 1653 567 1687 601
rect 1653 495 1687 529
rect 4610 588 4644 622
rect 4610 516 4644 550
rect 4763 588 4797 622
rect 4763 516 4797 550
rect 5393 1028 5427 1062
rect 5393 956 5427 990
rect 7050 1040 7084 1074
rect 7050 968 7084 1002
rect 5837 828 5871 862
rect 5837 779 5871 790
rect 5837 756 5871 779
rect 6013 586 6047 620
rect 6013 514 6047 548
rect 5642 120 5676 154
rect 5723 120 5757 154
rect 5837 381 5871 409
rect 5837 375 5871 381
rect 5837 313 5871 337
rect 5837 303 5871 313
rect 5837 231 5871 265
rect 834 -97 868 -63
rect 925 -97 959 -63
rect 1016 -97 1050 -63
rect 1107 -97 1141 -63
rect 3517 -60 3551 -26
rect 3589 -60 3623 -26
rect 8068 204 8102 238
rect 8142 204 8176 238
rect 8216 204 8250 238
rect 8290 204 8324 238
rect 8364 204 8398 238
rect 8438 204 8472 238
rect 8512 204 8546 238
rect 8586 204 8620 238
rect 8660 204 8694 238
rect 8734 204 8768 238
rect 8808 204 8842 238
rect 8882 204 8916 238
rect 8956 204 8990 238
rect 9030 204 9064 238
rect 9104 204 9138 238
rect 9178 204 9212 238
rect 9252 204 9286 238
rect 9326 204 9360 238
rect 9400 204 9434 238
rect 9475 204 9509 238
rect 9550 204 9584 238
rect 9625 204 9659 238
rect 9700 204 9734 238
rect 9775 204 9809 238
rect 9850 204 9884 238
rect 9925 204 9959 238
rect 10000 204 10034 238
rect 10075 204 10109 238
rect 4303 -192 4337 -158
rect 4384 -192 4418 -158
rect 4647 -240 4681 -233
rect 4647 -267 4681 -240
rect 4719 -267 4753 -233
<< metal1 >>
rect -179 2033 -139 2235
rect 6041 2230 6762 2231
rect 6041 2178 6047 2230
rect 6099 2178 6112 2230
rect 6164 2178 6177 2230
rect 6229 2178 6242 2230
rect 6294 2178 6308 2230
rect 6360 2178 6374 2230
rect 6426 2178 6440 2230
rect 6492 2178 6506 2230
rect 6558 2178 6572 2230
rect 6624 2178 6638 2230
rect 6690 2178 6704 2230
rect 6756 2178 6762 2230
rect 6041 2160 6762 2178
rect 6041 2108 6047 2160
rect 6099 2108 6112 2160
rect 6164 2108 6177 2160
rect 6229 2108 6242 2160
rect 6294 2108 6308 2160
rect 6360 2108 6374 2160
rect 6426 2108 6440 2160
rect 6492 2108 6506 2160
rect 6558 2108 6572 2160
rect 6624 2108 6638 2160
rect 6690 2108 6704 2160
rect 6756 2108 6762 2160
rect 6041 2090 6762 2108
rect 6041 2038 6047 2090
rect 6099 2038 6112 2090
rect 6164 2038 6177 2090
rect 6229 2038 6242 2090
rect 6294 2038 6308 2090
rect 6360 2038 6374 2090
rect 6426 2038 6440 2090
rect 6492 2038 6506 2090
rect 6558 2038 6572 2090
rect 6624 2038 6638 2090
rect 6690 2038 6704 2090
rect 6756 2038 6762 2090
rect 6041 2037 6762 2038
rect 12524 2033 12564 2235
rect -179 1875 -139 2005
rect 104 1998 220 2004
rect 2734 1999 2814 2005
rect 2734 1965 2746 1999
rect 2780 1965 2814 1999
rect 2734 1959 2814 1965
rect 2936 1999 3016 2005
rect 2936 1965 2948 1999
rect 2982 1965 3016 1999
rect 2936 1959 3016 1965
rect 3117 1999 3197 2005
rect 3117 1965 3129 1999
rect 3163 1965 3197 1999
rect 3117 1959 3197 1965
rect 3302 1999 3382 2005
rect 3302 1965 3314 1999
rect 3348 1965 3382 1999
rect 3302 1959 3382 1965
rect 3501 1999 3581 2005
rect 3501 1965 3513 1999
rect 3547 1965 3581 1999
rect 3501 1959 3581 1965
rect 104 1876 220 1882
rect 3744 1953 3750 2005
rect 3802 1953 3822 2005
rect 3874 1953 3894 2005
rect 3946 1953 3966 2005
rect 4018 1953 4038 2005
rect 4090 1953 4110 2005
rect 4162 1953 4182 2005
rect 4234 1953 4253 2005
rect 4305 1953 4324 2005
rect 4376 1953 4382 2005
rect 3744 1927 4382 1953
rect 3744 1875 3750 1927
rect 3802 1875 3822 1927
rect 3874 1875 3894 1927
rect 3946 1875 3966 1927
rect 4018 1875 4038 1927
rect 4090 1875 4110 1927
rect 4162 1875 4182 1927
rect 4234 1875 4253 1927
rect 4305 1875 4324 1927
rect 4376 1875 4382 1927
rect 6678 1875 6718 2005
tri 6860 1959 6887 1986 se
rect 6887 1959 7866 1986
tri 6777 1876 6860 1959 se
rect 6860 1934 7866 1959
rect 6860 1876 6887 1934
tri 6887 1876 6945 1934 nw
tri 6776 1875 6777 1876 se
rect 6777 1875 6858 1876
tri 6748 1847 6776 1875 se
rect 6776 1847 6858 1875
tri 6858 1847 6887 1876 nw
rect 2094 1795 2100 1847
rect 2152 1795 2164 1847
rect 2216 1795 6806 1847
tri 6806 1795 6858 1847 nw
rect 1532 1706 1538 1758
rect 1590 1706 1602 1758
rect 1654 1706 1660 1758
tri 3953 1543 3999 1589 se
rect 3999 1583 6798 1589
rect 3999 1543 6746 1583
tri 3940 1530 3953 1543 se
rect 3953 1530 3999 1543
tri 3999 1530 4012 1543 nw
tri 6721 1530 6734 1543 ne
rect 6734 1531 6746 1543
rect 6734 1530 6798 1531
tri 3928 1518 3940 1530 se
rect 3940 1518 3987 1530
tri 3987 1518 3999 1530 nw
tri 6734 1518 6746 1530 ne
rect 6746 1519 6798 1530
tri 3905 1495 3928 1518 se
rect 3928 1495 3964 1518
tri 3964 1495 3987 1518 nw
tri 3881 1471 3905 1495 se
rect 3905 1471 3940 1495
tri 3940 1471 3964 1495 nw
tri 3853 1443 3881 1471 se
rect 3881 1443 3912 1471
tri 3912 1443 3940 1471 nw
rect 6226 1443 6232 1495
rect 6284 1443 6296 1495
rect 6348 1443 6368 1495
rect 6746 1461 6798 1467
tri 3825 1415 3853 1443 se
rect 3853 1415 3884 1443
tri 3884 1415 3912 1443 nw
tri 6240 1415 6268 1443 ne
tri 3822 1412 3825 1415 se
rect 3825 1412 3881 1415
tri 3881 1412 3884 1415 nw
tri 3798 1388 3822 1412 se
rect 3822 1388 3857 1412
tri 3857 1388 3881 1412 nw
tri 3591 1382 3597 1388 se
rect 3597 1382 3811 1388
tri 206 1361 227 1382 sw
tri 3570 1361 3591 1382 se
rect 3591 1361 3811 1382
tri 3531 1322 3570 1361 se
rect 3570 1342 3811 1361
tri 3811 1342 3857 1388 nw
rect 3570 1322 3597 1342
tri 3597 1322 3617 1342 nw
tri 3496 1287 3531 1322 se
rect 3531 1287 3562 1322
tri 3562 1287 3597 1322 nw
tri 6240 1287 6268 1315 se
rect 6268 1311 6368 1443
rect 7493 1432 7545 1484
tri 6368 1311 6372 1315 sw
rect 6268 1287 6372 1311
tri 6372 1287 6396 1311 sw
tri 6726 1287 6750 1311 se
rect 6750 1287 11121 1311
tri 3484 1275 3496 1287 se
rect 3496 1275 3531 1287
rect 2300 1256 2368 1275
tri 2368 1256 2387 1275 sw
tri 3465 1256 3484 1275 se
rect 3484 1256 3531 1275
tri 3531 1256 3562 1287 nw
rect 6267 1276 11121 1287
tri 11121 1276 11156 1311 sw
rect 6130 1268 11156 1276
rect 2300 1235 2387 1256
tri 2387 1235 2408 1256 sw
tri 3444 1235 3465 1256 se
rect 3465 1235 3510 1256
tri 3510 1235 3531 1256 nw
rect 6130 1235 6735 1268
tri 6735 1235 6768 1268 nw
tri 11107 1235 11140 1268 ne
rect 11140 1235 11156 1268
rect 2300 1219 2408 1235
tri 2408 1219 2424 1235 sw
tri 3428 1219 3444 1235 se
rect 3444 1219 3494 1235
tri 3494 1219 3510 1235 nw
tri 6130 1230 6135 1235 ne
rect 6135 1230 6267 1235
tri 6267 1230 6272 1235 nw
tri 11140 1230 11145 1235 ne
rect 11145 1230 11156 1235
tri 11145 1219 11156 1230 ne
tri 11156 1219 11213 1276 sw
rect 2300 1213 2424 1219
tri 2424 1213 2430 1219 sw
tri 3422 1213 3428 1219 se
rect 3428 1213 3488 1219
tri 3488 1213 3494 1219 nw
tri 11156 1213 11162 1219 ne
rect 11162 1213 12335 1219
rect 2300 1190 2430 1213
tri 2430 1190 2453 1213 sw
tri 3399 1190 3422 1213 se
rect 3422 1190 3465 1213
tri 3465 1190 3488 1213 nw
tri 11162 1190 11185 1213 ne
rect 11185 1190 11785 1213
rect 2300 1189 2453 1190
tri 2453 1189 2454 1190 sw
tri 3398 1189 3399 1190 se
rect 3399 1189 3464 1190
tri 3464 1189 3465 1190 nw
tri 11185 1189 11186 1190 ne
rect 11186 1189 11785 1190
rect 2300 1176 3451 1189
tri 3451 1176 3464 1189 nw
tri 11186 1176 11199 1189 ne
rect 11199 1176 11785 1189
rect 2300 1170 3445 1176
tri 3445 1170 3451 1176 nw
rect 5785 1170 6409 1176
rect 2300 1143 3418 1170
tri 3418 1143 3445 1170 nw
rect 5785 1136 5797 1170
rect 5831 1136 5869 1170
rect 5903 1136 6409 1170
rect 5785 1130 6409 1136
tri 6389 1116 6403 1130 ne
rect 6403 1116 6409 1130
tri 6409 1116 6469 1176 sw
tri 11748 1160 11764 1176 ne
rect 11764 1160 11785 1176
rect 6746 1154 6798 1160
tri 6403 1110 6409 1116 ne
rect 6409 1110 6469 1116
tri 6409 1107 6412 1110 ne
rect 6412 1107 6469 1110
tri 6469 1107 6478 1116 sw
tri 6412 1086 6433 1107 ne
rect 6433 1086 6478 1107
tri 6478 1086 6499 1107 sw
tri 11764 1151 11773 1160 ne
rect 6746 1090 6798 1102
rect 11773 1107 11785 1160
rect 12323 1107 12335 1213
rect 11773 1101 12335 1107
rect -179 884 -96 1086
rect 104 1080 220 1086
rect 156 1028 168 1080
rect 104 1011 220 1028
rect 156 959 168 1011
rect 104 942 220 959
rect 156 890 168 942
rect 104 884 220 890
rect 3744 1034 3750 1086
rect 3802 1034 3822 1086
rect 3874 1034 3894 1086
rect 3946 1034 3966 1086
rect 4018 1034 4038 1086
rect 4090 1034 4110 1086
rect 4162 1034 4182 1086
rect 4234 1034 4253 1086
rect 4305 1034 4324 1086
rect 4376 1034 4382 1086
tri 6433 1074 6445 1086 ne
rect 6445 1074 6499 1086
tri 6499 1074 6511 1086 sw
rect 3744 1011 4382 1034
rect 3744 959 3750 1011
rect 3802 959 3822 1011
rect 3874 959 3894 1011
rect 3946 959 3966 1011
rect 4018 959 4038 1011
rect 4090 959 4110 1011
rect 4162 959 4182 1011
rect 4234 959 4253 1011
rect 4305 959 4324 1011
rect 4376 959 4382 1011
rect 3744 936 4382 959
rect 5387 1062 5433 1074
rect 5387 1028 5393 1062
rect 5427 1028 5433 1062
tri 6445 1050 6469 1074 ne
rect 6469 1050 6511 1074
tri 6511 1050 6535 1074 sw
tri 6469 1040 6479 1050 ne
rect 6479 1040 6535 1050
tri 6535 1040 6545 1050 sw
rect 5387 990 5433 1028
tri 6479 1002 6517 1040 ne
rect 6517 1009 6545 1040
tri 6545 1009 6576 1040 sw
rect 6746 1032 6798 1038
rect 7044 1074 7090 1086
rect 7044 1040 7050 1074
rect 7084 1040 7090 1074
rect 6517 1002 6576 1009
tri 6576 1002 6583 1009 sw
tri 7037 1002 7044 1009 se
rect 7044 1002 7090 1040
rect 5387 956 5393 990
rect 5427 956 5433 990
tri 6517 984 6535 1002 ne
rect 6535 984 6583 1002
tri 6583 984 6601 1002 sw
tri 7019 984 7037 1002 se
rect 7037 984 7050 1002
tri 6535 968 6551 984 ne
rect 6551 968 7050 984
rect 7084 968 7090 1002
tri 6551 956 6563 968 ne
rect 6563 956 7090 968
rect 5387 944 5433 956
rect 3744 884 3750 936
rect 3802 884 3822 936
rect 3874 884 3894 936
rect 3946 884 3966 936
rect 4018 884 4038 936
rect 4090 884 4110 936
rect 4162 884 4182 936
rect 4234 884 4253 936
rect 4305 884 4324 936
rect 4376 884 4382 936
rect 5783 862 6114 942
rect 5783 828 5837 862
rect 5871 828 6114 862
rect 1703 756 1709 808
rect 1761 756 1773 808
rect 1825 756 2404 808
rect 2456 756 2468 808
rect 2520 756 2526 808
rect 5783 790 6114 828
rect 3746 726 5170 773
rect 5211 769 5257 780
rect 3746 717 3823 726
tri 3823 717 3832 726 nw
rect 5211 717 5217 769
rect 5269 717 5281 769
rect 5333 717 5339 769
rect 5783 756 5837 790
rect 5871 756 6114 790
rect 5783 727 6114 756
rect 7927 793 7933 845
rect 7985 793 8016 845
rect 8068 793 8099 845
rect 8151 793 8181 845
rect 8233 793 8263 845
rect 8315 793 8345 845
rect 8397 793 8403 845
rect 7927 770 8403 793
rect 7927 718 7933 770
rect 7985 718 8016 770
rect 8068 718 8099 770
rect 8151 718 8181 770
rect 8233 718 8263 770
rect 8315 718 8345 770
rect 8397 718 8403 770
rect 3746 696 3802 717
tri 3802 696 3823 717 nw
rect 5211 696 5257 717
rect 3746 625 3801 696
tri 3801 695 3802 696 nw
rect 5211 662 5217 696
rect 5251 662 5257 696
rect 5211 650 5257 662
rect 7927 695 8403 718
rect 7927 643 7933 695
rect 7985 643 8016 695
rect 8068 643 8099 695
rect 8151 643 8181 695
rect 8233 643 8263 695
rect 8315 643 8345 695
rect 8397 643 8403 695
rect 1492 601 1538 613
rect 1492 567 1498 601
rect 1532 567 1538 601
rect 1492 561 1538 567
rect 1590 561 1602 613
rect 1654 601 1693 613
rect 1687 567 1693 601
rect 1654 561 1693 567
rect 1492 535 1693 561
rect 1492 529 1538 535
rect 1492 495 1498 529
rect 1532 495 1538 529
rect 1492 483 1538 495
rect 1590 483 1602 535
rect 1654 529 1693 535
rect 1687 495 1693 529
rect 3746 573 3748 625
rect 3800 573 3801 625
rect 3746 561 3801 573
rect 3746 509 3748 561
rect 3800 509 3801 561
rect 3746 503 3801 509
rect 4333 629 4803 635
rect 6007 630 6053 632
rect 4385 622 4803 629
rect 4385 588 4610 622
rect 4644 588 4763 622
rect 4797 588 4803 622
rect 4385 577 4803 588
rect 4333 565 4803 577
rect 4385 550 4803 565
rect 4385 516 4610 550
rect 4644 516 4763 550
rect 4797 516 4803 550
rect 4385 513 4803 516
rect 4333 504 4803 513
rect 6004 624 6056 630
rect 6004 560 6056 572
rect 6004 502 6056 508
rect 1654 483 1693 495
rect 3065 239 3231 441
rect 5367 239 5434 441
tri 5823 413 5831 421 se
rect 5831 413 5878 421
tri 5878 413 5886 421 sw
rect 5782 412 6056 413
rect 5782 409 6180 412
rect 5782 375 5837 409
rect 5871 375 6180 409
rect 5782 358 6180 375
rect 5782 337 6050 358
rect 5782 303 5837 337
rect 5871 303 6050 337
rect 5782 265 6050 303
rect 738 211 5499 239
rect 5782 231 5837 265
rect 5871 242 6050 265
rect 6166 246 6180 358
rect 6166 242 6176 246
tri 6176 242 6180 246 nw
rect 8763 244 8841 643
tri 9777 281 9779 283 se
rect 9779 281 9934 643
tri 9740 244 9777 281 se
rect 9777 244 9934 281
tri 9934 244 9971 281 sw
rect 5871 239 6173 242
tri 6173 239 6176 242 nw
rect 5871 238 6172 239
tri 6172 238 6173 239 nw
rect 8056 238 10159 244
rect 5871 231 6153 238
rect 5782 219 6153 231
tri 6153 219 6172 238 nw
rect 5367 93 5434 211
rect 8056 204 8068 238
rect 8102 204 8142 238
rect 8176 204 8216 238
rect 8250 204 8290 238
rect 8324 204 8364 238
rect 8398 204 8438 238
rect 8472 204 8512 238
rect 8546 204 8586 238
rect 8620 204 8660 238
rect 8694 204 8734 238
rect 8768 204 8808 238
rect 8842 204 8882 238
rect 8916 204 8956 238
rect 8990 204 9030 238
rect 9064 204 9104 238
rect 9138 204 9178 238
rect 9212 204 9252 238
rect 9286 204 9326 238
rect 9360 204 9400 238
rect 9434 204 9475 238
rect 9509 204 9550 238
rect 9584 204 9625 238
rect 9659 204 9700 238
rect 9734 204 9775 238
rect 9809 204 9850 238
rect 9884 204 9925 238
rect 9959 204 10000 238
rect 10034 204 10075 238
rect 10109 223 10159 238
tri 10159 223 10180 244 sw
rect 10109 204 10180 223
rect 8056 198 10180 204
rect 5640 160 5646 166
rect 5630 154 5646 160
rect 5630 120 5642 154
rect 5630 114 5646 120
rect 5698 114 5710 166
rect 5762 160 5768 166
rect 5762 114 5769 160
tri 2748 10 2755 17 ne
rect 2755 10 2761 17
rect 3505 -23 3635 -20
tri 1939 -26 1942 -23 se
rect 1942 -26 3635 -23
tri 1908 -57 1939 -26 se
rect 1939 -57 3517 -26
rect 822 -60 1153 -57
tri 1905 -60 1908 -57 se
rect 1908 -60 3517 -57
rect 3551 -60 3589 -26
rect 3623 -60 3635 -26
rect 822 -63 3635 -60
rect 822 -97 834 -63
rect 868 -97 925 -63
rect 959 -97 1016 -63
rect 1050 -97 1107 -63
rect 1141 -66 1957 -63
tri 1957 -66 1960 -63 nw
rect 3505 -66 3635 -63
rect 1141 -97 1923 -66
rect 822 -100 1923 -97
tri 1923 -100 1957 -66 nw
rect 822 -103 1153 -100
tri 5626 -152 5640 -138 se
rect 5640 -152 5646 -138
rect 4291 -158 5646 -152
rect 4291 -192 4303 -158
rect 4337 -192 4384 -158
rect 4418 -190 5646 -158
rect 5698 -190 5710 -138
rect 5762 -190 5768 -138
rect 4418 -192 4430 -190
rect 4291 -198 4430 -192
rect 4291 -205 4329 -198
tri 3798 -221 3814 -205 se
rect 3814 -221 4329 -205
tri 3792 -227 3798 -221 se
rect 3798 -227 4329 -221
rect 4686 -227 4692 -221
tri 3786 -233 3792 -227 se
rect 3792 -233 4329 -227
tri 3770 -249 3786 -233 se
rect 3786 -243 4329 -233
rect 4635 -233 4692 -227
rect 4744 -233 4756 -221
rect 3786 -249 3814 -243
tri 3814 -249 3820 -243 nw
tri 3752 -267 3770 -249 se
rect 3770 -267 3796 -249
tri 3796 -267 3814 -249 nw
rect 4635 -267 4647 -233
rect 4681 -267 4692 -233
rect 4753 -267 4756 -233
tri 3746 -273 3752 -267 se
rect 3752 -273 3790 -267
tri 3790 -273 3796 -267 nw
rect 4635 -273 4692 -267
rect 4744 -273 4756 -267
rect 4808 -273 4814 -221
tri 3726 -293 3746 -273 se
rect 3746 -293 3770 -273
tri 3770 -293 3790 -273 nw
tri 3693 -326 3726 -293 se
rect 3084 -332 3136 -326
tri 3682 -337 3693 -326 se
rect 3693 -337 3726 -326
tri 3726 -337 3770 -293 nw
tri 3680 -339 3682 -337 se
rect 3682 -339 3724 -337
tri 3724 -339 3726 -337 nw
rect 3136 -377 3686 -339
tri 3686 -377 3724 -339 nw
rect 3084 -396 3136 -384
rect 3084 -454 3136 -448
<< via1 >>
rect 6047 2178 6099 2230
rect 6112 2178 6164 2230
rect 6177 2178 6229 2230
rect 6242 2178 6294 2230
rect 6308 2178 6360 2230
rect 6374 2178 6426 2230
rect 6440 2178 6492 2230
rect 6506 2178 6558 2230
rect 6572 2178 6624 2230
rect 6638 2178 6690 2230
rect 6704 2178 6756 2230
rect 6047 2108 6099 2160
rect 6112 2108 6164 2160
rect 6177 2108 6229 2160
rect 6242 2108 6294 2160
rect 6308 2108 6360 2160
rect 6374 2108 6426 2160
rect 6440 2108 6492 2160
rect 6506 2108 6558 2160
rect 6572 2108 6624 2160
rect 6638 2108 6690 2160
rect 6704 2108 6756 2160
rect 6047 2038 6099 2090
rect 6112 2038 6164 2090
rect 6177 2038 6229 2090
rect 6242 2038 6294 2090
rect 6308 2038 6360 2090
rect 6374 2038 6426 2090
rect 6440 2038 6492 2090
rect 6506 2038 6558 2090
rect 6572 2038 6624 2090
rect 6638 2038 6690 2090
rect 6704 2038 6756 2090
rect 104 1882 220 1998
rect 3750 1953 3802 2005
rect 3822 1953 3874 2005
rect 3894 1953 3946 2005
rect 3966 1953 4018 2005
rect 4038 1953 4090 2005
rect 4110 1953 4162 2005
rect 4182 1953 4234 2005
rect 4253 1953 4305 2005
rect 4324 1953 4376 2005
rect 3750 1875 3802 1927
rect 3822 1875 3874 1927
rect 3894 1875 3946 1927
rect 3966 1875 4018 1927
rect 4038 1875 4090 1927
rect 4110 1875 4162 1927
rect 4182 1875 4234 1927
rect 4253 1875 4305 1927
rect 4324 1875 4376 1927
rect 2100 1795 2152 1847
rect 2164 1795 2216 1847
rect 1538 1706 1590 1758
rect 1602 1706 1654 1758
rect 6746 1531 6798 1583
rect 6232 1443 6284 1495
rect 6296 1443 6348 1495
rect 6746 1467 6798 1519
rect 6746 1102 6798 1154
rect 104 1028 156 1080
rect 168 1028 220 1080
rect 104 959 156 1011
rect 168 959 220 1011
rect 104 890 156 942
rect 168 890 220 942
rect 3750 1034 3802 1086
rect 3822 1034 3874 1086
rect 3894 1034 3946 1086
rect 3966 1034 4018 1086
rect 4038 1034 4090 1086
rect 4110 1034 4162 1086
rect 4182 1034 4234 1086
rect 4253 1034 4305 1086
rect 4324 1034 4376 1086
rect 3750 959 3802 1011
rect 3822 959 3874 1011
rect 3894 959 3946 1011
rect 3966 959 4018 1011
rect 4038 959 4090 1011
rect 4110 959 4162 1011
rect 4182 959 4234 1011
rect 4253 959 4305 1011
rect 4324 959 4376 1011
rect 6746 1038 6798 1090
rect 3750 884 3802 936
rect 3822 884 3874 936
rect 3894 884 3946 936
rect 3966 884 4018 936
rect 4038 884 4090 936
rect 4110 884 4162 936
rect 4182 884 4234 936
rect 4253 884 4305 936
rect 4324 884 4376 936
rect 1709 756 1761 808
rect 1773 756 1825 808
rect 2404 756 2456 808
rect 2468 756 2520 808
rect 5217 768 5269 769
rect 5217 734 5251 768
rect 5251 734 5269 768
rect 5217 717 5269 734
rect 5281 717 5333 769
rect 7933 793 7985 845
rect 8016 793 8068 845
rect 8099 793 8151 845
rect 8181 793 8233 845
rect 8263 793 8315 845
rect 8345 793 8397 845
rect 7933 718 7985 770
rect 8016 718 8068 770
rect 8099 718 8151 770
rect 8181 718 8233 770
rect 8263 718 8315 770
rect 8345 718 8397 770
rect 7933 643 7985 695
rect 8016 643 8068 695
rect 8099 643 8151 695
rect 8181 643 8233 695
rect 8263 643 8315 695
rect 8345 643 8397 695
rect 1538 561 1590 613
rect 1602 601 1654 613
rect 1602 567 1653 601
rect 1653 567 1654 601
rect 1602 561 1654 567
rect 1538 483 1590 535
rect 1602 529 1654 535
rect 1602 495 1653 529
rect 1653 495 1654 529
rect 3748 573 3800 625
rect 3748 509 3800 561
rect 4333 577 4385 629
rect 4333 513 4385 565
rect 6004 620 6056 624
rect 6004 586 6013 620
rect 6013 586 6047 620
rect 6047 586 6056 620
rect 6004 572 6056 586
rect 6004 548 6056 560
rect 6004 514 6013 548
rect 6013 514 6047 548
rect 6047 514 6056 548
rect 6004 508 6056 514
rect 1602 483 1654 495
rect 6050 242 6166 358
rect 5646 154 5698 166
rect 5646 120 5676 154
rect 5676 120 5698 154
rect 5646 114 5698 120
rect 5710 154 5762 166
rect 5710 120 5723 154
rect 5723 120 5757 154
rect 5757 120 5762 154
rect 5710 114 5762 120
rect 5646 -190 5698 -138
rect 5710 -190 5762 -138
rect 4692 -233 4744 -221
rect 4692 -267 4719 -233
rect 4719 -267 4744 -233
rect 4692 -273 4744 -267
rect 4756 -273 4808 -221
rect 3084 -384 3136 -332
rect 3084 -448 3136 -396
<< metal2 >>
rect 6041 2230 6762 2231
rect 6041 2178 6047 2230
rect 6099 2228 6112 2230
rect 6164 2228 6177 2230
rect 6229 2228 6242 2230
rect 6294 2228 6308 2230
rect 6360 2228 6374 2230
rect 6426 2228 6440 2230
rect 6492 2228 6506 2230
rect 6558 2228 6572 2230
rect 6624 2228 6638 2230
rect 6690 2228 6704 2230
rect 6109 2178 6112 2228
rect 6360 2178 6373 2228
rect 6429 2178 6440 2228
rect 6690 2178 6694 2228
rect 6756 2178 6762 2230
rect 6041 2172 6053 2178
rect 6109 2172 6133 2178
rect 6189 2172 6213 2178
rect 6269 2172 6293 2178
rect 6349 2172 6373 2178
rect 6429 2172 6453 2178
rect 6509 2172 6533 2178
rect 6589 2172 6613 2178
rect 6669 2172 6694 2178
rect 6750 2172 6762 2178
rect 6041 2160 6762 2172
rect 6041 2108 6047 2160
rect 6099 2108 6112 2160
rect 6164 2108 6177 2160
rect 6229 2108 6242 2160
rect 6294 2108 6308 2160
rect 6360 2108 6374 2160
rect 6426 2108 6440 2160
rect 6492 2108 6506 2160
rect 6558 2108 6572 2160
rect 6624 2108 6638 2160
rect 6690 2108 6704 2160
rect 6756 2108 6762 2160
rect 6041 2096 6762 2108
rect 6041 2090 6053 2096
rect 6109 2090 6133 2096
rect 6189 2090 6213 2096
rect 6269 2090 6293 2096
rect 6349 2090 6373 2096
rect 6429 2090 6453 2096
rect 6509 2090 6533 2096
rect 6589 2090 6613 2096
rect 6669 2090 6694 2096
rect 6750 2090 6762 2096
rect 6041 2038 6047 2090
rect 6109 2040 6112 2090
rect 6360 2040 6373 2090
rect 6429 2040 6440 2090
rect 6690 2040 6694 2090
rect 6099 2038 6112 2040
rect 6164 2038 6177 2040
rect 6229 2038 6242 2040
rect 6294 2038 6308 2040
rect 6360 2038 6374 2040
rect 6426 2038 6440 2040
rect 6492 2038 6506 2040
rect 6558 2038 6572 2040
rect 6624 2038 6638 2040
rect 6690 2038 6704 2040
rect 6756 2038 6762 2090
rect 6041 2037 6762 2038
rect 104 1998 220 2004
rect 104 1080 220 1882
rect 3744 1953 3750 2005
rect 3802 1953 3822 2005
rect 3874 1953 3894 2005
rect 3946 1953 3966 2005
rect 4018 1953 4038 2005
rect 4090 1953 4110 2005
rect 4162 1953 4182 2005
rect 4234 1953 4253 2005
rect 4305 1953 4324 2005
rect 4376 1953 4382 2005
rect 3744 1927 4382 1953
rect 3744 1875 3750 1927
rect 3802 1875 3822 1927
rect 3874 1875 3894 1927
rect 3946 1875 3966 1927
rect 4018 1875 4038 1927
rect 4090 1875 4110 1927
rect 4162 1875 4182 1927
rect 4234 1875 4253 1927
rect 4305 1875 4324 1927
rect 4376 1875 4382 1927
rect 2094 1795 2100 1847
rect 2152 1795 2164 1847
rect 2216 1795 2222 1847
rect 156 1028 168 1080
rect 104 1011 220 1028
rect 156 959 168 1011
rect 104 942 220 959
rect 156 890 168 942
rect 104 884 220 890
rect 1532 1706 1538 1758
rect 1590 1706 1602 1758
rect 1654 1706 1660 1758
rect 1532 808 1660 1706
rect 3744 1086 4382 1875
rect 6746 1583 6798 1589
rect 6746 1519 6798 1531
rect 6226 1443 6232 1495
rect 6284 1443 6296 1495
rect 6348 1443 6354 1495
rect 3744 1034 3750 1086
rect 3802 1034 3822 1086
rect 3874 1034 3894 1086
rect 3946 1034 3966 1086
rect 4018 1034 4038 1086
rect 4090 1034 4110 1086
rect 4162 1034 4182 1086
rect 4234 1034 4253 1086
rect 4305 1034 4324 1086
rect 4376 1034 4382 1086
rect 3744 1011 4382 1034
rect 6746 1154 6798 1467
rect 6746 1090 6798 1102
rect 6746 1032 6798 1038
rect 3744 959 3750 1011
rect 3802 959 3822 1011
rect 3874 959 3894 1011
rect 3946 959 3966 1011
rect 4018 959 4038 1011
rect 4090 959 4110 1011
rect 4162 959 4182 1011
rect 4234 959 4253 1011
rect 4305 959 4324 1011
rect 4376 959 4382 1011
rect 3744 936 4382 959
rect 3744 884 3750 936
rect 3802 884 3822 936
rect 3874 884 3894 936
rect 3946 884 3966 936
rect 4018 884 4038 936
rect 4090 884 4110 936
rect 4162 884 4182 936
rect 4234 884 4253 936
rect 4305 884 4324 936
rect 4376 884 4382 936
tri 1660 808 1695 843 sw
rect 1532 756 1709 808
rect 1761 756 1773 808
rect 1825 756 1831 808
rect 2398 756 2404 808
rect 2456 756 2468 808
rect 2520 756 2526 808
rect 7927 793 7933 845
rect 7992 793 8016 845
rect 8091 793 8099 845
rect 8315 793 8332 845
rect 8397 793 8403 845
rect 7927 789 7936 793
rect 7992 789 8035 793
rect 8091 789 8134 793
rect 8190 789 8233 793
rect 8289 789 8332 793
rect 8388 789 8403 793
rect 7927 770 8403 789
rect 1532 717 1664 756
tri 1664 717 1703 756 nw
rect 1532 613 1660 717
tri 1660 713 1664 717 nw
rect 1532 561 1538 613
rect 1590 561 1602 613
rect 1654 561 1660 613
rect 1532 535 1660 561
rect 1532 483 1538 535
rect 1590 483 1602 535
rect 1654 483 1660 535
rect 2448 483 2500 756
rect 5211 717 5217 769
rect 5269 717 5281 769
rect 5333 756 5610 769
tri 5610 756 5623 769 sw
rect 5333 718 5623 756
tri 5623 718 5661 756 sw
rect 7927 718 7933 770
rect 7985 718 8016 770
rect 8068 718 8099 770
rect 8151 718 8181 770
rect 8233 718 8263 770
rect 8315 718 8345 770
rect 8397 718 8403 770
rect 5333 717 5661 718
tri 5588 713 5592 717 ne
rect 5592 713 5661 717
tri 5661 713 5666 718 sw
tri 5592 704 5601 713 ne
rect 5601 704 5666 713
tri 5666 704 5675 713 sw
tri 5601 695 5610 704 ne
rect 5610 695 5675 704
tri 5675 695 5684 704 sw
rect 7927 699 8403 718
rect 7927 695 7936 699
rect 7992 695 8035 699
rect 8091 695 8134 699
rect 8190 695 8233 699
rect 8289 695 8332 699
rect 8388 695 8403 699
tri 5610 643 5662 695 ne
rect 5662 643 5684 695
tri 5684 643 5736 695 sw
rect 7927 643 7933 695
rect 7992 643 8016 695
rect 8091 643 8099 695
rect 8315 643 8332 695
rect 8397 643 8403 695
tri 5662 635 5670 643 ne
rect 5670 635 5736 643
rect 3748 625 3800 631
tri 3732 573 3748 589 se
tri 3731 572 3732 573 se
rect 3732 572 3800 573
tri 3724 565 3731 572 se
rect 3731 565 3800 572
tri 3720 561 3724 565 se
rect 3724 561 3800 565
tri 3714 555 3720 561 se
rect 3720 555 3748 561
rect 3748 503 3800 509
rect 4333 629 4385 635
tri 5670 630 5675 635 ne
rect 5675 630 5736 635
tri 5736 630 5749 643 sw
tri 5675 624 5681 630 ne
rect 5681 624 6056 630
tri 5681 578 5727 624 ne
rect 5727 578 6004 624
rect 4333 565 4385 577
tri 5987 572 5993 578 ne
rect 5993 572 6004 578
tri 5993 561 6004 572 ne
tri 2500 483 2517 500 sw
tri 4316 483 4333 500 se
rect 4333 483 4385 513
rect 6004 560 6056 572
rect 6004 502 6056 508
rect 2448 478 2517 483
tri 2448 468 2458 478 ne
rect 2458 468 2517 478
tri 2517 468 2532 483 sw
tri 4301 468 4316 483 se
rect 4316 478 4385 483
rect 4316 468 4375 478
tri 4375 468 4385 478 nw
tri 2458 426 2500 468 ne
rect 2500 426 4333 468
tri 4333 426 4375 468 nw
tri 2500 423 2503 426 ne
rect 2503 423 4330 426
tri 4330 423 4333 426 nw
rect 6036 371 6190 375
rect 6036 280 6045 371
tri 4786 242 4824 280 se
rect 4824 242 6045 280
tri 4762 218 4786 242 se
rect 4786 235 6045 242
rect 6181 235 6190 371
rect 4786 221 6190 235
rect 4786 219 6042 221
rect 4786 218 4863 219
tri 4863 218 4864 219 nw
tri 2987 62 3004 79 se
rect 2987 10 3004 62
tri 2977 -17 3004 10 ne
rect 4762 -221 4822 218
tri 4822 177 4863 218 nw
rect 5640 114 5646 166
rect 5698 114 5710 166
rect 5762 114 5768 166
rect 5640 -138 5768 114
rect 5640 -190 5646 -138
rect 5698 -190 5710 -138
rect 5762 -190 5768 -138
rect 4686 -273 4692 -221
rect 4744 -273 4756 -221
rect 4808 -273 4822 -221
rect 3084 -332 3136 -326
rect 3084 -396 3136 -384
rect 2606 -493 2662 -430
tri 2662 -493 2672 -483 sw
rect 2606 -501 2672 -493
tri 2606 -537 2642 -501 ne
rect 2642 -537 2672 -501
tri 2672 -537 2716 -493 sw
tri 3040 -537 3084 -493 se
rect 3084 -515 3136 -448
rect 3084 -537 3114 -515
tri 3114 -537 3136 -515 nw
tri 2642 -557 2662 -537 ne
rect 2662 -557 3094 -537
tri 3094 -557 3114 -537 nw
tri 2662 -581 2686 -557 ne
rect 2686 -581 3070 -557
tri 3070 -581 3094 -557 nw
<< via2 >>
rect 6053 2178 6099 2228
rect 6099 2178 6109 2228
rect 6133 2178 6164 2228
rect 6164 2178 6177 2228
rect 6177 2178 6189 2228
rect 6213 2178 6229 2228
rect 6229 2178 6242 2228
rect 6242 2178 6269 2228
rect 6293 2178 6294 2228
rect 6294 2178 6308 2228
rect 6308 2178 6349 2228
rect 6373 2178 6374 2228
rect 6374 2178 6426 2228
rect 6426 2178 6429 2228
rect 6453 2178 6492 2228
rect 6492 2178 6506 2228
rect 6506 2178 6509 2228
rect 6533 2178 6558 2228
rect 6558 2178 6572 2228
rect 6572 2178 6589 2228
rect 6613 2178 6624 2228
rect 6624 2178 6638 2228
rect 6638 2178 6669 2228
rect 6694 2178 6704 2228
rect 6704 2178 6750 2228
rect 6053 2172 6109 2178
rect 6133 2172 6189 2178
rect 6213 2172 6269 2178
rect 6293 2172 6349 2178
rect 6373 2172 6429 2178
rect 6453 2172 6509 2178
rect 6533 2172 6589 2178
rect 6613 2172 6669 2178
rect 6694 2172 6750 2178
rect 6053 2090 6109 2096
rect 6133 2090 6189 2096
rect 6213 2090 6269 2096
rect 6293 2090 6349 2096
rect 6373 2090 6429 2096
rect 6453 2090 6509 2096
rect 6533 2090 6589 2096
rect 6613 2090 6669 2096
rect 6694 2090 6750 2096
rect 6053 2040 6099 2090
rect 6099 2040 6109 2090
rect 6133 2040 6164 2090
rect 6164 2040 6177 2090
rect 6177 2040 6189 2090
rect 6213 2040 6229 2090
rect 6229 2040 6242 2090
rect 6242 2040 6269 2090
rect 6293 2040 6294 2090
rect 6294 2040 6308 2090
rect 6308 2040 6349 2090
rect 6373 2040 6374 2090
rect 6374 2040 6426 2090
rect 6426 2040 6429 2090
rect 6453 2040 6492 2090
rect 6492 2040 6506 2090
rect 6506 2040 6509 2090
rect 6533 2040 6558 2090
rect 6558 2040 6572 2090
rect 6572 2040 6589 2090
rect 6613 2040 6624 2090
rect 6624 2040 6638 2090
rect 6638 2040 6669 2090
rect 6694 2040 6704 2090
rect 6704 2040 6750 2090
rect 7936 793 7985 845
rect 7985 793 7992 845
rect 8035 793 8068 845
rect 8068 793 8091 845
rect 8134 793 8151 845
rect 8151 793 8181 845
rect 8181 793 8190 845
rect 8233 793 8263 845
rect 8263 793 8289 845
rect 8332 793 8345 845
rect 8345 793 8388 845
rect 7936 789 7992 793
rect 8035 789 8091 793
rect 8134 789 8190 793
rect 8233 789 8289 793
rect 8332 789 8388 793
rect 7936 695 7992 699
rect 8035 695 8091 699
rect 8134 695 8190 699
rect 8233 695 8289 699
rect 8332 695 8388 699
rect 7936 643 7985 695
rect 7985 643 7992 695
rect 8035 643 8068 695
rect 8068 643 8091 695
rect 8134 643 8151 695
rect 8151 643 8181 695
rect 8181 643 8190 695
rect 8233 643 8263 695
rect 8263 643 8289 695
rect 8332 643 8345 695
rect 8345 643 8388 695
rect 6045 358 6181 371
rect 6045 242 6050 358
rect 6050 242 6166 358
rect 6166 242 6181 358
rect 6045 235 6181 242
<< metal3 >>
rect 6041 2233 6186 2235
rect 6041 2228 6755 2233
rect 6041 2172 6053 2228
rect 6109 2172 6133 2228
rect 6189 2172 6213 2228
rect 6269 2172 6293 2228
rect 6349 2172 6373 2228
rect 6429 2172 6453 2228
rect 6509 2172 6533 2228
rect 6589 2172 6613 2228
rect 6669 2172 6694 2228
rect 6750 2172 6755 2228
rect 6041 2096 6755 2172
rect 6041 2040 6053 2096
rect 6109 2040 6133 2096
rect 6189 2040 6213 2096
rect 6269 2040 6293 2096
rect 6349 2040 6373 2096
rect 6429 2040 6453 2096
rect 6509 2040 6533 2096
rect 6589 2040 6613 2096
rect 6669 2040 6694 2096
rect 6750 2040 6755 2096
rect 6041 2035 6755 2040
rect 6041 376 6186 2035
rect 7931 845 8393 850
rect 7931 789 7936 845
rect 7992 789 8035 845
rect 8091 789 8134 845
rect 8190 789 8233 845
rect 8289 789 8332 845
rect 8388 789 8393 845
rect 7931 699 8393 789
rect 7931 643 7936 699
rect 7992 643 8035 699
rect 8091 643 8134 699
rect 8190 643 8233 699
rect 8289 643 8332 699
rect 8388 643 8393 699
rect 7931 638 8393 643
rect 6040 371 6186 376
rect 6040 235 6045 371
rect 6181 235 6186 371
rect 6040 230 6186 235
use sky130_fd_io__gpio_dat_ls_ovtv2_i2c_fix  sky130_fd_io__gpio_dat_ls_ovtv2_i2c_fix_0
timestamp 1694700623
transform 1 0 0 0 -1 2339
box -179 23 3312 2414
use sky130_fd_io__gpio_dat_ls_ovtv2_i2c_fix_2  sky130_fd_io__gpio_dat_ls_ovtv2_i2c_fix_2_0
timestamp 1694700623
transform -1 0 6296 0 -1 2339
box -179 23 3312 2414
use sky130_fd_io__gpio_ovtv2_cclat_i2c_fix  sky130_fd_io__gpio_ovtv2_cclat_i2c_fix_0
timestamp 1694700623
transform 1 0 6330 0 1 0
box -133 145 6328 2367
use sky130_fd_io__hvsbt_inv_x1_i2c_fix  sky130_fd_io__hvsbt_inv_x1_i2c_fix_0
timestamp 1694700623
transform 1 0 5763 0 -1 983
box 107 226 240 751
use sky130_fd_io__hvsbt_inv_x1_i2c_fix_2  sky130_fd_io__hvsbt_inv_x1_i2c_fix_2_0
timestamp 1694700623
transform 0 1 3623 1 0 -368
box 118 283 240 751
use sky130_fd_pr__tpl1__example_55959141808367  sky130_fd_pr__tpl1__example_55959141808367_0
timestamp 1694700623
transform -1 0 6365 0 1 171
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1694700623
transform -1 0 5903 0 1 1136
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1694700623
transform 0 -1 7084 -1 0 1074
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808368  sky130_fd_pr__via_l1m1__example_55959141808368_0
timestamp 1694700623
transform -1 0 12323 0 1 1107
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1694700623
transform 0 -1 6798 -1 0 1160
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1694700623
transform 0 -1 6798 -1 0 1589
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1694700623
transform 0 -1 220 -1 0 2004
box 0 0 1 1
<< labels >>
flabel metal2 s 3084 -395 3136 -331 3 FreeSans 520 0 0 0 OD_I_H_N
port 1 nsew
flabel metal1 s 7816 1934 7866 1986 3 FreeSans 300 180 0 0 DRVHI_H
port 3 nsew
flabel metal1 s 7493 1432 7545 1484 3 FreeSans 300 180 0 0 DRVLO_H_N
port 4 nsew
flabel metal1 s 12524 2033 12564 2235 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 6678 1875 6718 2005 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s -179 1875 -139 2005 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s -179 2033 -139 2235 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s -179 884 -139 1086 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 4628 586 4661 624 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 7 nsew
flabel metal1 s 5367 93 5434 441 3 FreeSans 520 0 0 0 VPWR_KA
port 8 nsew
flabel metal1 s 11926 1134 12003 1187 3 FreeSans 520 0 0 0 PD_DIS_H
port 9 nsew
flabel locali s 413 1188 448 1234 3 FreeSans 300 0 0 0 OE_H
port 2 nsew
flabel comment s 5990 1188 5990 1188 0 FreeSans 300 0 0 0 PU_DIS_H
flabel comment s 6309 1264 6309 1264 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 8460 1291 8460 1291 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 10075 1294 10075 1294 0 FreeSans 300 0 0 0 PD_DIS_H
flabel comment s 6363 1491 6363 1491 0 FreeSans 300 0 0 0 OE_H_N
<< properties >>
string GDS_END 36840028
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36806626
<< end >>
