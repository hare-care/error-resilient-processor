magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal1 >>
rect 6867 95 7067 195
rect 5242 -7 5540 74
<< metal2 >>
rect 316 38458 2258 38490
rect 316 12482 339 38458
rect 2235 12482 2258 38458
rect 316 12450 2258 12482
rect 13868 14551 14780 14576
rect 13868 12495 13896 14551
rect 14752 12495 14780 14551
rect 13868 12470 14780 12495
rect 316 10913 2258 10944
rect 316 2297 339 10913
rect 2235 2297 2258 10913
rect 13868 10904 14780 10936
rect 316 2266 2258 2297
rect 11514 4085 13669 4095
rect 3372 1036 3526 2009
rect 3372 287 4215 1036
rect 100 0 4215 287
rect 10707 715 11164 1901
rect 11514 1069 11523 4085
rect 13659 1069 13669 4085
rect 11514 1059 13669 1069
rect 13868 1088 13896 10904
rect 14752 1088 14780 10904
rect 13868 1056 14780 1088
rect 3372 -7 4215 0
rect 6888 -7 8888 58
rect 10707 -7 14940 715
<< via2 >>
rect 339 12482 2235 38458
rect 13896 12495 14752 14551
rect 339 2297 2235 10913
rect 11523 1069 13659 4085
rect 13896 1088 14752 10904
<< metal3 >>
rect 316 38458 2258 38490
rect 316 12482 339 38458
rect 2235 12482 2258 38458
rect 4215 18474 4822 18525
rect 4215 17930 4286 18474
rect 4750 17930 4822 18474
rect 9498 18461 10372 18510
rect 9498 17997 9543 18461
rect 10327 17997 10372 18461
rect 4215 17880 4822 17930
rect 6994 17890 7723 17952
rect 9498 17949 10372 17997
rect 5193 17556 5929 17609
rect 5193 16932 5249 17556
rect 5873 16932 5929 17556
rect 5193 16880 5929 16932
rect 6994 16866 7046 17890
rect 7670 16866 7723 17890
rect 6994 16804 7723 16866
rect 8628 17627 9586 17685
rect 8628 16923 8675 17627
rect 9539 16923 9586 17627
rect 8628 16865 9586 16923
rect 5272 16652 7324 16704
rect 5272 13708 5346 16652
rect 7250 13708 7324 16652
rect 7696 16676 9748 16728
rect 7696 15434 7770 16676
rect 7526 14364 7770 15434
tri 7526 14214 7676 14364 ne
rect 7676 13890 7770 14364
rect 5272 13656 7324 13708
rect 7696 13732 7770 13890
rect 9674 15434 9748 16676
rect 9674 15358 9774 15434
tri 9774 15358 9850 15434 sw
rect 9674 13890 9850 15358
rect 13868 14551 14780 14576
rect 9674 13732 9748 13890
rect 7696 13680 9748 13732
rect 316 12450 2258 12482
rect 13868 12495 13896 14551
rect 14752 12495 14780 14551
rect 13868 12470 14780 12495
rect 316 10913 2258 10944
rect 316 2297 339 10913
rect 2235 2297 2258 10913
rect 13868 10904 14780 10936
rect 316 2266 2258 2297
rect 11514 4085 13669 4095
rect 11514 1069 11523 4085
rect 13659 1069 13669 4085
rect 11514 1059 13669 1069
rect 13868 1088 13896 10904
rect 14752 1088 14780 10904
rect 13868 1056 14780 1088
rect 98 339 4900 862
rect 100 -7 4900 339
rect 5200 -7 7374 918
rect 7676 -7 9850 918
rect 10151 -7 14940 862
<< via3 >>
rect 4286 17930 4750 18474
rect 9543 17997 10327 18461
rect 5249 16932 5873 17556
rect 7046 16866 7670 17890
rect 8675 16923 9539 17627
rect 5346 13708 7250 16652
rect 7770 13732 9674 16676
<< metal4 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 4255 18474 4782 18485
rect 4255 17930 4286 18474
rect 4750 17930 4782 18474
rect 9538 18461 10332 18470
rect 9538 17997 9543 18461
rect 10327 17997 10332 18461
rect 9538 17989 10332 17997
rect 4255 17920 4782 17930
rect 7034 17890 7683 17912
rect 5233 17556 5889 17569
rect 5233 16932 5249 17556
rect 5873 16932 5889 17556
rect 5233 16920 5889 16932
rect 7034 16866 7046 17890
rect 7670 16866 7683 17890
rect 8668 17627 9546 17645
rect 8668 16923 8675 17627
rect 9539 16923 9546 17627
rect 8668 16905 9546 16923
rect 7034 16844 7683 16866
rect 7736 16676 9708 16688
rect 5312 16652 7284 16664
rect 5312 13708 5346 16652
rect 7250 13708 7284 16652
rect 7736 13732 7770 16676
rect 9674 13732 9708 16676
rect 7736 13720 9708 13732
rect 5312 13696 7284 13708
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10874 254 10940
rect 14746 10874 15000 10940
rect 0 10218 254 10814
rect 14746 10218 15000 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 254 9862
rect 14746 9266 15000 9862
rect 0 9140 254 9206
rect 14746 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 254 3270
rect 14746 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 0 254 1090
rect 14746 0 15000 1090
<< metal5 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 6339 32546 10468 33417
rect 0 13600 254 18590
rect 14746 13600 15000 18590
rect 0 12430 254 13280
rect 14746 12430 15000 13280
rect 0 11260 254 12110
rect 14746 11260 15000 12110
rect 0 9140 254 10940
rect 14746 9140 15000 10940
rect 0 7930 254 8820
rect 14746 7930 15000 8820
rect 0 6960 254 7610
rect 14746 6960 15000 7610
rect 0 5990 254 6640
rect 14746 5990 15000 6640
rect 0 4780 254 5670
rect 14746 4780 15000 5670
rect 0 3570 254 4460
rect 14746 3570 15000 4460
rect 0 2600 254 3250
rect 14746 2600 15000 3250
rect 0 1390 254 2280
rect 14746 1390 15000 2280
rect 0 20 254 1070
rect 14746 20 15000 1070
use sky130_fd_io__overlay_vssio_lvc  sky130_fd_io__overlay_vssio_lvc_0
timestamp 1694700623
transform 1 0 0 0 1 -7
box 0 7 15000 39600
use sky130_fd_io__top_ground_lvc_wpad  sky130_fd_io__top_ground_lvc_wpad_2
timestamp 1694700623
transform 1 0 0 0 1 -7
box 0 0 15000 39600
<< labels >>
flabel metal4 s 0 10218 254 10814 3 FreeSans 650 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 14746 10218 15000 10814 3 FreeSans 650 180 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 0 9266 254 9862 3 FreeSans 650 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal4 s 14746 9266 15000 9862 3 FreeSans 650 180 0 0 AMUXBUS_B
port 2 nsew
flabel metal5 s 6339 32546 10468 33417 0 FreeSans 2500 0 0 0 VSSIO_PAD
port 3 nsew
flabel metal4 s 0 6940 254 7630 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal4 s 0 10874 254 10940 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal4 s 0 9922 254 10158 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal4 s 0 9140 254 9206 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal4 s 14746 6940 15000 7630 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal4 s 14746 9140 15000 9206 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal4 s 14746 10874 15000 10940 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal4 s 14746 9922 15000 10158 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal5 s 0 6961 254 7610 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal5 s 0 9140 254 10940 3 FreeSans 650 0 0 0 VSSA
port 4 nsew
flabel metal5 s 14746 6961 15000 7610 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal5 s 14746 9140 15000 10940 3 FreeSans 650 180 0 0 VSSA
port 4 nsew
flabel metal4 s 0 2580 193 3270 3 FreeSans 650 0 0 0 VDDA
port 5 nsew
flabel metal4 s 14807 2580 15000 3270 3 FreeSans 650 180 0 0 VDDA
port 5 nsew
flabel metal5 s 0 2600 193 3250 3 FreeSans 650 0 0 0 VDDA
port 5 nsew
flabel metal5 s 14807 2600 15000 3250 3 FreeSans 650 180 0 0 VDDA
port 5 nsew
flabel metal4 s 0 5970 254 6660 3 FreeSans 650 0 0 0 VSWITCH
port 6 nsew
flabel metal4 s 14746 5970 15000 6660 3 FreeSans 650 180 0 0 VSWITCH
port 6 nsew
flabel metal5 s 0 5990 254 6640 3 FreeSans 650 0 0 0 VSWITCH
port 6 nsew
flabel metal5 s 14746 5990 15000 6640 3 FreeSans 650 180 0 0 VSWITCH
port 6 nsew
flabel metal4 s 0 12410 254 13300 3 FreeSans 650 0 0 0 VDDIO_Q
port 7 nsew
flabel metal4 s 14746 12410 15000 13300 3 FreeSans 650 180 0 0 VDDIO_Q
port 7 nsew
flabel metal5 s 0 12430 254 13280 3 FreeSans 650 0 0 0 VDDIO_Q
port 7 nsew
flabel metal5 s 14746 12430 15000 13280 3 FreeSans 650 180 0 0 VDDIO_Q
port 7 nsew
flabel metal4 s 0 0 254 1090 3 FreeSans 650 0 0 0 VCCHIB
port 8 nsew
flabel metal4 s 14746 0 15000 1090 3 FreeSans 650 180 0 0 VCCHIB
port 8 nsew
flabel metal5 s 0 20 254 1070 3 FreeSans 650 0 0 0 VCCHIB
port 8 nsew
flabel metal5 s 14746 20 15000 1070 3 FreeSans 650 180 0 0 VCCHIB
port 8 nsew
flabel metal4 s 0 13600 254 18593 3 FreeSans 650 0 0 0 VDDIO
port 9 nsew
flabel metal4 s 0 3550 254 4480 3 FreeSans 650 0 0 0 VDDIO
port 9 nsew
flabel metal4 s 14746 13600 15000 18593 3 FreeSans 650 180 0 0 VDDIO
port 9 nsew
flabel metal4 s 14746 3550 15000 4480 3 FreeSans 650 180 0 0 VDDIO
port 9 nsew
flabel metal5 s 0 3570 254 4460 3 FreeSans 650 0 0 0 VDDIO
port 9 nsew
flabel metal5 s 0 13600 254 18590 3 FreeSans 650 0 0 0 VDDIO
port 9 nsew
flabel metal5 s 14746 3570 15000 4460 3 FreeSans 650 180 0 0 VDDIO
port 9 nsew
flabel metal5 s 14746 13600 15000 18590 3 FreeSans 650 180 0 0 VDDIO
port 9 nsew
flabel metal4 s 0 1370 254 2300 3 FreeSans 650 0 0 0 VCCD
port 10 nsew
flabel metal4 s 14746 1370 15000 2300 3 FreeSans 650 180 0 0 VCCD
port 10 nsew
flabel metal5 s 0 1390 254 2280 3 FreeSans 650 0 0 0 VCCD
port 10 nsew
flabel metal5 s 14746 1390 15000 2280 3 FreeSans 650 180 0 0 VCCD
port 10 nsew
flabel metal4 s 0 4760 254 5690 3 FreeSans 650 0 0 0 VSSIO
port 11 nsew
flabel metal4 s 0 34750 254 39593 3 FreeSans 650 0 0 0 VSSIO
port 11 nsew
flabel metal4 s 14746 34750 15000 39593 3 FreeSans 650 180 0 0 VSSIO
port 11 nsew
flabel metal4 s 14746 4760 15000 5690 3 FreeSans 650 180 0 0 VSSIO
port 11 nsew
flabel metal5 s 0 4780 254 5670 3 FreeSans 650 0 0 0 VSSIO
port 11 nsew
flabel metal5 s 14746 4780 15000 5670 3 FreeSans 650 180 0 0 VSSIO
port 11 nsew
flabel metal3 s 100 -7 4900 862 0 FreeSans 2500 0 0 0 VSSIO
port 11 nsew
flabel metal3 s 10151 -7 14940 862 0 FreeSans 5000 0 0 0 VSSIO
port 11 nsew
flabel metal4 s 0 7910 254 8840 3 FreeSans 650 0 0 0 VSSD
port 12 nsew
flabel metal4 s 14746 7910 15000 8840 3 FreeSans 650 180 0 0 VSSD
port 12 nsew
flabel metal5 s 0 7930 254 8820 3 FreeSans 650 0 0 0 VSSD
port 12 nsew
flabel metal5 s 14746 7930 15000 8820 3 FreeSans 650 180 0 0 VSSD
port 12 nsew
flabel metal4 s 0 11240 254 12130 3 FreeSans 650 0 0 0 VSSIO_Q
port 13 nsew
flabel metal4 s 14746 11240 15000 12130 3 FreeSans 650 180 0 0 VSSIO_Q
port 13 nsew
flabel metal5 s 0 11260 254 12110 3 FreeSans 650 0 0 0 VSSIO_Q
port 13 nsew
flabel metal5 s 14746 11260 15000 12110 3 FreeSans 650 180 0 0 VSSIO_Q
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 15000 39593
string GDS_END 2025834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 1037644
<< end >>
