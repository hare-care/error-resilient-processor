magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< locali >>
rect 199 1548 207 1582
rect 241 1548 279 1582
rect 313 1548 351 1582
rect 385 1548 423 1582
rect 457 1548 495 1582
rect 529 1548 567 1582
rect 601 1548 639 1582
rect 673 1548 711 1582
rect 745 1548 783 1582
rect 817 1548 855 1582
rect 889 1548 927 1582
rect 961 1548 999 1582
rect 1033 1548 1071 1582
rect 1105 1548 1143 1582
rect 1177 1548 1215 1582
rect 1249 1548 1287 1582
rect 1321 1548 1359 1582
rect 1393 1548 1431 1582
rect 1465 1548 1503 1582
rect 1537 1548 1575 1582
rect 1609 1548 1647 1582
rect 1681 1548 1719 1582
rect 1753 1548 1761 1582
rect 199 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1761 54
<< viali >>
rect 207 1548 241 1582
rect 279 1548 313 1582
rect 351 1548 385 1582
rect 423 1548 457 1582
rect 495 1548 529 1582
rect 567 1548 601 1582
rect 639 1548 673 1582
rect 711 1548 745 1582
rect 783 1548 817 1582
rect 855 1548 889 1582
rect 927 1548 961 1582
rect 999 1548 1033 1582
rect 1071 1548 1105 1582
rect 1143 1548 1177 1582
rect 1215 1548 1249 1582
rect 1287 1548 1321 1582
rect 1359 1548 1393 1582
rect 1431 1548 1465 1582
rect 1503 1548 1537 1582
rect 1575 1548 1609 1582
rect 1647 1548 1681 1582
rect 1719 1548 1753 1582
rect 207 20 241 54
rect 279 20 313 54
rect 351 20 385 54
rect 423 20 457 54
rect 495 20 529 54
rect 567 20 601 54
rect 639 20 673 54
rect 711 20 745 54
rect 783 20 817 54
rect 855 20 889 54
rect 927 20 961 54
rect 999 20 1033 54
rect 1071 20 1105 54
rect 1143 20 1177 54
rect 1215 20 1249 54
rect 1287 20 1321 54
rect 1359 20 1393 54
rect 1431 20 1465 54
rect 1503 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1681 54
rect 1719 20 1753 54
<< obsli1 >>
rect 48 1466 82 1514
rect 48 1394 82 1432
rect 48 1322 82 1360
rect 48 1250 82 1288
rect 48 1178 82 1216
rect 48 1106 82 1144
rect 48 1034 82 1072
rect 48 962 82 1000
rect 48 890 82 928
rect 48 818 82 856
rect 48 746 82 784
rect 48 674 82 712
rect 48 602 82 640
rect 48 530 82 568
rect 48 458 82 496
rect 48 386 82 424
rect 48 314 82 352
rect 48 242 82 280
rect 48 170 82 208
rect 48 88 82 136
rect 183 88 217 1514
rect 339 88 373 1514
rect 495 88 529 1514
rect 651 88 685 1514
rect 807 88 841 1514
rect 963 88 997 1514
rect 1119 88 1153 1514
rect 1275 88 1309 1514
rect 1431 88 1465 1514
rect 1587 88 1621 1514
rect 1743 88 1777 1514
rect 1878 1466 1912 1514
rect 1878 1394 1912 1432
rect 1878 1322 1912 1360
rect 1878 1250 1912 1288
rect 1878 1178 1912 1216
rect 1878 1106 1912 1144
rect 1878 1034 1912 1072
rect 1878 962 1912 1000
rect 1878 890 1912 928
rect 1878 818 1912 856
rect 1878 746 1912 784
rect 1878 674 1912 712
rect 1878 602 1912 640
rect 1878 530 1912 568
rect 1878 458 1912 496
rect 1878 386 1912 424
rect 1878 314 1912 352
rect 1878 242 1912 280
rect 1878 170 1912 208
rect 1878 88 1912 136
<< obsli1c >>
rect 48 1432 82 1466
rect 48 1360 82 1394
rect 48 1288 82 1322
rect 48 1216 82 1250
rect 48 1144 82 1178
rect 48 1072 82 1106
rect 48 1000 82 1034
rect 48 928 82 962
rect 48 856 82 890
rect 48 784 82 818
rect 48 712 82 746
rect 48 640 82 674
rect 48 568 82 602
rect 48 496 82 530
rect 48 424 82 458
rect 48 352 82 386
rect 48 280 82 314
rect 48 208 82 242
rect 48 136 82 170
rect 1878 1432 1912 1466
rect 1878 1360 1912 1394
rect 1878 1288 1912 1322
rect 1878 1216 1912 1250
rect 1878 1144 1912 1178
rect 1878 1072 1912 1106
rect 1878 1000 1912 1034
rect 1878 928 1912 962
rect 1878 856 1912 890
rect 1878 784 1912 818
rect 1878 712 1912 746
rect 1878 640 1912 674
rect 1878 568 1912 602
rect 1878 496 1912 530
rect 1878 424 1912 458
rect 1878 352 1912 386
rect 1878 280 1912 314
rect 1878 208 1912 242
rect 1878 136 1912 170
<< metal1 >>
rect 195 1582 1765 1602
rect 195 1548 207 1582
rect 241 1548 279 1582
rect 313 1548 351 1582
rect 385 1548 423 1582
rect 457 1548 495 1582
rect 529 1548 567 1582
rect 601 1548 639 1582
rect 673 1548 711 1582
rect 745 1548 783 1582
rect 817 1548 855 1582
rect 889 1548 927 1582
rect 961 1548 999 1582
rect 1033 1548 1071 1582
rect 1105 1548 1143 1582
rect 1177 1548 1215 1582
rect 1249 1548 1287 1582
rect 1321 1548 1359 1582
rect 1393 1548 1431 1582
rect 1465 1548 1503 1582
rect 1537 1548 1575 1582
rect 1609 1548 1647 1582
rect 1681 1548 1719 1582
rect 1753 1548 1765 1582
rect 195 1536 1765 1548
rect 36 1466 94 1497
rect 36 1432 48 1466
rect 82 1432 94 1466
rect 36 1394 94 1432
rect 36 1360 48 1394
rect 82 1360 94 1394
rect 36 1322 94 1360
rect 36 1288 48 1322
rect 82 1288 94 1322
rect 36 1250 94 1288
rect 36 1216 48 1250
rect 82 1216 94 1250
rect 36 1178 94 1216
rect 36 1144 48 1178
rect 82 1144 94 1178
rect 36 1106 94 1144
rect 36 1072 48 1106
rect 82 1072 94 1106
rect 36 1034 94 1072
rect 36 1000 48 1034
rect 82 1000 94 1034
rect 36 962 94 1000
rect 36 928 48 962
rect 82 928 94 962
rect 36 890 94 928
rect 36 856 48 890
rect 82 856 94 890
rect 36 818 94 856
rect 36 784 48 818
rect 82 784 94 818
rect 36 746 94 784
rect 36 712 48 746
rect 82 712 94 746
rect 36 674 94 712
rect 36 640 48 674
rect 82 640 94 674
rect 36 602 94 640
rect 36 568 48 602
rect 82 568 94 602
rect 36 530 94 568
rect 36 496 48 530
rect 82 496 94 530
rect 36 458 94 496
rect 36 424 48 458
rect 82 424 94 458
rect 36 386 94 424
rect 36 352 48 386
rect 82 352 94 386
rect 36 314 94 352
rect 36 280 48 314
rect 82 280 94 314
rect 36 242 94 280
rect 36 208 48 242
rect 82 208 94 242
rect 36 170 94 208
rect 36 136 48 170
rect 82 136 94 170
rect 36 105 94 136
rect 1866 1466 1924 1497
rect 1866 1432 1878 1466
rect 1912 1432 1924 1466
rect 1866 1394 1924 1432
rect 1866 1360 1878 1394
rect 1912 1360 1924 1394
rect 1866 1322 1924 1360
rect 1866 1288 1878 1322
rect 1912 1288 1924 1322
rect 1866 1250 1924 1288
rect 1866 1216 1878 1250
rect 1912 1216 1924 1250
rect 1866 1178 1924 1216
rect 1866 1144 1878 1178
rect 1912 1144 1924 1178
rect 1866 1106 1924 1144
rect 1866 1072 1878 1106
rect 1912 1072 1924 1106
rect 1866 1034 1924 1072
rect 1866 1000 1878 1034
rect 1912 1000 1924 1034
rect 1866 962 1924 1000
rect 1866 928 1878 962
rect 1912 928 1924 962
rect 1866 890 1924 928
rect 1866 856 1878 890
rect 1912 856 1924 890
rect 1866 818 1924 856
rect 1866 784 1878 818
rect 1912 784 1924 818
rect 1866 746 1924 784
rect 1866 712 1878 746
rect 1912 712 1924 746
rect 1866 674 1924 712
rect 1866 640 1878 674
rect 1912 640 1924 674
rect 1866 602 1924 640
rect 1866 568 1878 602
rect 1912 568 1924 602
rect 1866 530 1924 568
rect 1866 496 1878 530
rect 1912 496 1924 530
rect 1866 458 1924 496
rect 1866 424 1878 458
rect 1912 424 1924 458
rect 1866 386 1924 424
rect 1866 352 1878 386
rect 1912 352 1924 386
rect 1866 314 1924 352
rect 1866 280 1878 314
rect 1912 280 1924 314
rect 1866 242 1924 280
rect 1866 208 1878 242
rect 1912 208 1924 242
rect 1866 170 1924 208
rect 1866 136 1878 170
rect 1912 136 1924 170
rect 1866 105 1924 136
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< obsm1 >>
rect 174 105 226 1497
rect 330 105 382 1497
rect 486 105 538 1497
rect 642 105 694 1497
rect 798 105 850 1497
rect 954 105 1006 1497
rect 1110 105 1162 1497
rect 1266 105 1318 1497
rect 1422 105 1474 1497
rect 1578 105 1630 1497
rect 1734 105 1786 1497
<< metal2 >>
rect 10 1177 1950 1497
rect 10 481 1950 1121
rect 10 105 1950 425
<< labels >>
rlabel metal2 s 10 481 1950 1121 6 DRAIN
port 1 nsew
rlabel viali s 1719 1548 1753 1582 6 GATE
port 2 nsew
rlabel viali s 1719 20 1753 54 6 GATE
port 2 nsew
rlabel viali s 1647 1548 1681 1582 6 GATE
port 2 nsew
rlabel viali s 1647 20 1681 54 6 GATE
port 2 nsew
rlabel viali s 1575 1548 1609 1582 6 GATE
port 2 nsew
rlabel viali s 1575 20 1609 54 6 GATE
port 2 nsew
rlabel viali s 1503 1548 1537 1582 6 GATE
port 2 nsew
rlabel viali s 1503 20 1537 54 6 GATE
port 2 nsew
rlabel viali s 1431 1548 1465 1582 6 GATE
port 2 nsew
rlabel viali s 1431 20 1465 54 6 GATE
port 2 nsew
rlabel viali s 1359 1548 1393 1582 6 GATE
port 2 nsew
rlabel viali s 1359 20 1393 54 6 GATE
port 2 nsew
rlabel viali s 1287 1548 1321 1582 6 GATE
port 2 nsew
rlabel viali s 1287 20 1321 54 6 GATE
port 2 nsew
rlabel viali s 1215 1548 1249 1582 6 GATE
port 2 nsew
rlabel viali s 1215 20 1249 54 6 GATE
port 2 nsew
rlabel viali s 1143 1548 1177 1582 6 GATE
port 2 nsew
rlabel viali s 1143 20 1177 54 6 GATE
port 2 nsew
rlabel viali s 1071 1548 1105 1582 6 GATE
port 2 nsew
rlabel viali s 1071 20 1105 54 6 GATE
port 2 nsew
rlabel viali s 999 1548 1033 1582 6 GATE
port 2 nsew
rlabel viali s 999 20 1033 54 6 GATE
port 2 nsew
rlabel viali s 927 1548 961 1582 6 GATE
port 2 nsew
rlabel viali s 927 20 961 54 6 GATE
port 2 nsew
rlabel viali s 855 1548 889 1582 6 GATE
port 2 nsew
rlabel viali s 855 20 889 54 6 GATE
port 2 nsew
rlabel viali s 783 1548 817 1582 6 GATE
port 2 nsew
rlabel viali s 783 20 817 54 6 GATE
port 2 nsew
rlabel viali s 711 1548 745 1582 6 GATE
port 2 nsew
rlabel viali s 711 20 745 54 6 GATE
port 2 nsew
rlabel viali s 639 1548 673 1582 6 GATE
port 2 nsew
rlabel viali s 639 20 673 54 6 GATE
port 2 nsew
rlabel viali s 567 1548 601 1582 6 GATE
port 2 nsew
rlabel viali s 567 20 601 54 6 GATE
port 2 nsew
rlabel viali s 495 1548 529 1582 6 GATE
port 2 nsew
rlabel viali s 495 20 529 54 6 GATE
port 2 nsew
rlabel viali s 423 1548 457 1582 6 GATE
port 2 nsew
rlabel viali s 423 20 457 54 6 GATE
port 2 nsew
rlabel viali s 351 1548 385 1582 6 GATE
port 2 nsew
rlabel viali s 351 20 385 54 6 GATE
port 2 nsew
rlabel viali s 279 1548 313 1582 6 GATE
port 2 nsew
rlabel viali s 279 20 313 54 6 GATE
port 2 nsew
rlabel viali s 207 1548 241 1582 6 GATE
port 2 nsew
rlabel viali s 207 20 241 54 6 GATE
port 2 nsew
rlabel locali s 199 1548 1761 1582 6 GATE
port 2 nsew
rlabel locali s 199 20 1761 54 6 GATE
port 2 nsew
rlabel metal1 s 195 1536 1765 1602 6 GATE
port 2 nsew
rlabel metal1 s 195 0 1765 66 6 GATE
port 2 nsew
rlabel metal2 s 10 1177 1950 1497 6 SOURCE
port 3 nsew
rlabel metal2 s 10 105 1950 425 6 SOURCE
port 3 nsew
rlabel metal1 s 36 105 94 1497 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1866 105 1924 1497 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 0 1950 1602
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7790306
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7733854
<< end >>
