magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 1151 102 1251
rect -66 419 3079 1151
rect -66 377 102 419
rect 1883 341 3079 419
rect 3479 409 4339 1219
<< pwell >>
rect -26 1585 5018 1671
rect 449 1353 2439 1585
rect 2748 1353 3006 1585
rect 183 1217 3006 1353
rect 3534 1303 4297 1585
rect 183 43 1175 359
rect 3534 43 4012 325
rect -26 -43 5018 43
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2815 1645
rect 2849 1611 2911 1645
rect 2945 1611 3007 1645
rect 3041 1611 3103 1645
rect 3137 1611 3199 1645
rect 3233 1611 3295 1645
rect 3329 1611 3391 1645
rect 3425 1611 3487 1645
rect 3521 1611 3583 1645
rect 3617 1611 3679 1645
rect 3713 1611 3775 1645
rect 3809 1611 3871 1645
rect 3905 1611 3967 1645
rect 4001 1611 4063 1645
rect 4097 1611 4159 1645
rect 4193 1611 4255 1645
rect 4289 1611 4351 1645
rect 4385 1611 4447 1645
rect 4481 1611 4543 1645
rect 4577 1611 4639 1645
rect 4673 1611 4735 1645
rect 4769 1611 4831 1645
rect 4865 1611 4927 1645
rect 4961 1611 4992 1645
rect 72 831 106 1036
rect 0 797 31 831
rect 65 797 103 831
rect 212 428 256 1023
rect 524 428 568 1023
rect 212 384 568 428
rect 212 129 256 384
rect 524 129 568 384
rect 2863 1109 2997 1175
rect 1827 797 1853 831
rect 1887 797 1925 831
rect 1959 797 1985 831
rect 4214 1195 4280 1291
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 2815 1611 2849 1645
rect 2911 1611 2945 1645
rect 3007 1611 3041 1645
rect 3103 1611 3137 1645
rect 3199 1611 3233 1645
rect 3295 1611 3329 1645
rect 3391 1611 3425 1645
rect 3487 1611 3521 1645
rect 3583 1611 3617 1645
rect 3679 1611 3713 1645
rect 3775 1611 3809 1645
rect 3871 1611 3905 1645
rect 3967 1611 4001 1645
rect 4063 1611 4097 1645
rect 4159 1611 4193 1645
rect 4255 1611 4289 1645
rect 4351 1611 4385 1645
rect 4447 1611 4481 1645
rect 4543 1611 4577 1645
rect 4639 1611 4673 1645
rect 4735 1611 4769 1645
rect 4831 1611 4865 1645
rect 4927 1611 4961 1645
rect 31 797 65 831
rect 103 797 137 831
rect 1853 797 1887 831
rect 1925 797 1959 831
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
<< obsli1 >>
rect 212 1554 2977 1560
rect 212 1520 223 1554
rect 257 1520 319 1554
rect 353 1520 415 1554
rect 449 1520 511 1554
rect 545 1520 607 1554
rect 641 1520 703 1554
rect 737 1520 799 1554
rect 833 1520 895 1554
rect 929 1520 991 1554
rect 1025 1520 1087 1554
rect 1121 1520 1183 1554
rect 1217 1520 1279 1554
rect 1313 1520 1375 1554
rect 1409 1520 1471 1554
rect 1505 1520 1567 1554
rect 1601 1520 1663 1554
rect 1697 1520 1759 1554
rect 1793 1520 1855 1554
rect 1889 1520 1951 1554
rect 1985 1520 2047 1554
rect 2081 1520 2143 1554
rect 2177 1520 2239 1554
rect 2273 1520 2335 1554
rect 2369 1520 2431 1554
rect 2465 1520 2527 1554
rect 2561 1520 2623 1554
rect 2657 1520 2718 1554
rect 2752 1520 2815 1554
rect 2849 1520 2911 1554
rect 2945 1520 2977 1554
rect 212 1514 2977 1520
rect 212 1436 256 1514
rect 472 1441 516 1514
rect 212 1370 362 1436
rect 212 1239 256 1370
rect 368 1195 412 1305
rect 472 1239 517 1441
rect 714 1195 758 1441
rect 950 1239 994 1514
rect 1186 1195 1230 1441
rect 1422 1239 1466 1514
rect 1658 1195 1702 1441
rect 1894 1239 1938 1514
rect 2130 1195 2174 1441
rect 2366 1239 2410 1514
rect 2511 1195 2555 1305
rect 2667 1239 2711 1514
rect 368 1151 1304 1195
rect 367 925 413 1023
rect 331 919 449 925
rect 331 885 337 919
rect 371 885 409 919
rect 443 885 449 919
rect 331 879 449 885
rect 367 481 413 879
rect 679 925 725 1023
rect 643 919 761 925
rect 643 885 649 919
rect 683 885 721 919
rect 755 885 761 919
rect 643 879 761 885
rect 679 481 725 879
rect 790 439 834 751
rect 945 743 1062 751
rect 945 709 950 743
rect 984 709 1022 743
rect 1056 709 1062 743
rect 945 703 1062 709
rect 945 481 991 703
rect 367 97 413 331
rect 602 428 834 439
rect 1102 428 1146 751
rect 1260 503 1304 1151
rect 1572 1151 2555 1195
rect 2777 1151 2821 1373
rect 2933 1239 2977 1514
rect 3556 1543 4275 1549
rect 3556 1509 3564 1543
rect 3598 1509 3660 1543
rect 3694 1509 3756 1543
rect 3790 1509 3852 1543
rect 3886 1509 3948 1543
rect 3982 1509 4044 1543
rect 4078 1509 4140 1543
rect 4174 1509 4236 1543
rect 4270 1509 4275 1543
rect 3556 1503 4275 1509
rect 3556 1383 3622 1503
rect 3658 1349 3692 1469
rect 3738 1383 3804 1503
rect 3840 1349 3890 1469
rect 3558 1315 3890 1349
rect 3924 1325 3990 1503
rect 4037 1325 4087 1503
rect 4123 1325 4189 1469
rect 4225 1325 4275 1503
rect 1572 1047 1616 1151
rect 2618 1085 2821 1151
rect 3558 1171 3604 1315
rect 4123 1281 4180 1325
rect 3653 1237 4180 1281
rect 3653 1195 3988 1237
rect 3432 1161 3604 1171
rect 4034 1161 4084 1187
rect 3432 1127 3893 1161
rect 1469 981 1616 1047
rect 1415 613 1461 869
rect 1415 567 1487 613
rect 1572 567 1616 981
rect 2042 1007 2710 1051
rect 2042 749 2086 1007
rect 2005 743 2123 749
rect 2005 709 2011 743
rect 2045 709 2083 743
rect 2117 709 2123 743
rect 2005 703 2123 709
rect 1441 531 1487 567
rect 1260 437 1399 503
rect 1441 485 1561 531
rect 602 384 1146 428
rect 602 373 834 384
rect 679 97 725 331
rect 790 129 834 373
rect 945 97 991 331
rect 1102 129 1146 384
rect 1515 361 1561 485
rect 2042 403 2086 703
rect 2198 361 2242 945
rect 2354 749 2398 1007
rect 2317 743 2435 749
rect 2317 709 2323 743
rect 2357 709 2395 743
rect 2429 709 2435 743
rect 2317 703 2435 709
rect 2354 403 2398 703
rect 2510 361 2554 945
rect 2666 749 2710 1007
rect 2777 853 2821 1085
rect 2931 925 2977 1011
rect 2859 919 2977 925
rect 2859 885 2865 919
rect 2899 885 2937 919
rect 2971 885 2977 919
rect 2859 879 2977 885
rect 2931 853 2977 879
rect 2629 743 2747 749
rect 2629 709 2635 743
rect 2669 709 2707 743
rect 2741 709 2747 743
rect 2629 703 2747 709
rect 2666 403 2710 703
rect 1515 317 2554 361
rect 2793 313 2859 457
rect 3432 433 3476 1127
rect 3557 921 3607 1093
rect 3647 955 3713 1127
rect 3753 921 3787 1093
rect 3827 955 3893 1127
rect 3933 921 4084 1161
rect 4123 955 4180 1237
rect 4214 921 4280 1161
rect 3557 887 4280 921
rect 3933 847 4084 887
rect 3559 781 4084 847
rect 3933 741 4084 781
rect 3563 707 4084 741
rect 3563 467 3613 707
rect 3653 501 3719 673
rect 3759 535 3793 707
rect 3833 501 3899 673
rect 3939 648 4084 707
rect 3939 614 3960 648
rect 3994 614 4032 648
rect 4066 614 4084 648
rect 3939 604 4084 614
rect 3939 535 3989 604
rect 3653 467 3988 501
rect 3432 347 3893 433
rect 3942 313 3988 467
rect 2793 279 3988 313
rect 2793 269 3706 279
rect 3556 125 3622 235
rect 3656 159 3706 269
rect 3742 125 3808 245
rect 3854 159 3888 279
rect 3924 125 3990 245
rect 3556 119 3990 125
rect 367 91 485 97
rect 367 57 373 91
rect 407 57 445 91
rect 479 57 485 91
rect 367 51 485 57
rect 607 91 725 97
rect 607 57 613 91
rect 647 57 685 91
rect 719 57 725 91
rect 607 51 725 57
rect 909 91 1027 97
rect 909 57 915 91
rect 949 57 987 91
rect 1021 57 1027 91
rect 3556 85 3564 119
rect 3598 85 3660 119
rect 3694 85 3756 119
rect 3790 85 3852 119
rect 3886 85 3948 119
rect 3982 85 3990 119
rect 3556 79 3990 85
rect 909 51 1027 57
<< obsli1c >>
rect 223 1520 257 1554
rect 319 1520 353 1554
rect 415 1520 449 1554
rect 511 1520 545 1554
rect 607 1520 641 1554
rect 703 1520 737 1554
rect 799 1520 833 1554
rect 895 1520 929 1554
rect 991 1520 1025 1554
rect 1087 1520 1121 1554
rect 1183 1520 1217 1554
rect 1279 1520 1313 1554
rect 1375 1520 1409 1554
rect 1471 1520 1505 1554
rect 1567 1520 1601 1554
rect 1663 1520 1697 1554
rect 1759 1520 1793 1554
rect 1855 1520 1889 1554
rect 1951 1520 1985 1554
rect 2047 1520 2081 1554
rect 2143 1520 2177 1554
rect 2239 1520 2273 1554
rect 2335 1520 2369 1554
rect 2431 1520 2465 1554
rect 2527 1520 2561 1554
rect 2623 1520 2657 1554
rect 2718 1520 2752 1554
rect 2815 1520 2849 1554
rect 2911 1520 2945 1554
rect 337 885 371 919
rect 409 885 443 919
rect 649 885 683 919
rect 721 885 755 919
rect 950 709 984 743
rect 1022 709 1056 743
rect 3564 1509 3598 1543
rect 3660 1509 3694 1543
rect 3756 1509 3790 1543
rect 3852 1509 3886 1543
rect 3948 1509 3982 1543
rect 4044 1509 4078 1543
rect 4140 1509 4174 1543
rect 4236 1509 4270 1543
rect 2011 709 2045 743
rect 2083 709 2117 743
rect 2323 709 2357 743
rect 2395 709 2429 743
rect 2865 885 2899 919
rect 2937 885 2971 919
rect 2635 709 2669 743
rect 2707 709 2741 743
rect 3960 614 3994 648
rect 4032 614 4066 648
rect 373 57 407 91
rect 445 57 479 91
rect 613 57 647 91
rect 685 57 719 91
rect 915 57 949 91
rect 987 57 1021 91
rect 3564 85 3598 119
rect 3660 85 3694 119
rect 3756 85 3790 119
rect 3852 85 3886 119
rect 3948 85 3982 119
<< metal1 >>
rect 0 1645 4992 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2815 1645
rect 2849 1611 2911 1645
rect 2945 1611 3007 1645
rect 3041 1611 3103 1645
rect 3137 1611 3199 1645
rect 3233 1611 3295 1645
rect 3329 1611 3391 1645
rect 3425 1611 3487 1645
rect 3521 1611 3583 1645
rect 3617 1611 3679 1645
rect 3713 1611 3775 1645
rect 3809 1611 3871 1645
rect 3905 1611 3967 1645
rect 4001 1611 4063 1645
rect 4097 1611 4159 1645
rect 4193 1611 4255 1645
rect 4289 1611 4351 1645
rect 4385 1611 4447 1645
rect 4481 1611 4543 1645
rect 4577 1611 4639 1645
rect 4673 1611 4735 1645
rect 4769 1611 4831 1645
rect 4865 1611 4927 1645
rect 4961 1611 4992 1645
rect 0 1605 4992 1611
rect 0 1554 4992 1577
rect 0 1520 223 1554
rect 257 1520 319 1554
rect 353 1520 415 1554
rect 449 1520 511 1554
rect 545 1520 607 1554
rect 641 1520 703 1554
rect 737 1520 799 1554
rect 833 1520 895 1554
rect 929 1520 991 1554
rect 1025 1520 1087 1554
rect 1121 1520 1183 1554
rect 1217 1520 1279 1554
rect 1313 1520 1375 1554
rect 1409 1520 1471 1554
rect 1505 1520 1567 1554
rect 1601 1520 1663 1554
rect 1697 1520 1759 1554
rect 1793 1520 1855 1554
rect 1889 1520 1951 1554
rect 1985 1520 2047 1554
rect 2081 1520 2143 1554
rect 2177 1520 2239 1554
rect 2273 1520 2335 1554
rect 2369 1520 2431 1554
rect 2465 1520 2527 1554
rect 2561 1520 2623 1554
rect 2657 1520 2718 1554
rect 2752 1520 2815 1554
rect 2849 1520 2911 1554
rect 2945 1543 4992 1554
rect 2945 1520 3564 1543
rect 0 1509 3564 1520
rect 3598 1509 3660 1543
rect 3694 1509 3756 1543
rect 3790 1509 3852 1543
rect 3886 1509 3948 1543
rect 3982 1509 4044 1543
rect 4078 1509 4140 1543
rect 4174 1509 4236 1543
rect 4270 1509 4992 1543
rect 0 1503 4992 1509
rect 0 919 4992 939
rect 0 885 337 919
rect 371 885 409 919
rect 443 885 649 919
rect 683 885 721 919
rect 755 885 2865 919
rect 2899 885 2937 919
rect 2971 885 4992 919
rect 0 865 4992 885
rect 0 831 4992 837
rect 0 797 31 831
rect 65 797 103 831
rect 137 797 1853 831
rect 1887 797 1925 831
rect 1959 797 4992 831
rect 0 791 4992 797
rect 0 743 4992 763
rect 0 709 950 743
rect 984 709 1022 743
rect 1056 709 2011 743
rect 2045 709 2083 743
rect 2117 709 2323 743
rect 2357 709 2395 743
rect 2429 709 2635 743
rect 2669 709 2707 743
rect 2741 709 4992 743
rect 0 689 4992 709
rect 14 648 4978 661
rect 14 614 3960 648
rect 3994 614 4032 648
rect 4066 614 4978 648
rect 14 604 4978 614
rect 0 119 4992 125
rect 0 91 3564 119
rect 0 57 373 91
rect 407 57 445 91
rect 479 57 613 91
rect 647 57 685 91
rect 719 57 915 91
rect 949 57 987 91
rect 1021 85 3564 91
rect 3598 85 3660 119
rect 3694 85 3756 119
rect 3790 85 3852 119
rect 3886 85 3948 119
rect 3982 85 4992 119
rect 1021 57 4992 85
rect 0 51 4992 57
rect 0 17 4992 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
rect 0 -23 4992 -17
<< labels >>
rlabel locali s 4214 1195 4280 1291 6 A
port 1 nsew signal input
rlabel locali s 2863 1109 2997 1175 6 SLEEP_B
port 2 nsew signal input
rlabel metal1 s 14 604 4978 661 6 LVPWR
port 3 nsew power bidirectional
rlabel nwell s 3479 409 4339 1219 6 LVPWR
port 3 nsew power bidirectional
rlabel metal1 s 0 51 4992 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 1503 4992 1577 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 1605 4992 1651 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 3534 1303 4297 1585 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 183 1217 3006 1353 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2748 1353 3006 1585 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 449 1353 2439 1585 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 1585 5018 1671 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 4992 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 5018 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 3534 43 4012 325 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 183 43 1175 359 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4927 1611 4961 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4831 1611 4865 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4735 1611 4769 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4639 1611 4673 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4543 1611 4577 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4447 1611 4481 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4351 1611 4385 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4255 1611 4289 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4159 1611 4193 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4063 1611 4097 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3967 1611 4001 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3871 1611 3905 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3775 1611 3809 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3679 1611 3713 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3583 1611 3617 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3487 1611 3521 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3391 1611 3425 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3295 1611 3329 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3199 1611 3233 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3103 1611 3137 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 3007 1611 3041 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2911 1611 2945 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2815 1611 2849 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 1611 2753 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 1611 2657 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 1611 2561 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 1611 2465 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 1611 2369 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 1611 2273 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 1611 2177 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 1611 2081 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 1611 1985 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 1611 1889 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 1611 1793 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 1611 1697 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 1611 1601 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 1611 1505 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 1611 1409 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 1611 1313 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 1611 1217 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 1611 1121 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 1611 1025 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 1611 929 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 1611 833 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 1611 737 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 1611 641 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 1611 545 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 1611 449 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 1611 353 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 1611 257 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 1611 161 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 1611 65 1645 6 VNB
port 5 nsew ground bidirectional
rlabel locali s 0 1611 4992 1645 6 VNB
port 5 nsew ground bidirectional
rlabel viali s 4927 -17 4961 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4831 -17 4865 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4735 -17 4769 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4639 -17 4673 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4543 -17 4577 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4447 -17 4481 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4351 -17 4385 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4255 -17 4289 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4159 -17 4193 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 4063 -17 4097 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3967 -17 4001 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3871 -17 3905 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3775 -17 3809 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3679 -17 3713 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3583 -17 3617 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3487 -17 3521 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3391 -17 3425 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3295 -17 3329 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3199 -17 3233 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3103 -17 3137 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 3007 -17 3041 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2911 -17 2945 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2815 -17 2849 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 -17 2753 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 -17 2657 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 -17 2561 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 -17 2465 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 -17 2369 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 -17 2273 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 -17 2177 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 -17 929 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 -17 833 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 -17 737 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 -17 641 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 -17 545 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 -17 449 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 -17 353 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 -17 257 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 -17 161 17 8 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 -17 65 17 8 VNB
port 5 nsew ground bidirectional
rlabel locali s 0 -17 4992 17 8 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 4992 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s 1883 341 3079 419 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 102 419 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 419 3079 1151 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 1151 102 1251 6 VPB
port 6 nsew power bidirectional
rlabel viali s 1925 797 1959 831 6 VPB
port 6 nsew power bidirectional
rlabel viali s 1853 797 1887 831 6 VPB
port 6 nsew power bidirectional
rlabel locali s 1827 797 1985 831 6 VPB
port 6 nsew power bidirectional
rlabel viali s 103 797 137 831 6 VPB
port 6 nsew power bidirectional
rlabel viali s 31 797 65 831 6 VPB
port 6 nsew power bidirectional
rlabel locali s 0 797 137 831 6 VPB
port 6 nsew power bidirectional
rlabel locali s 72 831 106 1036 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 865 4992 939 6 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 689 4992 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 524 129 568 384 6 X
port 8 nsew signal output
rlabel locali s 212 129 256 384 6 X
port 8 nsew signal output
rlabel locali s 212 384 568 428 6 X
port 8 nsew signal output
rlabel locali s 524 428 568 1023 6 X
port 8 nsew signal output
rlabel locali s 212 428 256 1023 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 4992 1628
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 531566
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 478572
<< end >>
