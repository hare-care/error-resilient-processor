magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -36 679 514 1471
<< pwell >>
rect 128 25 330 225
<< scnmos >>
rect 214 51 244 199
<< ndiff >>
rect 154 51 214 199
rect 244 51 304 199
<< poly >>
rect 114 303 144 1113
rect 214 427 244 1113
rect 314 551 344 1113
rect 314 535 395 551
rect 314 501 345 535
rect 379 501 395 535
rect 314 485 395 501
rect 196 411 262 427
rect 196 377 212 411
rect 246 377 262 411
rect 196 361 262 377
rect 63 287 144 303
rect 63 253 79 287
rect 113 253 144 287
rect 63 237 144 253
rect 114 225 144 237
rect 214 199 244 361
rect 314 225 344 485
rect 214 25 244 51
<< polycont >>
rect 345 501 379 535
rect 212 377 246 411
rect 79 253 113 287
<< locali >>
rect 0 1397 478 1431
rect 62 1218 96 1397
rect 162 1184 196 1251
rect 262 1218 296 1397
rect 362 1184 396 1251
rect 162 1150 464 1184
rect 345 535 379 551
rect 345 485 379 501
rect 212 411 246 427
rect 212 361 246 377
rect 79 287 113 303
rect 79 237 113 253
rect 430 158 464 1150
rect 379 92 464 158
rect 62 17 96 92
rect 0 -17 478 17
use contact_12  contact_12_0
timestamp 1694700623
transform 1 0 329 0 1 485
box 0 0 1 1
use contact_12  contact_12_1
timestamp 1694700623
transform 1 0 196 0 1 361
box 0 0 1 1
use contact_12  contact_12_2
timestamp 1694700623
transform 1 0 63 0 1 237
box 0 0 1 1
use nmos_m1_w0_740_sactive_dactive  nmos_m1_w0_740_sactive_dactive_0
timestamp 1694700623
transform 1 0 154 0 1 51
box 0 0 1 1
use nmos_m1_w0_740_sactive_dli  nmos_m1_w0_740_sactive_dli_0
timestamp 1694700623
transform 1 0 254 0 1 51
box -26 -26 176 174
use nmos_m1_w0_740_sli_dactive  nmos_m1_w0_740_sli_dactive_0
timestamp 1694700623
transform 1 0 54 0 1 51
box -26 -26 176 174
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_0
timestamp 1694700623
transform 1 0 254 0 1 1139
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_1
timestamp 1694700623
transform 1 0 154 0 1 1139
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_2
timestamp 1694700623
transform 1 0 54 0 1 1139
box -59 -54 209 278
<< labels >>
rlabel locali s 447 1167 447 1167 4 Z
port 4 nsew
rlabel locali s 239 1414 239 1414 4 vdd
port 5 nsew
rlabel locali s 239 0 239 0 4 gnd
port 6 nsew
rlabel locali s 96 270 96 270 4 A
port 1 nsew
rlabel locali s 362 518 362 518 4 C
port 3 nsew
rlabel locali s 229 394 229 394 4 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 478 1414
string GDS_END 4086642
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4083920
<< end >>
