magic
tech sky130B
timestamp 1694700623
<< properties >>
string GDS_END 3204570
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3204310
<< end >>
