magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal2 >>
rect -7432 33185 -987 33506
rect -7432 32929 -7331 33185
rect -7075 32929 -6807 33185
rect -6551 32929 -6253 33185
rect -5997 32929 -5699 33185
rect -5443 32929 -5175 33185
rect -4919 32929 -4561 33185
rect -4305 32929 -4037 33185
rect -3781 32929 -3483 33185
rect -3227 32929 -2929 33185
rect -2673 32929 -2405 33185
rect -2149 32929 -987 33185
rect -7432 32691 -987 32929
rect -7432 32435 -7331 32691
rect -7075 32435 -6807 32691
rect -6551 32435 -6253 32691
rect -5997 32435 -5699 32691
rect -5443 32435 -5175 32691
rect -4919 32435 -4561 32691
rect -4305 32435 -4037 32691
rect -3781 32435 -3483 32691
rect -3227 32435 -2929 32691
rect -2673 32435 -2405 32691
rect -2149 32435 -987 32691
rect -7432 32077 -987 32435
rect -7432 31821 -7331 32077
rect -7075 31821 -6807 32077
rect -6551 31821 -6253 32077
rect -5997 31821 -5699 32077
rect -5443 31821 -5175 32077
rect -4919 31821 -4561 32077
rect -4305 31821 -4037 32077
rect -3781 31821 -3483 32077
rect -3227 31821 -2929 32077
rect -2673 31821 -2405 32077
rect -2149 31821 -987 32077
rect -7432 31583 -987 31821
rect -7432 31327 -7331 31583
rect -7075 31327 -6807 31583
rect -6551 31327 -6253 31583
rect -5997 31327 -5699 31583
rect -5443 31327 -5175 31583
rect -4919 31327 -4561 31583
rect -4305 31327 -4037 31583
rect -3781 31327 -3483 31583
rect -3227 31327 -2929 31583
rect -2673 31327 -2405 31583
rect -2149 31327 -987 31583
rect -7432 31006 -987 31327
tri -987 31006 1513 33506 sw
tri -2023 28004 979 31006 ne
rect 979 30504 1513 31006
tri 1513 30504 2015 31006 sw
rect 979 30183 7787 30504
rect 979 29927 2504 30183
rect 2760 29927 3028 30183
rect 3284 29927 3582 30183
rect 3838 29927 4136 30183
rect 4392 29927 4660 30183
rect 4916 29927 5274 30183
rect 5530 29927 5798 30183
rect 6054 29927 6352 30183
rect 6608 29927 6906 30183
rect 7162 29927 7430 30183
rect 7686 29927 7787 30183
rect 979 29689 7787 29927
rect 979 29433 2504 29689
rect 2760 29433 3028 29689
rect 3284 29433 3582 29689
rect 3838 29433 4136 29689
rect 4392 29433 4660 29689
rect 4916 29433 5274 29689
rect 5530 29433 5798 29689
rect 6054 29433 6352 29689
rect 6608 29433 6906 29689
rect 7162 29433 7430 29689
rect 7686 29433 7787 29689
rect 979 29075 7787 29433
rect 979 28819 2504 29075
rect 2760 28819 3028 29075
rect 3284 28819 3582 29075
rect 3838 28819 4136 29075
rect 4392 28819 4660 29075
rect 4916 28819 5274 29075
rect 5530 28819 5798 29075
rect 6054 28819 6352 29075
rect 6608 28819 6906 29075
rect 7162 28819 7430 29075
rect 7686 28819 7787 29075
rect 979 28581 7787 28819
rect 979 28325 2504 28581
rect 2760 28325 3028 28581
rect 3284 28325 3582 28581
rect 3838 28325 4136 28581
rect 4392 28325 4660 28581
rect 4916 28325 5274 28581
rect 5530 28325 5798 28581
rect 6054 28325 6352 28581
rect 6608 28325 6906 28581
rect 7162 28325 7430 28581
rect 7686 28325 7787 28581
rect 979 28004 7787 28325
rect -7432 27181 -987 27502
rect -7432 26925 -7331 27181
rect -7075 26925 -6807 27181
rect -6551 26925 -6253 27181
rect -5997 26925 -5699 27181
rect -5443 26925 -5175 27181
rect -4919 26925 -4561 27181
rect -4305 26925 -4037 27181
rect -3781 26925 -3483 27181
rect -3227 26925 -2929 27181
rect -2673 26925 -2405 27181
rect -2149 26925 -987 27181
rect -7432 26687 -987 26925
rect -7432 26431 -7331 26687
rect -7075 26431 -6807 26687
rect -6551 26431 -6253 26687
rect -5997 26431 -5699 26687
rect -5443 26431 -5175 26687
rect -4919 26431 -4561 26687
rect -4305 26431 -4037 26687
rect -3781 26431 -3483 26687
rect -3227 26431 -2929 26687
rect -2673 26431 -2405 26687
rect -2149 26431 -987 26687
rect -7432 26073 -987 26431
rect -7432 25817 -7331 26073
rect -7075 25817 -6807 26073
rect -6551 25817 -6253 26073
rect -5997 25817 -5699 26073
rect -5443 25817 -5175 26073
rect -4919 25817 -4561 26073
rect -4305 25817 -4037 26073
rect -3781 25817 -3483 26073
rect -3227 25817 -2929 26073
rect -2673 25817 -2405 26073
rect -2149 25817 -987 26073
rect -7432 25579 -987 25817
rect -7432 25323 -7331 25579
rect -7075 25323 -6807 25579
rect -6551 25323 -6253 25579
rect -5997 25323 -5699 25579
rect -5443 25323 -5175 25579
rect -4919 25323 -4561 25579
rect -4305 25323 -4037 25579
rect -3781 25323 -3483 25579
rect -3227 25323 -2929 25579
rect -2673 25323 -2405 25579
rect -2149 25323 -987 25579
rect -7432 25002 -987 25323
tri -987 25002 1513 27502 sw
tri -2023 22000 979 25002 ne
rect 979 24500 1513 25002
tri 1513 24500 2015 25002 sw
rect 979 24179 7787 24500
rect 979 23923 2504 24179
rect 2760 23923 3028 24179
rect 3284 23923 3582 24179
rect 3838 23923 4136 24179
rect 4392 23923 4660 24179
rect 4916 23923 5274 24179
rect 5530 23923 5798 24179
rect 6054 23923 6352 24179
rect 6608 23923 6906 24179
rect 7162 23923 7430 24179
rect 7686 23923 7787 24179
rect 979 23685 7787 23923
rect 979 23429 2504 23685
rect 2760 23429 3028 23685
rect 3284 23429 3582 23685
rect 3838 23429 4136 23685
rect 4392 23429 4660 23685
rect 4916 23429 5274 23685
rect 5530 23429 5798 23685
rect 6054 23429 6352 23685
rect 6608 23429 6906 23685
rect 7162 23429 7430 23685
rect 7686 23429 7787 23685
rect 979 23071 7787 23429
rect 979 22815 2504 23071
rect 2760 22815 3028 23071
rect 3284 22815 3582 23071
rect 3838 22815 4136 23071
rect 4392 22815 4660 23071
rect 4916 22815 5274 23071
rect 5530 22815 5798 23071
rect 6054 22815 6352 23071
rect 6608 22815 6906 23071
rect 7162 22815 7430 23071
rect 7686 22815 7787 23071
rect 979 22577 7787 22815
rect 979 22321 2504 22577
rect 2760 22321 3028 22577
rect 3284 22321 3582 22577
rect 3838 22321 4136 22577
rect 4392 22321 4660 22577
rect 4916 22321 5274 22577
rect 5530 22321 5798 22577
rect 6054 22321 6352 22577
rect 6608 22321 6906 22577
rect 7162 22321 7430 22577
rect 7686 22321 7787 22577
rect 979 22000 7787 22321
rect 19408 929 37508 1250
rect 19408 673 19552 929
rect 19808 673 20076 929
rect 20332 673 20630 929
rect 20886 673 37508 929
rect 19408 435 37508 673
rect 19408 179 19552 435
rect 19808 179 20076 435
rect 20332 179 20630 435
rect 20886 179 37508 435
rect 19408 -179 37508 179
rect 19408 -435 19552 -179
rect 19808 -435 20076 -179
rect 20332 -435 20630 -179
rect 20886 -435 37508 -179
rect 19408 -673 37508 -435
rect 19408 -929 19552 -673
rect 19808 -929 20076 -673
rect 20332 -929 20630 -673
rect 20886 -929 37508 -673
rect 19408 -1250 37508 -929
tri -2023 -28004 979 -25002 se
rect 979 -25324 7675 -25002
rect 979 -25580 2393 -25324
rect 2649 -25580 2917 -25324
rect 3173 -25580 3471 -25324
rect 3727 -25580 4025 -25324
rect 4281 -25580 4549 -25324
rect 4805 -25580 5163 -25324
rect 5419 -25580 5687 -25324
rect 5943 -25580 6241 -25324
rect 6497 -25580 6795 -25324
rect 7051 -25580 7319 -25324
rect 7575 -25580 7675 -25324
rect 979 -25818 7675 -25580
rect 979 -26074 2393 -25818
rect 2649 -26074 2917 -25818
rect 3173 -26074 3471 -25818
rect 3727 -26074 4025 -25818
rect 4281 -26074 4549 -25818
rect 4805 -26074 5163 -25818
rect 5419 -26074 5687 -25818
rect 5943 -26074 6241 -25818
rect 6497 -26074 6795 -25818
rect 7051 -26074 7319 -25818
rect 7575 -26074 7675 -25818
rect 979 -26432 7675 -26074
rect 979 -26688 2393 -26432
rect 2649 -26688 2917 -26432
rect 3173 -26688 3471 -26432
rect 3727 -26688 4025 -26432
rect 4281 -26688 4549 -26432
rect 4805 -26688 5163 -26432
rect 5419 -26688 5687 -26432
rect 5943 -26688 6241 -26432
rect 6497 -26688 6795 -26432
rect 7051 -26688 7319 -26432
rect 7575 -26688 7675 -26432
rect 979 -26926 7675 -26688
rect 979 -27182 2393 -26926
rect 2649 -27182 2917 -26926
rect 3173 -27182 3471 -26926
rect 3727 -27182 4025 -26926
rect 4281 -27182 4549 -26926
rect 4805 -27182 5163 -26926
rect 5419 -27182 5687 -26926
rect 5943 -27182 6241 -26926
rect 6497 -27182 6795 -26926
rect 7051 -27182 7319 -26926
rect 7575 -27182 7675 -26926
rect 979 -27502 7675 -27182
rect 979 -28004 1513 -27502
tri 1513 -28004 2015 -27502 nw
rect -7544 -28325 -987 -28004
rect -7544 -28581 -7444 -28325
rect -7188 -28581 -6920 -28325
rect -6664 -28581 -6366 -28325
rect -6110 -28581 -5812 -28325
rect -5556 -28581 -5288 -28325
rect -5032 -28581 -4674 -28325
rect -4418 -28581 -4150 -28325
rect -3894 -28581 -3596 -28325
rect -3340 -28581 -3042 -28325
rect -2786 -28581 -2518 -28325
rect -2262 -28581 -987 -28325
rect -7544 -28819 -987 -28581
rect -7544 -29075 -7444 -28819
rect -7188 -29075 -6920 -28819
rect -6664 -29075 -6366 -28819
rect -6110 -29075 -5812 -28819
rect -5556 -29075 -5288 -28819
rect -5032 -29075 -4674 -28819
rect -4418 -29075 -4150 -28819
rect -3894 -29075 -3596 -28819
rect -3340 -29075 -3042 -28819
rect -2786 -29075 -2518 -28819
rect -2262 -29075 -987 -28819
rect -7544 -29433 -987 -29075
rect -7544 -29689 -7444 -29433
rect -7188 -29689 -6920 -29433
rect -6664 -29689 -6366 -29433
rect -6110 -29689 -5812 -29433
rect -5556 -29689 -5288 -29433
rect -5032 -29689 -4674 -29433
rect -4418 -29689 -4150 -29433
rect -3894 -29689 -3596 -29433
rect -3340 -29689 -3042 -29433
rect -2786 -29689 -2518 -29433
rect -2262 -29689 -987 -29433
rect -7544 -29927 -987 -29689
rect -7544 -30183 -7444 -29927
rect -7188 -30183 -6920 -29927
rect -6664 -30183 -6366 -29927
rect -6110 -30183 -5812 -29927
rect -5556 -30183 -5288 -29927
rect -5032 -30183 -4674 -29927
rect -4418 -30183 -4150 -29927
rect -3894 -30183 -3596 -29927
rect -3340 -30183 -3042 -29927
rect -2786 -30183 -2518 -29927
rect -2262 -30183 -987 -29927
rect -7544 -30504 -987 -30183
tri -987 -30504 1513 -28004 nw
tri -2023 -34008 979 -31006 se
rect 979 -31326 7675 -31006
rect 979 -31582 2393 -31326
rect 2649 -31582 2917 -31326
rect 3173 -31582 3471 -31326
rect 3727 -31582 4025 -31326
rect 4281 -31582 4549 -31326
rect 4805 -31582 5163 -31326
rect 5419 -31582 5687 -31326
rect 5943 -31582 6241 -31326
rect 6497 -31582 6795 -31326
rect 7051 -31582 7319 -31326
rect 7575 -31582 7675 -31326
rect 979 -31820 7675 -31582
rect 979 -32076 2393 -31820
rect 2649 -32076 2917 -31820
rect 3173 -32076 3471 -31820
rect 3727 -32076 4025 -31820
rect 4281 -32076 4549 -31820
rect 4805 -32076 5163 -31820
rect 5419 -32076 5687 -31820
rect 5943 -32076 6241 -31820
rect 6497 -32076 6795 -31820
rect 7051 -32076 7319 -31820
rect 7575 -32076 7675 -31820
rect 979 -32434 7675 -32076
rect 979 -32690 2393 -32434
rect 2649 -32690 2917 -32434
rect 3173 -32690 3471 -32434
rect 3727 -32690 4025 -32434
rect 4281 -32690 4549 -32434
rect 4805 -32690 5163 -32434
rect 5419 -32690 5687 -32434
rect 5943 -32690 6241 -32434
rect 6497 -32690 6795 -32434
rect 7051 -32690 7319 -32434
rect 7575 -32690 7675 -32434
rect 979 -32928 7675 -32690
rect 979 -33184 2393 -32928
rect 2649 -33184 2917 -32928
rect 3173 -33184 3471 -32928
rect 3727 -33184 4025 -32928
rect 4281 -33184 4549 -32928
rect 4805 -33184 5163 -32928
rect 5419 -33184 5687 -32928
rect 5943 -33184 6241 -32928
rect 6497 -33184 6795 -32928
rect 7051 -33184 7319 -32928
rect 7575 -33184 7675 -32928
rect 979 -33506 7675 -33184
rect 979 -34008 1513 -33506
tri 1513 -34008 2015 -33506 nw
rect -7544 -34329 -987 -34008
rect -7544 -34585 -7444 -34329
rect -7188 -34585 -6920 -34329
rect -6664 -34585 -6366 -34329
rect -6110 -34585 -5812 -34329
rect -5556 -34585 -5288 -34329
rect -5032 -34585 -4674 -34329
rect -4418 -34585 -4150 -34329
rect -3894 -34585 -3596 -34329
rect -3340 -34585 -3042 -34329
rect -2786 -34585 -2518 -34329
rect -2262 -34585 -987 -34329
rect -7544 -34823 -987 -34585
rect -7544 -35079 -7444 -34823
rect -7188 -35079 -6920 -34823
rect -6664 -35079 -6366 -34823
rect -6110 -35079 -5812 -34823
rect -5556 -35079 -5288 -34823
rect -5032 -35079 -4674 -34823
rect -4418 -35079 -4150 -34823
rect -3894 -35079 -3596 -34823
rect -3340 -35079 -3042 -34823
rect -2786 -35079 -2518 -34823
rect -2262 -35079 -987 -34823
rect -7544 -35437 -987 -35079
rect -7544 -35693 -7444 -35437
rect -7188 -35693 -6920 -35437
rect -6664 -35693 -6366 -35437
rect -6110 -35693 -5812 -35437
rect -5556 -35693 -5288 -35437
rect -5032 -35693 -4674 -35437
rect -4418 -35693 -4150 -35437
rect -3894 -35693 -3596 -35437
rect -3340 -35693 -3042 -35437
rect -2786 -35693 -2518 -35437
rect -2262 -35693 -987 -35437
rect -7544 -35931 -987 -35693
rect -7544 -36187 -7444 -35931
rect -7188 -36187 -6920 -35931
rect -6664 -36187 -6366 -35931
rect -6110 -36187 -5812 -35931
rect -5556 -36187 -5288 -35931
rect -5032 -36187 -4674 -35931
rect -4418 -36187 -4150 -35931
rect -3894 -36187 -3596 -35931
rect -3340 -36187 -3042 -35931
rect -2786 -36187 -2518 -35931
rect -2262 -36187 -987 -35931
rect -7544 -36508 -987 -36187
tri -987 -36508 1513 -34008 nw
<< via2 >>
rect -7331 32929 -7075 33185
rect -6807 32929 -6551 33185
rect -6253 32929 -5997 33185
rect -5699 32929 -5443 33185
rect -5175 32929 -4919 33185
rect -4561 32929 -4305 33185
rect -4037 32929 -3781 33185
rect -3483 32929 -3227 33185
rect -2929 32929 -2673 33185
rect -2405 32929 -2149 33185
rect -7331 32435 -7075 32691
rect -6807 32435 -6551 32691
rect -6253 32435 -5997 32691
rect -5699 32435 -5443 32691
rect -5175 32435 -4919 32691
rect -4561 32435 -4305 32691
rect -4037 32435 -3781 32691
rect -3483 32435 -3227 32691
rect -2929 32435 -2673 32691
rect -2405 32435 -2149 32691
rect -7331 31821 -7075 32077
rect -6807 31821 -6551 32077
rect -6253 31821 -5997 32077
rect -5699 31821 -5443 32077
rect -5175 31821 -4919 32077
rect -4561 31821 -4305 32077
rect -4037 31821 -3781 32077
rect -3483 31821 -3227 32077
rect -2929 31821 -2673 32077
rect -2405 31821 -2149 32077
rect -7331 31327 -7075 31583
rect -6807 31327 -6551 31583
rect -6253 31327 -5997 31583
rect -5699 31327 -5443 31583
rect -5175 31327 -4919 31583
rect -4561 31327 -4305 31583
rect -4037 31327 -3781 31583
rect -3483 31327 -3227 31583
rect -2929 31327 -2673 31583
rect -2405 31327 -2149 31583
rect 2504 29927 2760 30183
rect 3028 29927 3284 30183
rect 3582 29927 3838 30183
rect 4136 29927 4392 30183
rect 4660 29927 4916 30183
rect 5274 29927 5530 30183
rect 5798 29927 6054 30183
rect 6352 29927 6608 30183
rect 6906 29927 7162 30183
rect 7430 29927 7686 30183
rect 2504 29433 2760 29689
rect 3028 29433 3284 29689
rect 3582 29433 3838 29689
rect 4136 29433 4392 29689
rect 4660 29433 4916 29689
rect 5274 29433 5530 29689
rect 5798 29433 6054 29689
rect 6352 29433 6608 29689
rect 6906 29433 7162 29689
rect 7430 29433 7686 29689
rect 2504 28819 2760 29075
rect 3028 28819 3284 29075
rect 3582 28819 3838 29075
rect 4136 28819 4392 29075
rect 4660 28819 4916 29075
rect 5274 28819 5530 29075
rect 5798 28819 6054 29075
rect 6352 28819 6608 29075
rect 6906 28819 7162 29075
rect 7430 28819 7686 29075
rect 2504 28325 2760 28581
rect 3028 28325 3284 28581
rect 3582 28325 3838 28581
rect 4136 28325 4392 28581
rect 4660 28325 4916 28581
rect 5274 28325 5530 28581
rect 5798 28325 6054 28581
rect 6352 28325 6608 28581
rect 6906 28325 7162 28581
rect 7430 28325 7686 28581
rect -7331 26925 -7075 27181
rect -6807 26925 -6551 27181
rect -6253 26925 -5997 27181
rect -5699 26925 -5443 27181
rect -5175 26925 -4919 27181
rect -4561 26925 -4305 27181
rect -4037 26925 -3781 27181
rect -3483 26925 -3227 27181
rect -2929 26925 -2673 27181
rect -2405 26925 -2149 27181
rect -7331 26431 -7075 26687
rect -6807 26431 -6551 26687
rect -6253 26431 -5997 26687
rect -5699 26431 -5443 26687
rect -5175 26431 -4919 26687
rect -4561 26431 -4305 26687
rect -4037 26431 -3781 26687
rect -3483 26431 -3227 26687
rect -2929 26431 -2673 26687
rect -2405 26431 -2149 26687
rect -7331 25817 -7075 26073
rect -6807 25817 -6551 26073
rect -6253 25817 -5997 26073
rect -5699 25817 -5443 26073
rect -5175 25817 -4919 26073
rect -4561 25817 -4305 26073
rect -4037 25817 -3781 26073
rect -3483 25817 -3227 26073
rect -2929 25817 -2673 26073
rect -2405 25817 -2149 26073
rect -7331 25323 -7075 25579
rect -6807 25323 -6551 25579
rect -6253 25323 -5997 25579
rect -5699 25323 -5443 25579
rect -5175 25323 -4919 25579
rect -4561 25323 -4305 25579
rect -4037 25323 -3781 25579
rect -3483 25323 -3227 25579
rect -2929 25323 -2673 25579
rect -2405 25323 -2149 25579
rect 2504 23923 2760 24179
rect 3028 23923 3284 24179
rect 3582 23923 3838 24179
rect 4136 23923 4392 24179
rect 4660 23923 4916 24179
rect 5274 23923 5530 24179
rect 5798 23923 6054 24179
rect 6352 23923 6608 24179
rect 6906 23923 7162 24179
rect 7430 23923 7686 24179
rect 2504 23429 2760 23685
rect 3028 23429 3284 23685
rect 3582 23429 3838 23685
rect 4136 23429 4392 23685
rect 4660 23429 4916 23685
rect 5274 23429 5530 23685
rect 5798 23429 6054 23685
rect 6352 23429 6608 23685
rect 6906 23429 7162 23685
rect 7430 23429 7686 23685
rect 2504 22815 2760 23071
rect 3028 22815 3284 23071
rect 3582 22815 3838 23071
rect 4136 22815 4392 23071
rect 4660 22815 4916 23071
rect 5274 22815 5530 23071
rect 5798 22815 6054 23071
rect 6352 22815 6608 23071
rect 6906 22815 7162 23071
rect 7430 22815 7686 23071
rect 2504 22321 2760 22577
rect 3028 22321 3284 22577
rect 3582 22321 3838 22577
rect 4136 22321 4392 22577
rect 4660 22321 4916 22577
rect 5274 22321 5530 22577
rect 5798 22321 6054 22577
rect 6352 22321 6608 22577
rect 6906 22321 7162 22577
rect 7430 22321 7686 22577
rect 19552 673 19808 929
rect 20076 673 20332 929
rect 20630 673 20886 929
rect 19552 179 19808 435
rect 20076 179 20332 435
rect 20630 179 20886 435
rect 19552 -435 19808 -179
rect 20076 -435 20332 -179
rect 20630 -435 20886 -179
rect 19552 -929 19808 -673
rect 20076 -929 20332 -673
rect 20630 -929 20886 -673
rect 2393 -25580 2649 -25324
rect 2917 -25580 3173 -25324
rect 3471 -25580 3727 -25324
rect 4025 -25580 4281 -25324
rect 4549 -25580 4805 -25324
rect 5163 -25580 5419 -25324
rect 5687 -25580 5943 -25324
rect 6241 -25580 6497 -25324
rect 6795 -25580 7051 -25324
rect 7319 -25580 7575 -25324
rect 2393 -26074 2649 -25818
rect 2917 -26074 3173 -25818
rect 3471 -26074 3727 -25818
rect 4025 -26074 4281 -25818
rect 4549 -26074 4805 -25818
rect 5163 -26074 5419 -25818
rect 5687 -26074 5943 -25818
rect 6241 -26074 6497 -25818
rect 6795 -26074 7051 -25818
rect 7319 -26074 7575 -25818
rect 2393 -26688 2649 -26432
rect 2917 -26688 3173 -26432
rect 3471 -26688 3727 -26432
rect 4025 -26688 4281 -26432
rect 4549 -26688 4805 -26432
rect 5163 -26688 5419 -26432
rect 5687 -26688 5943 -26432
rect 6241 -26688 6497 -26432
rect 6795 -26688 7051 -26432
rect 7319 -26688 7575 -26432
rect 2393 -27182 2649 -26926
rect 2917 -27182 3173 -26926
rect 3471 -27182 3727 -26926
rect 4025 -27182 4281 -26926
rect 4549 -27182 4805 -26926
rect 5163 -27182 5419 -26926
rect 5687 -27182 5943 -26926
rect 6241 -27182 6497 -26926
rect 6795 -27182 7051 -26926
rect 7319 -27182 7575 -26926
rect -7444 -28581 -7188 -28325
rect -6920 -28581 -6664 -28325
rect -6366 -28581 -6110 -28325
rect -5812 -28581 -5556 -28325
rect -5288 -28581 -5032 -28325
rect -4674 -28581 -4418 -28325
rect -4150 -28581 -3894 -28325
rect -3596 -28581 -3340 -28325
rect -3042 -28581 -2786 -28325
rect -2518 -28581 -2262 -28325
rect -7444 -29075 -7188 -28819
rect -6920 -29075 -6664 -28819
rect -6366 -29075 -6110 -28819
rect -5812 -29075 -5556 -28819
rect -5288 -29075 -5032 -28819
rect -4674 -29075 -4418 -28819
rect -4150 -29075 -3894 -28819
rect -3596 -29075 -3340 -28819
rect -3042 -29075 -2786 -28819
rect -2518 -29075 -2262 -28819
rect -7444 -29689 -7188 -29433
rect -6920 -29689 -6664 -29433
rect -6366 -29689 -6110 -29433
rect -5812 -29689 -5556 -29433
rect -5288 -29689 -5032 -29433
rect -4674 -29689 -4418 -29433
rect -4150 -29689 -3894 -29433
rect -3596 -29689 -3340 -29433
rect -3042 -29689 -2786 -29433
rect -2518 -29689 -2262 -29433
rect -7444 -30183 -7188 -29927
rect -6920 -30183 -6664 -29927
rect -6366 -30183 -6110 -29927
rect -5812 -30183 -5556 -29927
rect -5288 -30183 -5032 -29927
rect -4674 -30183 -4418 -29927
rect -4150 -30183 -3894 -29927
rect -3596 -30183 -3340 -29927
rect -3042 -30183 -2786 -29927
rect -2518 -30183 -2262 -29927
rect 2393 -31582 2649 -31326
rect 2917 -31582 3173 -31326
rect 3471 -31582 3727 -31326
rect 4025 -31582 4281 -31326
rect 4549 -31582 4805 -31326
rect 5163 -31582 5419 -31326
rect 5687 -31582 5943 -31326
rect 6241 -31582 6497 -31326
rect 6795 -31582 7051 -31326
rect 7319 -31582 7575 -31326
rect 2393 -32076 2649 -31820
rect 2917 -32076 3173 -31820
rect 3471 -32076 3727 -31820
rect 4025 -32076 4281 -31820
rect 4549 -32076 4805 -31820
rect 5163 -32076 5419 -31820
rect 5687 -32076 5943 -31820
rect 6241 -32076 6497 -31820
rect 6795 -32076 7051 -31820
rect 7319 -32076 7575 -31820
rect 2393 -32690 2649 -32434
rect 2917 -32690 3173 -32434
rect 3471 -32690 3727 -32434
rect 4025 -32690 4281 -32434
rect 4549 -32690 4805 -32434
rect 5163 -32690 5419 -32434
rect 5687 -32690 5943 -32434
rect 6241 -32690 6497 -32434
rect 6795 -32690 7051 -32434
rect 7319 -32690 7575 -32434
rect 2393 -33184 2649 -32928
rect 2917 -33184 3173 -32928
rect 3471 -33184 3727 -32928
rect 4025 -33184 4281 -32928
rect 4549 -33184 4805 -32928
rect 5163 -33184 5419 -32928
rect 5687 -33184 5943 -32928
rect 6241 -33184 6497 -32928
rect 6795 -33184 7051 -32928
rect 7319 -33184 7575 -32928
rect -7444 -34585 -7188 -34329
rect -6920 -34585 -6664 -34329
rect -6366 -34585 -6110 -34329
rect -5812 -34585 -5556 -34329
rect -5288 -34585 -5032 -34329
rect -4674 -34585 -4418 -34329
rect -4150 -34585 -3894 -34329
rect -3596 -34585 -3340 -34329
rect -3042 -34585 -2786 -34329
rect -2518 -34585 -2262 -34329
rect -7444 -35079 -7188 -34823
rect -6920 -35079 -6664 -34823
rect -6366 -35079 -6110 -34823
rect -5812 -35079 -5556 -34823
rect -5288 -35079 -5032 -34823
rect -4674 -35079 -4418 -34823
rect -4150 -35079 -3894 -34823
rect -3596 -35079 -3340 -34823
rect -3042 -35079 -2786 -34823
rect -2518 -35079 -2262 -34823
rect -7444 -35693 -7188 -35437
rect -6920 -35693 -6664 -35437
rect -6366 -35693 -6110 -35437
rect -5812 -35693 -5556 -35437
rect -5288 -35693 -5032 -35437
rect -4674 -35693 -4418 -35437
rect -4150 -35693 -3894 -35437
rect -3596 -35693 -3340 -35437
rect -3042 -35693 -2786 -35437
rect -2518 -35693 -2262 -35437
rect -7444 -36187 -7188 -35931
rect -6920 -36187 -6664 -35931
rect -6366 -36187 -6110 -35931
rect -5812 -36187 -5556 -35931
rect -5288 -36187 -5032 -35931
rect -4674 -36187 -4418 -35931
rect -4150 -36187 -3894 -35931
rect -3596 -36187 -3340 -35931
rect -3042 -36187 -2786 -35931
rect -2518 -36187 -2262 -35931
<< metal3 >>
tri -17624 34008 -15124 36508 se
rect -15124 36340 15124 36508
tri 15124 36340 15292 36508 sw
rect -15124 34008 15292 36340
tri 15292 34008 17624 36340 sw
tri -18447 33185 -17624 34008 se
rect -17624 33506 -14590 34008
tri -14590 33506 -14088 34008 nw
tri 14088 33506 14590 34008 ne
rect 14590 33506 17624 34008
rect -17624 33185 -14911 33506
tri -14911 33185 -14590 33506 nw
tri -14202 33185 -13881 33506 se
rect -13881 33286 -2268 33506
tri -2268 33286 -2048 33506 sw
rect -13881 33185 -2048 33286
tri -18660 32972 -18447 33185 se
rect -18447 32972 -15124 33185
tri -15124 32972 -14911 33185 nw
tri -14415 32972 -14202 33185 se
rect -14202 32972 -7331 33185
tri -18703 32929 -18660 32972 se
rect -18660 32929 -15167 32972
tri -15167 32929 -15124 32972 nw
tri -14458 32929 -14415 32972 se
rect -14415 32929 -7331 32972
rect -7075 32929 -6807 33185
rect -6551 32929 -6253 33185
rect -5997 32929 -5699 33185
rect -5443 32929 -5175 33185
rect -4919 32929 -4561 33185
rect -4305 32929 -4037 33185
rect -3781 32929 -3483 33185
rect -3227 32929 -2929 33185
rect -2673 32929 -2405 33185
rect -2149 32929 -2048 33185
tri 453 32972 987 33506 se
rect 987 32972 13881 33506
tri 13881 32972 14415 33506 sw
tri 14590 32972 15124 33506 ne
rect 15124 32972 17624 33506
tri -18828 32804 -18703 32929 se
rect -18703 32804 -15292 32929
tri -15292 32804 -15167 32929 nw
tri -14583 32804 -14458 32929 se
rect -14458 32804 -2048 32929
tri 285 32804 453 32972 se
rect 453 32804 14415 32972
tri 14415 32804 14583 32972 sw
tri 15124 32804 15292 32972 ne
rect 15292 32804 17624 32972
tri 17624 32804 18828 34008 sw
tri -18941 32691 -18828 32804 se
rect -18828 32691 -15405 32804
tri -15405 32691 -15292 32804 nw
tri -14696 32691 -14583 32804 se
rect -14583 32691 -2048 32804
tri -19197 32435 -18941 32691 se
rect -18941 32435 -15661 32691
tri -15661 32435 -15405 32691 nw
tri -14952 32435 -14696 32691 se
rect -14696 32435 -7331 32691
rect -7075 32435 -6807 32691
rect -6551 32435 -6253 32691
rect -5997 32435 -5699 32691
rect -5443 32435 -5175 32691
rect -4919 32435 -4561 32691
rect -4305 32435 -4037 32691
rect -3781 32435 -3483 32691
rect -3227 32435 -2929 32691
rect -2673 32435 -2405 32691
rect -2149 32435 -2048 32691
tri -19555 32077 -19197 32435 se
rect -19197 32095 -16001 32435
tri -16001 32095 -15661 32435 nw
tri -15292 32095 -14952 32435 se
rect -14952 32095 -2048 32435
rect -19197 32077 -16019 32095
tri -16019 32077 -16001 32095 nw
tri -15310 32077 -15292 32095 se
rect -15292 32077 -2048 32095
tri -19811 31821 -19555 32077 se
rect -19555 31821 -16275 32077
tri -16275 31821 -16019 32077 nw
tri -15566 31821 -15310 32077 se
rect -15310 31821 -7331 32077
rect -7075 31821 -6807 32077
rect -6551 31821 -6253 32077
rect -5997 31821 -5699 32077
rect -5443 31821 -5175 32077
rect -4919 31821 -4561 32077
rect -4305 31821 -4037 32077
rect -3781 31821 -3483 32077
rect -3227 31821 -2929 32077
rect -2673 31821 -2405 32077
rect -2149 31821 -2048 32077
tri -20049 31583 -19811 31821 se
rect -19811 31583 -16513 31821
tri -16513 31583 -16275 31821 nw
tri -15804 31583 -15566 31821 se
rect -15566 31583 -2048 31821
tri -20305 31327 -20049 31583 se
rect -20049 31388 -16708 31583
tri -16708 31388 -16513 31583 nw
tri -15999 31388 -15804 31583 se
rect -15804 31388 -7331 31583
rect -20049 31327 -16769 31388
tri -16769 31327 -16708 31388 nw
tri -16060 31327 -15999 31388 se
rect -15999 31327 -7331 31388
rect -7075 31327 -6807 31583
rect -6551 31327 -6253 31583
rect -5997 31327 -5699 31583
rect -5443 31327 -5175 31583
rect -4919 31327 -4561 31583
rect -4305 31327 -4037 31583
rect -3781 31327 -3483 31583
rect -3227 31327 -2929 31583
rect -2673 31327 -2405 31583
rect -2149 31327 -2048 31583
tri -958 31561 285 32804 se
rect 285 32270 14583 32804
tri 14583 32270 15117 32804 sw
tri 15292 32270 15826 32804 ne
rect 15826 32270 18828 32804
rect 285 31561 15117 32270
tri 15117 31561 15826 32270 sw
tri 15826 31561 16535 32270 ne
rect 16535 31561 18828 32270
tri 18828 31561 20071 32804 sw
tri -21449 30183 -20305 31327 se
rect -20305 30679 -17417 31327
tri -17417 30679 -16769 31327 nw
tri -16708 30679 -16060 31327 se
rect -16060 31226 -2048 31327
rect -16060 31006 -2268 31226
tri -2268 31006 -2048 31226 nw
tri -1513 31006 -958 31561 se
rect -958 31006 15826 31561
rect -16060 30679 -13347 31006
rect -20305 30183 -17913 30679
tri -17913 30183 -17417 30679 nw
tri -17204 30183 -16708 30679 se
rect -16708 30504 -13347 30679
tri -13347 30504 -12845 31006 nw
tri -2015 30504 -1513 31006 se
rect -1513 30504 1521 31006
tri 1521 30504 2023 31006 nw
tri 12845 30504 13347 31006 ne
rect 13347 30852 15826 31006
tri 15826 30852 16535 31561 sw
tri 16535 30852 17244 31561 ne
rect 17244 30852 20071 31561
rect 13347 30504 16535 30852
rect -16708 30183 -13668 30504
tri -13668 30183 -13347 30504 nw
tri -12824 30317 -12637 30504 se
rect -12637 30317 1334 30504
tri 1334 30317 1521 30504 nw
tri 2436 30317 2623 30504 se
rect 2623 30317 12637 30504
tri 12637 30317 12824 30504 sw
tri 13347 30317 13534 30504 ne
rect 13534 30317 16535 30504
tri -12958 30183 -12824 30317 se
rect -12824 30183 1200 30317
tri 1200 30183 1334 30317 nw
tri 2403 30284 2436 30317 se
rect 2436 30284 12824 30317
rect 2403 30183 12824 30284
tri -21662 29970 -21449 30183 se
rect -21449 29970 -18126 30183
tri -18126 29970 -17913 30183 nw
tri -17417 29970 -17204 30183 se
rect -17204 29970 -13881 30183
tri -13881 29970 -13668 30183 nw
tri -13171 29970 -12958 30183 se
rect -12958 29970 987 30183
tri 987 29970 1200 30183 nw
tri -21705 29927 -21662 29970 se
rect -21662 29927 -18169 29970
tri -18169 29927 -18126 29970 nw
tri -17460 29927 -17417 29970 se
rect -17417 29927 -13924 29970
tri -13924 29927 -13881 29970 nw
tri -13214 29927 -13171 29970 se
rect -13171 29927 944 29970
tri 944 29927 987 29970 nw
rect 2403 29927 2504 30183
rect 2760 29927 3028 30183
rect 3284 29927 3582 30183
rect 3838 29927 4136 30183
rect 4392 29927 4660 30183
rect 4916 29927 5274 30183
rect 5530 29927 5798 30183
rect 6054 29927 6352 30183
rect 6608 29927 6906 30183
rect 7162 29927 7430 30183
rect 7686 29970 12824 30183
tri 12824 29970 13171 30317 sw
tri 13534 29970 13881 30317 ne
rect 13881 30143 16535 30317
tri 16535 30143 17244 30852 sw
tri 17244 30143 17953 30852 ne
rect 17953 30143 20071 30852
rect 13881 29977 17244 30143
tri 17244 29977 17410 30143 sw
tri 17953 29977 18119 30143 ne
rect 18119 29977 20071 30143
rect 13881 29970 17410 29977
rect 7686 29927 13171 29970
tri -21943 29689 -21705 29927 se
rect -21705 29689 -18407 29927
tri -18407 29689 -18169 29927 nw
tri -17698 29689 -17460 29927 se
rect -17460 29689 -14162 29927
tri -14162 29689 -13924 29927 nw
tri -13452 29689 -13214 29927 se
rect -13214 29689 706 29927
tri 706 29689 944 29927 nw
rect 2403 29689 13171 29927
tri -22196 29436 -21943 29689 se
rect -21943 29436 -18660 29689
tri -18660 29436 -18407 29689 nw
tri -17951 29436 -17698 29689 se
rect -17698 29436 -14415 29689
tri -14415 29436 -14162 29689 nw
tri -13705 29436 -13452 29689 se
rect -13452 29436 453 29689
tri 453 29436 706 29689 nw
tri -22199 29433 -22196 29436 se
rect -22196 29433 -18663 29436
tri -18663 29433 -18660 29436 nw
tri -17954 29433 -17951 29436 se
rect -17951 29433 -14418 29436
tri -14418 29433 -14415 29436 nw
tri -13708 29433 -13705 29436 se
rect -13705 29433 450 29436
tri 450 29433 453 29436 nw
rect 2403 29433 2504 29689
rect 2760 29433 3028 29689
rect 3284 29433 3582 29689
rect 3838 29433 4136 29689
rect 4392 29433 4660 29689
rect 4916 29433 5274 29689
rect 5530 29433 5798 29689
rect 6054 29433 6352 29689
rect 6608 29433 6906 29689
rect 7162 29433 7430 29689
rect 7686 29436 13171 29689
tri 13171 29436 13705 29970 sw
tri 13881 29436 14415 29970 ne
rect 14415 29436 17410 29970
tri 17410 29436 17951 29977 sw
tri 18119 29436 18660 29977 ne
rect 18660 29436 20071 29977
rect 7686 29433 13705 29436
tri -22364 29268 -22199 29433 se
rect -22199 29268 -18828 29433
tri -18828 29268 -18663 29433 nw
tri -18119 29268 -17954 29433 se
rect -17954 29268 -14583 29433
tri -14583 29268 -14418 29433 nw
tri -13873 29268 -13708 29433 se
rect -13708 29268 285 29433
tri 285 29268 450 29433 nw
rect 2403 29268 13705 29433
tri 13705 29268 13873 29436 sw
tri 14415 29268 14583 29436 ne
rect 14583 29268 17951 29436
tri 17951 29268 18119 29436 sw
tri 18660 29268 18828 29436 ne
rect 18828 29268 20071 29436
tri 20071 29268 22364 31561 sw
tri -22557 29075 -22364 29268 se
rect -22364 29075 -19021 29268
tri -19021 29075 -18828 29268 nw
tri -18312 29075 -18119 29268 se
rect -18119 29075 -14776 29268
tri -14776 29075 -14583 29268 nw
tri -14066 29075 -13873 29268 se
rect -13873 29075 92 29268
tri 92 29075 285 29268 nw
rect 2403 29075 13873 29268
tri -22813 28819 -22557 29075 se
rect -22557 28819 -19277 29075
tri -19277 28819 -19021 29075 nw
tri -18568 28819 -18312 29075 se
rect -18312 28819 -15032 29075
tri -15032 28819 -14776 29075 nw
tri -14322 28819 -14066 29075 se
rect -14066 28819 -164 29075
tri -164 28819 92 29075 nw
rect 2403 28819 2504 29075
rect 2760 28819 3028 29075
rect 3284 28819 3582 29075
rect 3838 28819 4136 29075
rect 4392 28819 4660 29075
rect 4916 28819 5274 29075
rect 5530 28819 5798 29075
rect 6054 28819 6352 29075
rect 6608 28819 6906 29075
rect 7162 28819 7430 29075
rect 7686 28819 13873 29075
tri -23051 28581 -22813 28819 se
rect -22813 28581 -19515 28819
tri -19515 28581 -19277 28819 nw
tri -18806 28581 -18568 28819 se
rect -18568 28581 -15270 28819
tri -15270 28581 -15032 28819 nw
tri -14560 28581 -14322 28819 se
rect -14322 28581 -402 28819
tri -402 28581 -164 28819 nw
rect 2403 28581 13873 28819
tri -23307 28325 -23051 28581 se
rect -23051 28559 -19537 28581
tri -19537 28559 -19515 28581 nw
tri -18828 28559 -18806 28581 se
rect -18806 28559 -15293 28581
rect -23051 28325 -19771 28559
tri -19771 28325 -19537 28559 nw
tri -19062 28325 -18828 28559 se
rect -18828 28558 -15293 28559
tri -15293 28558 -15270 28581 nw
tri -14583 28558 -14560 28581 se
rect -14560 28558 -658 28581
rect -18828 28325 -15526 28558
tri -15526 28325 -15293 28558 nw
tri -14816 28325 -14583 28558 se
rect -14583 28325 -658 28558
tri -658 28325 -402 28581 nw
rect 2403 28325 2504 28581
rect 2760 28325 3028 28581
rect 3284 28325 3582 28581
rect 3838 28325 4136 28581
rect 4392 28325 4660 28581
rect 4916 28325 5274 28581
rect 5530 28325 5798 28581
rect 6054 28325 6352 28581
rect 6608 28325 6906 28581
rect 7162 28325 7430 28581
rect 7686 28558 13873 28581
tri 13873 28558 14583 29268 sw
tri 14583 28558 15293 29268 ne
rect 15293 28734 18119 29268
tri 18119 28734 18653 29268 sw
tri 18828 28734 19362 29268 ne
rect 19362 28734 22364 29268
rect 15293 28558 18653 28734
rect 7686 28325 14583 28558
tri -24451 27181 -23307 28325 se
rect -23307 27852 -20244 28325
tri -20244 27852 -19771 28325 nw
tri -19535 27852 -19062 28325 se
rect -19062 28025 -15826 28325
tri -15826 28025 -15526 28325 nw
tri -15116 28025 -14816 28325 se
rect -14816 28025 -958 28325
tri -958 28025 -658 28325 nw
rect 2403 28224 14583 28325
tri 2403 28025 2602 28224 ne
rect 2602 28025 14583 28224
tri 14583 28025 15116 28558 sw
tri 15293 28025 15826 28558 ne
rect 15826 28025 18653 28558
tri 18653 28025 19362 28734 sw
tri 19362 28025 20071 28734 ne
rect 20071 28025 22364 28734
tri 22364 28025 23607 29268 sw
rect -19062 27852 -16173 28025
rect -23307 27181 -20915 27852
tri -20915 27181 -20244 27852 nw
tri -20206 27181 -19535 27852 se
rect -19535 27678 -16173 27852
tri -16173 27678 -15826 28025 nw
tri -15463 27678 -15116 28025 se
rect -15116 28004 -979 28025
tri -979 28004 -958 28025 nw
tri 2602 28004 2623 28025 ne
rect 2623 28004 15116 28025
rect -15116 27678 -12103 28004
rect -19535 27181 -16670 27678
tri -16670 27181 -16173 27678 nw
tri -15960 27181 -15463 27678 se
rect -15463 27502 -12103 27678
tri -12103 27502 -11601 28004 nw
tri 11601 27502 12103 28004 ne
rect 12103 27502 15116 28004
rect -15463 27181 -12424 27502
tri -12424 27181 -12103 27502 nw
tri -11715 27181 -11394 27502 se
rect -11394 27282 -2268 27502
tri -2268 27282 -2048 27502 sw
rect -11394 27181 -2048 27282
tri -24707 26925 -24451 27181 se
rect -24451 27143 -20953 27181
tri -20953 27143 -20915 27181 nw
tri -20244 27143 -20206 27181 se
rect -20206 27143 -16883 27181
rect -24451 26925 -21171 27143
tri -21171 26925 -20953 27143 nw
tri -20462 26925 -20244 27143 se
rect -20244 26968 -16883 27143
tri -16883 26968 -16670 27181 nw
tri -16173 26968 -15960 27181 se
rect -15960 26968 -12637 27181
tri -12637 26968 -12424 27181 nw
tri -11928 26968 -11715 27181 se
rect -11715 26968 -7331 27181
rect -20244 26925 -16926 26968
tri -16926 26925 -16883 26968 nw
tri -16216 26925 -16173 26968 se
rect -16173 26925 -12680 26968
tri -12680 26925 -12637 26968 nw
tri -11971 26925 -11928 26968 se
rect -11928 26925 -7331 26968
rect -7075 26925 -6807 27181
rect -6551 26925 -6253 27181
rect -5997 26925 -5699 27181
rect -5443 26925 -5175 27181
rect -4919 26925 -4561 27181
rect -4305 26925 -4037 27181
rect -3781 26925 -3483 27181
rect -3227 26925 -2929 27181
rect -2673 26925 -2405 27181
rect -2149 26925 -2048 27181
tri 453 26968 987 27502 se
rect 987 26968 11394 27502
tri 11394 26968 11928 27502 sw
tri 12103 26968 12637 27502 ne
rect 12637 27491 15116 27502
tri 15116 27491 15650 28025 sw
tri 15826 27491 16360 28025 ne
rect 16360 27491 19362 28025
rect 12637 26968 15650 27491
tri -24945 26687 -24707 26925 se
rect -24707 26687 -21409 26925
tri -21409 26687 -21171 26925 nw
tri -20700 26687 -20462 26925 se
rect -20462 26687 -17164 26925
tri -17164 26687 -16926 26925 nw
tri -16360 26781 -16216 26925 se
rect -16216 26781 -12824 26925
tri -12824 26781 -12680 26925 nw
tri -12115 26781 -11971 26925 se
rect -11971 26781 -2048 26925
tri 266 26781 453 26968 se
rect 453 26793 11928 26968
tri 11928 26793 12103 26968 sw
tri 12637 26793 12812 26968 ne
rect 12812 26793 15650 26968
rect 453 26781 12103 26793
tri 12103 26781 12115 26793 sw
tri 12812 26781 12824 26793 ne
rect 12824 26781 15650 26793
tri 15650 26781 16360 27491 sw
tri 16360 26781 17070 27491 ne
rect 17070 27316 19362 27491
tri 19362 27316 20071 28025 sw
tri 20071 27316 20780 28025 ne
rect 20780 27316 23607 28025
rect 17070 26781 20071 27316
tri -16454 26687 -16360 26781 se
rect -16360 26687 -12918 26781
tri -12918 26687 -12824 26781 nw
tri -12209 26687 -12115 26781 se
rect -12115 26687 -2048 26781
tri -25198 26434 -24945 26687 se
rect -24945 26434 -21662 26687
tri -21662 26434 -21409 26687 nw
tri -20953 26434 -20700 26687 se
rect -20700 26434 -17417 26687
tri -17417 26434 -17164 26687 nw
tri -16707 26434 -16454 26687 se
rect -16454 26434 -13171 26687
tri -13171 26434 -12918 26687 nw
tri -12462 26434 -12209 26687 se
rect -12209 26434 -7331 26687
tri -25201 26431 -25198 26434 se
rect -25198 26431 -21665 26434
tri -21665 26431 -21662 26434 nw
tri -20956 26431 -20953 26434 se
rect -20953 26431 -17420 26434
tri -17420 26431 -17417 26434 nw
tri -16710 26431 -16707 26434 se
rect -16707 26431 -13174 26434
tri -13174 26431 -13171 26434 nw
tri -12465 26431 -12462 26434 se
rect -12462 26431 -7331 26434
rect -7075 26431 -6807 26687
rect -6551 26431 -6253 26687
rect -5997 26431 -5699 26687
rect -5443 26431 -5175 26687
rect -4919 26431 -4561 26687
rect -4305 26431 -4037 26687
rect -3781 26431 -3483 26687
rect -3227 26431 -2929 26687
rect -2673 26431 -2405 26687
rect -2149 26431 -2048 26687
tri -81 26434 266 26781 se
rect 266 26434 12115 26781
tri 12115 26434 12462 26781 sw
tri 12824 26434 13171 26781 ne
rect 13171 26434 16360 26781
tri 16360 26434 16707 26781 sw
tri 17070 26434 17417 26781 ne
rect 17417 26607 20071 26781
tri 20071 26607 20780 27316 sw
tri 20780 26607 21489 27316 ne
rect 21489 26607 23607 27316
rect 17417 26441 20780 26607
tri 20780 26441 20946 26607 sw
tri 21489 26441 21655 26607 ne
rect 21655 26441 23607 26607
rect 17417 26434 20946 26441
tri -25559 26073 -25201 26431 se
rect -25201 26073 -22023 26431
tri -22023 26073 -21665 26431 nw
tri -21314 26073 -20956 26431 se
rect -20956 26073 -17778 26431
tri -17778 26073 -17420 26431 nw
tri -17068 26073 -16710 26431 se
rect -16710 26073 -13532 26431
tri -13532 26073 -13174 26431 nw
tri -12823 26073 -12465 26431 se
rect -12465 26073 -2048 26431
tri -25732 25900 -25559 26073 se
rect -25559 25900 -22196 26073
tri -22196 25900 -22023 26073 nw
tri -21487 25900 -21314 26073 se
rect -21314 25900 -17951 26073
tri -17951 25900 -17778 26073 nw
tri -17241 25900 -17068 26073 se
rect -17068 25900 -13705 26073
tri -13705 25900 -13532 26073 nw
tri -12996 25900 -12823 26073 se
rect -12823 25900 -7331 26073
tri -25815 25817 -25732 25900 se
rect -25732 25817 -22279 25900
tri -22279 25817 -22196 25900 nw
tri -21570 25817 -21487 25900 se
rect -21487 25817 -18034 25900
tri -18034 25817 -17951 25900 nw
tri -17324 25817 -17241 25900 se
rect -17241 25817 -13788 25900
tri -13788 25817 -13705 25900 nw
tri -13079 25817 -12996 25900 se
rect -12996 25817 -7331 25900
rect -7075 25817 -6807 26073
rect -6551 25817 -6253 26073
rect -5997 25817 -5699 26073
rect -5443 25817 -5175 26073
rect -4919 25817 -4561 26073
rect -4305 25817 -4037 26073
rect -3781 25817 -3483 26073
rect -3227 25817 -2929 26073
rect -2673 25817 -2405 26073
rect -2149 25817 -2048 26073
tri -615 25900 -81 26434 se
rect -81 26247 12462 26434
tri 12462 26247 12649 26434 sw
tri 13171 26247 13358 26434 ne
rect 13358 26247 16707 26434
rect -81 25900 12649 26247
tri 12649 25900 12996 26247 sw
tri 13358 25900 13705 26247 ne
rect 13705 26071 16707 26247
tri 16707 26071 17070 26434 sw
tri 17417 26071 17780 26434 ne
rect 17780 26071 20946 26434
rect 13705 25900 17070 26071
tri 17070 25900 17241 26071 sw
tri 17780 25900 17951 26071 ne
rect 17951 25900 20946 26071
tri 20946 25900 21487 26441 sw
tri 21655 25900 22196 26441 ne
rect 22196 25900 23607 26441
tri -25900 25732 -25815 25817 se
rect -25815 25732 -22364 25817
tri -22364 25732 -22279 25817 nw
tri -21655 25732 -21570 25817 se
rect -21570 25732 -18119 25817
tri -18119 25732 -18034 25817 nw
tri -17409 25732 -17324 25817 se
rect -17324 25732 -13873 25817
tri -13873 25732 -13788 25817 nw
tri -13164 25732 -13079 25817 se
rect -13079 25732 -2048 25817
tri -783 25732 -615 25900 se
rect -615 25732 12996 25900
tri 12996 25732 13164 25900 sw
tri 13705 25732 13873 25900 ne
rect 13873 25732 17241 25900
tri 17241 25732 17409 25900 sw
tri 17951 25732 18119 25900 ne
rect 18119 25732 21487 25900
tri 21487 25732 21655 25900 sw
tri 22196 25732 22364 25900 ne
rect 22364 25732 23607 25900
tri 23607 25732 25900 28025 sw
tri -26053 25579 -25900 25732 se
rect -25900 25579 -22517 25732
tri -22517 25579 -22364 25732 nw
tri -21808 25579 -21655 25732 se
rect -21655 25579 -18272 25732
tri -18272 25579 -18119 25732 nw
tri -17562 25579 -17409 25732 se
rect -17409 25579 -14026 25732
tri -14026 25579 -13873 25732 nw
tri -13317 25579 -13164 25732 se
rect -13164 25579 -2048 25732
tri -26309 25323 -26053 25579 se
rect -26053 25323 -22773 25579
tri -22773 25323 -22517 25579 nw
tri -22064 25323 -21808 25579 se
rect -21808 25323 -18528 25579
tri -18528 25323 -18272 25579 nw
tri -17818 25323 -17562 25579 se
rect -17562 25323 -14282 25579
tri -14282 25323 -14026 25579 nw
tri -13358 25538 -13317 25579 se
rect -13317 25538 -7331 25579
tri -13573 25323 -13358 25538 se
rect -13358 25323 -7331 25538
rect -7075 25323 -6807 25579
rect -6551 25323 -6253 25579
rect -5997 25323 -5699 25579
rect -5443 25323 -5175 25579
rect -4919 25323 -4561 25579
rect -4305 25323 -4037 25579
rect -3781 25323 -3483 25579
rect -3227 25323 -2929 25579
rect -2673 25323 -2405 25579
rect -2149 25323 -2048 25579
tri -977 25538 -783 25732 se
rect -783 25538 13164 25732
tri 13164 25538 13358 25732 sw
tri 13873 25538 14067 25732 ne
rect 14067 25538 17409 25732
tri -27453 24179 -26309 25323 se
rect -26309 25023 -23073 25323
tri -23073 25023 -22773 25323 nw
tri -22364 25023 -22064 25323 se
rect -22064 25023 -18829 25323
rect -26309 24316 -23780 25023
tri -23780 24316 -23073 25023 nw
tri -23071 24316 -22364 25023 se
rect -22364 25022 -18829 25023
tri -18829 25022 -18528 25323 nw
tri -18119 25022 -17818 25323 se
rect -17818 25023 -14582 25323
tri -14582 25023 -14282 25323 nw
tri -13873 25023 -13573 25323 se
rect -13573 25222 -2048 25323
rect -13573 25023 -2268 25222
rect -17818 25022 -14930 25023
rect -22364 24489 -19362 25022
tri -19362 24489 -18829 25022 nw
tri -18652 24489 -18119 25022 se
rect -18119 24675 -14930 25022
tri -14930 24675 -14582 25023 nw
tri -14221 24675 -13873 25023 se
rect -13873 25002 -2268 25023
tri -2268 25002 -2048 25222 nw
tri -1513 25002 -977 25538 se
rect -977 25002 13358 25538
rect -13873 24675 -10860 25002
rect -18119 24489 -15116 24675
tri -15116 24489 -14930 24675 nw
tri -14407 24489 -14221 24675 se
rect -14221 24500 -10860 24675
tri -10860 24500 -10358 25002 nw
tri -2015 24500 -1513 25002 se
rect -1513 24500 1521 25002
tri 1521 24500 2023 25002 nw
tri 10358 24500 10860 25002 ne
rect 10860 24829 13358 25002
tri 13358 24829 14067 25538 sw
tri 14067 24829 14776 25538 ne
rect 14776 25022 17409 25538
tri 17409 25022 18119 25732 sw
tri 18119 25022 18829 25732 ne
rect 18829 25198 21655 25732
tri 21655 25198 22189 25732 sw
tri 22364 25198 22898 25732 ne
rect 22898 25198 25900 25732
rect 18829 25022 22189 25198
rect 14776 24829 18119 25022
rect 10860 24500 14067 24829
rect -14221 24489 -10871 24500
tri -10871 24489 -10860 24500 nw
tri -10161 24489 -10150 24500 se
rect -10150 24489 1510 24500
tri 1510 24489 1521 24500 nw
tri 2612 24489 2623 24500 se
rect 2623 24489 10150 24500
tri 10150 24489 10161 24500 sw
tri 10860 24489 10871 24500 ne
rect 10871 24489 14067 24500
tri 14067 24489 14407 24829 sw
tri 14776 24489 15116 24829 ne
rect 15116 24489 18119 24829
tri 18119 24489 18652 25022 sw
tri 18829 24489 19362 25022 ne
rect 19362 24489 22189 25022
tri 22189 24489 22898 25198 sw
tri 22898 24489 23607 25198 ne
rect 23607 24489 25900 25198
tri 25900 24489 27143 25732 sw
rect -22364 24316 -19672 24489
rect -26309 24179 -23917 24316
tri -23917 24179 -23780 24316 nw
tri -23208 24179 -23071 24316 se
rect -23071 24179 -19672 24316
tri -19672 24179 -19362 24489 nw
tri -18962 24179 -18652 24489 se
rect -18652 24179 -15426 24489
tri -15426 24179 -15116 24489 nw
tri -14717 24179 -14407 24489 se
rect -14407 24179 -11181 24489
tri -11181 24179 -10871 24489 nw
tri -10356 24294 -10161 24489 se
rect -10161 24294 1315 24489
tri 1315 24294 1510 24489 nw
tri 2417 24294 2612 24489 se
rect 2612 24294 10161 24489
tri 10161 24294 10356 24489 sw
tri 10871 24294 11066 24489 ne
rect 11066 24294 14407 24489
tri -10471 24179 -10356 24294 se
rect -10356 24179 1200 24294
tri 1200 24179 1315 24294 nw
tri 2403 24280 2417 24294 se
rect 2417 24280 10356 24294
rect 2403 24179 10356 24280
tri -27709 23923 -27453 24179 se
rect -27453 23923 -24173 24179
tri -24173 23923 -23917 24179 nw
tri -23464 23923 -23208 24179 se
rect -23208 24142 -19709 24179
tri -19709 24142 -19672 24179 nw
tri -18999 24142 -18962 24179 se
rect -18962 24142 -15639 24179
rect -23208 23923 -19928 24142
tri -19928 23923 -19709 24142 nw
tri -19218 23923 -18999 24142 se
rect -18999 23966 -15639 24142
tri -15639 23966 -15426 24179 nw
tri -14930 23966 -14717 24179 se
rect -14717 23966 -11394 24179
tri -11394 23966 -11181 24179 nw
tri -10684 23966 -10471 24179 se
rect -10471 23966 987 24179
tri 987 23966 1200 24179 nw
rect -18999 23923 -15682 23966
tri -15682 23923 -15639 23966 nw
tri -14973 23923 -14930 23966 se
rect -14930 23923 -11437 23966
tri -11437 23923 -11394 23966 nw
tri -10727 23923 -10684 23966 se
rect -10684 23923 944 23966
tri 944 23923 987 23966 nw
rect 2403 23923 2504 24179
rect 2760 23923 3028 24179
rect 3284 23923 3582 24179
rect 3838 23923 4136 24179
rect 4392 23923 4660 24179
rect 4916 23923 5274 24179
rect 5530 23923 5798 24179
rect 6054 23923 6352 24179
rect 6608 23923 6906 24179
rect 7162 23923 7430 24179
rect 7686 23966 10356 24179
tri 10356 23966 10684 24294 sw
tri 11066 23966 11394 24294 ne
rect 11394 23966 14407 24294
rect 7686 23923 10684 23966
tri -27947 23685 -27709 23923 se
rect -27709 23685 -24411 23923
tri -24411 23685 -24173 23923 nw
tri -23702 23685 -23464 23923 se
rect -23464 23685 -20166 23923
tri -20166 23685 -19928 23923 nw
tri -19456 23685 -19218 23923 se
rect -19218 23685 -15920 23923
tri -15920 23685 -15682 23923 nw
tri -15211 23685 -14973 23923 se
rect -14973 23685 -11675 23923
tri -11675 23685 -11437 23923 nw
tri -10965 23685 -10727 23923 se
rect -10727 23685 706 23923
tri 706 23685 944 23923 nw
rect 2403 23685 10684 23923
tri -28203 23429 -27947 23685 se
rect -27947 23607 -24489 23685
tri -24489 23607 -24411 23685 nw
tri -23780 23607 -23702 23685 se
rect -23702 23607 -20419 23685
rect -27947 23429 -24667 23607
tri -24667 23429 -24489 23607 nw
tri -23958 23429 -23780 23607 se
rect -23780 23432 -20419 23607
tri -20419 23432 -20166 23685 nw
tri -19709 23432 -19456 23685 se
rect -19456 23432 -16173 23685
tri -16173 23432 -15920 23685 nw
tri -15464 23432 -15211 23685 se
rect -15211 23432 -11928 23685
tri -11928 23432 -11675 23685 nw
tri -11218 23432 -10965 23685 se
rect -10965 23432 453 23685
tri 453 23432 706 23685 nw
rect -23780 23429 -20422 23432
tri -20422 23429 -20419 23432 nw
tri -19712 23429 -19709 23432 se
rect -19709 23429 -16176 23432
tri -16176 23429 -16173 23432 nw
tri -15467 23429 -15464 23432 se
rect -15464 23429 -11931 23432
tri -11931 23429 -11928 23432 nw
tri -11221 23429 -11218 23432 se
rect -11218 23429 450 23432
tri 450 23429 453 23432 nw
rect 2403 23429 2504 23685
rect 2760 23429 3028 23685
rect 3284 23429 3582 23685
rect 3838 23429 4136 23685
rect 4392 23429 4660 23685
rect 4916 23429 5274 23685
rect 5530 23429 5798 23685
rect 6054 23429 6352 23685
rect 6608 23429 6906 23685
rect 7162 23429 7430 23685
rect 7686 23432 10684 23685
tri 10684 23432 11218 23966 sw
tri 11394 23432 11928 23966 ne
rect 11928 23780 14407 23966
tri 14407 23780 15116 24489 sw
tri 15116 23780 15825 24489 ne
rect 15825 23955 18652 24489
tri 18652 23955 19186 24489 sw
tri 19362 23955 19896 24489 ne
rect 19896 23955 22898 24489
rect 15825 23780 19186 23955
rect 11928 23432 15116 23780
tri 15116 23432 15464 23780 sw
tri 15825 23432 16173 23780 ne
rect 16173 23432 19186 23780
rect 7686 23429 11218 23432
tri -28561 23071 -28203 23429 se
rect -28203 23071 -25025 23429
tri -25025 23071 -24667 23429 nw
tri -24316 23071 -23958 23429 se
rect -23958 23071 -20780 23429
tri -20780 23071 -20422 23429 nw
tri -19896 23245 -19712 23429 se
rect -19712 23245 -16360 23429
tri -16360 23245 -16176 23429 nw
tri -15651 23245 -15467 23429 se
rect -15467 23245 -12115 23429
tri -12115 23245 -11931 23429 nw
tri -11405 23245 -11221 23429 se
rect -11221 23245 266 23429
tri 266 23245 450 23429 nw
rect 2403 23245 11218 23429
tri 11218 23245 11405 23432 sw
tri 11928 23245 12115 23432 ne
rect 12115 23245 15464 23432
tri 15464 23245 15651 23432 sw
tri 16173 23245 16360 23432 ne
rect 16360 23245 19186 23432
tri 19186 23245 19896 23955 sw
tri 19896 23245 20606 23955 ne
rect 20606 23780 22898 23955
tri 22898 23780 23607 24489 sw
tri 23607 23780 24316 24489 ne
rect 24316 23780 27143 24489
rect 20606 23245 23607 23780
tri -20070 23071 -19896 23245 se
rect -19896 23071 -16534 23245
tri -16534 23071 -16360 23245 nw
tri -15825 23071 -15651 23245 se
rect -15651 23071 -12289 23245
tri -12289 23071 -12115 23245 nw
tri -11579 23071 -11405 23245 se
rect -11405 23071 92 23245
tri 92 23071 266 23245 nw
rect 2403 23071 11405 23245
tri -28734 22898 -28561 23071 se
rect -28561 22898 -25198 23071
tri -25198 22898 -25025 23071 nw
tri -24489 22898 -24316 23071 se
rect -24316 22898 -20953 23071
tri -20953 22898 -20780 23071 nw
tri -20243 22898 -20070 23071 se
rect -20070 22898 -16707 23071
tri -16707 22898 -16534 23071 nw
tri -15998 22898 -15825 23071 se
rect -15825 22898 -12462 23071
tri -12462 22898 -12289 23071 nw
tri -11752 22898 -11579 23071 se
rect -11579 22898 -81 23071
tri -81 22898 92 23071 nw
tri -28817 22815 -28734 22898 se
rect -28734 22815 -25281 22898
tri -25281 22815 -25198 22898 nw
tri -24572 22815 -24489 22898 se
rect -24489 22815 -21036 22898
tri -21036 22815 -20953 22898 nw
tri -20326 22815 -20243 22898 se
rect -20243 22815 -16790 22898
tri -16790 22815 -16707 22898 nw
tri -16081 22815 -15998 22898 se
rect -15998 22815 -12545 22898
tri -12545 22815 -12462 22898 nw
tri -11835 22815 -11752 22898 se
rect -11752 22815 -164 22898
tri -164 22815 -81 22898 nw
rect 2403 22815 2504 23071
rect 2760 22815 3028 23071
rect 3284 22815 3582 23071
rect 3838 22815 4136 23071
rect 4392 22815 4660 23071
rect 4916 22815 5274 23071
rect 5530 22815 5798 23071
rect 6054 22815 6352 23071
rect 6608 22815 6906 23071
rect 7162 22815 7430 23071
rect 7686 22898 11405 23071
tri 11405 22898 11752 23245 sw
tri 12115 22898 12462 23245 ne
rect 12462 22898 15651 23245
tri 15651 22898 15998 23245 sw
tri 16360 22898 16707 23245 ne
rect 16707 22898 19896 23245
tri 19896 22898 20243 23245 sw
tri 20606 22898 20953 23245 ne
rect 20953 23071 23607 23245
tri 23607 23071 24316 23780 sw
tri 24316 23071 25025 23780 ne
rect 25025 23071 27143 23780
rect 20953 22905 24316 23071
tri 24316 22905 24482 23071 sw
tri 25025 22905 25191 23071 ne
rect 25191 22905 27143 23071
rect 20953 22898 24482 22905
rect 7686 22815 11752 22898
tri -29055 22577 -28817 22815 se
rect -28817 22577 -25519 22815
tri -25519 22577 -25281 22815 nw
tri -24810 22577 -24572 22815 se
rect -24572 22577 -21274 22815
tri -21274 22577 -21036 22815 nw
tri -20564 22577 -20326 22815 se
rect -20326 22577 -17028 22815
tri -17028 22577 -16790 22815 nw
tri -16319 22577 -16081 22815 se
rect -16081 22577 -12783 22815
tri -12783 22577 -12545 22815 nw
tri -12073 22577 -11835 22815 se
rect -11835 22577 -402 22815
tri -402 22577 -164 22815 nw
rect 2403 22577 11752 22815
tri -29268 22364 -29055 22577 se
rect -29055 22364 -25732 22577
tri -25732 22364 -25519 22577 nw
tri -25023 22364 -24810 22577 se
rect -24810 22364 -21487 22577
tri -21487 22364 -21274 22577 nw
tri -20777 22364 -20564 22577 se
rect -20564 22364 -17241 22577
tri -17241 22364 -17028 22577 nw
tri -16532 22364 -16319 22577 se
rect -16319 22364 -12996 22577
tri -12996 22364 -12783 22577 nw
tri -12286 22364 -12073 22577 se
rect -12073 22364 -615 22577
tri -615 22364 -402 22577 nw
tri -29311 22321 -29268 22364 se
rect -29268 22321 -25775 22364
tri -25775 22321 -25732 22364 nw
tri -25066 22321 -25023 22364 se
rect -25023 22321 -21530 22364
tri -21530 22321 -21487 22364 nw
tri -20820 22321 -20777 22364 se
rect -20777 22321 -17284 22364
tri -17284 22321 -17241 22364 nw
tri -16575 22321 -16532 22364 se
rect -16532 22321 -13039 22364
tri -13039 22321 -12996 22364 nw
tri -12329 22321 -12286 22364 se
rect -12286 22321 -658 22364
tri -658 22321 -615 22364 nw
rect 2403 22321 2504 22577
rect 2760 22321 3028 22577
rect 3284 22321 3582 22577
rect 3838 22321 4136 22577
rect 4392 22321 4660 22577
rect 4916 22321 5274 22577
rect 5530 22321 5798 22577
rect 6054 22321 6352 22577
rect 6608 22321 6906 22577
rect 7162 22321 7430 22577
rect 7686 22364 11752 22577
tri 11752 22364 12286 22898 sw
tri 12462 22364 12996 22898 ne
rect 12996 22711 15998 22898
tri 15998 22711 16185 22898 sw
tri 16707 22711 16894 22898 ne
rect 16894 22711 20243 22898
rect 12996 22364 16185 22711
tri 16185 22364 16532 22711 sw
tri 16894 22364 17241 22711 ne
rect 17241 22535 20243 22711
tri 20243 22535 20606 22898 sw
tri 20953 22535 21316 22898 ne
rect 21316 22535 24482 22898
rect 17241 22364 20606 22535
tri 20606 22364 20777 22535 sw
tri 21316 22364 21487 22535 ne
rect 21487 22364 24482 22535
tri 24482 22364 25023 22905 sw
tri 25191 22364 25732 22905 ne
rect 25732 22364 27143 22905
rect 7686 22321 12286 22364
tri -29436 22196 -29311 22321 se
rect -29311 22196 -25900 22321
tri -25900 22196 -25775 22321 nw
tri -25191 22196 -25066 22321 se
rect -25066 22196 -21655 22321
tri -21655 22196 -21530 22321 nw
tri -20945 22196 -20820 22321 se
rect -20820 22196 -17409 22321
tri -17409 22196 -17284 22321 nw
tri -16700 22196 -16575 22321 se
rect -16575 22196 -13164 22321
tri -13164 22196 -13039 22321 nw
tri -12454 22196 -12329 22321 se
rect -12329 22196 -783 22321
tri -783 22196 -658 22321 nw
rect 2403 22220 12286 22321
tri 2403 22196 2427 22220 ne
rect 2427 22196 12286 22220
tri 12286 22196 12454 22364 sw
tri 12996 22196 13164 22364 ne
rect 13164 22196 16532 22364
tri 16532 22196 16700 22364 sw
tri 17241 22196 17409 22364 ne
rect 17409 22196 20777 22364
tri 20777 22196 20945 22364 sw
tri 21487 22196 21655 22364 ne
rect 21655 22196 25023 22364
tri 25023 22196 25191 22364 sw
tri 25732 22196 25900 22364 ne
rect 25900 22196 27143 22364
tri 27143 22196 29436 24489 sw
tri -32270 19362 -29436 22196 se
rect -29436 21487 -26609 22196
tri -26609 21487 -25900 22196 nw
tri -25900 21487 -25191 22196 se
rect -25191 21487 -22365 22196
rect -29436 20780 -27316 21487
tri -27316 20780 -26609 21487 nw
tri -26607 20780 -25900 21487 se
rect -25900 21486 -22365 21487
tri -22365 21486 -21655 22196 nw
tri -21655 21486 -20945 22196 se
rect -20945 21487 -18118 22196
tri -18118 21487 -17409 22196 nw
tri -16894 22002 -16700 22196 se
rect -16700 22002 -13358 22196
tri -13358 22002 -13164 22196 nw
tri -12648 22002 -12454 22196 se
rect -12454 22002 -977 22196
tri -977 22002 -783 22196 nw
tri 2427 22002 2621 22196 ne
rect 2621 22002 12454 22196
tri 12454 22002 12648 22196 sw
tri 13164 22002 13358 22196 ne
rect 13358 22002 16700 22196
tri 16700 22002 16894 22196 sw
tri 17409 22002 17603 22196 ne
rect 17603 22002 20945 22196
tri -17409 21487 -16894 22002 se
rect -16894 21674 -13686 22002
tri -13686 21674 -13358 22002 nw
tri -12976 21674 -12648 22002 se
rect -12648 22000 -979 22002
tri -979 22000 -977 22002 nw
tri 2621 22000 2623 22002 ne
rect 2623 22000 12648 22002
rect -12648 21674 -10150 22000
rect -16894 21487 -14396 21674
rect -20945 21486 -18466 21487
rect -25900 20953 -22898 21486
tri -22898 20953 -22365 21486 nw
tri -22188 20953 -21655 21486 se
rect -21655 21139 -18466 21486
tri -18466 21139 -18118 21487 nw
tri -17757 21139 -17409 21487 se
rect -17409 21139 -14396 21487
rect -21655 20953 -18652 21139
tri -18652 20953 -18466 21139 nw
tri -17943 20953 -17757 21139 se
rect -17757 20964 -14396 21139
tri -14396 20964 -13686 21674 nw
tri -13686 20964 -12976 21674 se
rect -12976 20964 -10150 21674
tri -10150 20964 -9114 22000 nw
tri 9114 20964 10150 22000 ne
rect 10150 21468 12648 22000
tri 12648 21468 13182 22002 sw
tri 13358 21468 13892 22002 ne
rect 13892 21468 16894 22002
rect 10150 20964 13182 21468
rect -17757 20953 -14407 20964
tri -14407 20953 -14396 20964 nw
tri -13697 20953 -13686 20964 se
rect -13686 20953 -10161 20964
tri -10161 20953 -10150 20964 nw
tri 10150 20953 10161 20964 ne
rect 10161 20953 13182 20964
tri 13182 20953 13697 21468 sw
tri 13892 20953 14407 21468 ne
rect 14407 21293 16894 21468
tri 16894 21293 17603 22002 sw
tri 17603 21293 18312 22002 ne
rect 18312 21486 20945 22002
tri 20945 21486 21655 22196 sw
tri 21655 21486 22365 22196 ne
rect 22365 21662 25191 22196
tri 25191 21662 25725 22196 sw
tri 25900 21662 26434 22196 ne
rect 26434 21662 29436 22196
rect 22365 21486 25725 21662
rect 18312 21293 21655 21486
rect 14407 20953 17603 21293
tri 17603 20953 17943 21293 sw
tri 18312 20953 18652 21293 ne
rect 18652 20953 21655 21293
tri 21655 20953 22188 21486 sw
tri 22365 20953 22898 21486 ne
rect 22898 20953 25725 21486
tri 25725 20953 26434 21662 sw
tri 26434 20953 27143 21662 ne
rect 27143 20953 29436 21662
tri 29436 20953 30679 22196 sw
rect -25900 20780 -23245 20953
rect -29436 20071 -28025 20780
tri -28025 20071 -27316 20780 nw
tri -27316 20071 -26607 20780 se
rect -26607 20606 -23245 20780
tri -23245 20606 -22898 20953 nw
tri -22535 20606 -22188 20953 se
rect -22188 20606 -19175 20953
rect -26607 20071 -23955 20606
rect -29436 19362 -28734 20071
tri -28734 19362 -28025 20071 nw
tri -28025 19362 -27316 20071 se
rect -27316 19896 -23955 20071
tri -23955 19896 -23245 20606 nw
tri -23245 19896 -22535 20606 se
rect -22535 20430 -19175 20606
tri -19175 20430 -18652 20953 nw
tri -18466 20430 -17943 20953 se
rect -17943 20430 -14930 20953
tri -14930 20430 -14407 20953 nw
tri -13892 20758 -13697 20953 se
rect -13697 20758 -10356 20953
tri -10356 20758 -10161 20953 nw
tri 10161 20758 10356 20953 ne
rect 10356 20758 13697 20953
tri 13697 20758 13892 20953 sw
tri 14407 20758 14602 20953 ne
rect 14602 20758 17943 20953
tri -14220 20430 -13892 20758 se
rect -13892 20430 -10684 20758
tri -10684 20430 -10356 20758 nw
tri 10356 20430 10684 20758 ne
rect 10684 20430 13892 20758
tri 13892 20430 14220 20758 sw
tri 14602 20430 14930 20758 ne
rect 14930 20430 17943 20758
rect -22535 19896 -19709 20430
tri -19709 19896 -19175 20430 nw
tri -19000 19896 -18466 20430 se
rect -18466 19896 -15464 20430
tri -15464 19896 -14930 20430 nw
tri -14754 19896 -14220 20430 se
rect -14220 19896 -11218 20430
tri -11218 19896 -10684 20430 nw
tri 10684 19896 11218 20430 ne
rect 11218 20048 14220 20430
tri 14220 20048 14602 20430 sw
tri 14930 20048 15312 20430 ne
rect 15312 20244 17943 20430
tri 17943 20244 18652 20953 sw
tri 18652 20244 19361 20953 ne
rect 19361 20419 22188 20953
tri 22188 20419 22722 20953 sw
tri 22898 20419 23432 20953 ne
rect 23432 20419 26434 20953
rect 19361 20244 22722 20419
rect 15312 20048 18652 20244
rect 11218 19896 14602 20048
tri 14602 19896 14754 20048 sw
tri 15312 19896 15464 20048 ne
rect 15464 19896 18652 20048
tri 18652 19896 19000 20244 sw
tri 19361 19896 19709 20244 ne
rect 19709 19896 22722 20244
rect -27316 19362 -24489 19896
tri -24489 19362 -23955 19896 nw
tri -23432 19709 -23245 19896 se
rect -23245 19709 -19896 19896
tri -19896 19709 -19709 19896 nw
tri -19187 19709 -19000 19896 se
rect -19000 19709 -15651 19896
tri -15651 19709 -15464 19896 nw
tri -14941 19709 -14754 19896 se
rect -14754 19709 -11405 19896
tri -11405 19709 -11218 19896 nw
tri 11218 19709 11405 19896 ne
rect 11405 19709 14754 19896
tri 14754 19709 14941 19896 sw
tri 15464 19709 15651 19896 ne
rect 15651 19709 19000 19896
tri 19000 19709 19187 19896 sw
tri 19709 19709 19896 19896 ne
rect 19896 19709 22722 19896
tri 22722 19709 23432 20419 sw
tri 23432 19709 24142 20419 ne
rect 24142 20244 26434 20419
tri 26434 20244 27143 20953 sw
tri 27143 20244 27852 20953 ne
rect 27852 20244 30679 20953
rect 24142 19709 27143 20244
tri -23779 19362 -23432 19709 se
rect -23432 19362 -20243 19709
tri -20243 19362 -19896 19709 nw
tri -19534 19362 -19187 19709 se
rect -19187 19362 -15998 19709
tri -15998 19362 -15651 19709 nw
tri -15288 19362 -14941 19709 se
rect -14941 19362 -11752 19709
tri -11752 19362 -11405 19709 nw
tri 11405 19362 11752 19709 ne
rect 11752 19362 14941 19709
tri 14941 19362 15288 19709 sw
tri 15651 19362 15998 19709 ne
rect 15998 19362 19187 19709
tri 19187 19362 19534 19709 sw
tri 19896 19362 20243 19709 ne
rect 20243 19362 23432 19709
tri 23432 19362 23779 19709 sw
tri 24142 19362 24489 19709 ne
rect 24489 19535 27143 19709
tri 27143 19535 27852 20244 sw
tri 27852 19535 28561 20244 ne
rect 28561 19535 30679 20244
rect 24489 19369 27852 19535
tri 27852 19369 28018 19535 sw
tri 28561 19369 28727 19535 ne
rect 28727 19369 30679 19535
rect 24489 19362 28018 19369
tri -32804 18828 -32270 19362 se
rect -32270 18828 -29268 19362
tri -29268 18828 -28734 19362 nw
tri -28559 18828 -28025 19362 se
rect -28025 18828 -25023 19362
tri -25023 18828 -24489 19362 nw
tri -24313 18828 -23779 19362 se
rect -23779 18828 -20777 19362
tri -20777 18828 -20243 19362 nw
tri -20068 18828 -19534 19362 se
rect -19534 18828 -16532 19362
tri -16532 18828 -15998 19362 nw
tri -15822 18828 -15288 19362 se
rect -15288 18828 -12286 19362
tri -12286 18828 -11752 19362 nw
tri 11752 18828 12286 19362 ne
rect 12286 18828 15288 19362
tri 15288 18828 15822 19362 sw
tri 15998 18828 16532 19362 ne
rect 16532 19175 19534 19362
tri 19534 19175 19721 19362 sw
tri 20243 19175 20430 19362 ne
rect 20430 19175 23779 19362
rect 16532 18828 19721 19175
tri 19721 18828 20068 19175 sw
tri 20430 18828 20777 19175 ne
rect 20777 18999 23779 19175
tri 23779 18999 24142 19362 sw
tri 24489 18999 24852 19362 ne
rect 24852 18999 28018 19362
rect 20777 18828 24142 18999
tri 24142 18828 24313 18999 sw
tri 24852 18828 25023 18999 ne
rect 25023 18828 28018 18999
tri 28018 18828 28559 19369 sw
tri 28727 18828 29268 19369 ne
rect 29268 18828 30679 19369
tri -32972 18660 -32804 18828 se
rect -32804 18660 -29436 18828
tri -29436 18660 -29268 18828 nw
tri -28727 18660 -28559 18828 se
rect -28559 18660 -25191 18828
tri -25191 18660 -25023 18828 nw
tri -24481 18660 -24313 18828 se
rect -24313 18660 -20945 18828
tri -20945 18660 -20777 18828 nw
tri -20236 18660 -20068 18828 se
rect -20068 18660 -16700 18828
tri -16700 18660 -16532 18828 nw
tri -15990 18660 -15822 18828 se
rect -15822 18660 -12454 18828
tri -12454 18660 -12286 18828 nw
tri 12286 18660 12454 18828 ne
rect 12454 18660 15822 18828
tri 15822 18660 15990 18828 sw
tri 16532 18660 16700 18828 ne
rect 16700 18660 20068 18828
tri 20068 18660 20236 18828 sw
tri 20777 18660 20945 18828 ne
rect 20945 18660 24313 18828
tri 24313 18660 24481 18828 sw
tri 25023 18660 25191 18828 ne
rect 25191 18660 28559 18828
tri 28559 18660 28727 18828 sw
tri 29268 18660 29436 18828 ne
rect 29436 18660 30679 18828
tri 30679 18660 32972 20953 sw
tri -35806 15826 -32972 18660 se
rect -32972 17951 -30145 18660
tri -30145 17951 -29436 18660 nw
tri -29436 17951 -28727 18660 se
rect -28727 17951 -25901 18660
rect -32972 17244 -30852 17951
tri -30852 17244 -30145 17951 nw
tri -30143 17244 -29436 17951 se
rect -29436 17950 -25901 17951
tri -25901 17950 -25191 18660 nw
tri -25191 17950 -24481 18660 se
rect -24481 17951 -21654 18660
tri -21654 17951 -20945 18660 nw
tri -20430 18466 -20236 18660 se
rect -20236 18466 -16894 18660
tri -16894 18466 -16700 18660 nw
tri -16184 18466 -15990 18660 se
rect -15990 18466 -12648 18660
tri -12648 18466 -12454 18660 nw
tri 12454 18466 12648 18660 ne
rect 12648 18466 15990 18660
tri 15990 18466 16184 18660 sw
tri 16700 18466 16894 18660 ne
rect 16894 18466 20236 18660
tri 20236 18466 20430 18660 sw
tri 20945 18466 21139 18660 ne
rect 21139 18466 24481 18660
tri -20945 17951 -20430 18466 se
rect -20430 18138 -17222 18466
tri -17222 18138 -16894 18466 nw
tri -16512 18138 -16184 18466 se
rect -16184 18138 -13686 18466
rect -20430 17951 -17932 18138
rect -24481 17950 -22002 17951
rect -29436 17417 -26434 17950
tri -26434 17417 -25901 17950 nw
tri -25724 17417 -25191 17950 se
rect -25191 17603 -22002 17950
tri -22002 17603 -21654 17951 nw
tri -21293 17603 -20945 17951 se
rect -20945 17603 -17932 17951
rect -25191 17417 -22188 17603
tri -22188 17417 -22002 17603 nw
tri -21479 17417 -21293 17603 se
rect -21293 17428 -17932 17603
tri -17932 17428 -17222 18138 nw
tri -17222 17428 -16512 18138 se
rect -16512 17428 -13686 18138
tri -13686 17428 -12648 18466 nw
tri 12648 17428 13686 18466 ne
rect 13686 17932 16184 18466
tri 16184 17932 16718 18466 sw
tri 16894 17932 17428 18466 ne
rect 17428 17932 20430 18466
rect 13686 17428 16718 17932
rect -21293 17417 -17943 17428
tri -17943 17417 -17932 17428 nw
tri -17233 17417 -17222 17428 se
rect -17222 17417 -13697 17428
tri -13697 17417 -13686 17428 nw
tri 13686 17417 13697 17428 ne
rect 13697 17417 16718 17428
tri 16718 17417 17233 17932 sw
tri 17428 17417 17943 17932 ne
rect 17943 17757 20430 17932
tri 20430 17757 21139 18466 sw
tri 21139 17757 21848 18466 ne
rect 21848 17950 24481 18466
tri 24481 17950 25191 18660 sw
tri 25191 17950 25901 18660 ne
rect 25901 18126 28727 18660
tri 28727 18126 29261 18660 sw
tri 29436 18126 29970 18660 ne
rect 29970 18126 32972 18660
rect 25901 17950 29261 18126
rect 21848 17757 25191 17950
rect 17943 17417 21139 17757
tri 21139 17417 21479 17757 sw
tri 21848 17417 22188 17757 ne
rect 22188 17417 25191 17757
tri 25191 17417 25724 17950 sw
tri 25901 17417 26434 17950 ne
rect 26434 17417 29261 17950
tri 29261 17417 29970 18126 sw
tri 29970 17417 30679 18126 ne
rect 30679 17417 32972 18126
tri 32972 17417 34215 18660 sw
rect -29436 17244 -26781 17417
rect -32972 16535 -31561 17244
tri -31561 16535 -30852 17244 nw
tri -30852 16535 -30143 17244 se
rect -30143 17070 -26781 17244
tri -26781 17070 -26434 17417 nw
tri -26071 17070 -25724 17417 se
rect -25724 17070 -22711 17417
rect -30143 16535 -27491 17070
rect -32972 15826 -32270 16535
tri -32270 15826 -31561 16535 nw
tri -31561 15826 -30852 16535 se
rect -30852 16360 -27491 16535
tri -27491 16360 -26781 17070 nw
tri -26781 16360 -26071 17070 se
rect -26071 16894 -22711 17070
tri -22711 16894 -22188 17417 nw
tri -22002 16894 -21479 17417 se
rect -21479 16894 -18466 17417
tri -18466 16894 -17943 17417 nw
tri -17428 17222 -17233 17417 se
rect -17233 17222 -13892 17417
tri -13892 17222 -13697 17417 nw
tri 13697 17222 13892 17417 ne
rect 13892 17222 17233 17417
tri 17233 17222 17428 17417 sw
tri 17943 17222 18138 17417 ne
rect 18138 17222 21479 17417
tri -17756 16894 -17428 17222 se
rect -17428 16894 -14220 17222
tri -14220 16894 -13892 17222 nw
tri 13892 16894 14220 17222 ne
rect 14220 16894 17428 17222
tri 17428 16894 17756 17222 sw
tri 18138 16894 18466 17222 ne
rect 18466 16894 21479 17222
rect -26071 16360 -23245 16894
tri -23245 16360 -22711 16894 nw
tri -22536 16360 -22002 16894 se
rect -22002 16360 -19000 16894
tri -19000 16360 -18466 16894 nw
tri -18290 16360 -17756 16894 se
rect -17756 16360 -14754 16894
tri -14754 16360 -14220 16894 nw
tri 14220 16360 14754 16894 ne
rect 14754 16512 17756 16894
tri 17756 16512 18138 16894 sw
tri 18466 16512 18848 16894 ne
rect 18848 16708 21479 16894
tri 21479 16708 22188 17417 sw
tri 22188 16708 22897 17417 ne
rect 22897 16883 25724 17417
tri 25724 16883 26258 17417 sw
tri 26434 16883 26968 17417 ne
rect 26968 16883 29970 17417
rect 22897 16708 26258 16883
rect 18848 16512 22188 16708
rect 14754 16360 18138 16512
tri 18138 16360 18290 16512 sw
tri 18848 16360 19000 16512 ne
rect 19000 16360 22188 16512
tri 22188 16360 22536 16708 sw
tri 22897 16360 23245 16708 ne
rect 23245 16360 26258 16708
rect -30852 15826 -28025 16360
tri -28025 15826 -27491 16360 nw
tri -26968 16173 -26781 16360 se
rect -26781 16173 -23432 16360
tri -23432 16173 -23245 16360 nw
tri -22723 16173 -22536 16360 se
rect -22536 16173 -19187 16360
tri -19187 16173 -19000 16360 nw
tri -18477 16173 -18290 16360 se
rect -18290 16173 -14941 16360
tri -14941 16173 -14754 16360 nw
tri 14754 16173 14941 16360 ne
rect 14941 16173 18290 16360
tri 18290 16173 18477 16360 sw
tri 19000 16173 19187 16360 ne
rect 19187 16173 22536 16360
tri 22536 16173 22723 16360 sw
tri 23245 16173 23432 16360 ne
rect 23432 16173 26258 16360
tri 26258 16173 26968 16883 sw
tri 26968 16173 27678 16883 ne
rect 27678 16708 29970 16883
tri 29970 16708 30679 17417 sw
tri 30679 16708 31388 17417 ne
rect 31388 16708 34215 17417
rect 27678 16173 30679 16708
tri -27315 15826 -26968 16173 se
rect -26968 15826 -23779 16173
tri -23779 15826 -23432 16173 nw
tri -23070 15826 -22723 16173 se
rect -22723 15826 -19534 16173
tri -19534 15826 -19187 16173 nw
tri -18824 15826 -18477 16173 se
rect -18477 15826 -15288 16173
tri -15288 15826 -14941 16173 nw
tri 14941 15826 15288 16173 ne
rect 15288 15826 18477 16173
tri 18477 15826 18824 16173 sw
tri 19187 15826 19534 16173 ne
rect 19534 15826 22723 16173
tri 22723 15826 23070 16173 sw
tri 23432 15826 23779 16173 ne
rect 23779 15826 26968 16173
tri 26968 15826 27315 16173 sw
tri 27678 15826 28025 16173 ne
rect 28025 15999 30679 16173
tri 30679 15999 31388 16708 sw
tri 31388 15999 32097 16708 ne
rect 32097 15999 34215 16708
rect 28025 15833 31388 15999
tri 31388 15833 31554 15999 sw
tri 32097 15833 32263 15999 ne
rect 32263 15833 34215 15999
rect 28025 15826 31554 15833
tri -36340 15292 -35806 15826 se
rect -35806 15292 -32804 15826
tri -32804 15292 -32270 15826 nw
tri -32095 15292 -31561 15826 se
rect -31561 15292 -28559 15826
tri -28559 15292 -28025 15826 nw
tri -27849 15292 -27315 15826 se
rect -27315 15292 -24313 15826
tri -24313 15292 -23779 15826 nw
tri -23604 15292 -23070 15826 se
rect -23070 15292 -20068 15826
tri -20068 15292 -19534 15826 nw
tri -19358 15292 -18824 15826 se
rect -18824 15292 -15822 15826
tri -15822 15292 -15288 15826 nw
tri 15288 15292 15822 15826 ne
rect 15822 15292 18824 15826
tri 18824 15292 19358 15826 sw
tri 19534 15292 20068 15826 ne
rect 20068 15639 23070 15826
tri 23070 15639 23257 15826 sw
tri 23779 15639 23966 15826 ne
rect 23966 15639 27315 15826
rect 20068 15292 23257 15639
tri 23257 15292 23604 15639 sw
tri 23966 15292 24313 15639 ne
rect 24313 15463 27315 15639
tri 27315 15463 27678 15826 sw
tri 28025 15463 28388 15826 ne
rect 28388 15463 31554 15826
rect 24313 15292 27678 15463
tri 27678 15292 27849 15463 sw
tri 28388 15292 28559 15463 ne
rect 28559 15292 31554 15463
tri 31554 15292 32095 15833 sw
tri 32263 15292 32804 15833 ne
rect 32804 15292 34215 15833
tri -36508 15124 -36340 15292 se
rect -36340 15124 -32972 15292
tri -32972 15124 -32804 15292 nw
tri -32263 15124 -32095 15292 se
rect -32095 15124 -28727 15292
tri -28727 15124 -28559 15292 nw
tri -28017 15124 -27849 15292 se
rect -27849 15124 -24481 15292
tri -24481 15124 -24313 15292 nw
tri -23772 15124 -23604 15292 se
rect -23604 15124 -20236 15292
tri -20236 15124 -20068 15292 nw
tri -19526 15124 -19358 15292 se
rect -19358 15124 -15990 15292
tri -15990 15124 -15822 15292 nw
tri 15822 15124 15990 15292 ne
rect 15990 15124 19358 15292
tri 19358 15124 19526 15292 sw
tri 20068 15124 20236 15292 ne
rect 20236 15124 23604 15292
tri 23604 15124 23772 15292 sw
tri 24313 15124 24481 15292 ne
rect 24481 15124 27849 15292
tri 27849 15124 28017 15292 sw
tri 28559 15124 28727 15292 ne
rect 28727 15124 32095 15292
tri 32095 15124 32263 15292 sw
tri 32804 15124 32972 15292 ne
rect 32972 15124 34215 15292
tri 34215 15124 36508 17417 sw
rect -36508 14590 -33506 15124
tri -33506 14590 -32972 15124 nw
tri -32797 14590 -32263 15124 se
rect -32263 14590 -29437 15124
rect -36508 -14590 -34008 14590
tri -34008 14088 -33506 14590 nw
tri -33299 14088 -32797 14590 se
rect -32797 14414 -29437 14590
tri -29437 14414 -28727 15124 nw
tri -28727 14414 -28017 15124 se
rect -28017 14415 -25190 15124
tri -25190 14415 -24481 15124 nw
tri -23966 14930 -23772 15124 se
rect -23772 14930 -20430 15124
tri -20430 14930 -20236 15124 nw
tri -19720 14930 -19526 15124 se
rect -19526 14930 -16184 15124
tri -16184 14930 -15990 15124 nw
tri 15990 14930 16184 15124 ne
rect 16184 14930 19526 15124
tri 19526 14930 19720 15124 sw
tri 20236 14930 20430 15124 ne
rect 20430 14930 23772 15124
tri 23772 14930 23966 15124 sw
tri 24481 14930 24675 15124 ne
rect 24675 14930 28017 15124
tri -24481 14415 -23966 14930 se
rect -23966 14602 -20758 14930
tri -20758 14602 -20430 14930 nw
tri -20048 14602 -19720 14930 se
rect -19720 14602 -17026 14930
rect -23966 14415 -21272 14602
rect -28017 14414 -25517 14415
rect -32797 14088 -29763 14414
tri -29763 14088 -29437 14414 nw
tri -29053 14088 -28727 14414 se
rect -28727 14088 -25517 14414
tri -25517 14088 -25190 14415 nw
tri -24808 14088 -24481 14415 se
rect -24481 14088 -21272 14415
tri -21272 14088 -20758 14602 nw
tri -20562 14088 -20048 14602 se
rect -20048 14088 -17026 14602
tri -17026 14088 -16184 14930 nw
tri 16184 14088 17026 14930 ne
rect 17026 14396 19720 14930
tri 19720 14396 20254 14930 sw
tri 20430 14396 20964 14930 ne
rect 20964 14396 23966 14930
rect 17026 14088 20254 14396
tri 20254 14088 20562 14396 sw
tri 20964 14088 21272 14396 ne
rect 21272 14221 23966 14396
tri 23966 14221 24675 14930 sw
tri 24675 14221 25384 14930 ne
rect 25384 14414 28017 14930
tri 28017 14414 28727 15124 sw
tri 28727 14414 29437 15124 ne
rect 29437 14590 32263 15124
tri 32263 14590 32797 15124 sw
tri 32972 14590 33506 15124 ne
rect 33506 14590 36508 15124
rect 29437 14414 32797 14590
rect 25384 14221 28727 14414
rect 21272 14088 24675 14221
tri 24675 14088 24808 14221 sw
tri 25384 14088 25517 14221 ne
rect 25517 14088 28727 14221
tri 28727 14088 29053 14414 sw
tri 29437 14088 29763 14414 ne
rect 29763 14088 32797 14414
tri 32797 14088 33299 14590 sw
tri 33506 14088 34008 14590 ne
tri -33506 13881 -33299 14088 se
rect -33299 13881 -29970 14088
tri -29970 13881 -29763 14088 nw
tri -29260 13881 -29053 14088 se
rect -29053 14067 -25538 14088
tri -25538 14067 -25517 14088 nw
tri -24829 14067 -24808 14088 se
rect -24808 14067 -21468 14088
rect -29053 13881 -25724 14067
tri -25724 13881 -25538 14067 nw
tri -25015 13881 -24829 14067 se
rect -24829 13892 -21468 14067
tri -21468 13892 -21272 14088 nw
tri -20758 13892 -20562 14088 se
rect -20562 13892 -17222 14088
tri -17222 13892 -17026 14088 nw
tri 17026 13892 17222 14088 ne
rect 17222 13892 20562 14088
rect -24829 13881 -21479 13892
tri -21479 13881 -21468 13892 nw
tri -20769 13881 -20758 13892 se
rect -20758 13881 -17233 13892
tri -17233 13881 -17222 13892 nw
tri 17222 13881 17233 13892 ne
rect 17233 13881 20562 13892
tri 20562 13881 20769 14088 sw
tri 21272 13881 21479 14088 ne
rect 21479 13881 24808 14088
tri 24808 13881 25015 14088 sw
tri 25517 13881 25724 14088 ne
rect 25724 13881 29053 14088
tri 29053 13881 29260 14088 sw
tri 29763 13881 29970 14088 ne
rect 29970 13881 33299 14088
tri 33299 13881 33506 14088 sw
rect -33506 13534 -30317 13881
tri -30317 13534 -29970 13881 nw
tri -29607 13534 -29260 13881 se
rect -29260 13534 -26247 13881
rect -33506 -13347 -31006 13534
tri -31006 12845 -30317 13534 nw
tri -30296 12845 -29607 13534 se
rect -29607 13358 -26247 13534
tri -26247 13358 -25724 13881 nw
tri -25538 13358 -25015 13881 se
rect -25015 13358 -22002 13881
tri -22002 13358 -21479 13881 nw
tri -20964 13686 -20769 13881 se
rect -20769 13686 -17428 13881
tri -17428 13686 -17233 13881 nw
tri 17233 13686 17428 13881 ne
rect 17428 13686 20769 13881
tri 20769 13686 20964 13881 sw
tri 21479 13686 21674 13881 ne
rect 21674 13686 25015 13881
tri -21292 13358 -20964 13686 se
rect -20964 13358 -17756 13686
tri -17756 13358 -17428 13686 nw
tri 17428 13358 17756 13686 ne
rect 17756 13358 20964 13686
tri 20964 13358 21292 13686 sw
tri 21674 13358 22002 13686 ne
rect 22002 13358 25015 13686
rect -29607 12845 -26760 13358
tri -26760 12845 -26247 13358 nw
tri -26051 12845 -25538 13358 se
rect -25538 12845 -22515 13358
tri -22515 12845 -22002 13358 nw
tri -21805 12845 -21292 13358 se
rect -21292 12845 -18269 13358
tri -18269 12845 -17756 13358 nw
tri 17756 12845 18269 13358 ne
rect 18269 12976 21292 13358
tri 21292 12976 21674 13358 sw
tri 22002 12976 22384 13358 ne
rect 22384 13172 25015 13358
tri 25015 13172 25724 13881 sw
tri 25724 13172 26433 13881 ne
rect 26433 13347 29260 13881
tri 29260 13347 29794 13881 sw
tri 29970 13347 30504 13881 ne
rect 30504 13347 33506 13881
rect 26433 13172 29794 13347
rect 22384 12976 25724 13172
rect 18269 12845 21674 12976
tri 21674 12845 21805 12976 sw
tri 22384 12845 22515 12976 ne
rect 22515 12845 25724 12976
tri 25724 12845 26051 13172 sw
tri 26433 12845 26760 13172 ne
rect 26760 12845 29794 13172
tri 29794 12845 30296 13347 sw
tri 30504 12845 31006 13347 ne
tri -30317 12824 -30296 12845 se
rect -30296 12824 -26781 12845
tri -26781 12824 -26760 12845 nw
tri -26072 12824 -26051 12845 se
rect -26051 12824 -22536 12845
tri -22536 12824 -22515 12845 nw
tri -21826 12824 -21805 12845 se
rect -21805 12824 -18290 12845
tri -18290 12824 -18269 12845 nw
tri 18269 12824 18290 12845 ne
rect 18290 12824 21805 12845
tri 21805 12824 21826 12845 sw
tri 22515 12824 22536 12845 ne
rect 22536 12824 26051 12845
tri 26051 12824 26072 12845 sw
tri 26760 12824 26781 12845 ne
rect 26781 12824 30296 12845
tri -30504 12637 -30317 12824 se
rect -30317 12637 -26968 12824
tri -26968 12637 -26781 12824 nw
tri -26259 12637 -26072 12824 se
rect -26072 12637 -22723 12824
tri -22723 12637 -22536 12824 nw
tri -22013 12637 -21826 12824 se
rect -21826 12637 -18477 12824
tri -18477 12637 -18290 12824 nw
tri 18290 12637 18477 12824 ne
rect 18477 12637 21826 12824
tri 21826 12637 22013 12824 sw
tri 22536 12637 22723 12824 ne
rect 22723 12637 26072 12824
tri 26072 12637 26259 12824 sw
tri 26781 12637 26968 12824 ne
rect 26968 12637 30296 12824
tri 30296 12637 30504 12845 sw
rect -30504 12103 -27502 12637
tri -27502 12103 -26968 12637 nw
tri -26793 12103 -26259 12637 se
rect -26259 12103 -23433 12637
rect -30504 -12103 -28004 12103
tri -28004 11601 -27502 12103 nw
tri -27295 11601 -26793 12103 se
rect -26793 11927 -23433 12103
tri -23433 11927 -22723 12637 nw
tri -22723 11927 -22013 12637 se
rect -22013 11927 -19513 12637
rect -26793 11601 -23759 11927
tri -23759 11601 -23433 11927 nw
tri -23049 11601 -22723 11927 se
rect -22723 11601 -19513 11927
tri -19513 11601 -18477 12637 nw
tri 18477 11601 19513 12637 ne
rect 19513 11927 22013 12637
tri 22013 11927 22723 12637 sw
tri 22723 11927 23433 12637 ne
rect 23433 12103 26259 12637
tri 26259 12103 26793 12637 sw
tri 26968 12103 27502 12637 ne
rect 27502 12103 30504 12637
rect 23433 11927 26793 12103
rect 19513 11601 22723 11927
tri 22723 11601 23049 11927 sw
tri 23433 11601 23759 11927 ne
rect 23759 11601 26793 11927
tri 26793 11601 27295 12103 sw
tri 27502 11601 28004 12103 ne
tri -27502 11394 -27295 11601 se
rect -27295 11394 -23966 11601
tri -23966 11394 -23759 11601 nw
tri -23256 11394 -23049 11601 se
rect -23049 11394 -19720 11601
tri -19720 11394 -19513 11601 nw
tri 19513 11394 19720 11601 ne
rect 19720 11394 23049 11601
tri 23049 11394 23256 11601 sw
tri 23759 11394 23966 11601 ne
rect 23966 11394 27295 11601
tri 27295 11394 27502 11601 sw
rect -27502 11066 -24294 11394
tri -24294 11066 -23966 11394 nw
tri -23584 11066 -23256 11394 se
rect -23256 11066 -20756 11394
rect -27502 -10860 -25002 11066
tri -25002 10358 -24294 11066 nw
tri -24292 10358 -23584 11066 se
rect -23584 10358 -20756 11066
tri -20756 10358 -19720 11394 nw
tri 19720 10358 20756 11394 ne
rect 20756 10860 23256 11394
tri 23256 10860 23790 11394 sw
tri 23966 10860 24500 11394 ne
rect 24500 10860 27502 11394
rect 20756 10358 23790 10860
tri 23790 10358 24292 10860 sw
tri 24500 10358 25002 10860 ne
tri -24294 10356 -24292 10358 se
rect -24292 10356 -20758 10358
tri -20758 10356 -20756 10358 nw
tri 20756 10356 20758 10358 ne
rect 20758 10356 24292 10358
tri -24500 10150 -24294 10356 se
rect -24294 10150 -20964 10356
tri -20964 10150 -20758 10356 nw
tri 20758 10150 20964 10356 ne
rect 20964 10150 24292 10356
tri 24292 10150 24500 10358 sw
rect -24500 1250 -22000 10150
tri -22000 9114 -20964 10150 nw
tri 20964 9114 22000 10150 ne
rect -24500 929 21000 1250
rect -24500 673 19552 929
rect 19808 673 20076 929
rect 20332 673 20630 929
rect 20886 673 21000 929
rect -24500 435 21000 673
rect -24500 179 19552 435
rect 19808 179 20076 435
rect 20332 179 20630 435
rect 20886 179 21000 435
rect -24500 -179 21000 179
rect -24500 -435 19552 -179
rect 19808 -435 20076 -179
rect 20332 -435 20630 -179
rect 20886 -435 21000 -179
rect -24500 -673 21000 -435
rect -24500 -929 19552 -673
rect 19808 -929 20076 -673
rect 20332 -929 20630 -673
rect 20886 -929 21000 -673
rect -24500 -1250 21000 -929
rect -24500 -10150 -22000 -1250
tri -22000 -10150 -20964 -9114 sw
tri 20964 -10150 22000 -9114 se
rect 22000 -10150 24500 10150
tri -24500 -10356 -24294 -10150 ne
rect -24294 -10356 -20964 -10150
tri -20964 -10356 -20758 -10150 sw
tri 20758 -10356 20964 -10150 se
rect 20964 -10356 24294 -10150
tri 24294 -10356 24500 -10150 nw
tri -24294 -10358 -24292 -10356 ne
rect -24292 -10358 -20758 -10356
tri -20758 -10358 -20756 -10356 sw
tri 20756 -10358 20758 -10356 se
rect 20758 -10358 24292 -10356
tri 24292 -10358 24294 -10356 nw
tri -25002 -10860 -24500 -10358 sw
tri -24292 -10860 -23790 -10358 ne
rect -23790 -10860 -20756 -10358
rect -27502 -11394 -24500 -10860
tri -24500 -11394 -23966 -10860 sw
tri -23790 -11394 -23256 -10860 ne
rect -23256 -11394 -20756 -10860
tri -20756 -11394 -19720 -10358 sw
tri 19720 -11394 20756 -10358 se
rect 20756 -11066 23584 -10358
tri 23584 -11066 24292 -10358 nw
tri 24294 -11066 25002 -10358 se
rect 25002 -11066 27502 10860
rect 20756 -11394 23256 -11066
tri 23256 -11394 23584 -11066 nw
tri 23966 -11394 24294 -11066 se
rect 24294 -11394 27502 -11066
tri -27502 -11601 -27295 -11394 ne
rect -27295 -11601 -23966 -11394
tri -23966 -11601 -23759 -11394 sw
tri -23256 -11601 -23049 -11394 ne
rect -23049 -11601 -19720 -11394
tri -19720 -11601 -19513 -11394 sw
tri 19513 -11601 19720 -11394 se
rect 19720 -11601 23049 -11394
tri 23049 -11601 23256 -11394 nw
tri 23759 -11601 23966 -11394 se
rect 23966 -11601 27295 -11394
tri 27295 -11601 27502 -11394 nw
tri -28004 -12103 -27502 -11601 sw
tri -27295 -12103 -26793 -11601 ne
rect -26793 -11927 -23759 -11601
tri -23759 -11927 -23433 -11601 sw
tri -23049 -11927 -22723 -11601 ne
rect -22723 -11927 -19513 -11601
rect -26793 -12103 -23433 -11927
rect -30504 -12637 -27502 -12103
tri -27502 -12637 -26968 -12103 sw
tri -26793 -12637 -26259 -12103 ne
rect -26259 -12637 -23433 -12103
tri -23433 -12637 -22723 -11927 sw
tri -22723 -12637 -22013 -11927 ne
rect -22013 -12637 -19513 -11927
tri -19513 -12637 -18477 -11601 sw
tri 18477 -12637 19513 -11601 se
rect 19513 -11927 22723 -11601
tri 22723 -11927 23049 -11601 nw
tri 23433 -11927 23759 -11601 se
rect 23759 -11927 26793 -11601
rect 19513 -12637 22013 -11927
tri 22013 -12637 22723 -11927 nw
tri 22723 -12637 23433 -11927 se
rect 23433 -12103 26793 -11927
tri 26793 -12103 27295 -11601 nw
tri 27502 -12103 28004 -11601 se
rect 28004 -12103 30504 12103
rect 23433 -12637 26259 -12103
tri 26259 -12637 26793 -12103 nw
tri 26968 -12637 27502 -12103 se
rect 27502 -12637 30504 -12103
tri -30504 -12824 -30317 -12637 ne
rect -30317 -12824 -26968 -12637
tri -26968 -12824 -26781 -12637 sw
tri -26259 -12824 -26072 -12637 ne
rect -26072 -12824 -22723 -12637
tri -22723 -12824 -22536 -12637 sw
tri -22013 -12824 -21826 -12637 ne
rect -21826 -12824 -18477 -12637
tri -18477 -12824 -18290 -12637 sw
tri 18290 -12824 18477 -12637 se
rect 18477 -12824 21826 -12637
tri 21826 -12824 22013 -12637 nw
tri 22536 -12824 22723 -12637 se
rect 22723 -12824 26072 -12637
tri 26072 -12824 26259 -12637 nw
tri 26781 -12824 26968 -12637 se
rect 26968 -12824 30317 -12637
tri 30317 -12824 30504 -12637 nw
tri -30317 -12845 -30296 -12824 ne
rect -30296 -12845 -26781 -12824
tri -26781 -12845 -26760 -12824 sw
tri -26072 -12845 -26051 -12824 ne
rect -26051 -12845 -22536 -12824
tri -22536 -12845 -22515 -12824 sw
tri -21826 -12845 -21805 -12824 ne
rect -21805 -12845 -18290 -12824
tri -18290 -12845 -18269 -12824 sw
tri 18269 -12845 18290 -12824 se
rect 18290 -12845 21805 -12824
tri 21805 -12845 21826 -12824 nw
tri 22515 -12845 22536 -12824 se
rect 22536 -12845 26051 -12824
tri 26051 -12845 26072 -12824 nw
tri 26760 -12845 26781 -12824 se
rect 26781 -12845 30296 -12824
tri 30296 -12845 30317 -12824 nw
tri -31006 -13347 -30504 -12845 sw
tri -30296 -13347 -29794 -12845 ne
rect -29794 -13172 -26760 -12845
tri -26760 -13172 -26433 -12845 sw
tri -26051 -13172 -25724 -12845 ne
rect -25724 -13172 -22515 -12845
rect -29794 -13347 -26433 -13172
rect -33506 -13881 -30504 -13347
tri -30504 -13881 -29970 -13347 sw
tri -29794 -13881 -29260 -13347 ne
rect -29260 -13881 -26433 -13347
tri -26433 -13881 -25724 -13172 sw
tri -25724 -13358 -25538 -13172 ne
rect -25538 -13358 -22515 -13172
tri -22515 -13358 -22002 -12845 sw
tri -21805 -13358 -21292 -12845 ne
rect -21292 -13358 -18269 -12845
tri -18269 -13358 -17756 -12845 sw
tri 17756 -13358 18269 -12845 se
rect 18269 -13358 21292 -12845
tri 21292 -13358 21805 -12845 nw
tri 22002 -13358 22515 -12845 se
rect 22515 -13358 25538 -12845
tri 25538 -13358 26051 -12845 nw
tri 26247 -13358 26760 -12845 se
rect 26760 -13358 29607 -12845
tri -25538 -13881 -25015 -13358 ne
rect -25015 -13686 -22002 -13358
tri -22002 -13686 -21674 -13358 sw
tri -21292 -13686 -20964 -13358 ne
rect -20964 -13686 -17756 -13358
tri -17756 -13686 -17428 -13358 sw
tri 17428 -13686 17756 -13358 se
rect 17756 -13686 20769 -13358
rect -25015 -13881 -21674 -13686
tri -21674 -13881 -21479 -13686 sw
tri -20964 -13881 -20769 -13686 ne
rect -20769 -13881 -17428 -13686
tri -17428 -13881 -17233 -13686 sw
tri 17233 -13881 17428 -13686 se
rect 17428 -13881 20769 -13686
tri 20769 -13881 21292 -13358 nw
tri 21479 -13881 22002 -13358 se
rect 22002 -13881 25015 -13358
tri 25015 -13881 25538 -13358 nw
tri 25724 -13881 26247 -13358 se
rect 26247 -13534 29607 -13358
tri 29607 -13534 30296 -12845 nw
tri 30317 -13534 31006 -12845 se
rect 31006 -13534 33506 13347
rect 34008 5500 36508 14590
rect 34008 3000 37508 5500
rect 26247 -13881 29260 -13534
tri 29260 -13881 29607 -13534 nw
tri 29970 -13881 30317 -13534 se
rect 30317 -13881 33506 -13534
tri -33506 -14088 -33299 -13881 ne
rect -33299 -14088 -29970 -13881
tri -29970 -14088 -29763 -13881 sw
tri -29260 -14088 -29053 -13881 ne
rect -29053 -14088 -25724 -13881
tri -25724 -14088 -25517 -13881 sw
tri -25015 -14088 -24808 -13881 ne
rect -24808 -14088 -21479 -13881
tri -21479 -14088 -21272 -13881 sw
tri -20769 -13892 -20758 -13881 ne
rect -20758 -13892 -17233 -13881
tri -17233 -13892 -17222 -13881 sw
tri 17222 -13892 17233 -13881 se
rect 17233 -13892 20758 -13881
tri 20758 -13892 20769 -13881 nw
tri 21468 -13892 21479 -13881 se
rect 21479 -13892 24829 -13881
tri -20758 -14088 -20562 -13892 ne
rect -20562 -14088 -17222 -13892
tri -17222 -14088 -17026 -13892 sw
tri 17026 -14088 17222 -13892 se
rect 17222 -14088 20562 -13892
tri 20562 -14088 20758 -13892 nw
tri 21272 -14088 21468 -13892 se
rect 21468 -14067 24829 -13892
tri 24829 -14067 25015 -13881 nw
tri 25538 -14067 25724 -13881 se
rect 25724 -14067 29053 -13881
rect 21468 -14088 24808 -14067
tri 24808 -14088 24829 -14067 nw
tri 25517 -14088 25538 -14067 se
rect 25538 -14088 29053 -14067
tri 29053 -14088 29260 -13881 nw
tri 29763 -14088 29970 -13881 se
rect 29970 -14088 33299 -13881
tri 33299 -14088 33506 -13881 nw
rect 34008 -5500 37508 -3000
tri -34008 -14590 -33506 -14088 sw
tri -33299 -14590 -32797 -14088 ne
rect -32797 -14414 -29763 -14088
tri -29763 -14414 -29437 -14088 sw
tri -29053 -14414 -28727 -14088 ne
rect -28727 -14221 -25517 -14088
tri -25517 -14221 -25384 -14088 sw
tri -24808 -14221 -24675 -14088 ne
rect -24675 -14221 -21272 -14088
rect -28727 -14414 -25384 -14221
rect -32797 -14590 -29437 -14414
rect -36508 -15124 -33506 -14590
tri -33506 -15124 -32972 -14590 sw
tri -32797 -15124 -32263 -14590 ne
rect -32263 -15124 -29437 -14590
tri -29437 -15124 -28727 -14414 sw
tri -28727 -15124 -28017 -14414 ne
rect -28017 -14930 -25384 -14414
tri -25384 -14930 -24675 -14221 sw
tri -24675 -14930 -23966 -14221 ne
rect -23966 -14396 -21272 -14221
tri -21272 -14396 -20964 -14088 sw
tri -20562 -14396 -20254 -14088 ne
rect -20254 -14396 -17026 -14088
rect -23966 -14930 -20964 -14396
tri -20964 -14930 -20430 -14396 sw
tri -20254 -14930 -19720 -14396 ne
rect -19720 -14930 -17026 -14396
tri -17026 -14930 -16184 -14088 sw
tri 16184 -14930 17026 -14088 se
rect 17026 -14602 20048 -14088
tri 20048 -14602 20562 -14088 nw
tri 20758 -14602 21272 -14088 se
rect 21272 -14415 24481 -14088
tri 24481 -14415 24808 -14088 nw
tri 25190 -14415 25517 -14088 se
rect 25517 -14414 28727 -14088
tri 28727 -14414 29053 -14088 nw
tri 29437 -14414 29763 -14088 se
rect 29763 -14414 32797 -14088
rect 25517 -14415 28017 -14414
rect 21272 -14602 23772 -14415
rect 17026 -14930 19720 -14602
tri 19720 -14930 20048 -14602 nw
tri 20430 -14930 20758 -14602 se
rect 20758 -14930 23772 -14602
rect -28017 -15124 -24675 -14930
tri -24675 -15124 -24481 -14930 sw
tri -23966 -15124 -23772 -14930 ne
rect -23772 -15124 -20430 -14930
tri -20430 -15124 -20236 -14930 sw
tri -19720 -15124 -19526 -14930 ne
rect -19526 -15124 -16184 -14930
tri -16184 -15124 -15990 -14930 sw
tri 15990 -15124 16184 -14930 se
rect 16184 -15124 19526 -14930
tri 19526 -15124 19720 -14930 nw
tri 20236 -15124 20430 -14930 se
rect 20430 -15124 23772 -14930
tri 23772 -15124 24481 -14415 nw
tri 24481 -15124 25190 -14415 se
rect 25190 -15124 28017 -14415
tri 28017 -15124 28727 -14414 nw
tri 28727 -15124 29437 -14414 se
rect 29437 -14590 32797 -14414
tri 32797 -14590 33299 -14088 nw
tri 33506 -14590 34008 -14088 se
rect 34008 -14590 36508 -5500
rect 29437 -15124 32263 -14590
tri 32263 -15124 32797 -14590 nw
tri 32972 -15124 33506 -14590 se
rect 33506 -15124 36508 -14590
tri -36508 -15292 -36340 -15124 ne
rect -36340 -15292 -32972 -15124
tri -32972 -15292 -32804 -15124 sw
tri -32263 -15292 -32095 -15124 ne
rect -32095 -15292 -28727 -15124
tri -28727 -15292 -28559 -15124 sw
tri -28017 -15292 -27849 -15124 ne
rect -27849 -15292 -24481 -15124
tri -24481 -15292 -24313 -15124 sw
tri -23772 -15292 -23604 -15124 ne
rect -23604 -15292 -20236 -15124
tri -20236 -15292 -20068 -15124 sw
tri -19526 -15292 -19358 -15124 ne
rect -19358 -15292 -15990 -15124
tri -15990 -15292 -15822 -15124 sw
tri 15822 -15292 15990 -15124 se
rect 15990 -15292 19358 -15124
tri 19358 -15292 19526 -15124 nw
tri 20068 -15292 20236 -15124 se
rect 20236 -15292 23604 -15124
tri 23604 -15292 23772 -15124 nw
tri 24313 -15292 24481 -15124 se
rect 24481 -15292 27849 -15124
tri 27849 -15292 28017 -15124 nw
tri 28559 -15292 28727 -15124 se
rect 28727 -15292 32095 -15124
tri 32095 -15292 32263 -15124 nw
tri 32804 -15292 32972 -15124 se
rect 32972 -15292 36340 -15124
tri 36340 -15292 36508 -15124 nw
tri -36340 -17417 -34215 -15292 ne
rect -34215 -16001 -32804 -15292
tri -32804 -16001 -32095 -15292 sw
tri -32095 -16001 -31386 -15292 ne
rect -31386 -15826 -28559 -15292
tri -28559 -15826 -28025 -15292 sw
tri -27849 -15826 -27315 -15292 ne
rect -27315 -15639 -24313 -15292
tri -24313 -15639 -23966 -15292 sw
tri -23604 -15639 -23257 -15292 ne
rect -23257 -15639 -20068 -15292
rect -27315 -15826 -23966 -15639
tri -23966 -15826 -23779 -15639 sw
tri -23257 -15826 -23070 -15639 ne
rect -23070 -15826 -20068 -15639
tri -20068 -15826 -19534 -15292 sw
tri -19358 -15826 -18824 -15292 ne
rect -18824 -15826 -15822 -15292
tri -15822 -15826 -15288 -15292 sw
tri 15288 -15826 15822 -15292 se
rect 15822 -15826 18824 -15292
tri 18824 -15826 19358 -15292 nw
tri 19534 -15826 20068 -15292 se
rect 20068 -15826 23070 -15292
tri 23070 -15826 23604 -15292 nw
tri 23779 -15826 24313 -15292 se
rect 24313 -15826 27315 -15292
tri 27315 -15826 27849 -15292 nw
tri 28025 -15826 28559 -15292 se
rect 28559 -15826 31561 -15292
tri 31561 -15826 32095 -15292 nw
tri 32270 -15826 32804 -15292 se
rect 32804 -15826 35806 -15292
tri 35806 -15826 36340 -15292 nw
rect -31386 -16001 -28025 -15826
rect -34215 -16708 -32095 -16001
tri -32095 -16708 -31388 -16001 sw
tri -31386 -16708 -30679 -16001 ne
rect -30679 -16173 -28025 -16001
tri -28025 -16173 -27678 -15826 sw
tri -27315 -16173 -26968 -15826 ne
rect -26968 -16173 -23779 -15826
tri -23779 -16173 -23432 -15826 sw
tri -23070 -16173 -22723 -15826 ne
rect -22723 -16173 -19534 -15826
tri -19534 -16173 -19187 -15826 sw
tri -18824 -16173 -18477 -15826 ne
rect -18477 -16173 -15288 -15826
tri -15288 -16173 -14941 -15826 sw
tri 14941 -16173 15288 -15826 se
rect 15288 -16173 18477 -15826
tri 18477 -16173 18824 -15826 nw
tri 19187 -16173 19534 -15826 se
rect 19534 -16173 22723 -15826
tri 22723 -16173 23070 -15826 nw
tri 23432 -16173 23779 -15826 se
rect 23779 -16173 26781 -15826
rect -30679 -16708 -27678 -16173
rect -34215 -17417 -31388 -16708
tri -31388 -17417 -30679 -16708 sw
tri -30679 -17417 -29970 -16708 ne
rect -29970 -16883 -27678 -16708
tri -27678 -16883 -26968 -16173 sw
tri -26968 -16360 -26781 -16173 ne
rect -26781 -16360 -23432 -16173
tri -23432 -16360 -23245 -16173 sw
tri -22723 -16360 -22536 -16173 ne
rect -22536 -16360 -19187 -16173
tri -19187 -16360 -19000 -16173 sw
tri -18477 -16360 -18290 -16173 ne
rect -18290 -16360 -14941 -16173
tri -14941 -16360 -14754 -16173 sw
tri 14754 -16360 14941 -16173 se
rect 14941 -16360 18290 -16173
tri 18290 -16360 18477 -16173 nw
tri 19000 -16360 19187 -16173 se
rect 19187 -16360 22536 -16173
tri 22536 -16360 22723 -16173 nw
tri 23245 -16360 23432 -16173 se
rect 23432 -16360 26781 -16173
tri 26781 -16360 27315 -15826 nw
tri 27491 -16360 28025 -15826 se
rect 28025 -16360 30852 -15826
tri -26781 -16883 -26258 -16360 ne
rect -26258 -16708 -23245 -16360
tri -23245 -16708 -22897 -16360 sw
tri -22536 -16708 -22188 -16360 ne
rect -22188 -16708 -19000 -16360
rect -26258 -16883 -22897 -16708
rect -29970 -17417 -26968 -16883
tri -26968 -17417 -26434 -16883 sw
tri -26258 -17417 -25724 -16883 ne
rect -25724 -17417 -22897 -16883
tri -22897 -17417 -22188 -16708 sw
tri -22188 -16894 -22002 -16708 ne
rect -22002 -16894 -19000 -16708
tri -19000 -16894 -18466 -16360 sw
tri -18290 -16894 -17756 -16360 ne
rect -17756 -16894 -14754 -16360
tri -14754 -16894 -14220 -16360 sw
tri 14220 -16894 14754 -16360 se
rect 14754 -16894 17756 -16360
tri 17756 -16894 18290 -16360 nw
tri 18466 -16894 19000 -16360 se
rect 19000 -16894 22002 -16360
tri 22002 -16894 22536 -16360 nw
tri 22711 -16894 23245 -16360 se
rect 23245 -16894 26071 -16360
tri -22002 -17417 -21479 -16894 ne
rect -21479 -17222 -18466 -16894
tri -18466 -17222 -18138 -16894 sw
tri -17756 -17222 -17428 -16894 ne
rect -17428 -17222 -14220 -16894
tri -14220 -17222 -13892 -16894 sw
tri 13892 -17222 14220 -16894 se
rect 14220 -17222 17233 -16894
rect -21479 -17417 -18138 -17222
tri -18138 -17417 -17943 -17222 sw
tri -17428 -17417 -17233 -17222 ne
rect -17233 -17417 -13892 -17222
tri -13892 -17417 -13697 -17222 sw
tri 13697 -17417 13892 -17222 se
rect 13892 -17417 17233 -17222
tri 17233 -17417 17756 -16894 nw
tri 17943 -17417 18466 -16894 se
rect 18466 -17417 21479 -16894
tri 21479 -17417 22002 -16894 nw
tri 22188 -17417 22711 -16894 se
rect 22711 -17070 26071 -16894
tri 26071 -17070 26781 -16360 nw
tri 26781 -17070 27491 -16360 se
rect 27491 -16535 30852 -16360
tri 30852 -16535 31561 -15826 nw
tri 31561 -16535 32270 -15826 se
rect 32270 -16535 32804 -15826
rect 27491 -17070 30143 -16535
rect 22711 -17417 25724 -17070
tri 25724 -17417 26071 -17070 nw
tri 26434 -17417 26781 -17070 se
rect 26781 -17244 30143 -17070
tri 30143 -17244 30852 -16535 nw
tri 30852 -17244 31561 -16535 se
rect 31561 -17244 32804 -16535
rect 26781 -17410 29977 -17244
tri 29977 -17410 30143 -17244 nw
tri 30686 -17410 30852 -17244 se
rect 30852 -17410 32804 -17244
rect 26781 -17417 29268 -17410
tri -34215 -18660 -32972 -17417 ne
rect -32972 -18126 -30679 -17417
tri -30679 -18126 -29970 -17417 sw
tri -29970 -18126 -29261 -17417 ne
rect -29261 -17950 -26434 -17417
tri -26434 -17950 -25901 -17417 sw
tri -25724 -17950 -25191 -17417 ne
rect -25191 -17757 -22188 -17417
tri -22188 -17757 -21848 -17417 sw
tri -21479 -17757 -21139 -17417 ne
rect -21139 -17757 -17943 -17417
rect -25191 -17950 -21848 -17757
rect -29261 -18126 -25901 -17950
rect -32972 -18660 -29970 -18126
tri -29970 -18660 -29436 -18126 sw
tri -29261 -18660 -28727 -18126 ne
rect -28727 -18660 -25901 -18126
tri -25901 -18660 -25191 -17950 sw
tri -25191 -18660 -24481 -17950 ne
rect -24481 -18466 -21848 -17950
tri -21848 -18466 -21139 -17757 sw
tri -21139 -18466 -20430 -17757 ne
rect -20430 -17932 -17943 -17757
tri -17943 -17932 -17428 -17417 sw
tri -17233 -17428 -17222 -17417 ne
rect -17222 -17428 -13697 -17417
tri -13697 -17428 -13686 -17417 sw
tri 13686 -17428 13697 -17417 se
rect 13697 -17428 17222 -17417
tri 17222 -17428 17233 -17417 nw
tri 17932 -17428 17943 -17417 se
rect 17943 -17428 21293 -17417
tri -17222 -17932 -16718 -17428 ne
rect -16718 -17932 -13686 -17428
rect -20430 -18466 -17428 -17932
tri -17428 -18466 -16894 -17932 sw
tri -16718 -18466 -16184 -17932 ne
rect -16184 -18466 -13686 -17932
tri -13686 -18466 -12648 -17428 sw
tri 12648 -18466 13686 -17428 se
rect 13686 -18138 16512 -17428
tri 16512 -18138 17222 -17428 nw
tri 17222 -18138 17932 -17428 se
rect 17932 -17603 21293 -17428
tri 21293 -17603 21479 -17417 nw
tri 22002 -17603 22188 -17417 se
rect 22188 -17603 25361 -17417
rect 17932 -17951 20945 -17603
tri 20945 -17951 21293 -17603 nw
tri 21654 -17951 22002 -17603 se
rect 22002 -17780 25361 -17603
tri 25361 -17780 25724 -17417 nw
tri 26071 -17780 26434 -17417 se
rect 26434 -17780 29268 -17417
rect 22002 -17950 25191 -17780
tri 25191 -17950 25361 -17780 nw
tri 25901 -17950 26071 -17780 se
rect 26071 -17950 29268 -17780
rect 22002 -17951 24481 -17950
rect 17932 -18138 20236 -17951
rect 13686 -18466 16184 -18138
tri 16184 -18466 16512 -18138 nw
tri 16894 -18466 17222 -18138 se
rect 17222 -18466 20236 -18138
rect -24481 -18660 -21139 -18466
tri -21139 -18660 -20945 -18466 sw
tri -20430 -18660 -20236 -18466 ne
rect -20236 -18660 -16894 -18466
tri -16894 -18660 -16700 -18466 sw
tri -16184 -18660 -15990 -18466 ne
rect -15990 -18660 -12648 -18466
tri -12648 -18660 -12454 -18466 sw
tri 12454 -18660 12648 -18466 se
rect 12648 -18660 15990 -18466
tri 15990 -18660 16184 -18466 nw
tri 16700 -18660 16894 -18466 se
rect 16894 -18660 20236 -18466
tri 20236 -18660 20945 -17951 nw
tri 20945 -18660 21654 -17951 se
rect 21654 -18660 24481 -17951
tri 24481 -18660 25191 -17950 nw
tri 25191 -18660 25901 -17950 se
rect 25901 -18119 29268 -17950
tri 29268 -18119 29977 -17410 nw
tri 29977 -18119 30686 -17410 se
rect 30686 -18119 32804 -17410
rect 25901 -18660 28727 -18119
tri 28727 -18660 29268 -18119 nw
tri 29436 -18660 29977 -18119 se
rect 29977 -18660 32804 -18119
tri -32972 -18828 -32804 -18660 ne
rect -32804 -18828 -29436 -18660
tri -29436 -18828 -29268 -18660 sw
tri -28727 -18828 -28559 -18660 ne
rect -28559 -18828 -25191 -18660
tri -25191 -18828 -25023 -18660 sw
tri -24481 -18828 -24313 -18660 ne
rect -24313 -18828 -20945 -18660
tri -20945 -18828 -20777 -18660 sw
tri -20236 -18828 -20068 -18660 ne
rect -20068 -18828 -16700 -18660
tri -16700 -18828 -16532 -18660 sw
tri -15990 -18828 -15822 -18660 ne
rect -15822 -18828 -12454 -18660
tri -12454 -18828 -12286 -18660 sw
tri 12286 -18828 12454 -18660 se
rect 12454 -18828 15822 -18660
tri 15822 -18828 15990 -18660 nw
tri 16532 -18828 16700 -18660 se
rect 16700 -18828 20068 -18660
tri 20068 -18828 20236 -18660 nw
tri 20777 -18828 20945 -18660 se
rect 20945 -18828 24313 -18660
tri 24313 -18828 24481 -18660 nw
tri 25023 -18828 25191 -18660 se
rect 25191 -18828 28559 -18660
tri 28559 -18828 28727 -18660 nw
tri 29268 -18828 29436 -18660 se
rect 29436 -18828 32804 -18660
tri 32804 -18828 35806 -15826 nw
tri -32804 -20953 -30679 -18828 ne
rect -30679 -19537 -29268 -18828
tri -29268 -19537 -28559 -18828 sw
tri -28559 -19537 -27850 -18828 ne
rect -27850 -19362 -25023 -18828
tri -25023 -19362 -24489 -18828 sw
tri -24313 -19362 -23779 -18828 ne
rect -23779 -19175 -20777 -18828
tri -20777 -19175 -20430 -18828 sw
tri -20068 -19175 -19721 -18828 ne
rect -19721 -19175 -16532 -18828
rect -23779 -19362 -20430 -19175
tri -20430 -19362 -20243 -19175 sw
tri -19721 -19362 -19534 -19175 ne
rect -19534 -19362 -16532 -19175
tri -16532 -19362 -15998 -18828 sw
tri -15822 -19362 -15288 -18828 ne
rect -15288 -19362 -12286 -18828
tri -12286 -19362 -11752 -18828 sw
tri 11752 -19362 12286 -18828 se
rect 12286 -19362 15288 -18828
tri 15288 -19362 15822 -18828 nw
tri 15998 -19362 16532 -18828 se
rect 16532 -19362 19534 -18828
tri 19534 -19362 20068 -18828 nw
tri 20243 -19362 20777 -18828 se
rect 20777 -19362 23779 -18828
tri 23779 -19362 24313 -18828 nw
tri 24489 -19362 25023 -18828 se
rect 25023 -19362 28025 -18828
tri 28025 -19362 28559 -18828 nw
tri 28734 -19362 29268 -18828 se
rect 29268 -19362 32270 -18828
tri 32270 -19362 32804 -18828 nw
rect -27850 -19537 -24489 -19362
rect -30679 -20244 -28559 -19537
tri -28559 -20244 -27852 -19537 sw
tri -27850 -20244 -27143 -19537 ne
rect -27143 -19709 -24489 -19537
tri -24489 -19709 -24142 -19362 sw
tri -23779 -19709 -23432 -19362 ne
rect -23432 -19709 -20243 -19362
tri -20243 -19709 -19896 -19362 sw
tri -19534 -19709 -19187 -19362 ne
rect -19187 -19709 -15998 -19362
tri -15998 -19709 -15651 -19362 sw
tri -15288 -19709 -14941 -19362 ne
rect -14941 -19709 -11752 -19362
tri -11752 -19709 -11405 -19362 sw
tri 11405 -19709 11752 -19362 se
rect 11752 -19709 14941 -19362
tri 14941 -19709 15288 -19362 nw
tri 15651 -19709 15998 -19362 se
rect 15998 -19709 19187 -19362
tri 19187 -19709 19534 -19362 nw
tri 19896 -19709 20243 -19362 se
rect 20243 -19709 23245 -19362
rect -27143 -20244 -24142 -19709
rect -30679 -20953 -27852 -20244
tri -27852 -20953 -27143 -20244 sw
tri -27143 -20953 -26434 -20244 ne
rect -26434 -20419 -24142 -20244
tri -24142 -20419 -23432 -19709 sw
tri -23432 -19896 -23245 -19709 ne
rect -23245 -19896 -19896 -19709
tri -19896 -19896 -19709 -19709 sw
tri -19187 -19896 -19000 -19709 ne
rect -19000 -19896 -15651 -19709
tri -15651 -19896 -15464 -19709 sw
tri -14941 -19896 -14754 -19709 ne
rect -14754 -19896 -11405 -19709
tri -11405 -19896 -11218 -19709 sw
tri 11218 -19896 11405 -19709 se
rect 11405 -19896 14754 -19709
tri 14754 -19896 14941 -19709 nw
tri 15464 -19896 15651 -19709 se
rect 15651 -19896 19000 -19709
tri 19000 -19896 19187 -19709 nw
tri 19709 -19896 19896 -19709 se
rect 19896 -19896 23245 -19709
tri 23245 -19896 23779 -19362 nw
tri 23955 -19896 24489 -19362 se
rect 24489 -19896 27316 -19362
tri -23245 -20419 -22722 -19896 ne
rect -22722 -20244 -19709 -19896
tri -19709 -20244 -19361 -19896 sw
tri -19000 -20244 -18652 -19896 ne
rect -18652 -20244 -15464 -19896
rect -22722 -20419 -19361 -20244
rect -26434 -20953 -23432 -20419
tri -23432 -20953 -22898 -20419 sw
tri -22722 -20953 -22188 -20419 ne
rect -22188 -20953 -19361 -20419
tri -19361 -20953 -18652 -20244 sw
tri -18652 -20430 -18466 -20244 ne
rect -18466 -20430 -15464 -20244
tri -15464 -20430 -14930 -19896 sw
tri -14754 -20430 -14220 -19896 ne
rect -14220 -20430 -11218 -19896
tri -11218 -20430 -10684 -19896 sw
tri 10684 -20430 11218 -19896 se
rect 11218 -20430 14220 -19896
tri 14220 -20430 14754 -19896 nw
tri 14930 -20430 15464 -19896 se
rect 15464 -20430 18466 -19896
tri 18466 -20430 19000 -19896 nw
tri 19175 -20430 19709 -19896 se
rect 19709 -20430 22535 -19896
tri -18466 -20953 -17943 -20430 ne
rect -17943 -20758 -14930 -20430
tri -14930 -20758 -14602 -20430 sw
tri -14220 -20758 -13892 -20430 ne
rect -13892 -20758 -10684 -20430
tri -10684 -20758 -10356 -20430 sw
tri 10356 -20758 10684 -20430 se
rect 10684 -20758 13697 -20430
rect -17943 -20953 -14602 -20758
tri -14602 -20953 -14407 -20758 sw
tri -13892 -20953 -13697 -20758 ne
rect -13697 -20953 -10356 -20758
tri -10356 -20953 -10161 -20758 sw
tri 10161 -20953 10356 -20758 se
rect 10356 -20953 13697 -20758
tri 13697 -20953 14220 -20430 nw
tri 14407 -20953 14930 -20430 se
rect 14930 -20953 17943 -20430
tri 17943 -20953 18466 -20430 nw
tri 18652 -20953 19175 -20430 se
rect 19175 -20606 22535 -20430
tri 22535 -20606 23245 -19896 nw
tri 23245 -20606 23955 -19896 se
rect 23955 -20071 27316 -19896
tri 27316 -20071 28025 -19362 nw
tri 28025 -20071 28734 -19362 se
rect 28734 -20071 29268 -19362
rect 23955 -20606 26607 -20071
rect 19175 -20953 22188 -20606
tri 22188 -20953 22535 -20606 nw
tri 22898 -20953 23245 -20606 se
rect 23245 -20780 26607 -20606
tri 26607 -20780 27316 -20071 nw
tri 27316 -20780 28025 -20071 se
rect 28025 -20780 29268 -20071
rect 23245 -20946 26441 -20780
tri 26441 -20946 26607 -20780 nw
tri 27150 -20946 27316 -20780 se
rect 27316 -20946 29268 -20780
rect 23245 -20953 25732 -20946
tri -30679 -22196 -29436 -20953 ne
rect -29436 -21662 -27143 -20953
tri -27143 -21662 -26434 -20953 sw
tri -26434 -21662 -25725 -20953 ne
rect -25725 -21486 -22898 -20953
tri -22898 -21486 -22365 -20953 sw
tri -22188 -21486 -21655 -20953 ne
rect -21655 -21293 -18652 -20953
tri -18652 -21293 -18312 -20953 sw
tri -17943 -21293 -17603 -20953 ne
rect -17603 -21293 -14407 -20953
rect -21655 -21486 -18312 -21293
rect -25725 -21662 -22365 -21486
rect -29436 -22196 -26434 -21662
tri -26434 -22196 -25900 -21662 sw
tri -25725 -22196 -25191 -21662 ne
rect -25191 -22196 -22365 -21662
tri -22365 -22196 -21655 -21486 sw
tri -21655 -22196 -20945 -21486 ne
rect -20945 -22002 -18312 -21486
tri -18312 -22002 -17603 -21293 sw
tri -17603 -22002 -16894 -21293 ne
rect -16894 -21468 -14407 -21293
tri -14407 -21468 -13892 -20953 sw
tri -13697 -20964 -13686 -20953 ne
rect -13686 -20964 -10161 -20953
tri -10161 -20964 -10150 -20953 sw
tri 10150 -20964 10161 -20953 se
rect 10161 -20964 13686 -20953
tri 13686 -20964 13697 -20953 nw
tri 14396 -20964 14407 -20953 se
rect 14407 -20964 17757 -20953
tri -13686 -21468 -13182 -20964 ne
rect -13182 -21468 -10150 -20964
rect -16894 -22002 -13892 -21468
tri -13892 -22002 -13358 -21468 sw
tri -13182 -22002 -12648 -21468 ne
rect -12648 -22000 -10150 -21468
tri -10150 -22000 -9114 -20964 sw
tri 9114 -22000 10150 -20964 se
rect 10150 -21674 12976 -20964
tri 12976 -21674 13686 -20964 nw
tri 13686 -21674 14396 -20964 se
rect 14396 -21139 17757 -20964
tri 17757 -21139 17943 -20953 nw
tri 18466 -21139 18652 -20953 se
rect 18652 -21139 21825 -20953
rect 14396 -21487 17409 -21139
tri 17409 -21487 17757 -21139 nw
tri 18118 -21487 18466 -21139 se
rect 18466 -21316 21825 -21139
tri 21825 -21316 22188 -20953 nw
tri 22535 -21316 22898 -20953 se
rect 22898 -21316 25732 -20953
rect 18466 -21486 21655 -21316
tri 21655 -21486 21825 -21316 nw
tri 22365 -21486 22535 -21316 se
rect 22535 -21486 25732 -21316
rect 18466 -21487 20945 -21486
rect 14396 -21674 16700 -21487
rect 10150 -22000 12648 -21674
rect -12648 -22002 12648 -22000
tri 12648 -22002 12976 -21674 nw
tri 13358 -22002 13686 -21674 se
rect 13686 -22002 16700 -21674
rect -20945 -22196 -17603 -22002
tri -17603 -22196 -17409 -22002 sw
tri -16894 -22196 -16700 -22002 ne
rect -16700 -22196 -13358 -22002
tri -13358 -22196 -13164 -22002 sw
tri -12648 -22196 -12454 -22002 ne
rect -12454 -22196 12454 -22002
tri 12454 -22196 12648 -22002 nw
tri 13164 -22196 13358 -22002 se
rect 13358 -22196 16700 -22002
tri 16700 -22196 17409 -21487 nw
tri 17409 -22196 18118 -21487 se
rect 18118 -22196 20945 -21487
tri 20945 -22196 21655 -21486 nw
tri 21655 -22196 22365 -21486 se
rect 22365 -21655 25732 -21486
tri 25732 -21655 26441 -20946 nw
tri 26441 -21655 27150 -20946 se
rect 27150 -21655 29268 -20946
rect 22365 -22196 25191 -21655
tri 25191 -22196 25732 -21655 nw
tri 25900 -22196 26441 -21655 se
rect 26441 -22196 29268 -21655
tri -29436 -22364 -29268 -22196 ne
rect -29268 -22364 -25900 -22196
tri -25900 -22364 -25732 -22196 sw
tri -25191 -22364 -25023 -22196 ne
rect -25023 -22364 -21655 -22196
tri -21655 -22364 -21487 -22196 sw
tri -20945 -22364 -20777 -22196 ne
rect -20777 -22364 -17409 -22196
tri -17409 -22364 -17241 -22196 sw
tri -16700 -22364 -16532 -22196 ne
rect -16532 -22364 -13164 -22196
tri -13164 -22364 -12996 -22196 sw
tri -12454 -22364 -12286 -22196 ne
rect -12286 -22364 12286 -22196
tri 12286 -22364 12454 -22196 nw
tri 12996 -22364 13164 -22196 se
rect 13164 -22364 16532 -22196
tri 16532 -22364 16700 -22196 nw
tri 17241 -22364 17409 -22196 se
rect 17409 -22364 20777 -22196
tri 20777 -22364 20945 -22196 nw
tri 21487 -22364 21655 -22196 se
rect 21655 -22364 25023 -22196
tri 25023 -22364 25191 -22196 nw
tri 25732 -22364 25900 -22196 se
rect 25900 -22364 29268 -22196
tri 29268 -22364 32270 -19362 nw
tri -29268 -24489 -27143 -22364 ne
rect -27143 -23073 -25732 -22364
tri -25732 -23073 -25023 -22364 sw
tri -25023 -23073 -24314 -22364 ne
rect -24314 -22898 -21487 -22364
tri -21487 -22898 -20953 -22364 sw
tri -20777 -22898 -20243 -22364 ne
rect -20243 -22711 -17241 -22364
tri -17241 -22711 -16894 -22364 sw
tri -16532 -22711 -16185 -22364 ne
rect -16185 -22711 -12996 -22364
rect -20243 -22898 -16894 -22711
tri -16894 -22898 -16707 -22711 sw
tri -16185 -22898 -15998 -22711 ne
rect -15998 -22898 -12996 -22711
tri -12996 -22898 -12462 -22364 sw
tri -12286 -22898 -11752 -22364 ne
rect -11752 -22898 11752 -22364
tri 11752 -22898 12286 -22364 nw
tri 12462 -22898 12996 -22364 se
rect 12996 -22898 15998 -22364
tri 15998 -22898 16532 -22364 nw
tri 16707 -22898 17241 -22364 se
rect 17241 -22898 20243 -22364
tri 20243 -22898 20777 -22364 nw
tri 20953 -22898 21487 -22364 se
rect 21487 -22898 24489 -22364
tri 24489 -22898 25023 -22364 nw
tri 25198 -22898 25732 -22364 se
rect 25732 -22898 28734 -22364
tri 28734 -22898 29268 -22364 nw
rect -24314 -23073 -20953 -22898
rect -27143 -23780 -25023 -23073
tri -25023 -23780 -24316 -23073 sw
tri -24314 -23780 -23607 -23073 ne
rect -23607 -23245 -20953 -23073
tri -20953 -23245 -20606 -22898 sw
tri -20243 -23245 -19896 -22898 ne
rect -19896 -23245 -16707 -22898
tri -16707 -23245 -16360 -22898 sw
tri -15998 -23245 -15651 -22898 ne
rect -15651 -23245 -12462 -22898
tri -12462 -23245 -12115 -22898 sw
tri -11752 -23245 -11405 -22898 ne
rect -11405 -23245 11405 -22898
tri 11405 -23245 11752 -22898 nw
tri 12115 -23245 12462 -22898 se
rect 12462 -23245 15651 -22898
tri 15651 -23245 15998 -22898 nw
tri 16360 -23245 16707 -22898 se
rect 16707 -23245 19709 -22898
rect -23607 -23780 -20606 -23245
rect -27143 -24489 -24316 -23780
tri -24316 -24489 -23607 -23780 sw
tri -23607 -24489 -22898 -23780 ne
rect -22898 -23955 -20606 -23780
tri -20606 -23955 -19896 -23245 sw
tri -19896 -23432 -19709 -23245 ne
rect -19709 -23432 -16360 -23245
tri -16360 -23432 -16173 -23245 sw
tri -15651 -23432 -15464 -23245 ne
rect -15464 -23432 -12115 -23245
tri -12115 -23432 -11928 -23245 sw
tri -11405 -23432 -11218 -23245 ne
rect -11218 -23432 11218 -23245
tri 11218 -23432 11405 -23245 nw
tri 11928 -23432 12115 -23245 se
rect 12115 -23432 15464 -23245
tri 15464 -23432 15651 -23245 nw
tri 16173 -23432 16360 -23245 se
rect 16360 -23432 19709 -23245
tri 19709 -23432 20243 -22898 nw
tri 20419 -23432 20953 -22898 se
rect 20953 -23432 23780 -22898
tri -19709 -23955 -19186 -23432 ne
rect -19186 -23780 -16173 -23432
tri -16173 -23780 -15825 -23432 sw
tri -15464 -23780 -15116 -23432 ne
rect -15116 -23780 -11928 -23432
rect -19186 -23955 -15825 -23780
rect -22898 -24489 -19896 -23955
tri -19896 -24489 -19362 -23955 sw
tri -19186 -24489 -18652 -23955 ne
rect -18652 -24489 -15825 -23955
tri -15825 -24489 -15116 -23780 sw
tri -15116 -23966 -14930 -23780 ne
rect -14930 -23966 -11928 -23780
tri -11928 -23966 -11394 -23432 sw
tri -11218 -23966 -10684 -23432 ne
rect -10684 -23966 10684 -23432
tri 10684 -23966 11218 -23432 nw
tri 11394 -23966 11928 -23432 se
rect 11928 -23966 14930 -23432
tri 14930 -23966 15464 -23432 nw
tri 15639 -23966 16173 -23432 se
rect 16173 -23966 18999 -23432
tri -14930 -24489 -14407 -23966 ne
rect -14407 -24294 -11394 -23966
tri -11394 -24294 -11066 -23966 sw
tri -10684 -24294 -10356 -23966 ne
rect -10356 -24294 10161 -23966
rect -14407 -24489 -11066 -24294
tri -11066 -24489 -10871 -24294 sw
tri -10356 -24489 -10161 -24294 ne
rect -10161 -24489 10161 -24294
tri 10161 -24489 10684 -23966 nw
tri 10871 -24489 11394 -23966 se
rect 11394 -24489 14407 -23966
tri 14407 -24489 14930 -23966 nw
tri 15116 -24489 15639 -23966 se
rect 15639 -24142 18999 -23966
tri 18999 -24142 19709 -23432 nw
tri 19709 -24142 20419 -23432 se
rect 20419 -23607 23780 -23432
tri 23780 -23607 24489 -22898 nw
tri 24489 -23607 25198 -22898 se
rect 25198 -23607 25732 -22898
rect 20419 -24142 23071 -23607
rect 15639 -24489 18652 -24142
tri 18652 -24489 18999 -24142 nw
tri 19362 -24489 19709 -24142 se
rect 19709 -24316 23071 -24142
tri 23071 -24316 23780 -23607 nw
tri 23780 -24316 24489 -23607 se
rect 24489 -24316 25732 -23607
rect 19709 -24482 22905 -24316
tri 22905 -24482 23071 -24316 nw
tri 23614 -24482 23780 -24316 se
rect 23780 -24482 25732 -24316
rect 19709 -24489 22196 -24482
tri -27143 -25324 -26308 -24489 ne
rect -26308 -25198 -23607 -24489
tri -23607 -25198 -22898 -24489 sw
tri -22898 -25198 -22189 -24489 ne
rect -22189 -25022 -19362 -24489
tri -19362 -25022 -18829 -24489 sw
tri -18652 -25022 -18119 -24489 ne
rect -18119 -25002 -15116 -24489
tri -15116 -25002 -14603 -24489 sw
tri -14407 -25002 -13894 -24489 ne
rect -13894 -25002 -10871 -24489
tri -10871 -25002 -10358 -24489 sw
tri -10161 -24500 -10150 -24489 ne
rect -10150 -24500 10150 -24489
tri 10150 -24500 10161 -24489 nw
tri 10860 -24500 10871 -24489 se
rect 10871 -24500 14221 -24489
tri 10358 -25002 10860 -24500 se
rect 10860 -24675 14221 -24500
tri 14221 -24675 14407 -24489 nw
tri 14930 -24675 15116 -24489 se
rect 15116 -24675 18289 -24489
rect 10860 -25002 13894 -24675
tri 13894 -25002 14221 -24675 nw
tri 14603 -25002 14930 -24675 se
rect 14930 -24852 18289 -24675
tri 18289 -24852 18652 -24489 nw
tri 18999 -24852 19362 -24489 se
rect 19362 -24852 22196 -24489
rect 14930 -25002 18139 -24852
tri 18139 -25002 18289 -24852 nw
tri 18849 -25002 18999 -24852 se
rect 18999 -25002 22196 -24852
rect -18119 -25022 -14603 -25002
rect -22189 -25198 -18829 -25022
rect -26308 -25324 -22898 -25198
tri -22898 -25324 -22772 -25198 sw
tri -22189 -25324 -22063 -25198 ne
rect -22063 -25324 -18829 -25198
tri -18829 -25324 -18527 -25022 sw
tri -18119 -25324 -17817 -25022 ne
rect -17817 -25324 -14603 -25022
tri -14603 -25324 -14281 -25002 sw
tri -13894 -25324 -13572 -25002 ne
rect -13572 -25324 -979 -25002
tri -979 -25324 -657 -25002 sw
tri 2291 -25222 2511 -25002 se
rect 2511 -25023 13873 -25002
tri 13873 -25023 13894 -25002 nw
tri 14582 -25023 14603 -25002 se
rect 14603 -25022 18119 -25002
tri 18119 -25022 18139 -25002 nw
tri 18829 -25022 18849 -25002 se
rect 18849 -25022 22196 -25002
rect 14603 -25023 17409 -25022
rect 2511 -25222 13164 -25023
rect 2291 -25324 13164 -25222
tri -26308 -25580 -26052 -25324 ne
rect -26052 -25580 -22772 -25324
tri -22772 -25580 -22516 -25324 sw
tri -22063 -25580 -21807 -25324 ne
rect -21807 -25580 -18527 -25324
tri -18527 -25580 -18271 -25324 sw
tri -17817 -25580 -17561 -25324 ne
rect -17561 -25538 -14281 -25324
tri -14281 -25538 -14067 -25324 sw
tri -13572 -25538 -13358 -25324 ne
rect -13358 -25538 -657 -25324
rect -17561 -25580 -14067 -25538
tri -14067 -25580 -14025 -25538 sw
tri -13358 -25580 -13316 -25538 ne
rect -13316 -25580 -657 -25538
tri -657 -25580 -401 -25324 sw
rect 2291 -25580 2393 -25324
rect 2649 -25580 2917 -25324
rect 3173 -25580 3471 -25324
rect 3727 -25580 4025 -25324
rect 4281 -25580 4549 -25324
rect 4805 -25580 5163 -25324
rect 5419 -25580 5687 -25324
rect 5943 -25580 6241 -25324
rect 6497 -25580 6795 -25324
rect 7051 -25580 7319 -25324
rect 7575 -25580 13164 -25324
tri -26052 -25732 -25900 -25580 ne
rect -25900 -25732 -22516 -25580
tri -22516 -25732 -22364 -25580 sw
tri -21807 -25732 -21655 -25580 ne
rect -21655 -25732 -18271 -25580
tri -18271 -25732 -18119 -25580 sw
tri -17561 -25732 -17409 -25580 ne
rect -17409 -25732 -14025 -25580
tri -25900 -25818 -25814 -25732 ne
rect -25814 -25818 -22364 -25732
tri -22364 -25818 -22278 -25732 sw
tri -21655 -25818 -21569 -25732 ne
rect -21569 -25818 -18119 -25732
tri -18119 -25818 -18033 -25732 sw
tri -17409 -25818 -17323 -25732 ne
rect -17323 -25818 -14025 -25732
tri -14025 -25818 -13787 -25580 sw
tri -13316 -25818 -13078 -25580 ne
rect -13078 -25732 -401 -25580
tri -401 -25732 -249 -25580 sw
rect 2291 -25732 13164 -25580
tri 13164 -25732 13873 -25023 nw
tri 13873 -25732 14582 -25023 se
rect 14582 -25732 17409 -25023
tri 17409 -25732 18119 -25022 nw
tri 18119 -25732 18829 -25022 se
rect 18829 -25191 22196 -25022
tri 22196 -25191 22905 -24482 nw
tri 22905 -25191 23614 -24482 se
rect 23614 -25191 25732 -24482
rect 18829 -25732 21655 -25191
tri 21655 -25732 22196 -25191 nw
tri 22364 -25732 22905 -25191 se
rect 22905 -25732 25732 -25191
rect -13078 -25818 -249 -25732
tri -249 -25818 -163 -25732 sw
rect 2291 -25818 12996 -25732
tri -25814 -25900 -25732 -25818 ne
rect -25732 -25900 -22278 -25818
tri -22278 -25900 -22196 -25818 sw
tri -21569 -25900 -21487 -25818 ne
rect -21487 -25900 -18033 -25818
tri -18033 -25900 -17951 -25818 sw
tri -17323 -25900 -17241 -25818 ne
rect -17241 -25900 -13787 -25818
tri -25732 -26074 -25558 -25900 ne
rect -25558 -26074 -22196 -25900
tri -22196 -26074 -22022 -25900 sw
tri -21487 -26074 -21313 -25900 ne
rect -21313 -26074 -17951 -25900
tri -17951 -26074 -17777 -25900 sw
tri -17241 -26074 -17067 -25900 ne
rect -17067 -26074 -13787 -25900
tri -13787 -26074 -13531 -25818 sw
tri -13078 -26074 -12822 -25818 ne
rect -12822 -25900 -163 -25818
tri -163 -25900 -81 -25818 sw
rect -12822 -26074 -81 -25900
tri -81 -26074 93 -25900 sw
rect 2291 -26074 2393 -25818
rect 2649 -26074 2917 -25818
rect 3173 -26074 3471 -25818
rect 3727 -26074 4025 -25818
rect 4281 -26074 4549 -25818
rect 4805 -26074 5163 -25818
rect 5419 -26074 5687 -25818
rect 5943 -26074 6241 -25818
rect 6497 -26074 6795 -25818
rect 7051 -26074 7319 -25818
rect 7575 -25900 12996 -25818
tri 12996 -25900 13164 -25732 nw
tri 13705 -25900 13873 -25732 se
rect 13873 -25900 17241 -25732
tri 17241 -25900 17409 -25732 nw
tri 17951 -25900 18119 -25732 se
rect 18119 -25900 21487 -25732
tri 21487 -25900 21655 -25732 nw
tri 22196 -25900 22364 -25732 se
rect 22364 -25900 25732 -25732
tri 25732 -25900 28734 -22898 nw
rect 7575 -26074 12462 -25900
tri -25558 -26432 -25200 -26074 ne
rect -25200 -26432 -22022 -26074
tri -22022 -26432 -21664 -26074 sw
tri -21313 -26432 -20955 -26074 ne
rect -20955 -26432 -17777 -26074
tri -17777 -26432 -17419 -26074 sw
tri -17067 -26432 -16709 -26074 ne
rect -16709 -26247 -13531 -26074
tri -13531 -26247 -13358 -26074 sw
tri -12822 -26247 -12649 -26074 ne
rect -12649 -26247 93 -26074
rect -16709 -26432 -13358 -26247
tri -13358 -26432 -13173 -26247 sw
tri -12649 -26432 -12464 -26247 ne
rect -12464 -26432 93 -26247
tri 93 -26432 451 -26074 sw
rect 2291 -26432 12462 -26074
tri -25200 -26688 -24944 -26432 ne
rect -24944 -26609 -21664 -26432
tri -21664 -26609 -21487 -26432 sw
tri -20955 -26609 -20778 -26432 ne
rect -20778 -26434 -17419 -26432
tri -17419 -26434 -17417 -26432 sw
tri -16709 -26434 -16707 -26432 ne
rect -16707 -26434 -13173 -26432
rect -20778 -26609 -17417 -26434
rect -24944 -26688 -21487 -26609
tri -21487 -26688 -21408 -26609 sw
tri -20778 -26688 -20699 -26609 ne
rect -20699 -26688 -17417 -26609
tri -17417 -26688 -17163 -26434 sw
tri -16707 -26688 -16453 -26434 ne
rect -16453 -26688 -13173 -26434
tri -13173 -26688 -12917 -26432 sw
tri -12464 -26688 -12208 -26432 ne
rect -12208 -26434 451 -26432
tri 451 -26434 453 -26432 sw
rect -12208 -26688 453 -26434
tri 453 -26688 707 -26434 sw
rect 2291 -26688 2393 -26432
rect 2649 -26688 2917 -26432
rect 3173 -26688 3471 -26432
rect 3727 -26688 4025 -26432
rect 4281 -26688 4549 -26432
rect 4805 -26688 5163 -26432
rect 5419 -26688 5687 -26432
rect 5943 -26688 6241 -26432
rect 6497 -26688 6795 -26432
rect 7051 -26688 7319 -26432
rect 7575 -26434 12462 -26432
tri 12462 -26434 12996 -25900 nw
tri 13171 -26434 13705 -25900 se
rect 13705 -26434 16707 -25900
tri 16707 -26434 17241 -25900 nw
tri 17417 -26434 17951 -25900 se
rect 17951 -26434 20953 -25900
tri 20953 -26434 21487 -25900 nw
tri 21662 -26434 22196 -25900 se
rect 22196 -26434 25198 -25900
tri 25198 -26434 25732 -25900 nw
rect 7575 -26688 11928 -26434
tri -24944 -26926 -24706 -26688 ne
rect -24706 -26926 -21408 -26688
tri -21408 -26926 -21170 -26688 sw
tri -20699 -26926 -20461 -26688 ne
rect -20461 -26781 -17163 -26688
tri -17163 -26781 -17070 -26688 sw
tri -16453 -26781 -16360 -26688 ne
rect -16360 -26781 -12917 -26688
tri -12917 -26781 -12824 -26688 sw
tri -12208 -26781 -12115 -26688 ne
rect -12115 -26781 707 -26688
rect -20461 -26926 -17070 -26781
tri -17070 -26926 -16925 -26781 sw
tri -16360 -26926 -16215 -26781 ne
rect -16215 -26793 -12824 -26781
tri -12824 -26793 -12812 -26781 sw
tri -12115 -26793 -12103 -26781 ne
rect -12103 -26793 707 -26781
rect -16215 -26926 -12812 -26793
tri -12812 -26926 -12679 -26793 sw
tri -12103 -26926 -11970 -26793 ne
rect -11970 -26926 707 -26793
tri 707 -26926 945 -26688 sw
rect 2291 -26926 11928 -26688
tri -24706 -27182 -24450 -26926 ne
rect -24450 -27182 -21170 -26926
tri -21170 -27182 -20914 -26926 sw
tri -20461 -27182 -20205 -26926 ne
rect -20205 -27182 -16925 -26926
tri -16925 -27182 -16669 -26926 sw
tri -16215 -27182 -15959 -26926 ne
rect -15959 -27182 -12679 -26926
tri -12679 -27182 -12423 -26926 sw
tri -11970 -27182 -11714 -26926 ne
rect -11714 -27182 945 -26926
tri 945 -27182 1201 -26926 sw
rect 2291 -27182 2393 -26926
rect 2649 -27182 2917 -26926
rect 3173 -27182 3471 -26926
rect 3727 -27182 4025 -26926
rect 4281 -27182 4549 -26926
rect 4805 -27182 5163 -26926
rect 5419 -27182 5687 -26926
rect 5943 -27182 6241 -26926
rect 6497 -27182 6795 -26926
rect 7051 -27182 7319 -26926
rect 7575 -26968 11928 -26926
tri 11928 -26968 12462 -26434 nw
tri 12637 -26968 13171 -26434 se
rect 13171 -26968 16173 -26434
tri 16173 -26968 16707 -26434 nw
tri 16883 -26968 17417 -26434 se
rect 17417 -26968 20244 -26434
rect 7575 -27182 11394 -26968
tri -24450 -28025 -23607 -27182 ne
rect -23607 -27316 -20914 -27182
tri -20914 -27316 -20780 -27182 sw
tri -20205 -27316 -20071 -27182 ne
rect -20071 -27316 -16669 -27182
rect -23607 -28025 -20780 -27316
tri -20780 -28025 -20071 -27316 sw
tri -20071 -28025 -19362 -27316 ne
rect -19362 -27491 -16669 -27316
tri -16669 -27491 -16360 -27182 sw
tri -15959 -27491 -15650 -27182 ne
rect -15650 -27491 -12423 -27182
rect -19362 -28025 -16360 -27491
tri -16360 -28025 -15826 -27491 sw
tri -15650 -27502 -15639 -27491 ne
rect -15639 -27502 -12423 -27491
tri -12423 -27502 -12103 -27182 sw
tri -11714 -27502 -11394 -27182 ne
rect -11394 -27502 1201 -27182
tri 1201 -27502 1521 -27182 sw
rect 2291 -27282 11394 -27182
tri 2291 -27502 2511 -27282 ne
rect 2511 -27502 11394 -27282
tri 11394 -27502 11928 -26968 nw
tri 12103 -27502 12637 -26968 se
rect 12637 -27502 15639 -26968
tri 15639 -27502 16173 -26968 nw
tri 16349 -27502 16883 -26968 se
rect 16883 -27143 20244 -26968
tri 20244 -27143 20953 -26434 nw
tri 20953 -27143 21662 -26434 se
rect 21662 -27143 22196 -26434
rect 16883 -27502 19535 -27143
tri -15639 -28025 -15116 -27502 ne
rect -15116 -28004 -12103 -27502
tri -12103 -28004 -11601 -27502 sw
tri -2015 -28004 -1513 -27502 ne
rect -1513 -28004 1521 -27502
tri 1521 -28004 2023 -27502 sw
tri 11601 -28004 12103 -27502 se
rect 12103 -27678 15463 -27502
tri 15463 -27678 15639 -27502 nw
tri 16173 -27678 16349 -27502 se
rect 16349 -27678 19535 -27502
rect 12103 -28004 15137 -27678
tri 15137 -28004 15463 -27678 nw
tri 15847 -28004 16173 -27678 se
rect 16173 -27852 19535 -27678
tri 19535 -27852 20244 -27143 nw
tri 20244 -27852 20953 -27143 se
rect 20953 -27852 22196 -27143
rect 16173 -28004 19369 -27852
rect -15116 -28025 -2380 -28004
tri -2380 -28025 -2359 -28004 sw
tri -1513 -28025 -1492 -28004 ne
rect -1492 -28025 14753 -28004
tri -23607 -28325 -23307 -28025 ne
rect -23307 -28325 -20071 -28025
tri -20071 -28325 -19771 -28025 sw
tri -19362 -28325 -19062 -28025 ne
rect -19062 -28325 -15826 -28025
tri -15826 -28325 -15526 -28025 sw
tri -15116 -28325 -14816 -28025 ne
rect -14816 -28224 -2359 -28025
tri -2359 -28224 -2160 -28025 sw
rect -14816 -28325 -2160 -28224
tri -23307 -28581 -23051 -28325 ne
rect -23051 -28581 -19771 -28325
tri -19771 -28581 -19515 -28325 sw
tri -19062 -28581 -18806 -28325 ne
rect -18806 -28558 -15526 -28325
tri -15526 -28558 -15293 -28325 sw
tri -14816 -28558 -14583 -28325 ne
rect -14583 -28558 -7444 -28325
rect -18806 -28581 -15293 -28558
tri -15293 -28581 -15270 -28558 sw
tri -14583 -28581 -14560 -28558 ne
rect -14560 -28581 -7444 -28558
rect -7188 -28581 -6920 -28325
rect -6664 -28581 -6366 -28325
rect -6110 -28581 -5812 -28325
rect -5556 -28581 -5288 -28325
rect -5032 -28581 -4674 -28325
rect -4418 -28581 -4150 -28325
rect -3894 -28581 -3596 -28325
rect -3340 -28581 -3042 -28325
rect -2786 -28581 -2518 -28325
rect -2262 -28581 -2160 -28325
tri -23051 -28819 -22813 -28581 ne
rect -22813 -28734 -19515 -28581
tri -19515 -28734 -19362 -28581 sw
tri -18806 -28734 -18653 -28581 ne
rect -18653 -28734 -15270 -28581
rect -22813 -28819 -19362 -28734
tri -19362 -28819 -19277 -28734 sw
tri -18653 -28819 -18568 -28734 ne
rect -18568 -28819 -15270 -28734
tri -15270 -28819 -15032 -28581 sw
tri -14560 -28819 -14322 -28581 ne
rect -14322 -28819 -2160 -28581
tri -22813 -29075 -22557 -28819 ne
rect -22557 -29075 -19277 -28819
tri -19277 -29075 -19021 -28819 sw
tri -18568 -29075 -18312 -28819 ne
rect -18312 -29075 -15032 -28819
tri -15032 -29075 -14776 -28819 sw
tri -14322 -29075 -14066 -28819 ne
rect -14066 -29075 -7444 -28819
rect -7188 -29075 -6920 -28819
rect -6664 -29075 -6366 -28819
rect -6110 -29075 -5812 -28819
rect -5556 -29075 -5288 -28819
rect -5032 -29075 -4674 -28819
rect -4418 -29075 -4150 -28819
rect -3894 -29075 -3596 -28819
rect -3340 -29075 -3042 -28819
rect -2786 -29075 -2518 -28819
rect -2262 -29075 -2160 -28819
tri -22557 -29268 -22364 -29075 ne
rect -22364 -29268 -19021 -29075
tri -19021 -29268 -18828 -29075 sw
tri -18312 -29268 -18119 -29075 ne
rect -18119 -29268 -14776 -29075
tri -14776 -29268 -14583 -29075 sw
tri -14066 -29268 -13873 -29075 ne
rect -13873 -29268 -2160 -29075
tri -1492 -29268 -249 -28025 ne
rect -249 -28388 14753 -28025
tri 14753 -28388 15137 -28004 nw
tri 15463 -28388 15847 -28004 se
rect 15847 -28018 19369 -28004
tri 19369 -28018 19535 -27852 nw
tri 20078 -28018 20244 -27852 se
rect 20244 -28018 22196 -27852
rect 15847 -28388 18660 -28018
rect -249 -28558 14583 -28388
tri 14583 -28558 14753 -28388 nw
tri 15293 -28558 15463 -28388 se
rect 15463 -28558 18660 -28388
rect -249 -29268 13873 -28558
tri 13873 -29268 14583 -28558 nw
tri 14583 -29268 15293 -28558 se
rect 15293 -28727 18660 -28558
tri 18660 -28727 19369 -28018 nw
tri 19369 -28727 20078 -28018 se
rect 20078 -28727 22196 -28018
rect 15293 -29268 18119 -28727
tri 18119 -29268 18660 -28727 nw
tri 18828 -29268 19369 -28727 se
rect 19369 -29268 22196 -28727
tri -22364 -29433 -22199 -29268 ne
rect -22199 -29433 -18828 -29268
tri -18828 -29433 -18663 -29268 sw
tri -18119 -29433 -17954 -29268 ne
rect -17954 -29433 -14583 -29268
tri -14583 -29433 -14418 -29268 sw
tri -13873 -29433 -13708 -29268 ne
rect -13708 -29433 -2160 -29268
tri -22199 -29436 -22196 -29433 ne
rect -22196 -29436 -18663 -29433
tri -18663 -29436 -18660 -29433 sw
tri -17954 -29436 -17951 -29433 ne
rect -17951 -29436 -14418 -29433
tri -14418 -29436 -14415 -29433 sw
tri -13708 -29436 -13705 -29433 ne
rect -13705 -29436 -7444 -29433
tri -22196 -29689 -21943 -29436 ne
rect -21943 -29689 -18660 -29436
tri -18660 -29689 -18407 -29436 sw
tri -17951 -29689 -17698 -29436 ne
rect -17698 -29689 -14415 -29436
tri -14415 -29689 -14162 -29436 sw
tri -13705 -29689 -13452 -29436 ne
rect -13452 -29689 -7444 -29436
rect -7188 -29689 -6920 -29433
rect -6664 -29689 -6366 -29433
rect -6110 -29689 -5812 -29433
rect -5556 -29689 -5288 -29433
rect -5032 -29689 -4674 -29433
rect -4418 -29689 -4150 -29433
rect -3894 -29689 -3596 -29433
rect -3340 -29689 -3042 -29433
rect -2786 -29689 -2518 -29433
rect -2262 -29689 -2160 -29433
tri -249 -29436 -81 -29268 ne
rect -81 -29436 13705 -29268
tri 13705 -29436 13873 -29268 nw
tri 14415 -29436 14583 -29268 se
rect 14583 -29436 17951 -29268
tri 17951 -29436 18119 -29268 nw
tri 18660 -29436 18828 -29268 se
rect 18828 -29436 22196 -29268
tri 22196 -29436 25198 -26434 nw
tri -21943 -29927 -21705 -29689 ne
rect -21705 -29927 -18407 -29689
tri -18407 -29927 -18169 -29689 sw
tri -17698 -29927 -17460 -29689 ne
rect -17460 -29927 -14162 -29689
tri -14162 -29927 -13924 -29689 sw
tri -13452 -29927 -13214 -29689 ne
rect -13214 -29927 -2160 -29689
tri -21705 -30183 -21449 -29927 ne
rect -21449 -30145 -18169 -29927
tri -18169 -30145 -17951 -29927 sw
tri -17460 -30145 -17242 -29927 ne
rect -17242 -29970 -13924 -29927
tri -13924 -29970 -13881 -29927 sw
tri -13214 -29970 -13171 -29927 ne
rect -13171 -29970 -7444 -29927
rect -17242 -30145 -13881 -29970
rect -21449 -30183 -17951 -30145
tri -17951 -30183 -17913 -30145 sw
tri -17242 -30183 -17204 -30145 ne
rect -17204 -30183 -13881 -30145
tri -13881 -30183 -13668 -29970 sw
tri -13171 -30183 -12958 -29970 ne
rect -12958 -30183 -7444 -29970
rect -7188 -30183 -6920 -29927
rect -6664 -30183 -6366 -29927
rect -6110 -30183 -5812 -29927
rect -5556 -30183 -5288 -29927
rect -5032 -30183 -4674 -29927
rect -4418 -30183 -4150 -29927
rect -3894 -30183 -3596 -29927
rect -3340 -30183 -3042 -29927
rect -2786 -30183 -2518 -29927
rect -2262 -30183 -2160 -29927
tri -81 -29970 453 -29436 ne
rect 453 -29970 13171 -29436
tri 13171 -29970 13705 -29436 nw
tri 13881 -29970 14415 -29436 se
rect 14415 -29970 17417 -29436
tri 17417 -29970 17951 -29436 nw
tri 18126 -29970 18660 -29436 se
rect 18660 -29970 21662 -29436
tri 21662 -29970 22196 -29436 nw
tri -21449 -31326 -20306 -30183 ne
rect -20306 -30852 -17913 -30183
tri -17913 -30852 -17244 -30183 sw
tri -17204 -30852 -16535 -30183 ne
rect -16535 -30317 -13668 -30183
tri -13668 -30317 -13534 -30183 sw
tri -12958 -30317 -12824 -30183 ne
rect -12824 -30284 -2160 -30183
rect -12824 -30317 -2193 -30284
tri -2193 -30317 -2160 -30284 nw
tri 453 -30317 800 -29970 ne
rect 800 -30317 12637 -29970
rect -16535 -30852 -13534 -30317
rect -20306 -31326 -17244 -30852
tri -17244 -31326 -16770 -30852 sw
tri -16535 -31326 -16061 -30852 ne
rect -16061 -31006 -13534 -30852
tri -13534 -31006 -12845 -30317 sw
tri -12824 -30504 -12637 -30317 ne
rect -12637 -30504 -2380 -30317
tri -2380 -30504 -2193 -30317 nw
tri 800 -30504 987 -30317 ne
rect 987 -30504 12637 -30317
tri 12637 -30504 13171 -29970 nw
tri 13347 -30504 13881 -29970 se
rect 13881 -30504 16708 -29970
tri 12845 -31006 13347 -30504 se
rect 13347 -30679 16708 -30504
tri 16708 -30679 17417 -29970 nw
tri 17417 -30679 18126 -29970 se
rect 18126 -30679 18660 -29970
rect 13347 -31006 15999 -30679
rect -16061 -31326 -979 -31006
tri -979 -31326 -659 -31006 sw
tri 2291 -31226 2511 -31006 se
rect 2511 -31226 15999 -31006
rect 2291 -31326 15999 -31226
tri -20306 -31561 -20071 -31326 ne
rect -20071 -31561 -16770 -31326
tri -16770 -31561 -16535 -31326 sw
tri -16061 -31561 -15826 -31326 ne
rect -15826 -31561 -659 -31326
tri -659 -31561 -424 -31326 sw
tri -20071 -31582 -20050 -31561 ne
rect -20050 -31582 -16535 -31561
tri -16535 -31582 -16514 -31561 sw
tri -15826 -31582 -15805 -31561 ne
rect -15805 -31582 -424 -31561
tri -424 -31582 -403 -31561 sw
rect 2291 -31582 2393 -31326
rect 2649 -31582 2917 -31326
rect 3173 -31582 3471 -31326
rect 3727 -31582 4025 -31326
rect 4281 -31582 4549 -31326
rect 4805 -31582 5163 -31326
rect 5419 -31582 5687 -31326
rect 5943 -31582 6241 -31326
rect 6497 -31582 6795 -31326
rect 7051 -31582 7319 -31326
rect 7575 -31388 15999 -31326
tri 15999 -31388 16708 -30679 nw
tri 16708 -31388 17417 -30679 se
rect 17417 -31388 18660 -30679
rect 7575 -31554 15833 -31388
tri 15833 -31554 15999 -31388 nw
tri 16542 -31554 16708 -31388 se
rect 16708 -31554 18660 -31388
rect 7575 -31582 15124 -31554
tri -20050 -31820 -19812 -31582 ne
rect -19812 -31820 -16514 -31582
tri -16514 -31820 -16276 -31582 sw
tri -15805 -31820 -15567 -31582 ne
rect -15567 -31820 -403 -31582
tri -403 -31820 -165 -31582 sw
rect 2291 -31820 15124 -31582
tri -19812 -32076 -19556 -31820 ne
rect -19556 -32076 -16276 -31820
tri -16276 -32076 -16020 -31820 sw
tri -15567 -32076 -15311 -31820 ne
rect -15311 -32076 -165 -31820
tri -165 -32076 91 -31820 sw
rect 2291 -32076 2393 -31820
rect 2649 -32076 2917 -31820
rect 3173 -32076 3471 -31820
rect 3727 -32076 4025 -31820
rect 4281 -32076 4549 -31820
rect 4805 -32076 5163 -31820
rect 5419 -32076 5687 -31820
rect 5943 -32076 6241 -31820
rect 6497 -32076 6795 -31820
rect 7051 -32076 7319 -31820
rect 7575 -32076 15124 -31820
tri -19556 -32434 -19198 -32076 ne
rect -19198 -32270 -16020 -32076
tri -16020 -32270 -15826 -32076 sw
tri -15311 -32270 -15117 -32076 ne
rect -15117 -32270 91 -32076
rect -19198 -32434 -15826 -32270
tri -15826 -32434 -15662 -32270 sw
tri -15117 -32434 -14953 -32270 ne
rect -14953 -32434 91 -32270
tri 91 -32434 449 -32076 sw
rect 2291 -32263 15124 -32076
tri 15124 -32263 15833 -31554 nw
tri 15833 -32263 16542 -31554 se
rect 16542 -32263 18660 -31554
rect 2291 -32434 14583 -32263
tri -19198 -32690 -18942 -32434 ne
rect -18942 -32690 -15662 -32434
tri -15662 -32690 -15406 -32434 sw
tri -14953 -32690 -14697 -32434 ne
rect -14697 -32690 449 -32434
tri 449 -32690 705 -32434 sw
rect 2291 -32690 2393 -32434
rect 2649 -32690 2917 -32434
rect 3173 -32690 3471 -32434
rect 3727 -32690 4025 -32434
rect 4281 -32690 4549 -32434
rect 4805 -32690 5163 -32434
rect 5419 -32690 5687 -32434
rect 5943 -32690 6241 -32434
rect 6497 -32690 6795 -32434
rect 7051 -32690 7319 -32434
rect 7575 -32690 14583 -32434
tri -18942 -32804 -18828 -32690 ne
rect -18828 -32804 -15406 -32690
tri -15406 -32804 -15292 -32690 sw
tri -14697 -32804 -14583 -32690 ne
rect -14583 -32804 705 -32690
tri 705 -32804 819 -32690 sw
rect 2291 -32804 14583 -32690
tri 14583 -32804 15124 -32263 nw
tri 15292 -32804 15833 -32263 se
rect 15833 -32804 18660 -32263
tri -18828 -32928 -18704 -32804 ne
rect -18704 -32928 -15292 -32804
tri -15292 -32928 -15168 -32804 sw
tri -14583 -32928 -14459 -32804 ne
rect -14459 -32928 819 -32804
tri 819 -32928 943 -32804 sw
rect 2291 -32928 14415 -32804
tri -18704 -32972 -18660 -32928 ne
rect -18660 -32972 -15168 -32928
tri -15168 -32972 -15124 -32928 sw
tri -14459 -32972 -14415 -32928 ne
rect -14415 -32972 943 -32928
tri 943 -32972 987 -32928 sw
tri -18660 -33184 -18448 -32972 ne
rect -18448 -33184 -15124 -32972
tri -15124 -33184 -14912 -32972 sw
tri -14415 -33184 -14203 -32972 ne
rect -14203 -33184 987 -32972
tri 987 -33184 1199 -32972 sw
rect 2291 -33184 2393 -32928
rect 2649 -33184 2917 -32928
rect 3173 -33184 3471 -32928
rect 3727 -33184 4025 -32928
rect 4281 -33184 4549 -32928
rect 4805 -33184 5163 -32928
rect 5419 -33184 5687 -32928
rect 5943 -33184 6241 -32928
rect 6497 -33184 6795 -32928
rect 7051 -33184 7319 -32928
rect 7575 -32972 14415 -32928
tri 14415 -32972 14583 -32804 nw
tri 15124 -32972 15292 -32804 se
rect 15292 -32972 18660 -32804
tri 18660 -32972 21662 -29970 nw
rect 7575 -33184 13881 -32972
tri -18448 -33506 -18126 -33184 ne
rect -18126 -33506 -14912 -33184
tri -14912 -33506 -14590 -33184 sw
tri -14203 -33506 -13881 -33184 ne
rect -13881 -33506 1199 -33184
tri 1199 -33506 1521 -33184 sw
rect 2291 -33286 13881 -33184
tri 2291 -33506 2511 -33286 ne
rect 2511 -33506 13881 -33286
tri 13881 -33506 14415 -32972 nw
tri 14590 -33506 15124 -32972 se
rect 15124 -33506 18126 -32972
tri 18126 -33506 18660 -32972 nw
tri -18126 -34329 -17303 -33506 ne
rect -17303 -34008 -14590 -33506
tri -14590 -34008 -14088 -33506 sw
tri -2015 -34008 -1513 -33506 ne
rect -1513 -34008 1521 -33506
tri 1521 -34008 2023 -33506 sw
tri 14088 -34008 14590 -33506 se
rect 14590 -34008 15124 -33506
rect -17303 -34228 -2380 -34008
tri -2380 -34228 -2160 -34008 sw
rect -17303 -34329 -2160 -34228
tri -17303 -34585 -17047 -34329 ne
rect -17047 -34585 -7444 -34329
rect -7188 -34585 -6920 -34329
rect -6664 -34585 -6366 -34329
rect -6110 -34585 -5812 -34329
rect -5556 -34585 -5288 -34329
rect -5032 -34585 -4674 -34329
rect -4418 -34585 -4150 -34329
rect -3894 -34585 -3596 -34329
rect -3340 -34585 -3042 -34329
rect -2786 -34585 -2518 -34329
rect -2262 -34585 -2160 -34329
tri -17047 -34823 -16809 -34585 ne
rect -16809 -34823 -2160 -34585
tri -16809 -35079 -16553 -34823 ne
rect -16553 -35079 -7444 -34823
rect -7188 -35079 -6920 -34823
rect -6664 -35079 -6366 -34823
rect -6110 -35079 -5812 -34823
rect -5556 -35079 -5288 -34823
rect -5032 -35079 -4674 -34823
rect -4418 -35079 -4150 -34823
rect -3894 -35079 -3596 -34823
rect -3340 -35079 -3042 -34823
rect -2786 -35079 -2518 -34823
rect -2262 -35079 -2160 -34823
tri -16553 -35437 -16195 -35079 ne
rect -16195 -35437 -2160 -35079
tri -16195 -35693 -15939 -35437 ne
rect -15939 -35693 -7444 -35437
rect -7188 -35693 -6920 -35437
rect -6664 -35693 -6366 -35437
rect -6110 -35693 -5812 -35437
rect -5556 -35693 -5288 -35437
rect -5032 -35693 -4674 -35437
rect -4418 -35693 -4150 -35437
rect -3894 -35693 -3596 -35437
rect -3340 -35693 -3042 -35437
rect -2786 -35693 -2518 -35437
rect -2262 -35693 -2160 -35437
tri -15939 -35931 -15701 -35693 ne
rect -15701 -35931 -2160 -35693
tri -15701 -36187 -15445 -35931 ne
rect -15445 -36187 -7444 -35931
rect -7188 -36187 -6920 -35931
rect -6664 -36187 -6366 -35931
rect -6110 -36187 -5812 -35931
rect -5556 -36187 -5288 -35931
rect -5032 -36187 -4674 -35931
rect -4418 -36187 -4150 -35931
rect -3894 -36187 -3596 -35931
rect -3340 -36187 -3042 -35931
rect -2786 -36187 -2518 -35931
rect -2262 -36187 -2160 -35931
tri -15445 -36340 -15292 -36187 ne
rect -15292 -36288 -2160 -36187
rect -15292 -36340 -2212 -36288
tri -2212 -36340 -2160 -36288 nw
tri -1513 -36340 819 -34008 ne
rect 819 -36340 15124 -34008
tri -15292 -36508 -15124 -36340 ne
rect -15124 -36508 -2380 -36340
tri -2380 -36508 -2212 -36340 nw
tri 819 -36508 987 -36340 ne
rect 987 -36508 15124 -36340
tri 15124 -36508 18126 -33506 nw
<< comment >>
tri -15125 15125 -6266 36508 ne
rect -6266 15125 6266 36508
tri 6266 15125 15125 36508 nw
tri -36508 2596 -6266 15125 sw
tri -6266 2596 -1075 15125 ne
rect -1075 2596 1075 15125
tri 1075 2596 6266 15125 nw
tri 6266 2596 36508 15125 se
rect -36508 445 -6266 2596
tri -6266 445 -1075 2596 sw
tri -1075 445 -185 2596 ne
rect -185 446 185 2596
tri 185 446 1075 2596 nw
tri 1076 446 6266 2596 se
rect 6266 446 36508 2596
rect -185 445 32 446
rect -36508 76 -1075 445
tri -1075 76 -185 445 sw
tri -185 76 -32 445 ne
rect -32 76 32 445
tri 32 76 185 446 nw
tri 185 76 1075 446 se
rect 1075 76 36508 446
rect -36508 13 -185 76
tri -185 13 -32 76 sw
tri -32 13 -5 76 ne
rect -5 13 5 76
tri 5 13 32 76 nw
tri 32 13 184 76 se
rect 184 13 36508 76
rect -36508 2 -32 13
tri -32 2 -5 13 sw
tri -5 2 -1 13 ne
rect -1 2 1 13
tri 1 2 5 13 nw
tri 5 2 31 13 se
rect 31 2 36508 13
rect -36508 -2 -5 2
tri -5 0 -1 2 sw
tri -1 0 0 2 ne
tri 0 0 1 2 nw
tri 1 0 5 2 se
rect 5 0 36508 2
tri -5 -2 -1 0 nw
tri -1 -2 0 0 se
tri 0 -1 2 0 ne
rect 2 -1 36508 0
rect -36508 -13 -31 -2
tri -31 -13 -5 -2 nw
tri -5 -13 -1 -2 se
rect -1 -5 0 -2
tri 0 -5 2 -1 sw
tri 2 -5 13 -1 ne
rect 13 -5 36508 -1
rect -1 -13 2 -5
rect -36508 -76 -184 -13
tri -184 -76 -32 -13 nw
tri -32 -76 -5 -13 se
rect -5 -32 2 -13
tri 2 -32 13 -5 sw
tri 13 -32 76 -5 ne
rect 76 -32 36508 -5
rect -5 -76 13 -32
rect -36508 -446 -1075 -76
tri -1075 -446 -185 -76 nw
tri -185 -446 -32 -76 se
rect -32 -185 13 -76
tri 13 -185 76 -32 sw
tri 76 -185 445 -32 ne
rect 445 -185 36508 -32
rect -32 -446 76 -185
rect -36508 -2596 -6266 -446
tri -6266 -2596 -1076 -446 nw
tri -1075 -2596 -185 -446 se
rect -185 -1075 76 -446
tri 76 -1075 445 -185 sw
tri 445 -1075 2595 -185 ne
rect 2595 -1075 36508 -185
rect -185 -2596 445 -1075
tri -36508 -15125 -6266 -2596 nw
tri -6266 -15125 -1075 -2596 se
rect -1075 -6266 445 -2596
tri 445 -6266 2596 -1075 sw
tri 2596 -6266 15124 -1075 ne
rect 15124 -6266 36508 -1075
rect -1075 -15125 2596 -6266
tri 2596 -15125 6266 -6266 sw
tri 15125 -15125 36508 -6266 ne
tri -15125 -36508 -6266 -15125 se
rect -6266 -36508 6266 -15125
tri 6266 -36508 15125 -15125 sw
<< properties >>
string GDS_END 10411016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10379748
string gencell sky130_fd_pr__rf_test_coil3
string library sky130
string parameter m=1
string path 881.450 -378.100 881.450 -75.000 
<< end >>
