magic
tech sky130A
timestamp 1694700623
<< properties >>
string GDS_END 37256190
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37255674
<< end >>
