magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 11409 32865 11575 33597
rect 20086 31917 20191 33171
<< pwell >>
rect 20703 30227 20797 30315
<< pdiff >>
rect 24027 100 24059 338
rect 25279 100 25317 338
<< poly >>
rect 17794 31703 18050 31729
rect 17794 31669 17810 31703
rect 17844 31669 17905 31703
rect 17939 31669 18000 31703
rect 18034 31669 18050 31703
rect 17794 31653 18050 31669
rect 18278 31703 18534 31729
rect 18278 31669 18294 31703
rect 18328 31669 18389 31703
rect 18423 31669 18484 31703
rect 18518 31669 18534 31703
rect 18278 31653 18534 31669
rect 18740 31703 18996 31729
rect 18740 31669 18756 31703
rect 18790 31669 18851 31703
rect 18885 31669 18946 31703
rect 18980 31669 18996 31703
rect 18740 31653 18996 31669
<< polycont >>
rect 17810 31669 17844 31703
rect 17905 31669 17939 31703
rect 18000 31669 18034 31703
rect 18294 31669 18328 31703
rect 18389 31669 18423 31703
rect 18484 31669 18518 31703
rect 18756 31669 18790 31703
rect 18851 31669 18885 31703
rect 18946 31669 18980 31703
<< locali >>
rect 11905 32815 11943 32849
rect 18106 32832 18143 32883
rect 18072 32798 18110 32832
rect 18106 32781 18143 32798
rect 18420 32730 18486 32781
rect 18414 32696 18452 32730
rect 19219 32745 19253 32783
rect 18420 32693 18486 32696
rect 17794 31669 17810 31703
rect 17844 31669 17905 31703
rect 17939 31669 18000 31703
rect 18034 31669 18050 31703
rect 18278 31669 18294 31703
rect 18328 31669 18389 31703
rect 18423 31669 18484 31703
rect 18518 31669 18534 31703
rect 18740 31669 18756 31703
rect 18790 31669 18851 31703
rect 18885 31669 18946 31703
rect 18980 31669 18996 31703
rect 21039 31431 21141 31442
rect 21073 31397 21111 31431
rect 20858 31347 20965 31355
rect 20858 31313 20859 31347
rect 20893 31313 20931 31347
rect 20858 31229 20965 31313
rect 20855 31163 20965 31229
rect 21039 31196 21141 31397
rect 21555 31164 21733 31229
rect 20495 30803 20529 30841
rect 21276 30803 21310 30841
rect 21555 30560 21645 31164
rect 22011 31163 22085 31229
rect 22031 30803 22065 30841
rect 20319 30493 20353 30527
rect 20671 30493 20705 30539
rect 21175 30493 21209 30527
rect 21855 30493 21889 30527
rect 22207 30493 22241 30527
rect 20705 30427 20795 30493
rect 22633 30443 22671 30477
rect 21467 30347 21505 30381
rect 21641 30344 21679 30378
rect 21903 30344 21941 30378
rect 22495 30336 22533 30370
rect 20705 30271 20815 30303
rect 20705 30237 20795 30271
rect 20319 30191 20353 30237
rect 20671 29981 20829 30237
rect 21175 30191 21209 30237
rect 21555 30191 21589 30237
rect 21855 30191 21889 30237
rect 21935 30191 21969 30237
rect 22207 30183 22241 30237
rect 20419 29894 20493 29928
rect 20527 29894 20600 29928
rect 20855 29881 20929 29947
rect 22011 29881 22121 29947
rect 23494 1124 23532 1158
rect 25810 1124 25848 1158
rect 27356 1129 27394 1163
rect 27110 1060 27180 1063
rect 27132 1026 27170 1060
rect 27110 940 27180 1026
rect 23494 799 23532 833
rect 25923 -2 25961 32
<< viali >>
rect 11871 32815 11905 32849
rect 11943 32815 11977 32849
rect 18038 32798 18072 32832
rect 18110 32798 18144 32832
rect 19219 32783 19253 32817
rect 18380 32696 18414 32730
rect 18452 32696 18486 32730
rect 19219 32711 19253 32745
rect 21039 31397 21073 31431
rect 21111 31397 21145 31431
rect 20859 31313 20893 31347
rect 20931 31313 20965 31347
rect 20495 30841 20529 30875
rect 20495 30769 20529 30803
rect 21276 30841 21310 30875
rect 21276 30769 21310 30803
rect 22031 30841 22065 30875
rect 22031 30769 22065 30803
rect 22599 30443 22633 30477
rect 22671 30443 22705 30477
rect 21433 30347 21467 30381
rect 21505 30347 21539 30381
rect 21607 30344 21641 30378
rect 21679 30344 21713 30378
rect 21869 30344 21903 30378
rect 21941 30344 21975 30378
rect 22461 30336 22495 30370
rect 22533 30336 22567 30370
rect 20671 30237 20705 30271
rect 20795 30237 20829 30271
rect 20385 29894 20419 29928
rect 20493 29894 20527 29928
rect 20600 29894 20634 29928
rect 23460 1124 23494 1158
rect 23532 1124 23566 1158
rect 25776 1124 25810 1158
rect 25848 1124 25882 1158
rect 27322 1129 27356 1163
rect 27394 1129 27428 1163
rect 27098 1026 27132 1060
rect 27170 1026 27204 1060
rect 23460 799 23494 833
rect 23532 799 23566 833
rect 25889 -2 25923 32
rect 25961 -2 25995 32
<< metal1 >>
rect 13706 33704 14081 33705
rect 13706 33652 13712 33704
rect 13764 33652 13790 33704
rect 13842 33652 13868 33704
rect 13920 33652 13946 33704
rect 13998 33652 14023 33704
rect 14075 33652 14081 33704
rect 13706 33636 14081 33652
rect 13706 33584 13712 33636
rect 13764 33584 13790 33636
rect 13842 33584 13868 33636
rect 13920 33584 13946 33636
rect 13998 33584 14023 33636
rect 14075 33584 14081 33636
rect 13706 33568 14081 33584
rect 13706 33516 13712 33568
rect 13764 33516 13790 33568
rect 13842 33516 13868 33568
rect 13920 33516 13946 33568
rect 13998 33516 14023 33568
rect 14075 33516 14081 33568
rect 13706 33500 14081 33516
rect 13706 33448 13712 33500
rect 13764 33448 13790 33500
rect 13842 33448 13868 33500
rect 13920 33448 13946 33500
rect 13998 33448 14023 33500
rect 14075 33448 14081 33500
rect 18821 33497 19162 33656
rect 20137 33591 21700 33592
rect 20137 33539 21391 33591
rect 21443 33539 21473 33591
rect 21525 33539 21555 33591
rect 21607 33539 21636 33591
rect 21688 33539 21700 33591
tri 21700 33561 21731 33592 sw
rect 25522 33552 25809 33554
rect 20137 33527 21700 33539
rect 13706 33447 14081 33448
rect 20137 33475 21391 33527
rect 21443 33475 21473 33527
rect 21525 33475 21555 33527
rect 21607 33475 21636 33527
rect 21688 33478 21700 33527
rect 25453 33551 25809 33552
rect 25453 33499 25459 33551
rect 25511 33499 25548 33551
rect 25600 33499 25637 33551
rect 25689 33499 25726 33551
rect 25778 33499 25809 33551
rect 21688 33475 21694 33478
rect 20137 33463 21694 33475
rect 20137 33411 21391 33463
rect 21443 33411 21473 33463
rect 21525 33411 21555 33463
rect 21607 33411 21636 33463
rect 21688 33411 21694 33463
rect 20137 33399 21694 33411
rect 20137 33347 21391 33399
rect 21443 33347 21473 33399
rect 21525 33347 21555 33399
rect 21607 33347 21636 33399
rect 21688 33347 21694 33399
rect 25453 33471 25809 33499
rect 25453 33419 25459 33471
rect 25511 33419 25548 33471
rect 25600 33419 25637 33471
rect 25689 33419 25726 33471
rect 25778 33419 25809 33471
rect 25453 33391 25809 33419
tri 21694 33347 21725 33378 nw
rect 25453 33339 25459 33391
rect 25511 33339 25548 33391
rect 25600 33339 25637 33391
rect 25689 33339 25726 33391
rect 25778 33339 25809 33391
rect 25453 33338 25809 33339
tri 25529 33328 25539 33338 ne
rect 25539 33328 25809 33338
tri 25539 33274 25593 33328 ne
rect 25593 33322 25809 33328
rect 25593 33270 25595 33322
rect 25647 33270 25663 33322
rect 25715 33270 25731 33322
rect 25783 33270 25809 33322
rect 25593 33258 25809 33270
tri 22919 33189 22953 33223 se
rect 22953 33220 23005 33226
tri 21907 33123 21973 33189 se
rect 21973 33168 22953 33189
rect 21973 33156 23005 33168
rect 21973 33142 22953 33156
tri 21973 33123 21992 33142 nw
tri 22919 33123 22938 33142 ne
rect 22938 33123 22953 33142
tri 21882 33098 21907 33123 se
rect 21907 33098 21948 33123
tri 21948 33098 21973 33123 nw
tri 22938 33108 22953 33123 ne
rect 22953 33098 23005 33104
tri 21850 33066 21882 33098 se
rect 21882 33066 21907 33098
tri 12221 33020 12267 33066 se
rect 12267 33020 13460 33066
tri 12208 33007 12221 33020 se
rect 12221 33014 12281 33020
tri 12281 33014 12287 33020 nw
rect 13454 33014 13460 33020
rect 13512 33014 13524 33066
rect 13576 33014 13582 33066
tri 21841 33057 21850 33066 se
rect 21850 33057 21907 33066
tri 21907 33057 21948 33098 nw
tri 21833 33049 21841 33057 se
rect 20165 33043 20395 33049
rect 12221 33007 12274 33014
tri 12274 33007 12281 33014 nw
tri 12142 32941 12208 33007 se
tri 12208 32941 12274 33007 nw
rect 20217 32991 20395 33043
tri 21775 32991 21833 33049 se
rect 21833 32991 21841 33049
tri 21841 32991 21907 33057 nw
rect 22614 33023 22666 33029
rect 20165 32979 20395 32991
tri 12076 32875 12142 32941 se
tri 12142 32875 12208 32941 nw
rect 20217 32927 20395 32979
rect 20165 32919 20395 32927
tri 21709 32925 21775 32991 se
tri 21775 32925 21841 32991 nw
rect 22614 32959 22666 32971
tri 21703 32919 21709 32925 se
rect 21709 32919 21747 32925
tri 21690 32906 21703 32919 se
rect 21703 32906 21747 32919
tri 21132 32897 21141 32906 sw
tri 21681 32897 21690 32906 se
rect 21690 32897 21747 32906
tri 21747 32897 21775 32925 nw
tri 22666 32943 22700 32977 sw
tri 23275 32909 23309 32943 se
tri 23355 32909 23389 32943 sw
rect 22614 32901 22666 32907
rect 21132 32875 21725 32897
tri 21725 32875 21747 32897 nw
tri 12056 32855 12076 32875 se
rect 12076 32855 12099 32875
rect 11859 32849 12099 32855
rect 11859 32815 11871 32849
rect 11905 32815 11943 32849
rect 11977 32832 12099 32849
tri 12099 32832 12142 32875 nw
rect 21132 32851 21701 32875
tri 21701 32851 21725 32875 nw
rect 23270 32857 23276 32909
rect 23328 32857 23340 32909
rect 23392 32857 23398 32909
tri 23294 32851 23300 32857 ne
rect 23300 32851 23356 32857
rect 21132 32838 21153 32851
tri 21153 32838 21166 32851 nw
tri 23300 32842 23309 32851 ne
rect 23309 32842 23356 32851
tri 23356 32842 23371 32857 nw
rect 18026 32832 18156 32838
rect 11977 32815 12076 32832
rect 11859 32809 12076 32815
tri 12076 32809 12099 32832 nw
rect 18026 32798 18038 32832
rect 18098 32798 18110 32832
rect 18144 32798 18156 32832
rect 21132 32831 21146 32838
tri 21146 32831 21153 32838 nw
rect 18026 32792 18046 32798
rect 18098 32792 18156 32798
rect 19210 32825 19262 32831
tri 21132 32817 21146 32831 nw
rect 18046 32768 18098 32780
rect 19210 32761 19262 32773
rect 18046 32710 18098 32716
rect 18368 32730 18498 32736
rect 18368 32696 18380 32730
rect 18414 32696 18452 32730
rect 18486 32696 18498 32730
rect 18368 32690 18498 32696
rect 18533 32688 18539 32740
rect 18591 32688 18603 32740
rect 18655 32688 18661 32740
tri 25312 32727 25346 32761 se
rect 25346 32727 25398 33240
rect 25593 33206 25595 33258
rect 25647 33206 25663 33258
rect 25715 33206 25731 33258
rect 25783 33206 25809 33258
rect 25593 33194 25809 33206
rect 25593 33142 25595 33194
rect 25647 33142 25663 33194
rect 25715 33142 25731 33194
rect 25783 33142 25809 33194
rect 25593 33129 25809 33142
rect 27389 33256 27441 33262
rect 27389 33192 27441 33204
rect 27389 33134 27441 33140
tri 27441 33134 27515 33208 sw
tri 27390 33132 27392 33134 ne
rect 27392 33132 27515 33134
tri 27515 33132 27517 33134 sw
rect 25593 33077 25595 33129
rect 25647 33077 25663 33129
rect 25715 33077 25731 33129
rect 25783 33077 25809 33129
tri 27392 33103 27421 33132 ne
rect 27421 33103 27500 33132
tri 27421 33095 27429 33103 ne
rect 27429 33095 27500 33103
rect 25593 33064 25809 33077
rect 25593 33012 25595 33064
rect 25647 33012 25663 33064
rect 25715 33012 25731 33064
rect 25783 33012 25809 33064
rect 25593 32999 25809 33012
rect 25593 32947 25595 32999
rect 25647 32947 25663 32999
rect 25715 32947 25731 32999
rect 25783 32947 25809 32999
rect 25593 32934 25809 32947
rect 25593 32882 25595 32934
rect 25647 32882 25663 32934
rect 25715 32882 25731 32934
rect 25783 32882 25809 32934
rect 25593 32869 25809 32882
rect 25593 32817 25595 32869
rect 25647 32817 25663 32869
rect 25715 32817 25731 32869
rect 25783 32817 25809 32869
rect 25593 32804 25809 32817
rect 19210 32703 19262 32709
rect 19213 32699 19259 32703
rect 19964 32525 20257 32727
tri 25311 32726 25312 32727 se
rect 25312 32726 25398 32727
tri 25398 32726 25433 32761 sw
rect 25593 32752 25595 32804
rect 25647 32752 25663 32804
rect 25715 32752 25731 32804
rect 25783 32752 25809 32804
rect 25593 32739 25809 32752
rect 20979 32720 21285 32726
rect 20979 32668 20980 32720
rect 21032 32668 21064 32720
rect 21116 32668 21148 32720
rect 21200 32668 21232 32720
rect 21284 32668 21285 32720
tri 25304 32719 25311 32726 se
rect 25311 32719 25433 32726
tri 25433 32719 25440 32726 sw
rect 20979 32646 21285 32668
rect 20979 32594 20980 32646
rect 21032 32594 21064 32646
rect 21116 32594 21148 32646
rect 21200 32594 21232 32646
rect 21284 32594 21285 32646
rect 20979 32572 21285 32594
rect 14637 32447 14643 32499
rect 14695 32447 14710 32499
rect 14762 32447 14777 32499
rect 14829 32447 14844 32499
rect 14896 32447 14911 32499
rect 14963 32447 14978 32499
rect 15030 32447 15045 32499
rect 15097 32447 15112 32499
rect 15164 32447 15179 32499
rect 15231 32447 15246 32499
rect 15298 32447 15313 32499
rect 15365 32447 15379 32499
rect 15431 32447 15445 32499
rect 15497 32447 15511 32499
rect 15563 32447 15577 32499
rect 15629 32447 15635 32499
rect 14637 32427 15635 32447
rect 14637 32375 14643 32427
rect 14695 32375 14710 32427
rect 14762 32375 14777 32427
rect 14829 32375 14844 32427
rect 14896 32375 14911 32427
rect 14963 32375 14978 32427
rect 15030 32375 15045 32427
rect 15097 32375 15112 32427
rect 15164 32375 15179 32427
rect 15231 32375 15246 32427
rect 15298 32375 15313 32427
rect 15365 32375 15379 32427
rect 15431 32375 15445 32427
rect 15497 32375 15511 32427
rect 15563 32375 15577 32427
rect 15629 32375 15635 32427
rect 14637 32355 15635 32375
rect 19964 32362 20253 32525
rect 20979 32520 20980 32572
rect 21032 32520 21064 32572
rect 21116 32520 21148 32572
rect 21200 32520 21232 32572
rect 21284 32520 21285 32572
rect 20979 32498 21285 32520
rect 20979 32446 20980 32498
rect 21032 32446 21064 32498
rect 21116 32446 21148 32498
rect 21200 32446 21232 32498
rect 21284 32446 21285 32498
rect 20979 32423 21285 32446
rect 20979 32371 20980 32423
rect 21032 32371 21064 32423
rect 21116 32371 21148 32423
rect 21200 32371 21232 32423
rect 21284 32371 21285 32423
rect 20979 32365 21285 32371
rect 25593 32687 25595 32739
rect 25647 32687 25663 32739
rect 25715 32687 25731 32739
rect 25783 32687 25809 32739
rect 25593 32674 25809 32687
rect 25593 32622 25595 32674
rect 25647 32622 25663 32674
rect 25715 32622 25731 32674
rect 25783 32622 25809 32674
tri 25809 32653 25832 32676 nw
rect 25593 32616 25809 32622
rect 25593 32584 25755 32616
tri 25755 32585 25786 32616 nw
rect 25645 32532 25703 32584
rect 25593 32519 25755 32532
rect 25645 32467 25703 32519
rect 25593 32454 25755 32467
rect 25645 32402 25703 32454
rect 25593 32388 25755 32402
rect 14637 32303 14643 32355
rect 14695 32303 14710 32355
rect 14762 32303 14777 32355
rect 14829 32303 14844 32355
rect 14896 32303 14911 32355
rect 14963 32303 14978 32355
rect 15030 32303 15045 32355
rect 15097 32303 15112 32355
rect 15164 32303 15179 32355
rect 15231 32303 15246 32355
rect 15298 32303 15313 32355
rect 15365 32303 15379 32355
rect 15431 32303 15445 32355
rect 15497 32303 15511 32355
rect 15563 32303 15577 32355
rect 15629 32303 15635 32355
rect 25645 32336 25703 32388
rect 25593 32330 25755 32336
rect 23308 32309 23360 32318
rect 11529 32225 19054 32263
rect 19048 32211 19054 32225
rect 19106 32211 19118 32263
rect 19170 32211 19176 32263
rect 27140 32292 27192 32298
rect 23308 32245 23360 32257
rect 23037 32234 23089 32240
tri 23036 32211 23037 32212 se
tri 23003 32178 23036 32211 se
rect 23036 32182 23037 32211
rect 25001 32220 25007 32272
rect 25059 32220 25071 32272
rect 25123 32220 25129 32272
rect 23308 32187 23360 32193
rect 25611 32194 25881 32240
rect 27140 32228 27192 32240
rect 23036 32178 23089 32182
tri 21721 32170 21729 32178 se
rect 21729 32170 23089 32178
tri 21701 32150 21721 32170 se
rect 21721 32150 23037 32170
tri 21692 32141 21701 32150 se
rect 21701 32141 23037 32150
tri 21173 32101 21213 32141 se
rect 21213 32124 23037 32141
rect 21213 32101 21740 32124
tri 21740 32101 21763 32124 nw
tri 23025 32112 23037 32124 ne
rect 23037 32112 23089 32118
rect 21173 32094 21733 32101
tri 21733 32094 21740 32101 nw
tri 21078 31950 21079 31951 sw
rect 21078 31928 21079 31950
tri 21079 31928 21101 31950 sw
tri 21151 31928 21173 31950 se
rect 21173 31928 21233 32094
tri 21233 32060 21267 32094 nw
rect 19149 31924 19852 31928
rect 19149 31872 19337 31924
rect 19389 31872 19402 31924
rect 19454 31872 19467 31924
rect 19519 31872 19532 31924
rect 19584 31872 19597 31924
rect 19649 31872 19662 31924
rect 19714 31872 19726 31924
rect 19778 31872 19790 31924
rect 19842 31872 19852 31924
rect 19149 31852 19852 31872
rect 19149 31800 19337 31852
rect 19389 31800 19402 31852
rect 19454 31800 19467 31852
rect 19519 31800 19532 31852
rect 19584 31800 19597 31852
rect 19649 31800 19662 31852
rect 19714 31800 19726 31852
rect 19778 31800 19790 31852
rect 19842 31800 19852 31852
rect 21078 31925 21101 31928
tri 21101 31925 21104 31928 sw
tri 21148 31925 21151 31928 se
rect 21151 31925 21233 31928
rect 21078 31876 21233 31925
rect 21078 31827 21184 31876
tri 21184 31827 21233 31876 nw
rect 19149 31780 19852 31800
rect 19149 31728 19337 31780
rect 19389 31728 19402 31780
rect 19454 31728 19467 31780
rect 19519 31728 19532 31780
rect 19584 31728 19597 31780
rect 19649 31728 19662 31780
rect 19714 31728 19726 31780
rect 19778 31728 19790 31780
rect 19842 31728 19852 31780
rect 24327 31748 24980 31749
rect 25055 31748 25062 31749
rect 25357 31748 25535 31749
rect 24015 31743 25535 31748
rect 19149 31726 19852 31728
rect 21383 31739 21683 31741
rect 21383 31687 21389 31739
rect 21441 31687 21468 31739
rect 21520 31687 21547 31739
rect 21599 31687 21625 31739
rect 21677 31687 21683 31739
rect 21383 31671 21683 31687
rect 21383 31619 21389 31671
rect 21441 31619 21468 31671
rect 21520 31619 21547 31671
rect 21599 31619 21625 31671
rect 21677 31619 21683 31671
tri 21683 31644 21755 31716 sw
rect 24015 31691 25357 31743
rect 25409 31691 25483 31743
rect 24015 31668 25535 31691
rect 21383 31603 21683 31619
rect 21383 31551 21389 31603
rect 21441 31551 21468 31603
rect 21520 31551 21547 31603
rect 21599 31551 21625 31603
rect 21677 31551 21683 31603
rect 21383 31535 21683 31551
rect 21383 31483 21389 31535
rect 21441 31483 21468 31535
rect 21520 31483 21547 31535
rect 21599 31483 21625 31535
rect 21677 31483 21683 31535
rect 24015 31616 25357 31668
rect 25409 31616 25483 31668
rect 24015 31592 25535 31616
rect 24015 31540 25357 31592
rect 25409 31540 25483 31592
rect 24015 31534 25535 31540
rect 25611 31553 25663 32194
rect 27140 32170 27192 32176
rect 27698 32272 27750 32278
rect 27698 32208 27750 32220
rect 27698 32150 27750 32156
rect 27444 31986 27450 32038
rect 27502 31986 27529 32038
rect 27581 31986 27609 32038
rect 27661 31986 27689 32038
rect 27741 31986 27769 32038
rect 27821 31986 27827 32038
rect 27444 31962 27827 31986
rect 27444 31910 27450 31962
rect 27502 31910 27529 31962
rect 27581 31910 27609 31962
rect 27661 31910 27689 31962
rect 27741 31910 27769 31962
rect 27821 31910 27827 31962
rect 27134 31877 27480 31878
rect 27134 31825 27140 31877
rect 27192 31825 27211 31877
rect 27263 31825 27282 31877
rect 27334 31825 27352 31877
rect 27404 31825 27422 31877
rect 27474 31825 27480 31877
rect 27134 31805 27480 31825
rect 27134 31753 27140 31805
rect 27192 31753 27211 31805
rect 27263 31753 27282 31805
rect 27334 31753 27352 31805
rect 27404 31753 27422 31805
rect 27474 31753 27480 31805
rect 27134 31733 27480 31753
rect 27134 31681 27140 31733
rect 27192 31681 27211 31733
rect 27263 31681 27282 31733
rect 27334 31681 27352 31733
rect 27404 31681 27422 31733
rect 27474 31681 27480 31733
rect 27134 31680 27480 31681
rect 25611 31501 26320 31553
rect 26372 31501 26384 31553
rect 26436 31501 26442 31553
rect 21383 31481 21683 31483
rect 24787 31444 24839 31447
tri 24839 31444 24842 31447 sw
rect 24787 31441 24842 31444
tri 24842 31441 24845 31444 sw
tri 26543 31441 26546 31444 se
rect 26546 31441 26598 31444
rect 20715 31389 20721 31441
rect 20773 31389 20785 31441
rect 20837 31431 21157 31441
rect 20837 31397 21039 31431
rect 21073 31397 21111 31431
rect 21145 31397 21157 31431
rect 20837 31389 21157 31397
tri 21682 31389 21734 31441 se
rect 21734 31389 22575 31441
rect 22627 31389 22639 31441
rect 22691 31389 22697 31441
rect 24839 31439 24845 31441
tri 24845 31439 24847 31441 sw
tri 26541 31439 26543 31441 se
rect 26543 31439 26598 31441
rect 24839 31438 26598 31439
rect 24839 31389 26546 31438
tri 21660 31367 21682 31389 se
rect 21682 31367 21734 31389
tri 21734 31367 21756 31389 nw
rect 24787 31387 26546 31389
rect 24787 31377 24853 31387
tri 21648 31355 21660 31367 se
rect 21660 31355 21722 31367
tri 21722 31355 21734 31367 nw
rect 20828 31347 21670 31355
rect 20828 31313 20859 31347
rect 20893 31313 20931 31347
rect 20965 31313 21670 31347
rect 20828 31303 21670 31313
tri 21670 31303 21722 31355 nw
rect 24839 31367 24853 31377
tri 24853 31367 24873 31387 nw
tri 26512 31367 26532 31387 ne
rect 26532 31386 26546 31387
rect 26532 31374 26598 31386
rect 26532 31367 26546 31374
rect 24839 31355 24841 31367
tri 24841 31355 24853 31367 nw
tri 26532 31355 26544 31367 ne
rect 26544 31355 26546 31367
tri 24839 31353 24841 31355 nw
tri 26544 31353 26546 31355 ne
tri 26289 31347 26294 31352 se
rect 26294 31347 26346 31352
rect 24787 31319 24839 31325
rect 25041 31295 25047 31347
rect 25099 31295 25111 31347
rect 25163 31346 26346 31347
rect 25163 31295 26294 31346
tri 26257 31258 26294 31295 ne
rect 26546 31316 26598 31322
rect 27258 31316 27269 31339
tri 27269 31316 27292 31339 nw
tri 27544 31316 27567 31339 ne
rect 27567 31316 27578 31339
tri 27258 31305 27269 31316 nw
tri 27567 31305 27578 31316 ne
rect 26294 31282 26346 31294
rect 17900 31193 17906 31245
rect 17958 31193 17970 31245
rect 18022 31193 19127 31245
rect 19179 31193 19191 31245
rect 19243 31193 19249 31245
rect 26294 31224 26346 31230
rect 26798 31240 26850 31246
tri 26770 31163 26798 31191 se
rect 26798 31176 26850 31188
rect 24755 31124 26798 31163
tri 26850 31163 26861 31174 sw
rect 26850 31124 26861 31163
rect 24755 31111 26861 31124
tri 26893 31071 26924 31102 se
rect 26924 31096 26976 31102
rect 24844 31044 26924 31071
rect 24844 31032 26976 31044
rect 24844 31019 26924 31032
tri 26893 30988 26924 31019 ne
tri 27258 31024 27292 31058 sw
tri 27544 31024 27578 31058 se
rect 22930 30955 26736 30979
rect 26924 30974 26976 30980
rect 22930 30927 26672 30955
tri 26638 30893 26672 30927 ne
rect 26724 30927 26736 30955
tri 26724 30916 26735 30927 nw
rect 26672 30891 26724 30903
rect 20128 30875 20535 30887
rect 20128 30841 20495 30875
rect 20529 30841 20535 30875
rect 20128 30803 20535 30841
rect 20128 30769 20495 30803
rect 20529 30769 20535 30803
rect 20128 30757 20535 30769
rect 21025 30875 21316 30887
rect 21025 30841 21276 30875
rect 21310 30841 21316 30875
rect 21025 30803 21316 30841
rect 21025 30769 21276 30803
rect 21310 30769 21316 30803
rect 21025 30757 21316 30769
rect 22025 30875 22878 30887
rect 22025 30841 22031 30875
rect 22065 30841 22878 30875
rect 22025 30803 22878 30841
rect 24374 30868 26479 30887
rect 24374 30835 26420 30868
rect 22025 30769 22031 30803
rect 22065 30769 22878 30803
tri 26386 30801 26420 30835 ne
rect 26472 30835 26479 30868
rect 26472 30833 26477 30835
tri 26477 30833 26479 30835 nw
rect 26672 30833 26724 30839
tri 26472 30828 26477 30833 nw
rect 26420 30804 26472 30816
rect 22025 30757 22878 30769
rect 20128 30715 20258 30757
tri 20258 30722 20293 30757 nw
tri 22713 30729 22741 30757 ne
rect 22741 30729 22878 30757
rect 23685 30763 23737 30769
rect 20307 30727 22262 30729
rect 20128 30663 20134 30715
rect 20186 30663 20200 30715
rect 20252 30663 20258 30715
rect 14636 30441 14642 30493
rect 14694 30441 14709 30493
rect 14761 30441 14776 30493
rect 14828 30441 14843 30493
rect 14895 30441 14910 30493
rect 14962 30441 14977 30493
rect 15029 30441 15044 30493
rect 15096 30441 15111 30493
rect 15163 30441 15178 30493
rect 15230 30441 15245 30493
rect 15297 30441 15312 30493
rect 15364 30441 15378 30493
rect 15430 30441 15444 30493
rect 15496 30441 15510 30493
rect 15562 30441 15576 30493
rect 15628 30441 15634 30493
rect 14636 30409 15634 30441
rect 14636 30357 14642 30409
rect 14694 30357 14709 30409
rect 14761 30357 14776 30409
rect 14828 30357 14843 30409
rect 14895 30357 14910 30409
rect 14962 30357 14977 30409
rect 15029 30357 15044 30409
rect 15096 30357 15111 30409
rect 15163 30357 15178 30409
rect 15230 30357 15245 30409
rect 15297 30357 15312 30409
rect 15364 30357 15378 30409
rect 15430 30357 15444 30409
rect 15496 30357 15510 30409
rect 15562 30357 15576 30409
rect 15628 30357 15634 30409
rect 14636 30325 15634 30357
rect 20128 30387 20258 30663
rect 20307 30675 20985 30727
rect 21037 30675 21067 30727
rect 21119 30675 21149 30727
rect 21201 30675 21230 30727
rect 21282 30724 22262 30727
tri 22741 30724 22746 30729 ne
rect 22746 30724 22878 30729
rect 21282 30723 22623 30724
rect 21282 30675 22193 30723
rect 20307 30671 22193 30675
rect 22245 30671 22268 30723
rect 22320 30671 22343 30723
rect 22395 30671 22417 30723
rect 22469 30671 22491 30723
rect 22543 30671 22565 30723
rect 22617 30671 22623 30723
tri 22746 30722 22748 30724 ne
rect 20307 30655 22623 30671
rect 20307 30603 20985 30655
rect 21037 30603 21067 30655
rect 21119 30603 21149 30655
rect 21201 30603 21230 30655
rect 21282 30653 22623 30655
rect 21282 30603 22193 30653
rect 20307 30601 22193 30603
rect 22245 30601 22268 30653
rect 22320 30601 22343 30653
rect 22395 30601 22417 30653
rect 22469 30601 22491 30653
rect 22543 30601 22565 30653
rect 22617 30601 22623 30653
rect 20307 30583 22623 30601
rect 20307 30531 20985 30583
rect 21037 30531 21067 30583
rect 21119 30531 21149 30583
rect 21201 30531 21230 30583
rect 21282 30531 22193 30583
rect 22245 30531 22268 30583
rect 22320 30531 22343 30583
rect 22395 30531 22417 30583
rect 22469 30531 22491 30583
rect 22543 30531 22565 30583
rect 22617 30531 22623 30583
rect 20307 30530 22623 30531
rect 20307 30453 22262 30530
rect 22587 30431 22593 30483
rect 22645 30431 22657 30483
rect 22709 30437 22717 30483
rect 22709 30431 22715 30437
rect 22748 30427 22878 30724
rect 23445 30740 23497 30746
rect 23445 30676 23497 30688
tri 22878 30427 22913 30462 sw
tri 20258 30387 20293 30422 sw
rect 20128 30381 21551 30387
rect 20128 30347 21433 30381
rect 21467 30347 21505 30381
rect 21539 30347 21551 30381
rect 20128 30341 21551 30347
rect 21595 30378 21987 30384
rect 21595 30344 21607 30378
rect 21641 30344 21679 30378
rect 21713 30344 21869 30378
rect 21903 30344 21941 30378
rect 21975 30344 21987 30378
rect 21595 30338 21987 30344
rect 22449 30327 22455 30379
rect 22507 30327 22521 30379
rect 22573 30327 22579 30379
rect 14636 30273 14642 30325
rect 14694 30273 14709 30325
rect 14761 30273 14776 30325
rect 14828 30273 14843 30325
rect 14895 30273 14910 30325
rect 14962 30273 14977 30325
rect 15029 30273 15044 30325
rect 15096 30273 15111 30325
rect 15163 30273 15178 30325
rect 15230 30273 15245 30325
rect 15297 30273 15312 30325
rect 15364 30273 15378 30325
rect 15430 30273 15444 30325
rect 15496 30273 15510 30325
rect 15562 30273 15576 30325
rect 15628 30273 15634 30325
rect 22748 30297 23413 30427
tri 23322 30278 23341 30297 ne
rect 23341 30278 23413 30297
tri 20819 30277 20820 30278 sw
tri 23341 30277 23342 30278 ne
rect 23342 30277 23413 30278
rect 20298 30271 22705 30277
rect 20298 30237 20671 30271
rect 20705 30237 20795 30271
rect 20829 30237 22705 30271
tri 23342 30258 23361 30277 ne
rect 20298 30201 22705 30237
rect 20298 30149 21391 30201
rect 21443 30149 21473 30201
rect 21525 30149 21554 30201
rect 21606 30149 21635 30201
rect 21687 30149 22705 30201
rect 20298 30129 22705 30149
rect 20298 30077 21391 30129
rect 21443 30077 21473 30129
rect 21525 30077 21554 30129
rect 21606 30077 21635 30129
rect 21687 30077 22705 30129
rect 20298 30057 22705 30077
rect 20298 30005 21391 30057
rect 21443 30005 21473 30057
rect 21525 30005 21554 30057
rect 21606 30005 21635 30057
rect 21687 30005 22705 30057
rect 20298 30001 22705 30005
rect 20373 29882 20379 29934
rect 20431 29882 20449 29934
rect 20501 29928 20519 29934
rect 20501 29882 20519 29894
rect 20571 29882 20588 29934
rect 20640 29882 20646 29934
rect 23264 25131 23316 25137
rect 23264 25067 23316 25079
rect 23184 24637 23236 24643
rect 23184 24573 23236 24585
tri 23150 23396 23184 23430 se
rect 23184 23396 23236 24521
rect 22965 23380 23236 23396
rect 22965 23350 23206 23380
tri 23206 23350 23236 23380 nw
rect 22965 23344 23200 23350
tri 23200 23344 23206 23350 nw
tri 23258 23344 23264 23350 se
rect 23264 23344 23316 25015
rect 22965 23316 23023 23344
tri 23023 23316 23051 23344 nw
tri 23230 23316 23258 23344 se
rect 23258 23316 23316 23344
rect 22965 15957 23017 23316
tri 23017 23310 23023 23316 nw
tri 23074 23310 23080 23316 se
rect 23080 23310 23316 23316
tri 23045 23281 23074 23310 se
rect 23074 23281 23316 23310
rect 23045 23264 23316 23281
rect 23361 23341 23413 30277
rect 23445 30231 23497 30624
rect 23445 30167 23497 30179
rect 23445 30109 23497 30115
rect 23525 30740 23577 30746
rect 23525 30676 23577 30688
rect 23443 29837 23495 29843
rect 23443 29755 23495 29785
rect 23443 28484 23495 29703
rect 23443 28402 23495 28432
rect 23443 28336 23495 28350
rect 23361 23277 23413 23289
rect 23045 15957 23097 23264
tri 23097 23230 23131 23264 nw
rect 23361 23219 23413 23225
rect 23445 24063 23497 24082
rect 23445 23999 23497 24011
tri 23411 23156 23445 23190 se
rect 23445 23156 23497 23947
rect 23205 23104 23497 23156
rect 23125 20659 23177 20666
rect 23125 20595 23177 20607
rect 23125 15957 23177 20543
rect 23205 15957 23257 23104
tri 23257 23070 23291 23104 nw
rect 23525 22990 23577 30624
rect 23525 22926 23577 22938
rect 23525 22868 23577 22874
rect 23605 30740 23657 30746
rect 23605 30676 23657 30688
rect 23525 22824 23577 22830
rect 23525 22760 23577 22772
rect 23445 21995 23497 22052
rect 23445 21931 23497 21943
rect 23365 20822 23417 20865
rect 23365 20758 23417 20770
rect 23285 20108 23337 20125
rect 23285 20018 23337 20056
rect 23285 16019 23337 19966
rect 23365 16019 23417 20706
rect 23445 16019 23497 21879
rect 23525 16019 23577 22708
rect 23605 22417 23657 30624
rect 23685 30699 23737 30711
rect 23685 23507 23737 30647
rect 23685 23443 23737 23455
rect 23685 23385 23737 23391
rect 23767 30743 23773 30795
rect 23825 30743 23837 30795
rect 23889 30743 23895 30795
rect 26420 30746 26472 30752
rect 23605 22353 23657 22365
rect 23605 22295 23657 22301
rect 23685 23341 23737 23347
rect 23685 23277 23737 23289
tri 23626 21702 23685 21761 se
rect 23685 21739 23737 23225
rect 23685 21702 23700 21739
tri 23700 21702 23737 21739 nw
rect 23626 15958 23678 21702
tri 23678 21680 23700 21702 nw
tri 23759 20988 23767 20996 se
rect 23767 20989 23804 30743
tri 23804 30713 23834 30743 nw
rect 27973 30703 28028 30709
rect 23860 30632 23984 30638
rect 23912 30580 23932 30632
rect 27720 30625 27777 30660
rect 26861 30619 27063 30625
rect 23860 30560 23984 30580
rect 23912 30508 23932 30560
rect 23860 30488 23984 30508
rect 23912 30436 23932 30488
rect 23860 30430 23984 30436
rect 24018 30535 24024 30587
rect 24076 30535 24094 30587
rect 24146 30535 24164 30587
rect 24216 30535 24234 30587
rect 24286 30535 24304 30587
rect 24356 30535 24374 30587
rect 24426 30535 24444 30587
rect 24496 30535 24514 30587
rect 24566 30535 24584 30587
rect 24636 30535 24642 30587
rect 24018 30523 24642 30535
rect 24018 30471 24024 30523
rect 24076 30471 24094 30523
rect 24146 30471 24164 30523
rect 24216 30471 24234 30523
rect 24286 30471 24304 30523
rect 24356 30471 24374 30523
rect 24426 30471 24444 30523
rect 24496 30471 24514 30523
rect 24566 30471 24584 30523
rect 24636 30471 24642 30523
rect 24018 30459 24642 30471
rect 24018 30407 24024 30459
rect 24076 30407 24094 30459
rect 24146 30407 24164 30459
rect 24216 30407 24234 30459
rect 24286 30407 24304 30459
rect 24356 30407 24374 30459
rect 24426 30407 24444 30459
rect 24496 30407 24514 30459
rect 24566 30407 24584 30459
rect 24636 30407 24642 30459
rect 24018 30395 24642 30407
rect 24018 30343 24024 30395
rect 24076 30343 24094 30395
rect 24146 30343 24164 30395
rect 24216 30343 24234 30395
rect 24286 30343 24304 30395
rect 24356 30343 24374 30395
rect 24426 30343 24444 30395
rect 24496 30343 24514 30395
rect 24566 30343 24584 30395
rect 24636 30343 24642 30395
rect 26861 30567 26862 30619
rect 26914 30567 26936 30619
rect 26988 30567 27010 30619
rect 27062 30567 27063 30619
rect 26861 30547 27063 30567
rect 26861 30495 26862 30547
rect 26914 30495 26936 30547
rect 26988 30495 27010 30547
rect 27062 30495 27063 30547
rect 26861 30475 27063 30495
rect 26861 30423 26862 30475
rect 26914 30423 26936 30475
rect 26988 30423 27010 30475
rect 27062 30423 27063 30475
rect 26861 30402 27063 30423
rect 26861 30350 26862 30402
rect 26914 30350 26936 30402
rect 26988 30350 27010 30402
rect 27062 30350 27063 30402
rect 26861 30344 27063 30350
rect 27575 30619 27777 30625
tri 27777 30623 27811 30657 nw
rect 28025 30651 28028 30703
rect 27973 30623 28028 30651
rect 27575 30567 27576 30619
rect 27628 30567 27650 30619
rect 27702 30567 27724 30619
rect 27776 30567 27777 30619
rect 27575 30547 27777 30567
rect 27575 30495 27576 30547
rect 27628 30495 27650 30547
rect 27702 30495 27724 30547
rect 27776 30495 27777 30547
rect 27575 30474 27777 30495
rect 27575 30422 27576 30474
rect 27628 30422 27650 30474
rect 27702 30422 27724 30474
rect 27776 30422 27777 30474
rect 27575 30401 27777 30422
rect 27575 30349 27576 30401
rect 27628 30349 27650 30401
rect 27702 30349 27724 30401
rect 27776 30349 27777 30401
rect 28025 30571 28028 30623
rect 27973 30543 28028 30571
rect 28025 30491 28028 30543
rect 27973 30463 28028 30491
rect 28025 30411 28028 30463
rect 27973 30406 28028 30411
rect 27973 30405 28027 30406
tri 28027 30405 28028 30406 nw
rect 27973 30402 28024 30405
tri 28024 30402 28027 30405 nw
tri 27973 30399 27976 30402 ne
rect 27976 30399 28021 30402
tri 28021 30399 28024 30402 nw
rect 27575 30343 27777 30349
rect 27313 30021 27365 30027
rect 27313 29957 27365 29969
rect 27313 29899 27365 29905
rect 24184 28137 24386 28143
rect 24184 28085 24185 28137
rect 24237 28085 24259 28137
rect 24311 28085 24333 28137
rect 24385 28085 24386 28137
rect 24184 28067 24386 28085
rect 24184 28015 24185 28067
rect 24237 28015 24259 28067
rect 24311 28015 24333 28067
rect 24385 28015 24386 28067
rect 24184 27997 24386 28015
rect 24184 27945 24185 27997
rect 24237 27945 24259 27997
rect 24311 27945 24333 27997
rect 24385 27945 24386 27997
rect 24184 27927 24386 27945
rect 24184 27875 24185 27927
rect 24237 27875 24259 27927
rect 24311 27875 24333 27927
rect 24385 27875 24386 27927
rect 24184 27857 24386 27875
rect 24184 27805 24185 27857
rect 24237 27805 24259 27857
rect 24311 27805 24333 27857
rect 24385 27805 24386 27857
rect 24184 27786 24386 27805
rect 24184 27734 24185 27786
rect 24237 27734 24259 27786
rect 24311 27734 24333 27786
rect 24385 27734 24386 27786
rect 24184 27715 24386 27734
rect 24184 27663 24185 27715
rect 24237 27663 24259 27715
rect 24311 27663 24333 27715
rect 24385 27663 24386 27715
rect 24184 27657 24386 27663
rect 25307 28137 25437 28143
rect 25359 28085 25385 28137
rect 25307 28053 25437 28085
rect 25359 28001 25385 28053
rect 25307 27969 25437 28001
rect 25359 27917 25385 27969
rect 25307 27884 25437 27917
rect 25359 27832 25385 27884
rect 25307 27799 25437 27832
rect 25359 27747 25385 27799
rect 25307 27714 25437 27747
rect 25359 27662 25385 27714
rect 25307 27656 25437 27662
rect 25923 28137 26053 28143
rect 25975 28085 26001 28137
rect 25923 28053 26053 28085
rect 25975 28001 26001 28053
rect 25923 27969 26053 28001
rect 25975 27917 26001 27969
rect 25923 27884 26053 27917
rect 25975 27832 26001 27884
rect 25923 27799 26053 27832
rect 25975 27747 26001 27799
rect 25923 27714 26053 27747
rect 25975 27662 26001 27714
rect 25923 27656 26053 27662
rect 26335 28137 26537 28143
rect 26335 28085 26336 28137
rect 26388 28085 26410 28137
rect 26462 28085 26484 28137
rect 26536 28085 26537 28137
rect 26335 28067 26537 28085
rect 26335 28015 26336 28067
rect 26388 28015 26410 28067
rect 26462 28015 26484 28067
rect 26536 28015 26537 28067
rect 26335 27997 26537 28015
rect 26335 27945 26336 27997
rect 26388 27945 26410 27997
rect 26462 27945 26484 27997
rect 26536 27945 26537 27997
rect 26335 27927 26537 27945
rect 26335 27875 26336 27927
rect 26388 27875 26410 27927
rect 26462 27875 26484 27927
rect 26536 27875 26537 27927
rect 26335 27856 26537 27875
rect 26335 27804 26336 27856
rect 26388 27804 26410 27856
rect 26462 27804 26484 27856
rect 26536 27804 26537 27856
rect 26335 27785 26537 27804
rect 26335 27733 26336 27785
rect 26388 27733 26410 27785
rect 26462 27733 26484 27785
rect 26536 27733 26537 27785
rect 26335 27714 26537 27733
rect 26335 27662 26336 27714
rect 26388 27662 26410 27714
rect 26462 27662 26484 27714
rect 26536 27662 26537 27714
rect 26335 27656 26537 27662
rect 24184 26791 24386 26797
rect 24184 26739 24185 26791
rect 24237 26739 24259 26791
rect 24311 26739 24333 26791
rect 24385 26739 24386 26791
rect 24184 26721 24386 26739
rect 24184 26669 24185 26721
rect 24237 26669 24259 26721
rect 24311 26669 24333 26721
rect 24385 26669 24386 26721
rect 24184 26651 24386 26669
rect 24184 26599 24185 26651
rect 24237 26599 24259 26651
rect 24311 26599 24333 26651
rect 24385 26599 24386 26651
rect 24184 26581 24386 26599
rect 24184 26529 24185 26581
rect 24237 26529 24259 26581
rect 24311 26529 24333 26581
rect 24385 26529 24386 26581
rect 24184 26510 24386 26529
rect 24184 26458 24185 26510
rect 24237 26458 24259 26510
rect 24311 26458 24333 26510
rect 24385 26458 24386 26510
rect 24184 26439 24386 26458
rect 24184 26387 24185 26439
rect 24237 26387 24259 26439
rect 24311 26387 24333 26439
rect 24385 26387 24386 26439
rect 24184 26368 24386 26387
rect 24184 26316 24185 26368
rect 24237 26316 24259 26368
rect 24311 26316 24333 26368
rect 24385 26316 24386 26368
rect 24184 26310 24386 26316
rect 25413 26791 25543 26797
rect 25465 26739 25491 26791
rect 25413 26707 25543 26739
rect 25465 26655 25491 26707
rect 25413 26623 25543 26655
rect 25465 26571 25491 26623
rect 25413 26538 25543 26571
rect 25465 26486 25491 26538
rect 25413 26453 25543 26486
rect 25465 26401 25491 26453
rect 25413 26368 25543 26401
rect 25465 26316 25491 26368
rect 25413 26310 25543 26316
rect 25923 26791 26053 26797
rect 25975 26739 26001 26791
rect 25923 26707 26053 26739
rect 25975 26655 26001 26707
rect 25923 26623 26053 26655
rect 25975 26571 26001 26623
rect 25923 26538 26053 26571
rect 25975 26486 26001 26538
rect 25923 26453 26053 26486
rect 25975 26401 26001 26453
rect 25923 26368 26053 26401
rect 25975 26316 26001 26368
rect 25923 26310 26053 26316
rect 26335 26791 26537 26797
rect 26335 26739 26336 26791
rect 26388 26739 26410 26791
rect 26462 26739 26484 26791
rect 26536 26739 26537 26791
rect 26335 26721 26537 26739
rect 26335 26669 26336 26721
rect 26388 26669 26410 26721
rect 26462 26669 26484 26721
rect 26536 26669 26537 26721
rect 26335 26651 26537 26669
rect 26335 26599 26336 26651
rect 26388 26599 26410 26651
rect 26462 26599 26484 26651
rect 26536 26599 26537 26651
rect 26335 26581 26537 26599
rect 26335 26529 26336 26581
rect 26388 26529 26410 26581
rect 26462 26529 26484 26581
rect 26536 26529 26537 26581
rect 26335 26510 26537 26529
rect 26335 26458 26336 26510
rect 26388 26458 26410 26510
rect 26462 26458 26484 26510
rect 26536 26458 26537 26510
rect 26335 26439 26537 26458
rect 26335 26387 26336 26439
rect 26388 26387 26410 26439
rect 26462 26387 26484 26439
rect 26536 26387 26537 26439
rect 26335 26368 26537 26387
rect 26335 26316 26336 26368
rect 26388 26316 26410 26368
rect 26462 26316 26484 26368
rect 26536 26316 26537 26368
rect 26335 26310 26537 26316
rect 27171 24063 27223 24069
rect 27171 23999 27223 24011
rect 27171 23941 27223 23947
rect 25657 23437 25663 23489
rect 25715 23437 25727 23489
rect 25779 23437 25785 23489
tri 25691 23419 25709 23437 ne
rect 25709 23419 25720 23437
tri 25772 23424 25785 23437 nw
rect 27171 23419 27217 23941
tri 27217 23935 27223 23941 nw
tri 25709 23408 25720 23419 ne
rect 26707 23136 26759 23143
rect 26707 23072 26759 23084
rect 26707 23013 26759 23020
rect 27283 22813 27335 22823
rect 27283 22749 27335 22761
rect 27283 22691 27335 22697
rect 26633 22428 26685 22436
rect 26633 22364 26685 22376
rect 26633 22306 26685 22312
rect 24184 22263 24386 22269
rect 24184 22211 24185 22263
rect 24237 22211 24259 22263
rect 24311 22211 24333 22263
rect 24385 22211 24386 22263
rect 24184 22198 24386 22211
rect 24184 22146 24185 22198
rect 24237 22146 24259 22198
rect 24311 22146 24333 22198
rect 24385 22146 24386 22198
rect 24184 22133 24386 22146
rect 24184 22081 24185 22133
rect 24237 22081 24259 22133
rect 24311 22081 24333 22133
rect 24385 22081 24386 22133
rect 24184 22067 24386 22081
rect 24184 22015 24185 22067
rect 24237 22015 24259 22067
rect 24311 22015 24333 22067
rect 24385 22015 24386 22067
rect 24184 22009 24386 22015
rect 25307 22263 25437 22269
rect 25359 22211 25385 22263
rect 25307 22165 25437 22211
rect 25359 22113 25385 22165
rect 25307 22067 25437 22113
rect 25359 22015 25385 22067
rect 25307 22009 25437 22015
rect 25923 22263 26053 22269
rect 25975 22211 26001 22263
rect 25923 22165 26053 22211
rect 25975 22113 26001 22165
rect 25923 22067 26053 22113
rect 25975 22015 26001 22067
rect 25923 22009 26053 22015
rect 26335 22263 26537 22269
rect 26335 22211 26336 22263
rect 26388 22211 26410 22263
rect 26462 22211 26484 22263
rect 26536 22211 26537 22263
rect 26335 22198 26537 22211
rect 26335 22146 26336 22198
rect 26388 22146 26410 22198
rect 26462 22146 26484 22198
rect 26536 22146 26537 22198
rect 26335 22133 26537 22146
rect 26335 22081 26336 22133
rect 26388 22081 26410 22133
rect 26462 22081 26484 22133
rect 26536 22081 26537 22133
rect 26335 22067 26537 22081
rect 26335 22015 26336 22067
rect 26388 22015 26410 22067
rect 26462 22015 26484 22067
rect 26536 22015 26537 22067
rect 26335 22009 26537 22015
rect 27283 21984 27335 21990
rect 27283 21920 27335 21932
rect 27283 21862 27335 21868
tri 27283 21856 27289 21862 ne
rect 27289 21665 27335 21862
tri 27293 21048 27299 21054 sw
rect 27247 21042 27299 21048
tri 23804 20989 23811 20996 sw
rect 23767 20988 23811 20989
rect 23759 20982 23811 20988
rect 23759 20918 23811 20930
rect 23759 20860 23811 20866
tri 23759 20852 23767 20860 ne
rect 23767 19251 23804 20860
tri 23804 20853 23811 20860 nw
rect 25465 20961 25517 20986
rect 27247 20978 27299 20990
rect 27247 20920 27299 20926
tri 27293 20914 27299 20920 nw
rect 25465 20897 25517 20909
tri 27502 20854 27519 20871 se
rect 27519 20854 27547 23545
rect 27720 23166 27777 30343
tri 27710 23099 27777 23166 nw
rect 25465 20839 25517 20845
tri 26127 20847 26134 20854 sw
rect 26127 20717 26134 20847
tri 27495 20847 27502 20854 se
rect 27502 20847 27547 20854
rect 27495 20841 27547 20847
rect 27495 20777 27547 20789
rect 27495 20719 27547 20725
tri 26127 20710 26134 20717 nw
rect 25661 18956 25665 18961
rect 24184 18271 24386 18277
rect 24184 18219 24185 18271
rect 24237 18219 24259 18271
rect 24311 18219 24333 18271
rect 24385 18219 24386 18271
rect 24184 18206 24386 18219
rect 24184 18154 24185 18206
rect 24237 18154 24259 18206
rect 24311 18154 24333 18206
rect 24385 18154 24386 18206
rect 24184 18141 24386 18154
rect 24184 18089 24185 18141
rect 24237 18089 24259 18141
rect 24311 18089 24333 18141
rect 24385 18089 24386 18141
rect 24184 18075 24386 18089
rect 24184 18023 24185 18075
rect 24237 18023 24259 18075
rect 24311 18023 24333 18075
rect 24385 18023 24386 18075
rect 24184 18017 24386 18023
rect 25307 18271 25437 18277
rect 25359 18219 25385 18271
rect 25307 18173 25437 18219
rect 25359 18121 25385 18173
rect 25307 18075 25437 18121
rect 25359 18023 25385 18075
rect 25307 18017 25437 18023
rect 25923 18271 26053 18277
rect 25975 18219 26001 18271
rect 25923 18173 26053 18219
rect 25975 18121 26001 18173
rect 25923 18075 26053 18121
rect 25975 18023 26001 18075
rect 25923 18017 26053 18023
rect 26335 18271 26537 18277
rect 26335 18219 26336 18271
rect 26388 18219 26410 18271
rect 26462 18219 26484 18271
rect 26536 18219 26537 18271
rect 26335 18206 26537 18219
rect 26335 18154 26336 18206
rect 26388 18154 26410 18206
rect 26462 18154 26484 18206
rect 26536 18154 26537 18206
rect 26335 18141 26537 18154
rect 26335 18089 26336 18141
rect 26388 18089 26410 18141
rect 26462 18089 26484 18141
rect 26536 18089 26537 18141
rect 26335 18075 26537 18089
rect 26335 18023 26336 18075
rect 26388 18023 26410 18075
rect 26462 18023 26484 18075
rect 26536 18023 26537 18075
rect 26335 18017 26537 18023
rect 22370 1898 22620 2182
rect 23269 2133 23385 2139
rect 23321 2081 23333 2133
rect 23269 2019 23385 2081
rect 23321 1967 23333 2019
rect 23269 1961 23385 1967
rect 25764 1875 25770 1927
rect 25822 1875 25836 1927
rect 25888 1875 25894 1927
rect 23083 1691 23153 1780
rect 25138 1648 25144 1700
rect 25196 1648 25208 1700
rect 25260 1648 25390 1700
tri 25368 1641 25375 1648 ne
rect 25375 1641 25390 1648
tri 25390 1641 25449 1700 sw
tri 25375 1626 25390 1641 ne
rect 25390 1637 26545 1641
tri 26545 1637 26549 1641 sw
rect 25390 1626 26549 1637
tri 25390 1595 25421 1626 ne
rect 25421 1595 26549 1626
tri 25421 1589 25427 1595 ne
rect 25427 1589 26066 1595
tri 26066 1589 26072 1595 nw
tri 26525 1589 26531 1595 ne
rect 26531 1589 26549 1595
tri 26531 1571 26549 1589 ne
tri 26549 1577 26609 1637 sw
rect 26549 1571 26609 1577
tri 26609 1571 26615 1577 sw
tri 26851 1571 26857 1577 se
rect 26857 1571 26863 1577
tri 26549 1525 26595 1571 ne
rect 26595 1525 26863 1571
rect 26915 1525 26927 1577
rect 26979 1525 26985 1577
rect 27043 1420 27543 1421
rect 27043 1368 27049 1420
rect 27101 1368 27122 1420
rect 27174 1368 27195 1420
rect 27247 1368 27268 1420
rect 27320 1368 27341 1420
rect 27393 1368 27413 1420
rect 27465 1368 27485 1420
rect 27537 1368 27543 1420
rect 27043 1346 27543 1368
rect 27043 1294 27049 1346
rect 27101 1294 27122 1346
rect 27174 1294 27195 1346
rect 27247 1294 27268 1346
rect 27320 1294 27341 1346
rect 27393 1294 27413 1346
rect 27465 1294 27485 1346
rect 27537 1294 27543 1346
rect 27043 1272 27543 1294
rect 27043 1220 27049 1272
rect 27101 1220 27122 1272
rect 27174 1220 27195 1272
rect 27247 1220 27268 1272
rect 27320 1220 27341 1272
rect 27393 1220 27413 1272
rect 27465 1220 27485 1272
rect 27537 1220 27543 1272
rect 27043 1219 27543 1220
tri 27308 1167 27310 1169 se
rect 27310 1167 27440 1169
tri 27440 1167 27441 1168 sw
rect 23248 1115 23254 1167
rect 23306 1115 23320 1167
rect 23372 1158 23578 1167
rect 23372 1124 23460 1158
rect 23494 1124 23532 1158
rect 23566 1124 23578 1158
rect 23372 1115 23578 1124
rect 24138 1125 24190 1131
tri 24123 1085 24138 1100 se
tri 22828 1070 22843 1085 se
rect 22843 1073 24138 1085
rect 25505 1115 25511 1167
rect 25563 1115 25575 1167
rect 25627 1115 25633 1167
rect 25764 1115 25770 1167
rect 25822 1115 25836 1167
rect 25888 1115 25894 1167
tri 26611 1163 26615 1167 se
rect 26615 1163 27319 1167
tri 26577 1129 26611 1163 se
rect 26611 1129 27319 1163
tri 26563 1115 26577 1129 se
rect 26577 1115 27319 1129
rect 27371 1115 27383 1167
rect 27435 1115 27441 1167
rect 22843 1070 24190 1073
rect 22124 1061 24190 1070
rect 22124 1033 24138 1061
rect 22124 1026 22858 1033
tri 22858 1026 22865 1033 nw
tri 24108 1026 24115 1033 ne
rect 24115 1026 24138 1033
rect 22124 1018 22850 1026
tri 22850 1018 22858 1026 nw
tri 24115 1018 24123 1026 ne
rect 24123 1018 24138 1026
tri 24123 1003 24138 1018 ne
tri 24420 1060 24445 1085 se
rect 24445 1060 25303 1085
tri 25303 1060 25328 1085 sw
rect 25505 1082 25633 1115
tri 25633 1082 25666 1115 sw
tri 26530 1082 26563 1115 se
rect 26563 1082 26623 1115
tri 26623 1082 26656 1115 nw
rect 25505 1060 26601 1082
tri 26601 1060 26623 1082 nw
tri 24393 1033 24420 1060 se
rect 24420 1033 25328 1060
tri 25328 1033 25355 1060 sw
tri 24390 1030 24393 1033 se
rect 24393 1030 24464 1033
tri 24464 1030 24467 1033 nw
tri 25281 1030 25284 1033 ne
rect 25284 1030 25355 1033
rect 25505 1030 26571 1060
tri 26571 1030 26601 1060 nw
tri 24386 1026 24390 1030 se
rect 24390 1026 24460 1030
tri 24460 1026 24464 1030 nw
tri 25284 1026 25288 1030 ne
rect 25288 1026 25355 1030
tri 24371 1011 24386 1026 se
rect 24386 1011 24445 1026
tri 24445 1011 24460 1026 nw
tri 25288 1011 25303 1026 ne
rect 24138 1003 24190 1009
tri 24363 1003 24371 1011 se
tri 24297 937 24363 1003 se
rect 24363 937 24371 1003
tri 24371 937 24445 1011 nw
tri 24279 919 24297 937 se
rect 24297 919 24353 937
tri 24353 919 24371 937 nw
tri 24276 916 24279 919 se
rect 24279 916 24350 919
tri 24350 916 24353 919 nw
tri 24678 916 24681 919 se
rect 24681 916 24733 919
tri 24239 879 24276 916 se
rect 24276 879 24313 916
tri 24313 879 24350 916 nw
rect 24579 913 24733 916
tri 24027 873 24033 879 se
rect 24033 873 24304 879
rect 20327 870 20770 873
tri 20770 870 20773 873 sw
tri 24024 870 24027 873 se
rect 24027 870 24304 873
tri 24304 870 24313 879 nw
rect 24579 870 24681 913
rect 20327 833 20773 870
tri 20773 833 20810 870 sw
tri 23996 842 24024 870 se
rect 24024 842 24274 870
rect 20327 832 20810 833
tri 20810 832 20811 833 sw
rect 20327 823 20811 832
tri 20811 823 20820 832 sw
rect 20327 821 20820 823
tri 20748 799 20770 821 ne
rect 20770 799 20820 821
tri 20820 799 20844 823 sw
tri 20770 758 20811 799 ne
rect 20811 791 20844 799
tri 20844 791 20852 799 sw
rect 20811 767 20852 791
tri 20852 767 20876 791 sw
rect 23248 790 23254 842
rect 23306 790 23320 842
rect 23372 833 23578 842
rect 23372 799 23460 833
rect 23494 799 23532 833
rect 23566 799 23578 833
tri 23977 823 23996 842 se
rect 23996 840 24274 842
tri 24274 840 24304 870 nw
tri 24645 840 24675 870 ne
rect 24675 861 24681 870
rect 24675 849 24733 861
rect 24675 840 24681 849
rect 23996 823 24033 840
tri 24033 823 24050 840 nw
tri 24675 834 24681 840 ne
rect 23372 790 23578 799
tri 23945 791 23977 823 se
rect 23977 791 24001 823
tri 24001 791 24033 823 nw
rect 24681 791 24733 797
tri 23944 790 23945 791 se
rect 23945 790 23977 791
tri 23921 767 23944 790 se
rect 23944 767 23977 790
tri 23977 767 24001 791 nw
rect 20811 758 20876 767
tri 20876 758 20885 767 sw
tri 23912 758 23921 767 se
tri 20811 684 20885 758 ne
tri 20885 711 20932 758 sw
tri 23865 711 23912 758 se
rect 23912 711 23921 758
tri 23921 711 23977 767 nw
rect 20885 697 20932 711
tri 20932 697 20946 711 sw
tri 23851 697 23865 711 se
rect 23865 697 23907 711
tri 23907 697 23921 711 nw
rect 20885 684 20946 697
tri 20946 684 20959 697 sw
tri 23838 684 23851 697 se
rect 23851 684 23894 697
tri 23894 684 23907 697 nw
rect 25303 684 25355 1026
rect 27086 1020 27092 1072
rect 27144 1020 27156 1072
rect 27208 1066 27214 1072
rect 27208 1020 27216 1066
tri 25355 684 25368 697 sw
tri 20885 632 20937 684 ne
rect 20937 681 23891 684
tri 23891 681 23894 684 nw
rect 20937 632 23842 681
tri 23842 632 23891 681 nw
rect 23946 678 24152 681
rect 23946 626 23953 678
rect 24005 626 24018 678
rect 24070 626 24152 678
rect 25303 675 25377 684
tri 25303 632 25346 675 ne
rect 25346 632 25377 675
rect 25429 632 25441 684
rect 25493 632 25499 684
rect 23946 614 24152 626
rect 23946 562 23953 614
rect 24005 562 24018 614
rect 24070 562 24152 614
rect 23946 551 24152 562
rect 27043 378 27049 430
rect 27101 378 27158 430
rect 27210 378 27267 430
rect 27319 378 27376 430
rect 27428 378 27485 430
rect 27537 378 27543 430
rect 27043 352 27543 378
rect 27043 300 27049 352
rect 27101 300 27158 352
rect 27210 300 27267 352
rect 27319 300 27376 352
rect 27428 300 27485 352
rect 27537 300 27543 352
rect 18821 86 19162 245
rect 25877 -11 25883 41
rect 25935 -11 25949 41
rect 26001 -11 26007 41
<< via1 >>
rect 13712 33652 13764 33704
rect 13790 33652 13842 33704
rect 13868 33652 13920 33704
rect 13946 33652 13998 33704
rect 14023 33652 14075 33704
rect 13712 33584 13764 33636
rect 13790 33584 13842 33636
rect 13868 33584 13920 33636
rect 13946 33584 13998 33636
rect 14023 33584 14075 33636
rect 13712 33516 13764 33568
rect 13790 33516 13842 33568
rect 13868 33516 13920 33568
rect 13946 33516 13998 33568
rect 14023 33516 14075 33568
rect 13712 33448 13764 33500
rect 13790 33448 13842 33500
rect 13868 33448 13920 33500
rect 13946 33448 13998 33500
rect 14023 33448 14075 33500
rect 21391 33539 21443 33591
rect 21473 33539 21525 33591
rect 21555 33539 21607 33591
rect 21636 33539 21688 33591
rect 21391 33475 21443 33527
rect 21473 33475 21525 33527
rect 21555 33475 21607 33527
rect 21636 33475 21688 33527
rect 25459 33499 25511 33551
rect 25548 33499 25600 33551
rect 25637 33499 25689 33551
rect 25726 33499 25778 33551
rect 21391 33411 21443 33463
rect 21473 33411 21525 33463
rect 21555 33411 21607 33463
rect 21636 33411 21688 33463
rect 21391 33347 21443 33399
rect 21473 33347 21525 33399
rect 21555 33347 21607 33399
rect 21636 33347 21688 33399
rect 25459 33419 25511 33471
rect 25548 33419 25600 33471
rect 25637 33419 25689 33471
rect 25726 33419 25778 33471
rect 25459 33339 25511 33391
rect 25548 33339 25600 33391
rect 25637 33339 25689 33391
rect 25726 33339 25778 33391
rect 25595 33270 25647 33322
rect 25663 33270 25715 33322
rect 25731 33270 25783 33322
rect 22953 33168 23005 33220
rect 22953 33104 23005 33156
rect 13460 33014 13512 33066
rect 13524 33014 13576 33066
rect 20165 32991 20217 33043
rect 20165 32927 20217 32979
rect 22614 32971 22666 33023
rect 22614 32907 22666 32959
rect 23276 32857 23328 32909
rect 23340 32857 23392 32909
rect 18046 32798 18072 32832
rect 18072 32798 18098 32832
rect 18046 32780 18098 32798
rect 19210 32817 19262 32825
rect 18046 32716 18098 32768
rect 19210 32783 19219 32817
rect 19219 32783 19253 32817
rect 19253 32783 19262 32817
rect 19210 32773 19262 32783
rect 19210 32745 19262 32761
rect 18539 32688 18591 32740
rect 18603 32688 18655 32740
rect 19210 32711 19219 32745
rect 19219 32711 19253 32745
rect 19253 32711 19262 32745
rect 25595 33206 25647 33258
rect 25663 33206 25715 33258
rect 25731 33206 25783 33258
rect 25595 33142 25647 33194
rect 25663 33142 25715 33194
rect 25731 33142 25783 33194
rect 27389 33204 27441 33256
rect 27389 33140 27441 33192
rect 25595 33077 25647 33129
rect 25663 33077 25715 33129
rect 25731 33077 25783 33129
rect 25595 33012 25647 33064
rect 25663 33012 25715 33064
rect 25731 33012 25783 33064
rect 25595 32947 25647 32999
rect 25663 32947 25715 32999
rect 25731 32947 25783 32999
rect 25595 32882 25647 32934
rect 25663 32882 25715 32934
rect 25731 32882 25783 32934
rect 25595 32817 25647 32869
rect 25663 32817 25715 32869
rect 25731 32817 25783 32869
rect 19210 32709 19262 32711
rect 25595 32752 25647 32804
rect 25663 32752 25715 32804
rect 25731 32752 25783 32804
rect 20980 32668 21032 32720
rect 21064 32668 21116 32720
rect 21148 32668 21200 32720
rect 21232 32668 21284 32720
rect 20980 32594 21032 32646
rect 21064 32594 21116 32646
rect 21148 32594 21200 32646
rect 21232 32594 21284 32646
rect 14643 32447 14695 32499
rect 14710 32447 14762 32499
rect 14777 32447 14829 32499
rect 14844 32447 14896 32499
rect 14911 32447 14963 32499
rect 14978 32447 15030 32499
rect 15045 32447 15097 32499
rect 15112 32447 15164 32499
rect 15179 32447 15231 32499
rect 15246 32447 15298 32499
rect 15313 32447 15365 32499
rect 15379 32447 15431 32499
rect 15445 32447 15497 32499
rect 15511 32447 15563 32499
rect 15577 32447 15629 32499
rect 14643 32375 14695 32427
rect 14710 32375 14762 32427
rect 14777 32375 14829 32427
rect 14844 32375 14896 32427
rect 14911 32375 14963 32427
rect 14978 32375 15030 32427
rect 15045 32375 15097 32427
rect 15112 32375 15164 32427
rect 15179 32375 15231 32427
rect 15246 32375 15298 32427
rect 15313 32375 15365 32427
rect 15379 32375 15431 32427
rect 15445 32375 15497 32427
rect 15511 32375 15563 32427
rect 15577 32375 15629 32427
rect 20980 32520 21032 32572
rect 21064 32520 21116 32572
rect 21148 32520 21200 32572
rect 21232 32520 21284 32572
rect 20980 32446 21032 32498
rect 21064 32446 21116 32498
rect 21148 32446 21200 32498
rect 21232 32446 21284 32498
rect 20980 32371 21032 32423
rect 21064 32371 21116 32423
rect 21148 32371 21200 32423
rect 21232 32371 21284 32423
rect 25595 32687 25647 32739
rect 25663 32687 25715 32739
rect 25731 32687 25783 32739
rect 25595 32622 25647 32674
rect 25663 32622 25715 32674
rect 25731 32622 25783 32674
rect 25593 32532 25645 32584
rect 25703 32532 25755 32584
rect 25593 32467 25645 32519
rect 25703 32467 25755 32519
rect 25593 32402 25645 32454
rect 25703 32402 25755 32454
rect 14643 32303 14695 32355
rect 14710 32303 14762 32355
rect 14777 32303 14829 32355
rect 14844 32303 14896 32355
rect 14911 32303 14963 32355
rect 14978 32303 15030 32355
rect 15045 32303 15097 32355
rect 15112 32303 15164 32355
rect 15179 32303 15231 32355
rect 15246 32303 15298 32355
rect 15313 32303 15365 32355
rect 15379 32303 15431 32355
rect 15445 32303 15497 32355
rect 15511 32303 15563 32355
rect 15577 32303 15629 32355
rect 25593 32336 25645 32388
rect 25703 32336 25755 32388
rect 19054 32211 19106 32263
rect 19118 32211 19170 32263
rect 23308 32257 23360 32309
rect 23037 32182 23089 32234
rect 23308 32193 23360 32245
rect 25007 32220 25059 32272
rect 25071 32220 25123 32272
rect 27140 32240 27192 32292
rect 23037 32118 23089 32170
rect 19337 31872 19389 31924
rect 19402 31872 19454 31924
rect 19467 31872 19519 31924
rect 19532 31872 19584 31924
rect 19597 31872 19649 31924
rect 19662 31872 19714 31924
rect 19726 31872 19778 31924
rect 19790 31872 19842 31924
rect 19337 31800 19389 31852
rect 19402 31800 19454 31852
rect 19467 31800 19519 31852
rect 19532 31800 19584 31852
rect 19597 31800 19649 31852
rect 19662 31800 19714 31852
rect 19726 31800 19778 31852
rect 19790 31800 19842 31852
rect 19337 31728 19389 31780
rect 19402 31728 19454 31780
rect 19467 31728 19519 31780
rect 19532 31728 19584 31780
rect 19597 31728 19649 31780
rect 19662 31728 19714 31780
rect 19726 31728 19778 31780
rect 19790 31728 19842 31780
rect 21389 31687 21441 31739
rect 21468 31687 21520 31739
rect 21547 31687 21599 31739
rect 21625 31687 21677 31739
rect 21389 31619 21441 31671
rect 21468 31619 21520 31671
rect 21547 31619 21599 31671
rect 21625 31619 21677 31671
rect 25357 31691 25409 31743
rect 25483 31691 25535 31743
rect 21389 31551 21441 31603
rect 21468 31551 21520 31603
rect 21547 31551 21599 31603
rect 21625 31551 21677 31603
rect 21389 31483 21441 31535
rect 21468 31483 21520 31535
rect 21547 31483 21599 31535
rect 21625 31483 21677 31535
rect 25357 31616 25409 31668
rect 25483 31616 25535 31668
rect 25357 31540 25409 31592
rect 25483 31540 25535 31592
rect 27140 32176 27192 32228
rect 27698 32220 27750 32272
rect 27698 32156 27750 32208
rect 27450 31986 27502 32038
rect 27529 31986 27581 32038
rect 27609 31986 27661 32038
rect 27689 31986 27741 32038
rect 27769 31986 27821 32038
rect 27450 31910 27502 31962
rect 27529 31910 27581 31962
rect 27609 31910 27661 31962
rect 27689 31910 27741 31962
rect 27769 31910 27821 31962
rect 27140 31825 27192 31877
rect 27211 31825 27263 31877
rect 27282 31825 27334 31877
rect 27352 31825 27404 31877
rect 27422 31825 27474 31877
rect 27140 31753 27192 31805
rect 27211 31753 27263 31805
rect 27282 31753 27334 31805
rect 27352 31753 27404 31805
rect 27422 31753 27474 31805
rect 27140 31681 27192 31733
rect 27211 31681 27263 31733
rect 27282 31681 27334 31733
rect 27352 31681 27404 31733
rect 27422 31681 27474 31733
rect 26320 31501 26372 31553
rect 26384 31501 26436 31553
rect 20721 31389 20773 31441
rect 20785 31389 20837 31441
rect 22575 31389 22627 31441
rect 22639 31389 22691 31441
rect 24787 31389 24839 31441
rect 24787 31325 24839 31377
rect 26546 31386 26598 31438
rect 25047 31295 25099 31347
rect 25111 31295 25163 31347
rect 26294 31294 26346 31346
rect 26546 31322 26598 31374
rect 17906 31193 17958 31245
rect 17970 31193 18022 31245
rect 19127 31193 19179 31245
rect 19191 31193 19243 31245
rect 26294 31230 26346 31282
rect 26798 31188 26850 31240
rect 26798 31124 26850 31176
rect 26924 31044 26976 31096
rect 26924 30980 26976 31032
rect 26672 30903 26724 30955
rect 26420 30816 26472 30868
rect 26672 30839 26724 30891
rect 20134 30663 20186 30715
rect 20200 30663 20252 30715
rect 14642 30441 14694 30493
rect 14709 30441 14761 30493
rect 14776 30441 14828 30493
rect 14843 30441 14895 30493
rect 14910 30441 14962 30493
rect 14977 30441 15029 30493
rect 15044 30441 15096 30493
rect 15111 30441 15163 30493
rect 15178 30441 15230 30493
rect 15245 30441 15297 30493
rect 15312 30441 15364 30493
rect 15378 30441 15430 30493
rect 15444 30441 15496 30493
rect 15510 30441 15562 30493
rect 15576 30441 15628 30493
rect 14642 30357 14694 30409
rect 14709 30357 14761 30409
rect 14776 30357 14828 30409
rect 14843 30357 14895 30409
rect 14910 30357 14962 30409
rect 14977 30357 15029 30409
rect 15044 30357 15096 30409
rect 15111 30357 15163 30409
rect 15178 30357 15230 30409
rect 15245 30357 15297 30409
rect 15312 30357 15364 30409
rect 15378 30357 15430 30409
rect 15444 30357 15496 30409
rect 15510 30357 15562 30409
rect 15576 30357 15628 30409
rect 20985 30675 21037 30727
rect 21067 30675 21119 30727
rect 21149 30675 21201 30727
rect 21230 30675 21282 30727
rect 22193 30671 22245 30723
rect 22268 30671 22320 30723
rect 22343 30671 22395 30723
rect 22417 30671 22469 30723
rect 22491 30671 22543 30723
rect 22565 30671 22617 30723
rect 20985 30603 21037 30655
rect 21067 30603 21119 30655
rect 21149 30603 21201 30655
rect 21230 30603 21282 30655
rect 22193 30601 22245 30653
rect 22268 30601 22320 30653
rect 22343 30601 22395 30653
rect 22417 30601 22469 30653
rect 22491 30601 22543 30653
rect 22565 30601 22617 30653
rect 20985 30531 21037 30583
rect 21067 30531 21119 30583
rect 21149 30531 21201 30583
rect 21230 30531 21282 30583
rect 22193 30531 22245 30583
rect 22268 30531 22320 30583
rect 22343 30531 22395 30583
rect 22417 30531 22469 30583
rect 22491 30531 22543 30583
rect 22565 30531 22617 30583
rect 22593 30477 22645 30483
rect 22593 30443 22599 30477
rect 22599 30443 22633 30477
rect 22633 30443 22645 30477
rect 22593 30431 22645 30443
rect 22657 30477 22709 30483
rect 22657 30443 22671 30477
rect 22671 30443 22705 30477
rect 22705 30443 22709 30477
rect 22657 30431 22709 30443
rect 23445 30688 23497 30740
rect 23445 30624 23497 30676
rect 22455 30370 22507 30379
rect 22455 30336 22461 30370
rect 22461 30336 22495 30370
rect 22495 30336 22507 30370
rect 22455 30327 22507 30336
rect 22521 30370 22573 30379
rect 22521 30336 22533 30370
rect 22533 30336 22567 30370
rect 22567 30336 22573 30370
rect 22521 30327 22573 30336
rect 14642 30273 14694 30325
rect 14709 30273 14761 30325
rect 14776 30273 14828 30325
rect 14843 30273 14895 30325
rect 14910 30273 14962 30325
rect 14977 30273 15029 30325
rect 15044 30273 15096 30325
rect 15111 30273 15163 30325
rect 15178 30273 15230 30325
rect 15245 30273 15297 30325
rect 15312 30273 15364 30325
rect 15378 30273 15430 30325
rect 15444 30273 15496 30325
rect 15510 30273 15562 30325
rect 15576 30273 15628 30325
rect 21391 30149 21443 30201
rect 21473 30149 21525 30201
rect 21554 30149 21606 30201
rect 21635 30149 21687 30201
rect 21391 30077 21443 30129
rect 21473 30077 21525 30129
rect 21554 30077 21606 30129
rect 21635 30077 21687 30129
rect 21391 30005 21443 30057
rect 21473 30005 21525 30057
rect 21554 30005 21606 30057
rect 21635 30005 21687 30057
rect 20379 29928 20431 29934
rect 20379 29894 20385 29928
rect 20385 29894 20419 29928
rect 20419 29894 20431 29928
rect 20379 29882 20431 29894
rect 20449 29928 20501 29934
rect 20519 29928 20571 29934
rect 20449 29894 20493 29928
rect 20493 29894 20501 29928
rect 20519 29894 20527 29928
rect 20527 29894 20571 29928
rect 20449 29882 20501 29894
rect 20519 29882 20571 29894
rect 20588 29928 20640 29934
rect 20588 29894 20600 29928
rect 20600 29894 20634 29928
rect 20634 29894 20640 29928
rect 20588 29882 20640 29894
rect 23264 25079 23316 25131
rect 23264 25015 23316 25067
rect 23184 24585 23236 24637
rect 23184 24521 23236 24573
rect 23445 30179 23497 30231
rect 23445 30115 23497 30167
rect 23525 30688 23577 30740
rect 23525 30624 23577 30676
rect 23443 29785 23495 29837
rect 23443 29703 23495 29755
rect 23443 28432 23495 28484
rect 23443 28350 23495 28402
rect 23361 23289 23413 23341
rect 23361 23225 23413 23277
rect 23445 24011 23497 24063
rect 23445 23947 23497 23999
rect 23125 20607 23177 20659
rect 23125 20543 23177 20595
rect 23525 22938 23577 22990
rect 23525 22874 23577 22926
rect 23605 30688 23657 30740
rect 23605 30624 23657 30676
rect 23525 22772 23577 22824
rect 23525 22708 23577 22760
rect 23445 21943 23497 21995
rect 23445 21879 23497 21931
rect 23365 20770 23417 20822
rect 23365 20706 23417 20758
rect 23285 20056 23337 20108
rect 23285 19966 23337 20018
rect 23685 30711 23737 30763
rect 23685 30647 23737 30699
rect 23685 23455 23737 23507
rect 23685 23391 23737 23443
rect 23773 30743 23825 30795
rect 23837 30743 23889 30795
rect 26420 30752 26472 30804
rect 23605 22365 23657 22417
rect 23605 22301 23657 22353
rect 23685 23289 23737 23341
rect 23685 23225 23737 23277
rect 23860 30580 23912 30632
rect 23932 30580 23984 30632
rect 23860 30508 23912 30560
rect 23932 30508 23984 30560
rect 23860 30436 23912 30488
rect 23932 30436 23984 30488
rect 24024 30535 24076 30587
rect 24094 30535 24146 30587
rect 24164 30535 24216 30587
rect 24234 30535 24286 30587
rect 24304 30535 24356 30587
rect 24374 30535 24426 30587
rect 24444 30535 24496 30587
rect 24514 30535 24566 30587
rect 24584 30535 24636 30587
rect 24024 30471 24076 30523
rect 24094 30471 24146 30523
rect 24164 30471 24216 30523
rect 24234 30471 24286 30523
rect 24304 30471 24356 30523
rect 24374 30471 24426 30523
rect 24444 30471 24496 30523
rect 24514 30471 24566 30523
rect 24584 30471 24636 30523
rect 24024 30407 24076 30459
rect 24094 30407 24146 30459
rect 24164 30407 24216 30459
rect 24234 30407 24286 30459
rect 24304 30407 24356 30459
rect 24374 30407 24426 30459
rect 24444 30407 24496 30459
rect 24514 30407 24566 30459
rect 24584 30407 24636 30459
rect 24024 30343 24076 30395
rect 24094 30343 24146 30395
rect 24164 30343 24216 30395
rect 24234 30343 24286 30395
rect 24304 30343 24356 30395
rect 24374 30343 24426 30395
rect 24444 30343 24496 30395
rect 24514 30343 24566 30395
rect 24584 30343 24636 30395
rect 26862 30567 26914 30619
rect 26936 30567 26988 30619
rect 27010 30567 27062 30619
rect 26862 30495 26914 30547
rect 26936 30495 26988 30547
rect 27010 30495 27062 30547
rect 26862 30423 26914 30475
rect 26936 30423 26988 30475
rect 27010 30423 27062 30475
rect 26862 30350 26914 30402
rect 26936 30350 26988 30402
rect 27010 30350 27062 30402
rect 27973 30651 28025 30703
rect 27576 30567 27628 30619
rect 27650 30567 27702 30619
rect 27724 30567 27776 30619
rect 27576 30495 27628 30547
rect 27650 30495 27702 30547
rect 27724 30495 27776 30547
rect 27576 30422 27628 30474
rect 27650 30422 27702 30474
rect 27724 30422 27776 30474
rect 27576 30349 27628 30401
rect 27650 30349 27702 30401
rect 27724 30349 27776 30401
rect 27973 30571 28025 30623
rect 27973 30491 28025 30543
rect 27973 30411 28025 30463
rect 27313 29969 27365 30021
rect 27313 29905 27365 29957
rect 24185 28085 24237 28137
rect 24259 28085 24311 28137
rect 24333 28085 24385 28137
rect 24185 28015 24237 28067
rect 24259 28015 24311 28067
rect 24333 28015 24385 28067
rect 24185 27945 24237 27997
rect 24259 27945 24311 27997
rect 24333 27945 24385 27997
rect 24185 27875 24237 27927
rect 24259 27875 24311 27927
rect 24333 27875 24385 27927
rect 24185 27805 24237 27857
rect 24259 27805 24311 27857
rect 24333 27805 24385 27857
rect 24185 27734 24237 27786
rect 24259 27734 24311 27786
rect 24333 27734 24385 27786
rect 24185 27663 24237 27715
rect 24259 27663 24311 27715
rect 24333 27663 24385 27715
rect 25307 28085 25359 28137
rect 25385 28085 25437 28137
rect 25307 28001 25359 28053
rect 25385 28001 25437 28053
rect 25307 27917 25359 27969
rect 25385 27917 25437 27969
rect 25307 27832 25359 27884
rect 25385 27832 25437 27884
rect 25307 27747 25359 27799
rect 25385 27747 25437 27799
rect 25307 27662 25359 27714
rect 25385 27662 25437 27714
rect 25923 28085 25975 28137
rect 26001 28085 26053 28137
rect 25923 28001 25975 28053
rect 26001 28001 26053 28053
rect 25923 27917 25975 27969
rect 26001 27917 26053 27969
rect 25923 27832 25975 27884
rect 26001 27832 26053 27884
rect 25923 27747 25975 27799
rect 26001 27747 26053 27799
rect 25923 27662 25975 27714
rect 26001 27662 26053 27714
rect 26336 28085 26388 28137
rect 26410 28085 26462 28137
rect 26484 28085 26536 28137
rect 26336 28015 26388 28067
rect 26410 28015 26462 28067
rect 26484 28015 26536 28067
rect 26336 27945 26388 27997
rect 26410 27945 26462 27997
rect 26484 27945 26536 27997
rect 26336 27875 26388 27927
rect 26410 27875 26462 27927
rect 26484 27875 26536 27927
rect 26336 27804 26388 27856
rect 26410 27804 26462 27856
rect 26484 27804 26536 27856
rect 26336 27733 26388 27785
rect 26410 27733 26462 27785
rect 26484 27733 26536 27785
rect 26336 27662 26388 27714
rect 26410 27662 26462 27714
rect 26484 27662 26536 27714
rect 24185 26739 24237 26791
rect 24259 26739 24311 26791
rect 24333 26739 24385 26791
rect 24185 26669 24237 26721
rect 24259 26669 24311 26721
rect 24333 26669 24385 26721
rect 24185 26599 24237 26651
rect 24259 26599 24311 26651
rect 24333 26599 24385 26651
rect 24185 26529 24237 26581
rect 24259 26529 24311 26581
rect 24333 26529 24385 26581
rect 24185 26458 24237 26510
rect 24259 26458 24311 26510
rect 24333 26458 24385 26510
rect 24185 26387 24237 26439
rect 24259 26387 24311 26439
rect 24333 26387 24385 26439
rect 24185 26316 24237 26368
rect 24259 26316 24311 26368
rect 24333 26316 24385 26368
rect 25413 26739 25465 26791
rect 25491 26739 25543 26791
rect 25413 26655 25465 26707
rect 25491 26655 25543 26707
rect 25413 26571 25465 26623
rect 25491 26571 25543 26623
rect 25413 26486 25465 26538
rect 25491 26486 25543 26538
rect 25413 26401 25465 26453
rect 25491 26401 25543 26453
rect 25413 26316 25465 26368
rect 25491 26316 25543 26368
rect 25923 26739 25975 26791
rect 26001 26739 26053 26791
rect 25923 26655 25975 26707
rect 26001 26655 26053 26707
rect 25923 26571 25975 26623
rect 26001 26571 26053 26623
rect 25923 26486 25975 26538
rect 26001 26486 26053 26538
rect 25923 26401 25975 26453
rect 26001 26401 26053 26453
rect 25923 26316 25975 26368
rect 26001 26316 26053 26368
rect 26336 26739 26388 26791
rect 26410 26739 26462 26791
rect 26484 26739 26536 26791
rect 26336 26669 26388 26721
rect 26410 26669 26462 26721
rect 26484 26669 26536 26721
rect 26336 26599 26388 26651
rect 26410 26599 26462 26651
rect 26484 26599 26536 26651
rect 26336 26529 26388 26581
rect 26410 26529 26462 26581
rect 26484 26529 26536 26581
rect 26336 26458 26388 26510
rect 26410 26458 26462 26510
rect 26484 26458 26536 26510
rect 26336 26387 26388 26439
rect 26410 26387 26462 26439
rect 26484 26387 26536 26439
rect 26336 26316 26388 26368
rect 26410 26316 26462 26368
rect 26484 26316 26536 26368
rect 27171 24011 27223 24063
rect 27171 23947 27223 23999
rect 25663 23437 25715 23489
rect 25727 23437 25779 23489
rect 26707 23084 26759 23136
rect 26707 23020 26759 23072
rect 27283 22761 27335 22813
rect 27283 22697 27335 22749
rect 26633 22376 26685 22428
rect 26633 22312 26685 22364
rect 24185 22211 24237 22263
rect 24259 22211 24311 22263
rect 24333 22211 24385 22263
rect 24185 22146 24237 22198
rect 24259 22146 24311 22198
rect 24333 22146 24385 22198
rect 24185 22081 24237 22133
rect 24259 22081 24311 22133
rect 24333 22081 24385 22133
rect 24185 22015 24237 22067
rect 24259 22015 24311 22067
rect 24333 22015 24385 22067
rect 25307 22211 25359 22263
rect 25385 22211 25437 22263
rect 25307 22113 25359 22165
rect 25385 22113 25437 22165
rect 25307 22015 25359 22067
rect 25385 22015 25437 22067
rect 25923 22211 25975 22263
rect 26001 22211 26053 22263
rect 25923 22113 25975 22165
rect 26001 22113 26053 22165
rect 25923 22015 25975 22067
rect 26001 22015 26053 22067
rect 26336 22211 26388 22263
rect 26410 22211 26462 22263
rect 26484 22211 26536 22263
rect 26336 22146 26388 22198
rect 26410 22146 26462 22198
rect 26484 22146 26536 22198
rect 26336 22081 26388 22133
rect 26410 22081 26462 22133
rect 26484 22081 26536 22133
rect 26336 22015 26388 22067
rect 26410 22015 26462 22067
rect 26484 22015 26536 22067
rect 27283 21932 27335 21984
rect 27283 21868 27335 21920
rect 27247 20990 27299 21042
rect 23759 20930 23811 20982
rect 23759 20866 23811 20918
rect 25465 20909 25517 20961
rect 27247 20926 27299 20978
rect 25465 20845 25517 20897
rect 27495 20789 27547 20841
rect 27495 20725 27547 20777
rect 24185 18219 24237 18271
rect 24259 18219 24311 18271
rect 24333 18219 24385 18271
rect 24185 18154 24237 18206
rect 24259 18154 24311 18206
rect 24333 18154 24385 18206
rect 24185 18089 24237 18141
rect 24259 18089 24311 18141
rect 24333 18089 24385 18141
rect 24185 18023 24237 18075
rect 24259 18023 24311 18075
rect 24333 18023 24385 18075
rect 25307 18219 25359 18271
rect 25385 18219 25437 18271
rect 25307 18121 25359 18173
rect 25385 18121 25437 18173
rect 25307 18023 25359 18075
rect 25385 18023 25437 18075
rect 25923 18219 25975 18271
rect 26001 18219 26053 18271
rect 25923 18121 25975 18173
rect 26001 18121 26053 18173
rect 25923 18023 25975 18075
rect 26001 18023 26053 18075
rect 26336 18219 26388 18271
rect 26410 18219 26462 18271
rect 26484 18219 26536 18271
rect 26336 18154 26388 18206
rect 26410 18154 26462 18206
rect 26484 18154 26536 18206
rect 26336 18089 26388 18141
rect 26410 18089 26462 18141
rect 26484 18089 26536 18141
rect 26336 18023 26388 18075
rect 26410 18023 26462 18075
rect 26484 18023 26536 18075
rect 23269 2081 23321 2133
rect 23333 2081 23385 2133
rect 23269 1967 23321 2019
rect 23333 1967 23385 2019
rect 25770 1875 25822 1927
rect 25836 1875 25888 1927
rect 25144 1648 25196 1700
rect 25208 1648 25260 1700
rect 26863 1525 26915 1577
rect 26927 1525 26979 1577
rect 27049 1368 27101 1420
rect 27122 1368 27174 1420
rect 27195 1368 27247 1420
rect 27268 1368 27320 1420
rect 27341 1368 27393 1420
rect 27413 1368 27465 1420
rect 27485 1368 27537 1420
rect 27049 1294 27101 1346
rect 27122 1294 27174 1346
rect 27195 1294 27247 1346
rect 27268 1294 27320 1346
rect 27341 1294 27393 1346
rect 27413 1294 27465 1346
rect 27485 1294 27537 1346
rect 27049 1220 27101 1272
rect 27122 1220 27174 1272
rect 27195 1220 27247 1272
rect 27268 1220 27320 1272
rect 27341 1220 27393 1272
rect 27413 1220 27465 1272
rect 27485 1220 27537 1272
rect 23254 1115 23306 1167
rect 23320 1115 23372 1167
rect 24138 1073 24190 1125
rect 25511 1115 25563 1167
rect 25575 1115 25627 1167
rect 25770 1158 25822 1167
rect 25770 1124 25776 1158
rect 25776 1124 25810 1158
rect 25810 1124 25822 1158
rect 25770 1115 25822 1124
rect 25836 1158 25888 1167
rect 25836 1124 25848 1158
rect 25848 1124 25882 1158
rect 25882 1124 25888 1158
rect 25836 1115 25888 1124
rect 27319 1163 27371 1167
rect 27319 1129 27322 1163
rect 27322 1129 27356 1163
rect 27356 1129 27371 1163
rect 27319 1115 27371 1129
rect 27383 1163 27435 1167
rect 27383 1129 27394 1163
rect 27394 1129 27428 1163
rect 27428 1129 27435 1163
rect 27383 1115 27435 1129
rect 24138 1009 24190 1061
rect 23254 790 23306 842
rect 23320 790 23372 842
rect 24681 861 24733 913
rect 24681 797 24733 849
rect 27092 1060 27144 1072
rect 27092 1026 27098 1060
rect 27098 1026 27132 1060
rect 27132 1026 27144 1060
rect 27092 1020 27144 1026
rect 27156 1060 27208 1072
rect 27156 1026 27170 1060
rect 27170 1026 27204 1060
rect 27204 1026 27208 1060
rect 27156 1020 27208 1026
rect 23953 626 24005 678
rect 24018 626 24070 678
rect 25377 632 25429 684
rect 25441 632 25493 684
rect 23953 562 24005 614
rect 24018 562 24070 614
rect 27049 378 27101 430
rect 27158 378 27210 430
rect 27267 378 27319 430
rect 27376 378 27428 430
rect 27485 378 27537 430
rect 27049 300 27101 352
rect 27158 300 27210 352
rect 27267 300 27319 352
rect 27376 300 27428 352
rect 27485 300 27537 352
rect 25883 32 25935 41
rect 25883 -2 25889 32
rect 25889 -2 25923 32
rect 25923 -2 25935 32
rect 25883 -11 25935 -2
rect 25949 32 26001 41
rect 25949 -2 25961 32
rect 25961 -2 25995 32
rect 25995 -2 26001 32
rect 25949 -11 26001 -2
<< metal2 >>
rect 13706 33704 14081 33705
rect 13706 33652 13712 33704
rect 13764 33652 13790 33704
rect 13842 33652 13868 33704
rect 13920 33652 13946 33704
rect 13998 33652 14023 33704
rect 14075 33652 14081 33704
rect 13706 33636 14081 33652
rect 13706 33584 13712 33636
rect 13764 33584 13790 33636
rect 13842 33584 13868 33636
rect 13920 33584 13946 33636
rect 13998 33584 14023 33636
rect 14075 33584 14081 33636
rect 13706 33568 14081 33584
rect 13706 33516 13712 33568
rect 13764 33516 13790 33568
rect 13842 33516 13868 33568
rect 13920 33516 13946 33568
rect 13998 33516 14023 33568
rect 14075 33516 14081 33568
rect 13706 33500 14081 33516
rect 13706 33448 13712 33500
rect 13764 33448 13790 33500
rect 13842 33448 13868 33500
rect 13920 33448 13946 33500
rect 13998 33448 14023 33500
rect 14075 33448 14081 33500
rect 19975 33592 20911 33705
tri 20911 33592 21024 33705 sw
rect 19975 33591 21024 33592
tri 21024 33591 21025 33592 sw
rect 21383 33591 21695 33592
rect 19975 33539 21025 33591
tri 21025 33539 21077 33591 sw
rect 21383 33539 21391 33591
rect 21443 33539 21473 33591
rect 21525 33539 21555 33591
rect 21607 33539 21636 33591
rect 21688 33539 21695 33591
rect 19975 33527 21077 33539
tri 21077 33527 21089 33539 sw
rect 21383 33527 21695 33539
rect 19975 33475 21089 33527
tri 21089 33475 21141 33527 sw
rect 21383 33475 21391 33527
rect 21443 33475 21473 33527
rect 21525 33475 21555 33527
rect 21607 33475 21636 33527
rect 21688 33475 21695 33527
rect 19975 33471 21141 33475
tri 21141 33471 21145 33475 sw
rect 19975 33463 21145 33471
tri 21145 33463 21153 33471 sw
rect 21383 33463 21695 33475
rect 19975 33462 21153 33463
rect 13706 33447 14081 33448
tri 20712 33447 20727 33462 ne
rect 20727 33447 21153 33462
tri 21153 33447 21169 33463 sw
tri 20727 33411 20763 33447 ne
rect 20763 33411 21169 33447
tri 21169 33411 21205 33447 sw
rect 21383 33411 21391 33463
rect 21443 33411 21473 33463
rect 21525 33411 21555 33463
rect 21607 33411 21636 33463
rect 21688 33411 21695 33463
tri 20763 33399 20775 33411 ne
rect 20775 33399 21205 33411
tri 21205 33399 21217 33411 sw
rect 21383 33399 21695 33411
tri 20775 33347 20827 33399 ne
rect 20827 33347 21217 33399
tri 21217 33347 21269 33399 sw
rect 21383 33347 21391 33399
rect 21443 33347 21473 33399
rect 21525 33347 21555 33399
rect 21607 33347 21636 33399
rect 21688 33347 21695 33399
tri 20827 33339 20835 33347 ne
rect 20835 33339 21269 33347
tri 21269 33339 21277 33347 sw
tri 20835 33327 20847 33339 ne
rect 20847 33327 21277 33339
tri 21277 33327 21289 33339 sw
rect 18962 33322 18991 33327
tri 18991 33322 18996 33327 nw
tri 20847 33326 20848 33327 ne
rect 20848 33326 21289 33327
tri 21289 33326 21290 33327 sw
tri 20848 33322 20852 33326 ne
rect 20852 33322 21290 33326
tri 18962 33293 18991 33322 nw
tri 20852 33293 20881 33322 ne
rect 20881 33293 21290 33322
tri 20881 33270 20904 33293 ne
rect 20904 33270 21290 33293
tri 20904 33263 20911 33270 ne
rect 20911 33263 21290 33270
tri 20911 33258 20916 33263 ne
rect 20916 33258 21290 33263
tri 20916 33220 20954 33258 ne
rect 20954 33220 21290 33258
tri 20954 33196 20978 33220 ne
rect 13454 33014 13460 33066
rect 13512 33014 13524 33066
rect 13576 33014 13582 33066
tri 13442 32123 13454 32135 se
rect 13454 32123 13582 33014
rect 20165 33043 20217 33051
rect 20165 32979 20217 32991
rect 18046 32832 18098 32838
rect 19210 32825 19262 32831
rect 18046 32768 18098 32780
tri 18219 32773 18228 32782 se
rect 18228 32773 18283 32820
tri 18207 32761 18219 32773 se
rect 18219 32761 18283 32773
rect 14636 32499 15638 32500
rect 14636 32447 14643 32499
rect 14695 32447 14710 32499
rect 14762 32447 14777 32499
rect 14829 32447 14844 32499
rect 14896 32447 14911 32499
rect 14963 32447 14978 32499
rect 15030 32447 15045 32499
rect 15097 32447 15112 32499
rect 15164 32447 15179 32499
rect 15231 32447 15246 32499
rect 15298 32447 15313 32499
rect 15365 32447 15379 32499
rect 15431 32447 15445 32499
rect 15497 32447 15511 32499
rect 15563 32447 15577 32499
rect 15629 32447 15638 32499
rect 14636 32427 15638 32447
rect 14636 32375 14643 32427
rect 14695 32375 14710 32427
rect 14762 32375 14777 32427
rect 14829 32375 14844 32427
rect 14896 32375 14911 32427
rect 14963 32375 14978 32427
rect 15030 32375 15045 32427
rect 15097 32375 15112 32427
rect 15164 32375 15179 32427
rect 15231 32375 15246 32427
rect 15298 32375 15313 32427
rect 15365 32375 15379 32427
rect 15431 32375 15445 32427
rect 15497 32375 15511 32427
rect 15563 32375 15577 32427
rect 15629 32375 15638 32427
rect 14636 32355 15638 32375
rect 14636 32303 14643 32355
rect 14695 32303 14710 32355
rect 14762 32303 14777 32355
rect 14829 32303 14844 32355
rect 14896 32303 14911 32355
rect 14963 32303 14978 32355
rect 15030 32303 15045 32355
rect 15097 32303 15112 32355
rect 15164 32303 15179 32355
rect 15231 32303 15246 32355
rect 15298 32303 15313 32355
rect 15365 32303 15379 32355
rect 15431 32303 15445 32355
rect 15497 32303 15511 32355
rect 15563 32303 15577 32355
rect 15629 32303 15638 32355
tri 13582 32123 13596 32137 sw
rect 13442 32067 13451 32123
rect 13507 32067 13531 32123
rect 13587 32067 13596 32123
rect 3608 31960 3664 31969
tri 3589 31924 3608 31943 se
tri 3573 31908 3589 31924 se
rect 3589 31908 3608 31924
rect 3608 31880 3664 31904
rect 3608 31815 3664 31824
rect 2161 31730 3838 31745
rect 2161 31674 2170 31730
rect 2226 31674 2250 31730
rect 2306 31722 3838 31730
rect 2306 31674 3693 31722
rect 2161 31666 3693 31674
rect 3749 31666 3773 31722
rect 3829 31666 3838 31722
rect 2161 31651 3838 31666
rect 3899 31655 3955 31664
tri 3879 31619 3899 31639 se
tri 3876 31616 3879 31619 se
rect 3879 31616 3899 31619
tri 3864 31604 3876 31616 se
rect 3876 31604 3899 31616
rect 2165 31599 3899 31604
rect 2165 31593 3955 31599
rect 2165 31537 2174 31593
rect 2230 31537 2254 31593
rect 2310 31575 3955 31593
rect 2310 31537 3899 31575
rect 2165 31519 3899 31537
rect 2165 31510 3955 31519
rect 14636 31573 15638 32303
tri 18026 31986 18046 32006 se
rect 18046 31986 18098 32716
tri 18199 32753 18207 32761 se
rect 18207 32753 18283 32761
rect 18199 32697 18283 32753
rect 19210 32761 19262 32773
tri 18199 32692 18204 32697 ne
rect 18204 32692 18283 32697
rect 18533 32688 18539 32740
rect 18591 32688 18603 32740
rect 18655 32688 18661 32740
rect 18533 32249 18661 32688
rect 19210 32668 19262 32709
tri 19262 32668 19264 32670 sw
rect 19210 32648 19264 32668
tri 19210 32646 19212 32648 ne
rect 19212 32646 19264 32648
tri 19264 32646 19286 32668 sw
tri 19212 32596 19262 32646 ne
rect 19262 32596 19286 32646
tri 19286 32596 19336 32646 sw
tri 19262 32594 19264 32596 ne
rect 19264 32594 19336 32596
tri 19336 32594 19338 32596 sw
tri 19264 32584 19274 32594 ne
rect 19274 32584 19338 32594
tri 19338 32584 19348 32594 sw
tri 19274 32572 19286 32584 ne
rect 19286 32572 19348 32584
tri 19348 32572 19360 32584 sw
tri 19286 32522 19336 32572 ne
rect 19336 32522 19360 32572
tri 19360 32522 19410 32572 sw
rect 19704 32564 19713 32620
rect 19769 32564 19811 32620
rect 19867 32564 19910 32620
rect 19966 32564 19975 32620
tri 19336 32520 19338 32522 ne
rect 19338 32520 19410 32522
tri 19410 32520 19412 32522 sw
tri 19338 32519 19339 32520 ne
rect 19339 32519 19412 32520
tri 19412 32519 19413 32520 sw
tri 19339 32508 19350 32519 ne
rect 19350 32501 19413 32519
tri 19413 32501 19431 32519 sw
rect 19704 32516 19975 32564
rect 19350 32445 19359 32501
rect 19415 32445 19439 32501
rect 19495 32445 19504 32501
rect 19704 32460 19713 32516
rect 19769 32460 19811 32516
rect 19867 32460 19910 32516
rect 19966 32460 19975 32516
rect 18511 32193 18520 32249
rect 18576 32193 18600 32249
rect 18656 32193 18665 32249
rect 19048 32211 19054 32263
rect 19106 32211 19118 32263
rect 19170 32211 19176 32263
rect 18533 32187 18661 32193
tri 18002 31962 18026 31986 se
rect 18026 31976 18098 31986
rect 18026 31962 18084 31976
tri 18084 31962 18098 31976 nw
tri 17964 31924 18002 31962 se
rect 18002 31924 18046 31962
tri 18046 31924 18084 31962 nw
rect 14636 31517 14888 31573
rect 14944 31517 14970 31573
rect 15026 31517 15052 31573
rect 15108 31517 15134 31573
rect 15190 31517 15216 31573
rect 15272 31517 15298 31573
rect 15354 31517 15380 31573
rect 15436 31517 15638 31573
tri 4017 31483 4025 31491 se
rect 4025 31485 4081 31494
tri 3990 31456 4017 31483 se
rect 4017 31456 4025 31483
rect 2166 31400 2176 31456
rect 2232 31400 2256 31456
rect 2312 31429 4025 31456
rect 2312 31405 4081 31429
rect 2312 31400 4025 31405
rect 1971 31366 2027 31375
rect 2166 31356 4025 31400
tri 4009 31340 4025 31356 ne
rect 4025 31340 4081 31349
rect 14636 31492 15638 31517
rect 14636 31436 14888 31492
rect 14944 31436 14970 31492
rect 15026 31436 15052 31492
rect 15108 31436 15134 31492
rect 15190 31436 15216 31492
rect 15272 31436 15298 31492
rect 15354 31436 15380 31492
rect 15436 31436 15638 31492
rect 14636 31411 15638 31436
rect 14636 31355 14888 31411
rect 14944 31355 14970 31411
rect 15026 31355 15052 31411
rect 15108 31355 15134 31411
rect 15190 31355 15216 31411
rect 15272 31355 15298 31411
rect 15354 31355 15380 31411
rect 15436 31355 15638 31411
tri 2027 31325 2039 31337 sw
rect 14636 31330 15638 31355
rect 2027 31310 2039 31325
rect 1971 31295 2039 31310
tri 2039 31295 2069 31325 sw
rect 1971 31294 2069 31295
tri 2069 31294 2070 31295 sw
rect 1971 31286 4207 31294
rect 2027 31285 4207 31286
rect 2027 31230 4151 31285
rect 1971 31229 4151 31230
rect 1971 31221 4207 31229
tri 2741 31193 2769 31221 ne
rect 2769 31205 4207 31221
rect 2769 31193 4151 31205
tri 2769 31188 2774 31193 ne
rect 2774 31188 4151 31193
tri 2774 31176 2786 31188 ne
rect 2786 31176 4151 31188
tri 2786 31140 2822 31176 ne
rect 2822 31149 4151 31176
rect 2822 31140 4207 31149
rect 14636 31274 14888 31330
rect 14944 31274 14970 31330
rect 15026 31274 15052 31330
rect 15108 31274 15134 31330
rect 15190 31274 15216 31330
rect 15272 31274 15298 31330
rect 15354 31274 15380 31330
rect 15436 31274 15638 31330
rect 14636 31249 15638 31274
rect 14636 31193 14888 31249
rect 14944 31193 14970 31249
rect 15026 31193 15052 31249
rect 15108 31193 15134 31249
rect 15190 31193 15216 31249
rect 15272 31193 15298 31249
rect 15354 31193 15380 31249
rect 15436 31193 15638 31249
tri 17927 31887 17964 31924 se
rect 17964 31887 18009 31924
tri 18009 31887 18046 31924 nw
rect 17927 31872 17994 31887
tri 17994 31872 18009 31887 nw
rect 17927 31245 17979 31872
tri 17979 31857 17994 31872 nw
rect 19048 31738 19092 32211
tri 19092 32182 19121 32211 nw
rect 19329 31947 19975 31954
rect 19329 31924 19360 31947
rect 19416 31924 19468 31947
rect 19524 31924 19575 31947
rect 19631 31924 19682 31947
rect 19738 31924 19789 31947
rect 19329 31872 19337 31924
rect 19389 31872 19402 31891
rect 19454 31872 19467 31924
rect 19524 31891 19532 31924
rect 19519 31872 19532 31891
rect 19584 31872 19597 31891
rect 19649 31872 19662 31924
rect 19778 31891 19789 31924
rect 19845 31891 19896 31947
rect 19952 31891 19975 31947
rect 19714 31872 19726 31891
rect 19778 31872 19790 31891
rect 19842 31872 19975 31891
rect 19329 31852 19975 31872
rect 19329 31800 19337 31852
rect 19389 31800 19402 31852
rect 19454 31800 19467 31852
rect 19519 31800 19532 31852
rect 19584 31800 19597 31852
rect 19649 31800 19662 31852
rect 19714 31800 19726 31852
rect 19778 31800 19790 31852
rect 19842 31800 19975 31852
rect 19329 31789 19975 31800
rect 19329 31780 19360 31789
rect 19416 31780 19468 31789
rect 19524 31780 19575 31789
rect 19631 31780 19682 31789
rect 19738 31780 19789 31789
tri 19048 31728 19058 31738 ne
rect 19058 31728 19092 31738
tri 19092 31728 19135 31771 sw
tri 19058 31695 19091 31728 ne
tri 18380 31483 18397 31500 se
tri 18363 31466 18380 31483 se
rect 18380 31466 18397 31483
tri 18463 31495 18468 31500 sw
rect 18463 31483 18468 31495
tri 18468 31483 18480 31495 sw
tri 19079 31483 19091 31495 se
rect 19091 31483 19135 31728
rect 19329 31728 19337 31780
rect 19389 31728 19402 31733
rect 19454 31728 19467 31780
rect 19524 31733 19532 31780
rect 19519 31728 19532 31733
rect 19584 31728 19597 31733
rect 19649 31728 19662 31780
rect 19778 31733 19789 31780
rect 19845 31733 19896 31789
rect 19952 31733 19975 31789
rect 19714 31728 19726 31733
rect 19778 31728 19790 31733
rect 19842 31728 19975 31733
rect 19329 31724 19975 31728
rect 18463 31466 18480 31483
tri 18480 31466 18497 31483 sw
tri 19062 31466 19079 31483 se
rect 19079 31466 19135 31483
tri 19058 31462 19062 31466 se
rect 19062 31462 19135 31466
tri 19048 31452 19058 31462 se
rect 19058 31452 19114 31462
rect 19048 31441 19114 31452
tri 19114 31441 19135 31462 nw
tri 17979 31245 18014 31280 sw
rect 17900 31193 17906 31245
rect 17958 31193 17970 31245
rect 18022 31193 18028 31245
rect 14636 31168 15638 31193
rect 14636 31112 14888 31168
rect 14944 31112 14970 31168
rect 15026 31112 15052 31168
rect 15108 31112 15134 31168
rect 15190 31112 15216 31168
rect 15272 31112 15298 31168
rect 15354 31112 15380 31168
rect 15436 31112 15638 31168
rect 14636 31087 15638 31112
rect 14636 31031 14888 31087
rect 14944 31031 14970 31087
rect 15026 31031 15052 31087
rect 15108 31031 15134 31087
rect 15190 31031 15216 31087
rect 15272 31031 15298 31087
rect 15354 31031 15380 31087
rect 15436 31031 15638 31087
rect 14636 31006 15638 31031
rect 14636 30950 14888 31006
rect 14944 30950 14970 31006
rect 15026 30950 15052 31006
rect 15108 30950 15134 31006
rect 15190 30950 15216 31006
rect 15272 30950 15298 31006
rect 15354 30950 15380 31006
rect 15436 30950 15638 31006
rect 14636 30924 15638 30950
rect 14636 30868 14888 30924
rect 14944 30868 14970 30924
rect 15026 30868 15052 30924
rect 15108 30868 15134 30924
rect 15190 30868 15216 30924
rect 15272 30868 15298 30924
rect 15354 30868 15380 30924
rect 15436 30868 15638 30924
rect 14636 30842 15638 30868
rect 14636 30786 14888 30842
rect 14944 30786 14970 30842
rect 15026 30786 15052 30842
rect 15108 30786 15134 30842
rect 15190 30786 15216 30842
rect 15272 30786 15298 30842
rect 15354 30786 15380 30842
rect 15436 30786 15638 30842
rect 14636 30760 15638 30786
rect 14636 30704 14888 30760
rect 14944 30704 14970 30760
rect 15026 30704 15052 30760
rect 15108 30704 15134 30760
rect 15190 30704 15216 30760
rect 15272 30704 15298 30760
rect 15354 30704 15380 30760
rect 15436 30704 15638 30760
rect 14636 30678 15638 30704
rect 14636 30622 14888 30678
rect 14944 30622 14970 30678
rect 15026 30622 15052 30678
rect 15108 30622 15134 30678
rect 15190 30622 15216 30678
rect 15272 30622 15298 30678
rect 15354 30622 15380 30678
rect 15436 30622 15638 30678
rect 19048 30715 19092 31441
tri 19092 31419 19114 31441 nw
tri 20162 31282 20165 31285 se
rect 20165 31282 20217 32927
rect 20978 32720 21290 33220
rect 20978 32668 20980 32720
rect 21032 32668 21064 32720
rect 21116 32668 21148 32720
rect 21200 32668 21232 32720
rect 21284 32668 21290 32720
rect 20978 32646 21290 32668
rect 20978 32594 20980 32646
rect 21032 32620 21064 32646
rect 21116 32620 21148 32646
rect 21200 32620 21232 32646
rect 21043 32594 21064 32620
rect 21200 32594 21225 32620
rect 21284 32594 21290 32646
rect 20978 32572 20987 32594
rect 21043 32572 21106 32594
rect 21162 32572 21225 32594
rect 21281 32572 21290 32594
rect 20978 32520 20980 32572
rect 21043 32564 21064 32572
rect 21200 32564 21225 32572
rect 21032 32520 21064 32564
rect 21116 32520 21148 32564
rect 21200 32520 21232 32564
rect 21284 32520 21290 32572
rect 20978 32516 21290 32520
rect 20978 32498 20987 32516
rect 21043 32498 21106 32516
rect 21162 32498 21225 32516
rect 21281 32498 21290 32516
rect 20978 32446 20980 32498
rect 21043 32460 21064 32498
rect 21200 32460 21225 32498
rect 21032 32446 21064 32460
rect 21116 32446 21148 32460
rect 21200 32446 21232 32460
rect 21284 32446 21290 32498
rect 20978 32423 21290 32446
rect 20978 32371 20980 32423
rect 21032 32371 21064 32423
rect 21116 32371 21148 32423
rect 21200 32371 21232 32423
rect 21284 32371 21290 32423
tri 20715 31441 20732 31458 se
rect 20732 31441 20784 32185
rect 20978 31964 21290 32371
rect 21034 31908 21106 31964
rect 21162 31908 21234 31964
rect 20978 31854 21290 31908
rect 21034 31798 21106 31854
rect 21162 31798 21234 31854
rect 20978 31743 21290 31798
rect 21034 31687 21106 31743
rect 21162 31687 21234 31743
rect 20978 31632 21290 31687
rect 21034 31576 21106 31632
rect 21162 31576 21234 31632
tri 20784 31441 20809 31466 sw
rect 20715 31389 20721 31441
rect 20773 31389 20785 31441
rect 20837 31389 20843 31441
tri 20125 31245 20162 31282 se
rect 20162 31245 20217 31282
rect 19121 31193 19127 31245
rect 19179 31193 19191 31245
rect 19243 31233 20217 31245
rect 19243 31230 20214 31233
tri 20214 31230 20217 31233 nw
rect 19243 31193 20177 31230
tri 20177 31193 20214 31230 nw
rect 20978 30727 21290 31576
rect 19048 30663 20134 30715
rect 20186 30663 20200 30715
rect 20252 30663 20258 30715
rect 20978 30675 20985 30727
rect 21037 30675 21067 30727
rect 21119 30675 21149 30727
rect 21201 30675 21230 30727
rect 21282 30675 21290 30727
rect 14636 30596 15638 30622
rect 14636 30540 14888 30596
rect 14944 30540 14970 30596
rect 15026 30540 15052 30596
rect 15108 30540 15134 30596
rect 15190 30540 15216 30596
rect 15272 30540 15298 30596
rect 15354 30540 15380 30596
rect 15436 30540 15638 30596
rect 14636 30514 15638 30540
rect 20978 30655 21290 30675
rect 20978 30603 20985 30655
rect 21037 30603 21067 30655
rect 21119 30603 21149 30655
rect 21201 30603 21230 30655
rect 21282 30603 21290 30655
rect 20978 30583 21290 30603
rect 20978 30531 20985 30583
rect 21037 30531 21067 30583
rect 21119 30531 21149 30583
rect 21201 30531 21230 30583
rect 21282 30531 21290 30583
rect 20978 30527 21290 30531
rect 21383 31739 21695 33347
rect 25439 33551 25784 33552
rect 25439 33499 25459 33551
rect 25511 33499 25548 33551
rect 25600 33499 25637 33551
rect 25689 33499 25726 33551
rect 25778 33499 25784 33551
rect 25439 33471 25784 33499
rect 25439 33419 25459 33471
rect 25511 33419 25548 33471
rect 25600 33419 25637 33471
rect 25689 33419 25726 33471
rect 25778 33419 25784 33471
tri 26100 33433 26156 33489 se
rect 26156 33437 26442 33489
rect 26156 33433 26174 33437
tri 26174 33433 26178 33437 nw
tri 26429 33433 26433 33437 ne
rect 26433 33433 26442 33437
rect 26498 33433 26522 33489
rect 26578 33433 26587 33489
rect 26891 33433 26900 33489
rect 26956 33433 26980 33489
rect 27036 33437 27617 33489
rect 27036 33433 27045 33437
tri 27045 33433 27049 33437 nw
tri 27595 33433 27599 33437 ne
rect 27599 33433 27617 33437
tri 26097 33430 26100 33433 se
rect 26100 33430 26171 33433
tri 26171 33430 26174 33433 nw
tri 27599 33430 27602 33433 ne
rect 27602 33430 27617 33433
tri 27617 33430 27676 33489 sw
rect 25439 33391 25784 33419
tri 26082 33415 26097 33430 se
rect 26097 33415 26156 33430
tri 26156 33415 26171 33430 nw
tri 27602 33415 27617 33430 ne
rect 27617 33415 27676 33430
rect 25439 33339 25459 33391
rect 25511 33339 25548 33391
rect 25600 33339 25637 33391
rect 25689 33339 25726 33391
rect 25778 33339 25784 33391
tri 26051 33384 26082 33415 se
rect 26082 33384 26125 33415
tri 26125 33384 26156 33415 nw
tri 27617 33384 27648 33415 ne
rect 27648 33384 27676 33415
tri 27676 33384 27722 33430 sw
tri 26008 33341 26051 33384 se
rect 26051 33341 26082 33384
tri 26082 33341 26125 33384 nw
tri 26266 33341 26309 33384 se
rect 26309 33341 27377 33384
rect 25439 33322 25784 33339
rect 25439 33270 25595 33322
rect 25647 33270 25663 33322
rect 25715 33270 25731 33322
rect 25783 33270 25784 33322
rect 25439 33258 25784 33270
rect 22953 33220 23005 33226
rect 22953 33156 23005 33168
rect 21383 31687 21389 31739
rect 21441 31687 21468 31739
rect 21520 31687 21547 31739
rect 21599 31687 21625 31739
rect 21677 31687 21695 31739
rect 21383 31671 21695 31687
rect 21383 31619 21389 31671
rect 21441 31619 21468 31671
rect 21520 31619 21547 31671
rect 21599 31619 21625 31671
rect 21677 31619 21695 31671
rect 21383 31603 21695 31619
rect 21383 31551 21389 31603
rect 21441 31551 21468 31603
rect 21520 31551 21547 31603
rect 21599 31551 21625 31603
rect 21677 31551 21695 31603
rect 21383 31535 21695 31551
rect 21383 31483 21389 31535
rect 21441 31483 21468 31535
rect 21520 31483 21547 31535
rect 21599 31483 21625 31535
rect 21677 31483 21695 31535
rect 22614 33023 22666 33029
rect 22614 32959 22666 32971
rect 14636 30493 14888 30514
rect 14944 30493 14970 30514
rect 15026 30493 15052 30514
rect 15108 30493 15134 30514
rect 15190 30493 15216 30514
rect 15272 30493 15298 30514
rect 15354 30493 15380 30514
rect 15436 30493 15638 30514
rect 14636 30441 14642 30493
rect 14694 30441 14709 30493
rect 14761 30441 14776 30493
rect 14828 30441 14843 30493
rect 14962 30458 14970 30493
rect 14895 30441 14910 30458
rect 14962 30441 14977 30458
rect 15029 30441 15044 30493
rect 15108 30458 15111 30493
rect 15297 30458 15298 30493
rect 15096 30441 15111 30458
rect 15163 30441 15178 30458
rect 15230 30441 15245 30458
rect 15297 30441 15312 30458
rect 15364 30441 15378 30493
rect 15436 30458 15444 30493
rect 15430 30441 15444 30458
rect 15496 30441 15510 30493
rect 15562 30441 15576 30493
rect 15628 30441 15638 30493
rect 14636 30432 15638 30441
rect 14636 30409 14888 30432
rect 14944 30409 14970 30432
rect 15026 30409 15052 30432
rect 15108 30409 15134 30432
rect 15190 30409 15216 30432
rect 15272 30409 15298 30432
rect 15354 30409 15380 30432
rect 15436 30409 15638 30432
rect 14636 30357 14642 30409
rect 14694 30357 14709 30409
rect 14761 30357 14776 30409
rect 14828 30357 14843 30409
rect 14962 30376 14970 30409
rect 14895 30357 14910 30376
rect 14962 30357 14977 30376
rect 15029 30357 15044 30409
rect 15108 30376 15111 30409
rect 15297 30376 15298 30409
rect 15096 30357 15111 30376
rect 15163 30357 15178 30376
rect 15230 30357 15245 30376
rect 15297 30357 15312 30376
rect 15364 30357 15378 30409
rect 15436 30376 15444 30409
rect 15430 30357 15444 30376
rect 15496 30357 15510 30409
rect 15562 30357 15576 30409
rect 15628 30357 15638 30409
rect 14636 30350 15638 30357
rect 14636 30325 14888 30350
rect 14944 30325 14970 30350
rect 15026 30325 15052 30350
rect 15108 30325 15134 30350
rect 15190 30325 15216 30350
rect 15272 30325 15298 30350
rect 15354 30325 15380 30350
rect 15436 30325 15638 30350
rect 14636 30273 14642 30325
rect 14694 30273 14709 30325
rect 14761 30273 14776 30325
rect 14828 30273 14843 30325
rect 14962 30294 14970 30325
rect 14895 30273 14910 30294
rect 14962 30273 14977 30294
rect 15029 30273 15044 30325
rect 15108 30294 15111 30325
rect 15297 30294 15298 30325
rect 15096 30273 15111 30294
rect 15163 30273 15178 30294
rect 15230 30273 15245 30294
rect 15297 30273 15312 30294
rect 15364 30273 15378 30325
rect 15436 30294 15444 30325
rect 15430 30273 15444 30294
rect 15496 30273 15510 30325
rect 15562 30273 15576 30325
rect 15628 30273 15638 30325
rect 14636 30268 15638 30273
rect 14636 30212 14888 30268
rect 14944 30212 14970 30268
rect 15026 30212 15052 30268
rect 15108 30212 15134 30268
rect 15190 30212 15216 30268
rect 15272 30212 15298 30268
rect 15354 30212 15380 30268
rect 15436 30212 15638 30268
rect 14636 30187 15638 30212
rect 21383 30201 21695 31483
tri 22569 31441 22614 31486 se
rect 22614 31441 22666 32907
tri 22666 31441 22697 31472 sw
rect 22569 31389 22575 31441
rect 22627 31389 22639 31441
rect 22691 31389 22697 31441
rect 22953 31230 23005 33104
rect 25439 33206 25595 33258
rect 25647 33206 25663 33258
rect 25715 33206 25731 33258
rect 25783 33206 25784 33258
rect 25439 33194 25784 33206
rect 25439 33142 25595 33194
rect 25647 33142 25663 33194
rect 25715 33142 25731 33194
rect 25783 33142 25784 33194
rect 25439 33129 25784 33142
rect 25439 33077 25595 33129
rect 25647 33077 25663 33129
rect 25715 33077 25731 33129
rect 25783 33077 25784 33129
rect 25439 33064 25784 33077
rect 25439 33012 25595 33064
rect 25647 33012 25663 33064
rect 25715 33012 25731 33064
rect 25783 33012 25784 33064
rect 25439 32999 25784 33012
rect 25439 32947 25595 32999
rect 25647 32947 25663 32999
rect 25715 32947 25731 32999
rect 25783 32947 25784 32999
rect 25439 32934 25784 32947
rect 23266 32879 23276 32909
rect 23328 32879 23340 32909
rect 23392 32889 23457 32909
tri 23457 32889 23477 32909 sw
rect 23392 32882 23477 32889
tri 23477 32882 23484 32889 sw
tri 25432 32882 25439 32889 se
rect 25439 32882 25595 32934
rect 25647 32882 25663 32934
rect 25715 32882 25731 32934
rect 25783 32882 25784 32934
rect 23392 32879 23484 32882
rect 23266 32823 23275 32879
rect 23331 32857 23340 32879
rect 23413 32869 23484 32879
tri 23484 32869 23497 32882 sw
tri 25419 32869 25432 32882 se
rect 25432 32869 25784 32882
rect 23331 32823 23357 32857
rect 23413 32823 23497 32869
tri 23447 32821 23449 32823 ne
rect 23449 32821 23497 32823
tri 23497 32821 23545 32869 sw
tri 23449 32817 23453 32821 ne
rect 23453 32817 23545 32821
tri 25367 32817 25419 32869 se
rect 25419 32817 25595 32869
rect 25647 32817 25663 32869
rect 25715 32817 25731 32869
rect 25783 32817 25784 32869
tri 23453 32813 23457 32817 ne
rect 23457 32813 23545 32817
tri 23457 32804 23466 32813 ne
rect 23466 32804 23545 32813
tri 23466 32777 23493 32804 ne
rect 23308 32309 23360 32317
rect 23308 32245 23360 32257
rect 23037 32234 23089 32240
rect 23037 32170 23089 32182
rect 23037 31282 23089 32118
tri 23089 31282 23101 31294 sw
rect 23037 31272 23101 31282
tri 23037 31240 23069 31272 ne
rect 23069 31240 23101 31272
tri 23005 31230 23015 31240 sw
tri 23069 31230 23079 31240 ne
rect 23079 31230 23101 31240
tri 23101 31230 23153 31282 sw
rect 22953 31220 23015 31230
tri 23015 31220 23025 31230 sw
tri 23079 31220 23089 31230 ne
rect 23089 31229 23153 31230
tri 23153 31229 23154 31230 sw
rect 23089 31220 23154 31229
tri 23154 31220 23163 31229 sw
rect 22953 31218 23025 31220
tri 22953 31188 22983 31218 ne
rect 22983 31188 23025 31218
tri 23025 31188 23057 31220 sw
tri 23089 31188 23121 31220 ne
rect 23121 31188 23163 31220
tri 23163 31188 23195 31220 sw
tri 22983 31176 22995 31188 ne
rect 22995 31176 23057 31188
tri 23057 31176 23069 31188 sw
tri 23121 31176 23133 31188 ne
rect 23133 31176 23195 31188
tri 23195 31176 23207 31188 sw
tri 22995 31166 23005 31176 ne
rect 23005 31166 23069 31176
tri 23069 31166 23079 31176 sw
tri 23133 31166 23143 31176 ne
rect 23143 31166 23207 31176
tri 23005 31124 23047 31166 ne
rect 23047 31156 23079 31166
tri 23079 31156 23089 31166 sw
tri 23143 31156 23153 31166 ne
rect 23153 31156 23207 31166
rect 23047 31146 23089 31156
tri 23089 31146 23099 31156 sw
tri 23153 31146 23163 31156 ne
rect 23163 31155 23207 31156
tri 23207 31155 23228 31176 sw
rect 23163 31146 23228 31155
tri 23228 31146 23237 31155 sw
rect 23047 31124 23099 31146
tri 23099 31124 23121 31146 sw
tri 23163 31124 23185 31146 ne
rect 23185 31124 23237 31146
tri 23237 31124 23259 31146 sw
rect 23308 31139 23360 32193
tri 23360 31139 23361 31140 sw
rect 23308 31124 23361 31139
tri 23361 31124 23376 31139 sw
tri 23047 31096 23075 31124 ne
rect 23075 31096 23121 31124
tri 23121 31096 23149 31124 sw
tri 23185 31096 23213 31124 ne
rect 23213 31096 23259 31124
tri 23259 31096 23287 31124 sw
rect 23308 31118 23376 31124
tri 23308 31096 23330 31118 ne
rect 23330 31096 23376 31118
tri 23376 31096 23404 31124 sw
rect 23493 31096 23545 32804
tri 25364 32814 25367 32817 se
rect 25367 32814 25784 32817
rect 25364 32805 25784 32814
rect 25420 32749 25506 32805
rect 25562 32804 25648 32805
rect 25704 32804 25784 32805
rect 25562 32752 25595 32804
rect 25647 32752 25648 32804
rect 25715 32752 25731 32804
rect 25783 32752 25784 32804
rect 25562 32749 25648 32752
rect 25704 32749 25784 32752
rect 25364 32739 25784 32749
rect 25364 32687 25595 32739
rect 25647 32687 25663 32739
rect 25715 32687 25731 32739
rect 25783 32687 25784 32739
rect 25364 32686 25784 32687
rect 25420 32630 25506 32686
rect 25562 32674 25648 32686
rect 25704 32674 25784 32686
rect 25562 32630 25595 32674
rect 25364 32622 25595 32630
rect 25647 32630 25648 32674
rect 25647 32622 25663 32630
rect 25715 32622 25731 32674
rect 25783 32622 25784 32674
rect 25364 32584 25784 32622
rect 25364 32567 25593 32584
rect 25420 32511 25506 32567
rect 25562 32532 25593 32567
rect 25645 32567 25703 32584
rect 25645 32532 25648 32567
rect 25755 32532 25784 32584
rect 25562 32519 25648 32532
rect 25704 32519 25784 32532
rect 25562 32511 25593 32519
rect 25364 32467 25593 32511
rect 25645 32511 25648 32519
rect 25645 32467 25703 32511
rect 25755 32467 25784 32519
rect 25364 32454 25784 32467
rect 25364 32447 25593 32454
rect 25420 32391 25506 32447
rect 25562 32402 25593 32447
rect 25645 32447 25703 32454
rect 25645 32402 25648 32447
rect 25755 32402 25784 32454
tri 25998 33331 26008 33341 se
rect 26008 33331 26072 33341
tri 26072 33331 26082 33341 nw
tri 26256 33331 26266 33341 se
rect 26266 33332 27377 33341
rect 26266 33331 26319 33332
rect 25998 33320 26061 33331
tri 26061 33320 26072 33331 nw
tri 26245 33320 26256 33331 se
rect 26256 33320 26319 33331
tri 26319 33320 26331 33332 nw
tri 27355 33320 27367 33332 ne
rect 27367 33320 27377 33332
tri 27377 33320 27441 33384 sw
tri 27648 33356 27676 33384 ne
rect 27676 33356 27722 33384
tri 27722 33356 27750 33384 sw
tri 27676 33334 27698 33356 ne
rect 25998 33310 26051 33320
tri 26051 33310 26061 33320 nw
tri 26235 33310 26245 33320 se
rect 26245 33310 26309 33320
tri 26309 33310 26319 33320 nw
tri 27367 33310 27377 33320 ne
rect 27377 33310 27441 33320
rect 25562 32391 25648 32402
rect 25704 32391 25784 32402
rect 25364 32388 25784 32391
rect 25364 32336 25593 32388
rect 25645 32336 25703 32388
rect 25755 32336 25784 32388
tri 25924 32359 25998 32433 se
rect 25998 32411 26050 33310
tri 26050 33309 26051 33310 nw
tri 26234 33309 26235 33310 se
rect 26235 33309 26305 33310
tri 26231 33306 26234 33309 se
rect 26234 33306 26305 33309
tri 26305 33306 26309 33310 nw
tri 27377 33306 27381 33310 ne
rect 27381 33306 27441 33310
tri 26187 33262 26231 33306 se
rect 26231 33262 26261 33306
tri 26261 33262 26305 33306 nw
tri 27381 33298 27389 33306 ne
tri 26181 33256 26187 33262 se
rect 26187 33256 26255 33262
tri 26255 33256 26261 33262 nw
rect 27389 33256 27441 33306
tri 26161 33236 26181 33256 se
rect 26181 33236 26235 33256
tri 26235 33236 26255 33256 nw
tri 26147 33222 26161 33236 se
rect 26161 33222 26221 33236
tri 26221 33222 26235 33236 nw
tri 26136 33211 26147 33222 se
rect 26147 33211 26210 33222
tri 26210 33211 26221 33222 nw
tri 26417 33211 26428 33222 se
rect 26428 33211 27107 33222
tri 27107 33211 27118 33222 sw
tri 26129 33204 26136 33211 se
rect 26136 33204 26203 33211
tri 26203 33204 26210 33211 nw
tri 26410 33204 26417 33211 se
rect 26417 33204 27118 33211
tri 27118 33204 27125 33211 sw
tri 25998 32359 26050 32411 nw
tri 26118 33193 26129 33204 se
rect 26129 33193 26192 33204
tri 26192 33193 26203 33204 nw
tri 26399 33193 26410 33204 se
rect 26410 33193 27125 33204
rect 26118 33192 26191 33193
tri 26191 33192 26192 33193 nw
tri 26398 33192 26399 33193 se
rect 26399 33192 27125 33193
tri 27125 33192 27137 33204 sw
rect 27389 33192 27441 33204
rect 25364 32327 25784 32336
rect 25001 32220 25007 32272
rect 25059 32220 25071 32272
rect 25123 32220 25129 32272
rect 25420 32271 25506 32327
rect 25562 32271 25648 32327
rect 25704 32271 25784 32327
rect 25364 32262 25784 32271
tri 25364 32240 25386 32262 ne
rect 25386 32240 25784 32262
tri 25386 32228 25398 32240 ne
rect 25398 32228 25784 32240
tri 25398 32220 25406 32228 ne
rect 25406 32220 25784 32228
tri 25001 32180 25041 32220 ne
rect 25041 32211 25129 32220
rect 25041 32187 25105 32211
tri 25105 32187 25129 32211 nw
tri 25406 32187 25439 32220 ne
tri 24787 31793 24789 31795 se
rect 24789 31793 24841 31795
rect 24787 31441 24839 31793
tri 24839 31791 24841 31793 nw
rect 24787 31377 24839 31389
rect 24787 31319 24839 31325
rect 25041 31377 25097 32187
tri 25097 32179 25105 32187 nw
tri 25409 31753 25439 31783 se
rect 25439 31753 25784 32220
tri 25873 32308 25924 32359 se
rect 25924 32308 25947 32359
tri 25947 32308 25998 32359 nw
rect 25873 32292 25931 32308
tri 25931 32292 25947 32308 nw
tri 25869 32016 25873 32020 se
rect 25873 32016 25925 32292
tri 25925 32286 25931 32292 nw
tri 26075 32240 26118 32283 se
rect 26118 32257 26170 33192
tri 26170 33171 26191 33192 nw
tri 26377 33171 26398 33192 se
rect 26398 33171 27137 33192
tri 26354 33148 26377 33171 se
rect 26377 33170 27137 33171
rect 26377 33148 26428 33170
tri 26428 33148 26450 33170 nw
tri 27085 33148 27107 33170 ne
rect 27107 33148 27137 33170
tri 26346 33140 26354 33148 se
rect 26354 33140 26420 33148
tri 26420 33140 26428 33148 nw
tri 27107 33140 27115 33148 ne
rect 27115 33140 27137 33148
tri 27137 33140 27189 33192 sw
tri 26343 33137 26346 33140 se
rect 26346 33137 26417 33140
tri 26417 33137 26420 33140 nw
tri 27115 33137 27118 33140 ne
rect 27118 33137 27189 33140
tri 27189 33137 27192 33140 sw
rect 26118 32240 26153 32257
tri 26153 32240 26170 32257 nw
tri 26281 33075 26343 33137 se
rect 26343 33075 26355 33137
tri 26355 33075 26417 33137 nw
tri 27118 33115 27140 33137 ne
tri 26063 32228 26075 32240 se
rect 26075 32228 26141 32240
tri 26141 32228 26153 32240 nw
tri 26040 32205 26063 32228 se
rect 26063 32205 26118 32228
tri 26118 32205 26141 32228 nw
tri 26011 32176 26040 32205 se
rect 26040 32176 26089 32205
tri 26089 32176 26118 32205 nw
rect 25869 32007 25925 32016
rect 25869 31927 25925 31951
rect 25869 31862 25925 31871
tri 26001 32166 26011 32176 se
rect 26011 32166 26079 32176
tri 26079 32166 26089 32176 nw
rect 26001 32156 26069 32166
tri 26069 32156 26079 32166 nw
rect 26001 32007 26057 32156
tri 26057 32144 26069 32156 nw
tri 26234 32038 26281 32085 se
rect 26281 32038 26333 33075
tri 26333 33053 26355 33075 nw
rect 27140 32292 27192 33137
rect 27389 33134 27441 33140
rect 27525 33297 27654 33310
rect 27525 33241 27559 33297
rect 27615 33241 27654 33297
rect 27525 33232 27654 33241
rect 27525 33200 27649 33232
rect 27525 33144 27559 33200
rect 27615 33144 27649 33200
rect 27525 33103 27649 33144
rect 27525 33047 27559 33103
rect 27615 33047 27649 33103
rect 27525 33006 27649 33047
rect 27525 32950 27559 33006
rect 27615 32950 27649 33006
rect 27525 32941 27649 32950
tri 27525 32937 27529 32941 ne
rect 27529 32937 27654 32941
rect 27140 32228 27192 32240
rect 27140 32170 27192 32176
rect 27698 32272 27750 33356
rect 27698 32208 27750 32220
tri 27489 32113 27526 32150 se
rect 27526 32113 27654 32163
rect 27698 32150 27750 32156
tri 26212 32016 26234 32038 se
rect 26234 32016 26333 32038
rect 26001 31927 26057 31951
rect 26001 31862 26057 31871
rect 26142 32007 26333 32016
rect 26198 31951 26333 32007
tri 26490 32111 26492 32113 se
rect 26492 32111 26544 32113
tri 27487 32111 27489 32113 se
rect 27489 32111 27654 32113
tri 27654 32111 27693 32150 sw
tri 26483 31962 26490 31969 se
rect 26490 31962 26542 32111
tri 26542 32109 26544 32111 nw
tri 27485 32109 27487 32111 se
rect 27487 32109 27693 32111
rect 26142 31927 26333 31951
rect 26198 31919 26333 31927
tri 26445 31924 26483 31962 se
rect 26483 31947 26542 31962
rect 26483 31924 26505 31947
rect 26198 31910 26324 31919
tri 26324 31910 26333 31919 nw
tri 26431 31910 26445 31924 se
rect 26445 31910 26505 31924
tri 26505 31910 26542 31947 nw
tri 27444 32068 27485 32109 se
rect 27485 32068 27693 32109
tri 27693 32068 27736 32111 sw
rect 27444 32038 27660 32068
rect 27716 32038 27773 32068
rect 27444 31986 27450 32038
rect 27502 31986 27529 32038
rect 27581 31986 27609 32038
rect 27661 31986 27689 32012
rect 27741 31986 27769 32038
rect 27829 32012 27885 32068
rect 27941 32012 27950 32068
rect 27821 31986 27950 32012
rect 27444 31964 27950 31986
rect 27444 31962 27660 31964
rect 27716 31962 27773 31964
rect 27444 31910 27450 31962
rect 27502 31910 27529 31962
rect 27581 31910 27609 31962
rect 27741 31910 27769 31962
rect 26198 31908 26322 31910
tri 26322 31908 26324 31910 nw
tri 26429 31908 26431 31910 se
rect 26431 31908 26503 31910
tri 26503 31908 26505 31910 nw
rect 27444 31908 27660 31910
rect 27716 31908 27773 31910
rect 27829 31908 27885 31964
rect 27941 31908 27950 31964
rect 26198 31895 26309 31908
tri 26309 31895 26322 31908 nw
tri 26416 31895 26429 31908 se
rect 26429 31895 26490 31908
tri 26490 31895 26503 31908 nw
rect 26198 31877 26291 31895
tri 26291 31877 26309 31895 nw
tri 26398 31877 26416 31895 se
rect 26416 31877 26472 31895
tri 26472 31877 26490 31895 nw
rect 27132 31877 27482 31880
rect 26198 31871 26276 31877
rect 26142 31862 26276 31871
tri 26276 31862 26291 31877 nw
tri 26383 31862 26398 31877 se
rect 26398 31862 26420 31877
tri 26346 31825 26383 31862 se
rect 26383 31825 26420 31862
tri 26420 31825 26472 31877 nw
rect 27132 31825 27140 31877
rect 27192 31825 27211 31877
rect 27263 31825 27282 31877
rect 27334 31825 27352 31877
rect 27404 31825 27422 31877
rect 27474 31825 27482 31877
tri 26342 31821 26346 31825 se
rect 26346 31821 26416 31825
tri 26416 31821 26420 31825 nw
tri 26326 31805 26342 31821 se
rect 26342 31805 26400 31821
tri 26400 31805 26416 31821 nw
rect 27132 31805 27482 31825
tri 26274 31753 26326 31805 se
rect 26326 31753 26348 31805
tri 26348 31753 26400 31805 nw
rect 27132 31753 27140 31805
rect 27192 31753 27211 31805
rect 27263 31753 27282 31805
rect 27334 31753 27352 31805
rect 27404 31753 27422 31805
rect 27474 31753 27482 31805
tri 25405 31749 25409 31753 se
rect 25409 31749 25784 31753
rect 25357 31743 25784 31749
tri 26268 31747 26274 31753 se
rect 26274 31747 26342 31753
tri 26342 31747 26348 31753 nw
rect 25409 31691 25483 31743
rect 25535 31691 25784 31743
tri 26254 31733 26268 31747 se
rect 26268 31733 26328 31747
tri 26328 31733 26342 31747 nw
rect 27132 31733 27482 31753
tri 26249 31728 26254 31733 se
rect 26254 31728 26276 31733
tri 26243 31722 26249 31728 se
rect 26249 31722 26276 31728
rect 25357 31681 25784 31691
tri 25784 31681 25825 31722 sw
tri 26202 31681 26243 31722 se
rect 26243 31681 26276 31722
tri 26276 31681 26328 31733 nw
rect 27132 31681 27140 31733
rect 27192 31681 27211 31733
rect 27263 31681 27282 31733
rect 27334 31681 27352 31733
rect 27404 31681 27422 31733
rect 27474 31681 27482 31733
rect 25357 31673 25825 31681
tri 25825 31673 25833 31681 sw
tri 26194 31673 26202 31681 se
rect 26202 31673 26268 31681
tri 26268 31673 26276 31681 nw
rect 25357 31668 25833 31673
rect 25409 31616 25483 31668
rect 25535 31642 25833 31668
tri 25833 31642 25864 31673 sw
tri 26163 31642 26194 31673 se
rect 25535 31616 25849 31642
rect 25357 31599 25849 31616
tri 26120 31599 26163 31642 se
rect 26163 31599 26194 31642
tri 26194 31599 26268 31673 nw
rect 25357 31592 25803 31599
rect 25409 31540 25483 31592
rect 25535 31553 25803 31592
tri 25803 31553 25849 31599 nw
tri 26074 31553 26120 31599 se
rect 26120 31553 26148 31599
tri 26148 31553 26194 31599 nw
rect 25535 31540 25784 31553
rect 25357 31534 25784 31540
tri 25784 31534 25803 31553 nw
tri 26055 31534 26074 31553 se
rect 26074 31534 26120 31553
tri 26046 31525 26055 31534 se
rect 26055 31525 26120 31534
tri 26120 31525 26148 31553 nw
tri 26285 31525 26313 31553 se
rect 26313 31525 26320 31553
tri 26022 31501 26046 31525 se
rect 26046 31501 26096 31525
tri 26096 31501 26120 31525 nw
tri 26261 31501 26285 31525 se
rect 26285 31501 26320 31525
rect 26372 31501 26384 31553
rect 26436 31501 26442 31553
tri 25972 31451 26022 31501 se
rect 26022 31451 26046 31501
tri 26046 31451 26096 31501 nw
tri 26239 31479 26261 31501 se
rect 26261 31479 26313 31501
tri 26313 31479 26335 31501 nw
tri 26211 31451 26239 31479 se
rect 26239 31451 26272 31479
tri 25959 31438 25972 31451 se
rect 25972 31438 26033 31451
tri 26033 31438 26046 31451 nw
tri 26198 31438 26211 31451 se
rect 26211 31438 26272 31451
tri 26272 31438 26313 31479 nw
rect 26544 31454 26600 31463
tri 25907 31386 25959 31438 se
rect 25959 31386 25981 31438
tri 25981 31386 26033 31438 nw
tri 26165 31405 26198 31438 se
rect 26198 31405 26239 31438
tri 26239 31405 26272 31438 nw
tri 26146 31386 26165 31405 se
rect 26165 31386 26220 31405
tri 26220 31386 26239 31405 nw
rect 26544 31386 26546 31398
rect 26598 31386 26600 31398
tri 25902 31381 25907 31386 se
rect 25907 31381 25972 31386
tri 25097 31377 25101 31381 sw
tri 25898 31377 25902 31381 se
rect 25902 31377 25972 31381
tri 25972 31377 25981 31386 nw
tri 26137 31377 26146 31386 se
rect 26146 31377 26208 31386
rect 25041 31374 25101 31377
tri 25101 31374 25104 31377 sw
tri 25895 31374 25898 31377 se
rect 25898 31374 25969 31377
tri 25969 31374 25972 31377 nw
tri 26134 31374 26137 31377 se
rect 26137 31374 26208 31377
tri 26208 31374 26220 31386 nw
rect 26544 31374 26600 31386
rect 25041 31347 25104 31374
tri 25104 31347 25131 31374 sw
tri 25868 31347 25895 31374 se
rect 25895 31347 25941 31374
rect 25041 31295 25047 31347
rect 25099 31295 25111 31347
rect 25163 31295 25169 31347
tri 25867 31346 25868 31347 se
rect 25868 31346 25941 31347
tri 25941 31346 25969 31374 nw
tri 26106 31346 26134 31374 se
rect 26134 31346 26180 31374
tri 26180 31346 26208 31374 nw
rect 26292 31362 26348 31371
tri 25824 31303 25867 31346 se
rect 25867 31303 25898 31346
tri 25898 31303 25941 31346 nw
tri 26091 31331 26106 31346 se
rect 26106 31331 26165 31346
tri 26165 31331 26180 31346 nw
tri 26063 31303 26091 31331 se
rect 26091 31303 26128 31331
tri 25816 31295 25824 31303 se
rect 25824 31295 25889 31303
tri 25815 31294 25816 31295 se
rect 25816 31294 25889 31295
tri 25889 31294 25898 31303 nw
tri 26054 31294 26063 31303 se
rect 26063 31294 26128 31303
tri 26128 31294 26165 31331 nw
rect 26544 31309 26600 31318
rect 26292 31294 26294 31306
rect 26346 31294 26348 31306
tri 25803 31282 25815 31294 se
rect 25815 31282 25877 31294
tri 25877 31282 25889 31294 nw
tri 26042 31282 26054 31294 se
rect 26054 31282 26116 31294
tri 26116 31282 26128 31294 nw
rect 26292 31282 26348 31294
tri 25751 31230 25803 31282 se
rect 25803 31230 25825 31282
tri 25825 31230 25877 31282 nw
tri 26017 31257 26042 31282 se
rect 26042 31257 26091 31282
tri 26091 31257 26116 31282 nw
tri 25990 31230 26017 31257 se
rect 26017 31230 26064 31257
tri 26064 31230 26091 31257 nw
tri 25750 31229 25751 31230 se
rect 25751 31229 25824 31230
tri 25824 31229 25825 31230 nw
tri 25989 31229 25990 31230 se
rect 25990 31229 26022 31230
tri 25709 31188 25750 31229 se
rect 25750 31188 25783 31229
tri 25783 31188 25824 31229 nw
tri 25948 31188 25989 31229 se
rect 25989 31188 26022 31229
tri 26022 31188 26064 31230 nw
rect 26292 31217 26348 31226
rect 26796 31256 26852 31265
rect 26796 31188 26798 31200
rect 26850 31188 26852 31200
tri 25697 31176 25709 31188 se
rect 25709 31176 25771 31188
tri 25771 31176 25783 31188 nw
tri 25943 31183 25948 31188 se
rect 25948 31183 26017 31188
tri 26017 31183 26022 31188 nw
tri 25936 31176 25943 31183 se
rect 25943 31176 26010 31183
tri 26010 31176 26017 31183 nw
rect 26796 31176 26852 31188
tri 25676 31155 25697 31176 se
rect 25697 31155 25750 31176
tri 25750 31155 25771 31176 nw
tri 25915 31155 25936 31176 se
rect 25936 31155 25958 31176
tri 25645 31124 25676 31155 se
rect 25676 31124 25719 31155
tri 25719 31124 25750 31155 nw
tri 25884 31124 25915 31155 se
rect 25915 31124 25958 31155
tri 25958 31124 26010 31176 nw
tri 25629 31108 25645 31124 se
rect 25645 31108 25691 31124
tri 23545 31096 23557 31108 sw
tri 25617 31096 25629 31108 se
rect 25629 31096 25691 31108
tri 25691 31096 25719 31124 nw
tri 25869 31109 25884 31124 se
rect 25884 31109 25943 31124
tri 25943 31109 25958 31124 nw
rect 26796 31111 26852 31120
rect 26922 31112 26978 31121
tri 25856 31096 25869 31109 se
rect 25869 31096 25930 31109
tri 25930 31096 25943 31109 nw
tri 23075 31092 23079 31096 ne
rect 23079 31092 23149 31096
tri 23149 31092 23153 31096 sw
tri 23213 31092 23217 31096 ne
rect 23217 31092 23287 31096
tri 23079 31044 23127 31092 ne
rect 23127 31082 23153 31092
tri 23153 31082 23163 31092 sw
tri 23217 31082 23227 31092 ne
rect 23227 31082 23287 31092
rect 23127 31072 23163 31082
tri 23163 31072 23173 31082 sw
tri 23227 31072 23237 31082 ne
rect 23237 31081 23287 31082
tri 23287 31081 23302 31096 sw
tri 23330 31081 23345 31096 ne
rect 23345 31081 23404 31096
tri 23404 31081 23419 31096 sw
rect 23493 31086 23557 31096
tri 23493 31081 23498 31086 ne
rect 23498 31081 23557 31086
tri 23557 31081 23572 31096 sw
tri 25602 31081 25617 31096 se
rect 25617 31081 25676 31096
tri 25676 31081 25691 31096 nw
tri 25841 31081 25856 31096 se
rect 25856 31081 25878 31096
rect 23237 31075 23302 31081
tri 23302 31075 23308 31081 sw
tri 23345 31075 23351 31081 ne
rect 23351 31075 23419 31081
rect 23237 31072 23308 31075
tri 23308 31072 23311 31075 sw
tri 23351 31072 23354 31075 ne
rect 23354 31072 23419 31075
tri 23419 31072 23428 31081 sw
tri 23498 31072 23507 31081 ne
rect 23507 31072 23572 31081
tri 23572 31072 23581 31081 sw
tri 25593 31072 25602 31081 se
rect 25602 31072 25639 31081
rect 23127 31065 23173 31072
tri 23173 31065 23180 31072 sw
tri 23237 31065 23244 31072 ne
rect 23244 31065 23311 31072
tri 23311 31065 23318 31072 sw
tri 23354 31065 23361 31072 ne
rect 23361 31065 23428 31072
tri 23428 31065 23435 31072 sw
tri 23507 31065 23514 31072 ne
rect 23514 31065 23581 31072
rect 23127 31044 23180 31065
tri 23180 31044 23201 31065 sw
tri 23244 31044 23265 31065 ne
rect 23265 31044 23318 31065
tri 23318 31044 23339 31065 sw
tri 23361 31044 23382 31065 ne
rect 23382 31064 23435 31065
tri 23435 31064 23436 31065 sw
tri 23514 31064 23515 31065 ne
rect 23515 31064 23581 31065
tri 23581 31064 23589 31072 sw
tri 25585 31064 25593 31072 se
rect 25593 31064 25639 31072
rect 23382 31044 23436 31064
tri 23436 31044 23456 31064 sw
tri 23515 31044 23535 31064 ne
rect 23535 31044 23589 31064
tri 23589 31044 23609 31064 sw
tri 25581 31060 25585 31064 se
rect 25585 31060 25639 31064
rect 24402 31051 24458 31060
tri 23127 31032 23139 31044 ne
rect 23139 31032 23201 31044
tri 23201 31032 23213 31044 sw
tri 23265 31032 23277 31044 ne
rect 23277 31032 23339 31044
tri 23339 31032 23351 31044 sw
tri 23382 31032 23394 31044 ne
rect 23394 31034 23456 31044
tri 23456 31034 23466 31044 sw
tri 23535 31034 23545 31044 ne
rect 23545 31034 23609 31044
rect 23394 31032 23466 31034
tri 23466 31032 23468 31034 sw
tri 23545 31032 23547 31034 ne
rect 23547 31032 23609 31034
tri 23609 31032 23621 31044 sw
tri 23139 31018 23153 31032 ne
rect 23153 31018 23213 31032
tri 23213 31018 23227 31032 sw
tri 23277 31018 23291 31032 ne
rect 23291 31022 23351 31032
tri 23351 31022 23361 31032 sw
tri 23394 31022 23404 31032 ne
rect 23404 31022 23468 31032
rect 23291 31018 23361 31022
tri 23153 30980 23191 31018 ne
rect 23191 31008 23227 31018
tri 23227 31008 23237 31018 sw
tri 23291 31008 23301 31018 ne
rect 23301 31008 23361 31018
rect 23191 30998 23237 31008
tri 23237 30998 23247 31008 sw
tri 23301 30998 23311 31008 ne
rect 23311 31007 23361 31008
tri 23361 31007 23376 31022 sw
tri 23404 31007 23419 31022 ne
rect 23419 31007 23468 31022
tri 23468 31007 23493 31032 sw
tri 23547 31007 23572 31032 ne
rect 23572 31007 23621 31032
tri 23621 31007 23646 31032 sw
rect 23311 30998 23376 31007
tri 23376 30998 23385 31007 sw
tri 23419 30998 23428 31007 ne
rect 23428 30998 23493 31007
tri 23493 30998 23502 31007 sw
tri 23572 30998 23581 31007 ne
rect 23581 30998 23646 31007
tri 23646 30998 23655 31007 sw
rect 23191 30991 23247 30998
tri 23247 30991 23254 30998 sw
tri 23311 30991 23318 30998 ne
rect 23318 30991 23385 30998
tri 23385 30991 23392 30998 sw
tri 23428 30991 23435 30998 ne
rect 23435 30991 23502 30998
tri 23502 30991 23509 30998 sw
tri 23581 30991 23588 30998 ne
rect 23588 30991 23655 30998
rect 23191 30980 23254 30991
tri 23254 30980 23265 30991 sw
tri 23318 30980 23329 30991 ne
rect 23329 30980 23392 30991
tri 23392 30980 23403 30991 sw
tri 23435 30980 23446 30991 ne
rect 23446 30990 23509 30991
tri 23509 30990 23510 30991 sw
tri 23588 30990 23589 30991 ne
rect 23589 30990 23655 30991
tri 23655 30990 23663 30998 sw
tri 25565 31044 25581 31060 se
rect 25581 31044 25639 31060
tri 25639 31044 25676 31081 nw
tri 25804 31044 25841 31081 se
rect 25841 31044 25878 31081
tri 25878 31044 25930 31096 nw
rect 26922 31044 26924 31056
rect 26976 31044 26978 31056
tri 25553 31032 25565 31044 se
rect 25565 31032 25627 31044
tri 25627 31032 25639 31044 nw
tri 25795 31035 25804 31044 se
rect 25804 31035 25869 31044
tri 25869 31035 25878 31044 nw
tri 25792 31032 25795 31035 se
rect 25795 31032 25866 31035
tri 25866 31032 25869 31035 nw
rect 26922 31032 26978 31044
tri 24458 31007 24483 31032 sw
tri 25528 31007 25553 31032 se
rect 25553 31007 25602 31032
tri 25602 31007 25627 31032 nw
tri 25767 31007 25792 31032 se
rect 25792 31007 25814 31032
rect 24458 30995 24483 31007
rect 23446 30980 23510 30990
tri 23510 30980 23520 30990 sw
tri 23589 30980 23599 30990 ne
rect 23599 30980 23663 30990
tri 23663 30980 23673 30990 sw
rect 24402 30980 24483 30995
tri 24483 30980 24510 31007 sw
tri 25501 30980 25528 31007 se
rect 25528 30980 25575 31007
tri 25575 30980 25602 31007 nw
tri 25740 30980 25767 31007 se
rect 25767 30980 25814 31007
tri 25814 30980 25866 31032 nw
tri 23191 30955 23216 30980 ne
rect 23216 30955 23265 30980
tri 23265 30955 23290 30980 sw
tri 23329 30955 23354 30980 ne
rect 23354 30976 23403 30980
tri 23403 30976 23407 30980 sw
tri 23446 30976 23450 30980 ne
rect 23450 30976 23520 30980
tri 23520 30976 23524 30980 sw
tri 23599 30976 23603 30980 ne
rect 23603 30976 23673 30980
tri 23673 30976 23677 30980 sw
rect 24402 30976 24510 30980
tri 24510 30976 24514 30980 sw
tri 25497 30976 25501 30980 se
rect 25501 30976 25571 30980
tri 25571 30976 25575 30980 nw
tri 25736 30976 25740 30980 se
rect 25740 30976 25795 30980
rect 23354 30955 23407 30976
tri 23407 30955 23428 30976 sw
tri 23450 30955 23471 30976 ne
rect 23471 30955 23524 30976
tri 23524 30955 23545 30976 sw
tri 23603 30955 23624 30976 ne
rect 23624 30955 23677 30976
tri 23677 30955 23698 30976 sw
rect 24402 30971 25550 30976
tri 23216 30944 23227 30955 ne
rect 23227 30944 23290 30955
tri 23290 30944 23301 30955 sw
tri 23354 30944 23365 30955 ne
rect 23365 30948 23428 30955
tri 23428 30948 23435 30955 sw
tri 23471 30948 23478 30955 ne
rect 23478 30948 23545 30955
rect 23365 30944 23435 30948
tri 23227 30903 23268 30944 ne
rect 23268 30934 23301 30944
tri 23301 30934 23311 30944 sw
tri 23365 30934 23375 30944 ne
rect 23375 30934 23435 30944
rect 23268 30924 23311 30934
tri 23311 30924 23321 30934 sw
tri 23375 30924 23385 30934 ne
rect 23385 30924 23435 30934
tri 23435 30924 23459 30948 sw
tri 23478 30924 23502 30948 ne
rect 23502 30924 23545 30948
tri 23545 30924 23576 30955 sw
tri 23624 30924 23655 30955 ne
rect 23655 30924 23698 30955
tri 23698 30924 23729 30955 sw
rect 23268 30917 23321 30924
tri 23321 30917 23328 30924 sw
tri 23385 30917 23392 30924 ne
rect 23392 30917 23459 30924
tri 23459 30917 23466 30924 sw
tri 23502 30917 23509 30924 ne
rect 23509 30917 23576 30924
tri 23576 30917 23583 30924 sw
tri 23655 30917 23662 30924 ne
rect 23662 30917 23729 30924
rect 23268 30903 23328 30917
tri 23328 30903 23342 30917 sw
tri 23392 30903 23406 30917 ne
rect 23406 30903 23466 30917
tri 23466 30903 23480 30917 sw
tri 23509 30903 23523 30917 ne
rect 23523 30916 23583 30917
tri 23583 30916 23584 30917 sw
tri 23662 30916 23663 30917 ne
rect 23663 30916 23729 30917
tri 23729 30916 23737 30924 sw
rect 23523 30903 23584 30916
tri 23584 30903 23597 30916 sw
tri 23663 30903 23676 30916 ne
rect 23676 30903 23737 30916
rect 24458 30955 25550 30971
tri 25550 30955 25571 30976 nw
tri 25721 30961 25736 30976 se
rect 25736 30961 25795 30976
tri 25795 30961 25814 30980 nw
rect 26670 30971 26726 30980
tri 25715 30955 25721 30961 se
rect 25721 30955 25789 30961
tri 25789 30955 25795 30961 nw
rect 26922 30967 26978 30976
rect 24458 30924 25519 30955
tri 25519 30924 25550 30955 nw
tri 25691 30931 25715 30955 se
rect 25715 30931 25765 30955
tri 25765 30931 25789 30955 nw
tri 25684 30924 25691 30931 se
rect 25691 30924 25737 30931
rect 24402 30906 24458 30915
tri 24458 30906 24476 30924 nw
tri 25666 30906 25684 30924 se
rect 25684 30906 25737 30924
tri 25663 30903 25666 30906 se
rect 25666 30903 25737 30906
tri 25737 30903 25765 30931 nw
rect 25925 30924 25941 30931
tri 25941 30924 25948 30931 sw
rect 25925 30903 25948 30924
tri 25948 30903 25969 30924 sw
rect 26670 30903 26672 30915
rect 26724 30903 26726 30915
tri 23268 30891 23280 30903 ne
rect 23280 30891 23342 30903
tri 23342 30891 23354 30903 sw
tri 23406 30891 23418 30903 ne
rect 23418 30891 23480 30903
tri 23480 30891 23492 30903 sw
tri 23523 30891 23535 30903 ne
rect 23535 30894 23597 30903
tri 23597 30894 23606 30903 sw
tri 23676 30894 23685 30903 ne
rect 23535 30891 23606 30894
tri 23606 30891 23609 30894 sw
tri 23280 30870 23301 30891 ne
rect 23301 30870 23354 30891
tri 23354 30870 23375 30891 sw
tri 23418 30870 23439 30891 ne
rect 23439 30874 23492 30891
tri 23492 30874 23509 30891 sw
tri 23535 30874 23552 30891 ne
rect 23552 30874 23609 30891
rect 23439 30870 23509 30874
tri 23301 30868 23303 30870 ne
rect 23303 30868 23375 30870
tri 23375 30868 23377 30870 sw
tri 23439 30868 23441 30870 ne
rect 23441 30868 23509 30870
tri 23509 30868 23515 30874 sw
tri 23552 30868 23558 30874 ne
rect 23558 30868 23609 30874
tri 23609 30868 23632 30891 sw
tri 23303 30816 23355 30868 ne
rect 23355 30860 23377 30868
tri 23377 30860 23385 30868 sw
tri 23441 30860 23449 30868 ne
rect 23449 30860 23515 30868
rect 23355 30850 23385 30860
tri 23385 30850 23395 30860 sw
tri 23449 30850 23459 30860 ne
rect 23459 30850 23515 30860
tri 23515 30850 23533 30868 sw
tri 23558 30850 23576 30868 ne
rect 23576 30850 23632 30868
tri 23632 30850 23650 30868 sw
rect 23355 30816 23395 30850
tri 23395 30816 23429 30850 sw
tri 23459 30816 23493 30850 ne
rect 23493 30843 23533 30850
tri 23533 30843 23540 30850 sw
tri 23576 30843 23583 30850 ne
rect 23583 30843 23650 30850
tri 23650 30843 23657 30850 sw
rect 23493 30816 23540 30843
tri 23540 30816 23567 30843 sw
tri 23583 30821 23605 30843 ne
tri 23355 30804 23367 30816 ne
rect 23367 30806 23429 30816
tri 23429 30806 23439 30816 sw
tri 23493 30806 23503 30816 ne
rect 23503 30806 23567 30816
tri 23567 30806 23577 30816 sw
rect 23367 30804 23439 30806
tri 23439 30804 23441 30806 sw
tri 23503 30804 23505 30806 ne
rect 23505 30804 23577 30806
tri 23367 30796 23375 30804 ne
rect 23375 30796 23441 30804
tri 23441 30796 23449 30804 sw
tri 23505 30796 23513 30804 ne
rect 23513 30796 23577 30804
tri 23375 30795 23376 30796 ne
rect 23376 30795 23449 30796
tri 23449 30795 23450 30796 sw
tri 23513 30795 23514 30796 ne
rect 23514 30795 23577 30796
tri 23376 30763 23408 30795 ne
rect 23408 30784 23450 30795
tri 23450 30784 23461 30795 sw
tri 23514 30784 23525 30795 ne
rect 23408 30763 23461 30784
tri 23461 30763 23482 30784 sw
tri 23408 30748 23423 30763 ne
rect 23423 30748 23482 30763
tri 23482 30748 23497 30763 sw
tri 23423 30746 23425 30748 ne
rect 23425 30746 23497 30748
tri 23425 30740 23431 30746 ne
rect 23431 30740 23497 30746
tri 23431 30733 23438 30740 ne
rect 23438 30733 23445 30740
rect 22183 30723 22945 30733
rect 22183 30671 22193 30723
rect 22245 30671 22268 30723
rect 22320 30671 22343 30723
rect 22395 30671 22417 30723
rect 22469 30671 22491 30723
rect 22543 30671 22565 30723
rect 22617 30688 22945 30723
tri 22945 30688 22990 30733 sw
tri 23438 30726 23445 30733 ne
rect 22617 30676 22990 30688
tri 22990 30676 23002 30688 sw
rect 23445 30676 23497 30688
rect 22617 30671 23002 30676
rect 22183 30653 23002 30671
rect 22183 30601 22193 30653
rect 22245 30601 22268 30653
rect 22320 30601 22343 30653
rect 22395 30601 22417 30653
rect 22469 30601 22491 30653
rect 22543 30601 22565 30653
rect 22617 30624 23002 30653
tri 23002 30624 23054 30676 sw
rect 22617 30618 23054 30624
tri 23054 30618 23060 30624 sw
rect 23445 30618 23497 30624
rect 23525 30740 23577 30795
rect 23525 30676 23577 30688
rect 23525 30618 23577 30624
rect 23605 30740 23657 30843
rect 23605 30676 23657 30688
rect 23685 30763 23737 30903
tri 25651 30891 25663 30903 se
rect 25663 30891 25725 30903
tri 25725 30891 25737 30903 nw
rect 25925 30895 25969 30903
tri 25969 30895 25977 30903 sw
tri 25650 30890 25651 30891 se
rect 25651 30890 25724 30891
tri 25724 30890 25725 30891 nw
tri 24548 30868 24570 30890 se
rect 24570 30868 25702 30890
tri 25702 30868 25724 30890 nw
tri 24496 30816 24548 30868 se
rect 24548 30838 25672 30868
tri 25672 30838 25702 30868 nw
rect 24548 30816 24573 30838
tri 24573 30816 24595 30838 nw
rect 25925 30829 25977 30895
rect 25925 30816 25964 30829
tri 25964 30816 25977 30829 nw
rect 26418 30884 26474 30893
rect 26418 30816 26420 30828
rect 26472 30816 26474 30828
rect 26670 30891 26726 30903
rect 26670 30826 26726 30835
tri 27090 30826 27132 30868 se
rect 27132 30826 27482 31681
tri 24493 30813 24496 30816 se
rect 24496 30813 24570 30816
tri 24570 30813 24573 30816 nw
rect 25925 30813 25961 30816
tri 25961 30813 25964 30816 nw
tri 24484 30804 24493 30813 se
rect 24493 30804 24561 30813
tri 24561 30804 24570 30813 nw
rect 25925 30804 25952 30813
tri 25952 30804 25961 30813 nw
rect 26418 30804 26474 30816
tri 24475 30795 24484 30804 se
rect 24484 30795 24552 30804
tri 24552 30795 24561 30804 nw
rect 25925 30795 25943 30804
tri 25943 30795 25952 30804 nw
rect 23767 30743 23773 30795
rect 23825 30743 23837 30795
rect 23889 30777 24534 30795
tri 24534 30777 24552 30795 nw
tri 25925 30777 25943 30795 nw
rect 23889 30752 24509 30777
tri 24509 30752 24534 30777 nw
tri 27041 30777 27090 30826 se
rect 27090 30777 27482 30826
tri 27482 30777 27589 30884 sw
rect 23889 30743 24500 30752
tri 24500 30743 24509 30752 nw
rect 26418 30739 26474 30748
tri 27007 30743 27041 30777 se
rect 27041 30743 27589 30777
tri 27589 30743 27623 30777 sw
tri 27003 30739 27007 30743 se
rect 27007 30739 27623 30743
rect 23685 30699 23737 30711
tri 26973 30709 27003 30739 se
rect 27003 30709 27623 30739
tri 27623 30709 27657 30743 sw
tri 23859 30708 23860 30709 se
rect 23860 30708 28025 30709
tri 23858 30707 23859 30708 se
rect 23859 30707 28025 30708
tri 23854 30703 23858 30707 se
rect 23858 30703 28025 30707
tri 23802 30651 23854 30703 se
rect 23854 30695 27973 30703
rect 23854 30651 24164 30695
rect 23685 30641 23737 30647
tri 23792 30641 23802 30651 se
rect 23802 30641 24164 30651
tri 23783 30632 23792 30641 se
rect 23792 30639 24164 30641
rect 24220 30639 24268 30695
rect 24324 30651 27973 30695
rect 24324 30639 28025 30651
rect 23792 30632 28025 30639
rect 23605 30618 23657 30624
tri 23769 30618 23783 30632 se
rect 23783 30618 23860 30632
rect 22617 30601 23060 30618
rect 22183 30583 23060 30601
rect 22183 30531 22193 30583
rect 22245 30531 22268 30583
rect 22320 30531 22343 30583
rect 22395 30531 22417 30583
rect 22469 30531 22491 30583
rect 22543 30531 22565 30583
rect 22617 30580 23060 30583
tri 23060 30580 23098 30618 sw
tri 23731 30580 23769 30618 se
rect 23769 30580 23860 30618
rect 23912 30580 23932 30632
rect 23984 30623 28025 30632
rect 23984 30619 27973 30623
rect 23984 30600 26862 30619
rect 23984 30587 24164 30600
rect 24220 30587 24268 30600
rect 24324 30587 26862 30600
rect 23984 30580 24024 30587
rect 22617 30574 23098 30580
tri 23098 30574 23104 30580 sw
tri 23725 30574 23731 30580 se
rect 23731 30574 24024 30580
rect 22617 30560 24024 30574
rect 22617 30531 23860 30560
rect 22183 30525 23860 30531
tri 22859 30508 22876 30525 ne
rect 22876 30508 23860 30525
rect 23912 30508 23932 30560
rect 23984 30535 24024 30560
rect 24076 30535 24094 30587
rect 24146 30535 24164 30587
rect 24220 30544 24234 30587
rect 24216 30535 24234 30544
rect 24286 30535 24304 30544
rect 24356 30535 24374 30587
rect 24426 30535 24444 30587
rect 24496 30535 24514 30587
rect 24566 30535 24584 30587
rect 24636 30567 26862 30587
rect 26914 30567 26936 30619
rect 26988 30567 27010 30619
rect 27062 30567 27576 30619
rect 27628 30567 27650 30619
rect 27702 30567 27724 30619
rect 27776 30571 27973 30619
rect 27776 30567 28025 30571
rect 24636 30547 28025 30567
rect 24636 30535 26862 30547
rect 23984 30523 26862 30535
rect 23984 30508 24024 30523
tri 22876 30488 22896 30508 ne
rect 22896 30488 24024 30508
tri 22896 30483 22901 30488 ne
rect 22901 30483 23860 30488
rect 22587 30431 22593 30483
rect 22645 30431 22657 30483
rect 22709 30436 22843 30483
tri 22843 30436 22890 30483 sw
tri 22901 30436 22948 30483 ne
rect 22948 30436 23860 30483
rect 23912 30436 23932 30488
rect 23984 30471 24024 30488
rect 24076 30471 24094 30523
rect 24146 30471 24164 30523
rect 24216 30505 24234 30523
rect 24286 30505 24304 30523
rect 24220 30471 24234 30505
rect 24356 30471 24374 30523
rect 24426 30471 24444 30523
rect 24496 30471 24514 30523
rect 24566 30471 24584 30523
rect 24636 30495 26862 30523
rect 26914 30495 26936 30547
rect 26988 30495 27010 30547
rect 27062 30495 27576 30547
rect 27628 30495 27650 30547
rect 27702 30495 27724 30547
rect 27776 30543 28025 30547
rect 27776 30495 27973 30543
rect 24636 30491 27973 30495
rect 24636 30475 28025 30491
rect 24636 30471 26862 30475
rect 23984 30459 24164 30471
rect 24220 30459 24268 30471
rect 24324 30459 26862 30471
rect 23984 30436 24024 30459
rect 22709 30431 22890 30436
tri 22837 30425 22843 30431 ne
rect 22843 30425 22890 30431
tri 22890 30425 22901 30436 sw
tri 22948 30425 22959 30436 ne
rect 22959 30425 24024 30436
tri 22843 30407 22861 30425 ne
rect 22861 30407 22901 30425
tri 22901 30407 22919 30425 sw
tri 22959 30407 22977 30425 ne
rect 22977 30407 24024 30425
rect 24076 30407 24094 30459
rect 24146 30407 24164 30459
rect 24220 30449 24234 30459
rect 24216 30410 24234 30449
rect 24286 30410 24304 30449
rect 24220 30407 24234 30410
rect 24356 30407 24374 30459
rect 24426 30407 24444 30459
rect 24496 30407 24514 30459
rect 24566 30407 24584 30459
rect 24636 30423 26862 30459
rect 26914 30423 26936 30475
rect 26988 30423 27010 30475
rect 27062 30474 28025 30475
rect 27062 30423 27576 30474
rect 24636 30422 27576 30423
rect 27628 30422 27650 30474
rect 27702 30422 27724 30474
rect 27776 30463 28025 30474
rect 27776 30422 27973 30463
rect 24636 30411 27973 30422
rect 24636 30407 28025 30411
tri 22861 30402 22866 30407 ne
rect 22866 30402 22919 30407
tri 22919 30402 22924 30407 sw
tri 22977 30402 22982 30407 ne
rect 22982 30402 24164 30407
tri 22866 30395 22873 30402 ne
rect 22873 30395 22924 30402
tri 22924 30395 22931 30402 sw
tri 22982 30395 22989 30402 ne
rect 22989 30395 24164 30402
rect 24220 30395 24268 30407
rect 24324 30402 28025 30407
rect 24324 30395 26862 30402
tri 22873 30379 22889 30395 ne
rect 22889 30379 22931 30395
rect 22449 30327 22455 30379
rect 22507 30327 22521 30379
rect 22573 30367 22791 30379
tri 22791 30367 22803 30379 sw
tri 22889 30367 22901 30379 ne
rect 22901 30367 22931 30379
tri 22931 30367 22959 30395 sw
tri 22989 30367 23017 30395 ne
rect 23017 30367 24024 30395
rect 22573 30343 22803 30367
tri 22803 30343 22827 30367 sw
tri 22901 30343 22925 30367 ne
rect 22925 30343 22959 30367
tri 22959 30343 22983 30367 sw
tri 23017 30343 23041 30367 ne
rect 23041 30343 24024 30367
rect 24076 30343 24094 30395
rect 24146 30343 24164 30395
rect 24220 30354 24234 30395
rect 24216 30343 24234 30354
rect 24286 30343 24304 30354
rect 24356 30343 24374 30395
rect 24426 30343 24444 30395
rect 24496 30343 24514 30395
rect 24566 30343 24584 30395
rect 24636 30350 26862 30395
rect 26914 30350 26936 30402
rect 26988 30350 27010 30402
rect 27062 30401 28025 30402
rect 27062 30350 27576 30401
rect 24636 30349 27576 30350
rect 27628 30349 27650 30401
rect 27702 30349 27724 30401
rect 27776 30349 28025 30401
rect 24636 30343 28025 30349
rect 22573 30327 22827 30343
tri 22769 30269 22827 30327 ne
tri 22827 30309 22861 30343 sw
tri 22925 30309 22959 30343 ne
rect 22959 30309 22983 30343
tri 22983 30309 23017 30343 sw
rect 22827 30269 22861 30309
tri 22861 30269 22901 30309 sw
tri 22959 30269 22999 30309 ne
rect 22999 30284 23614 30309
tri 23614 30284 23639 30309 sw
rect 22999 30269 23639 30284
tri 22827 30231 22865 30269 ne
rect 22865 30267 22901 30269
tri 22901 30267 22903 30269 sw
tri 22999 30267 23001 30269 ne
rect 23001 30267 23639 30269
rect 22865 30248 22903 30267
tri 22903 30248 22922 30267 sw
tri 23593 30248 23612 30267 ne
rect 23612 30248 23639 30267
tri 23639 30248 23675 30284 sw
rect 25732 30275 25788 30284
rect 22865 30246 22922 30248
tri 22922 30246 22924 30248 sw
tri 23612 30246 23614 30248 ne
rect 23614 30246 23675 30248
rect 22865 30237 22924 30246
tri 22924 30237 22933 30246 sw
tri 23614 30237 23623 30246 ne
rect 23623 30237 23675 30246
tri 23675 30237 23686 30248 sw
rect 22865 30231 22933 30237
tri 22933 30231 22939 30237 sw
rect 23445 30231 23497 30237
rect 21383 30149 21391 30201
rect 21443 30149 21473 30201
rect 21525 30149 21554 30201
rect 21606 30149 21635 30201
rect 21687 30149 21695 30201
tri 22865 30195 22901 30231 ne
rect 22901 30195 22939 30231
tri 22939 30195 22975 30231 sw
tri 22901 30179 22917 30195 ne
rect 22917 30179 23314 30195
tri 23314 30179 23330 30195 sw
tri 23623 30185 23675 30237 ne
rect 23675 30194 23686 30237
tri 23686 30194 23729 30237 sw
rect 25732 30195 25788 30219
rect 23675 30185 23729 30194
tri 23729 30185 23738 30194 sw
tri 25723 30185 25732 30194 se
tri 22917 30171 22925 30179 ne
rect 22925 30171 23330 30179
tri 23330 30171 23338 30179 sw
tri 22925 30167 22929 30171 ne
rect 22929 30167 23338 30171
tri 23338 30167 23342 30171 sw
rect 23445 30167 23497 30179
rect 21383 30129 21695 30149
tri 22929 30143 22953 30167 ne
rect 22953 30143 23342 30167
rect 21383 30077 21391 30129
rect 21443 30077 21473 30129
rect 21525 30077 21554 30129
rect 21606 30077 21635 30129
rect 21687 30077 21695 30129
tri 23292 30115 23320 30143 ne
rect 23320 30115 23342 30143
tri 23342 30115 23394 30167 sw
tri 23675 30160 23700 30185 ne
rect 23700 30180 23738 30185
tri 23738 30180 23743 30185 sw
tri 25718 30180 25723 30185 se
rect 25723 30180 25732 30185
rect 23700 30160 23743 30180
rect 23497 30122 23573 30160
tri 23573 30122 23611 30160 sw
tri 23700 30122 23738 30160 ne
rect 23738 30130 23743 30160
tri 23743 30130 23793 30180 sw
tri 24073 30130 24123 30180 se
rect 24123 30139 25732 30180
rect 24123 30138 25788 30139
rect 24123 30130 24131 30138
tri 24131 30130 24139 30138 nw
tri 25724 30130 25732 30138 ne
rect 25732 30130 25788 30138
rect 23738 30122 23793 30130
tri 23793 30122 23801 30130 sw
tri 24065 30122 24073 30130 se
rect 24073 30122 24123 30130
tri 24123 30122 24131 30130 nw
rect 23497 30115 23611 30122
tri 23320 30097 23338 30115 ne
rect 23338 30109 23394 30115
tri 23394 30109 23400 30115 sw
rect 23445 30109 23611 30115
tri 23611 30109 23624 30122 sw
tri 23738 30109 23751 30122 ne
rect 23751 30109 24080 30122
rect 23338 30105 23400 30109
tri 23400 30105 23404 30109 sw
tri 23550 30105 23554 30109 ne
rect 23554 30105 23624 30109
tri 23624 30105 23628 30109 sw
tri 23751 30105 23755 30109 ne
rect 23755 30105 24080 30109
rect 23338 30097 23404 30105
tri 23404 30097 23412 30105 sw
tri 23554 30097 23562 30105 ne
rect 23562 30097 23628 30105
tri 23338 30088 23347 30097 ne
rect 23347 30088 23412 30097
tri 23412 30088 23421 30097 sw
tri 23562 30088 23571 30097 ne
rect 23571 30088 23628 30097
tri 23628 30088 23645 30105 sw
tri 23755 30088 23772 30105 ne
rect 23772 30088 24080 30105
rect 21383 30057 21695 30077
rect 21383 30005 21391 30057
rect 21443 30005 21473 30057
rect 21525 30005 21554 30057
rect 21606 30005 21635 30057
rect 21687 30005 21695 30057
tri 22634 30045 22677 30088 se
rect 22677 30046 23296 30088
tri 23296 30046 23338 30088 sw
tri 23347 30046 23389 30088 ne
rect 23389 30086 23421 30088
tri 23421 30086 23423 30088 sw
tri 23571 30086 23573 30088 ne
rect 23573 30086 23645 30088
rect 23389 30046 23423 30086
rect 22677 30045 23338 30046
tri 23338 30045 23339 30046 sw
tri 23389 30045 23390 30046 ne
rect 23390 30045 23423 30046
tri 23423 30045 23464 30086 sw
tri 23573 30045 23614 30086 ne
rect 23614 30079 23645 30086
tri 23645 30079 23654 30088 sw
tri 23772 30079 23781 30088 ne
rect 23781 30079 24080 30088
tri 24080 30079 24123 30122 nw
rect 23614 30045 23654 30079
tri 23654 30045 23688 30079 sw
tri 22610 30021 22634 30045 se
rect 22634 30036 23339 30045
rect 22634 30021 22684 30036
tri 22684 30021 22699 30036 nw
tri 23274 30021 23289 30036 ne
rect 23289 30027 23339 30036
tri 23339 30027 23357 30045 sw
tri 23390 30027 23408 30045 ne
rect 23408 30031 23464 30045
tri 23464 30031 23478 30045 sw
tri 23614 30031 23628 30045 ne
rect 23628 30031 23688 30045
tri 23688 30031 23702 30045 sw
rect 23408 30027 23478 30031
tri 23478 30027 23482 30031 sw
tri 23628 30027 23632 30031 ne
rect 23632 30027 23702 30031
tri 23702 30027 23706 30031 sw
rect 23289 30023 23357 30027
tri 23357 30023 23361 30027 sw
tri 23408 30023 23412 30027 ne
rect 23412 30023 23482 30027
tri 23482 30023 23486 30027 sw
tri 23632 30023 23636 30027 ne
rect 23636 30023 23706 30027
rect 23289 30021 23361 30023
tri 23361 30021 23363 30023 sw
tri 23412 30021 23414 30023 ne
rect 23414 30021 23486 30023
tri 23486 30021 23488 30023 sw
tri 23636 30021 23638 30023 ne
rect 23638 30021 23706 30023
tri 23706 30021 23712 30027 sw
tri 27307 30021 27313 30027 se
rect 27313 30021 27365 30027
tri 22603 30014 22610 30021 se
rect 22610 30014 22677 30021
tri 22677 30014 22684 30021 nw
tri 23289 30014 23296 30021 ne
rect 23296 30014 23363 30021
rect 21383 30001 21695 30005
tri 22590 30001 22603 30014 se
rect 22603 30001 22634 30014
tri 22560 29971 22590 30001 se
rect 22590 29971 22634 30001
tri 22634 29971 22677 30014 nw
tri 23296 29971 23339 30014 ne
rect 23339 30009 23363 30014
tri 23363 30009 23375 30021 sw
tri 23414 30009 23426 30021 ne
rect 23426 30009 23488 30021
tri 23488 30009 23500 30021 sw
tri 23638 30009 23650 30021 ne
rect 23650 30009 23712 30021
tri 23712 30009 23724 30021 sw
tri 27295 30009 27307 30021 se
rect 27307 30009 27313 30021
rect 23339 30001 23375 30009
tri 23375 30001 23383 30009 sw
tri 23426 30001 23434 30009 ne
rect 23434 30001 23500 30009
tri 23500 30001 23508 30009 sw
tri 23650 30001 23658 30009 ne
rect 23658 30001 23724 30009
tri 23724 30001 23732 30009 sw
tri 24275 30001 24283 30009 se
rect 24283 30001 27313 30009
rect 23339 29972 23383 30001
tri 23383 29972 23412 30001 sw
tri 23434 29972 23463 30001 ne
rect 23463 29972 23508 30001
rect 23339 29971 23412 29972
tri 23412 29971 23413 29972 sw
tri 22558 29969 22560 29971 se
rect 22560 29969 22632 29971
tri 22632 29969 22634 29971 nw
tri 23339 29969 23341 29971 ne
rect 23341 29969 23413 29971
tri 23463 29969 23466 29972 ne
rect 23466 29969 23508 29972
tri 23508 29969 23540 30001 sw
tri 23658 29969 23690 30001 ne
rect 23690 29969 23732 30001
tri 23732 29969 23764 30001 sw
tri 24243 29969 24275 30001 se
rect 24275 29969 27313 30001
tri 22546 29957 22558 29969 se
rect 22558 29957 22620 29969
tri 22620 29957 22632 29969 nw
tri 23341 29957 23353 29969 ne
rect 23353 29957 23413 29969
tri 23466 29957 23478 29969 ne
rect 23478 29957 23540 29969
tri 23540 29957 23552 29969 sw
tri 23690 29957 23702 29969 ne
rect 23702 29957 23764 29969
tri 23764 29957 23776 29969 sw
tri 24231 29957 24243 29969 se
rect 24243 29957 27365 29969
tri 22529 29940 22546 29957 se
rect 22546 29940 22603 29957
tri 22603 29940 22620 29957 nw
tri 23353 29949 23361 29957 ne
tri 22523 29934 22529 29940 se
rect 22529 29934 22597 29940
tri 22597 29934 22603 29940 nw
rect 20373 29882 20379 29934
rect 20431 29882 20449 29934
rect 20501 29882 20519 29934
rect 20571 29882 20588 29934
rect 20640 29925 22588 29934
tri 22588 29925 22597 29934 nw
rect 20640 29905 22568 29925
tri 22568 29905 22588 29925 nw
rect 20640 29882 22545 29905
tri 22545 29882 22568 29905 nw
rect 23361 29842 23413 29957
tri 23478 29949 23486 29957 ne
rect 23486 29949 23552 29957
tri 23552 29949 23560 29957 sw
tri 23702 29949 23710 29957 ne
rect 23710 29949 24300 29957
tri 23486 29905 23530 29949 ne
rect 23530 29905 23560 29949
tri 23560 29905 23604 29949 sw
tri 23710 29905 23754 29949 ne
rect 23754 29925 24300 29949
tri 24300 29925 24332 29957 nw
tri 27281 29925 27313 29957 ne
rect 23754 29905 24280 29925
tri 24280 29905 24300 29925 nw
tri 23530 29875 23560 29905 ne
rect 23560 29899 23604 29905
tri 23604 29899 23610 29905 sw
rect 27313 29899 27365 29905
rect 23560 29875 23610 29899
tri 23610 29875 23634 29899 sw
tri 23560 29843 23592 29875 ne
rect 23592 29843 23634 29875
tri 23634 29843 23666 29875 sw
rect 23443 29842 23495 29843
rect 23361 29837 23495 29842
rect 23361 29785 23443 29837
tri 23592 29801 23634 29843 ne
rect 23634 29801 23666 29843
tri 23666 29801 23708 29843 sw
rect 23443 29755 23495 29785
tri 23634 29727 23708 29801 ne
tri 23708 29727 23782 29801 sw
rect 25410 29727 25466 29731
rect 23443 29697 23495 29703
tri 23708 29697 23738 29727 ne
rect 23738 29722 25471 29727
rect 23738 29697 25410 29722
tri 23738 29675 23760 29697 ne
rect 23760 29675 25410 29697
rect 25466 29675 25471 29722
rect 25410 29642 25466 29666
rect 25410 29577 25466 29586
tri 18759 29210 18793 29244 se
tri 18885 29125 18919 29159 se
tri 18631 28947 18665 28981 ne
rect 8162 28590 8339 28887
rect 23758 28860 24317 28869
rect 23758 28804 23765 28860
rect 23821 28804 24261 28860
rect 23758 28780 24317 28804
rect 23758 28724 23765 28780
rect 23821 28724 24261 28780
rect 23758 28715 24317 28724
tri 25532 28490 25536 28494 se
rect 25536 28490 25593 28494
tri 25593 28490 25597 28494 sw
rect 23443 28485 25673 28490
rect 23443 28484 25536 28485
rect 23495 28432 25536 28484
rect 23443 28429 25536 28432
rect 25592 28429 25673 28485
rect 23443 28405 25673 28429
rect 23443 28402 25536 28405
rect 23495 28350 25536 28402
rect 23443 28349 25536 28350
rect 25592 28349 25673 28405
rect 23443 28344 25673 28349
tri 25532 28340 25536 28344 ne
rect 25536 28340 25593 28344
tri 25593 28340 25597 28344 nw
rect 24184 28137 26537 28143
rect 24184 28085 24185 28137
rect 24237 28085 24259 28137
rect 24311 28085 24333 28137
rect 24385 28085 25307 28137
rect 25359 28085 25385 28137
rect 25437 28085 25923 28137
rect 25975 28085 26001 28137
rect 26053 28085 26336 28137
rect 26388 28085 26410 28137
rect 26462 28085 26484 28137
rect 26536 28085 26537 28137
rect 24184 28067 26537 28085
rect 24184 28015 24185 28067
rect 24237 28015 24259 28067
rect 24311 28015 24333 28067
rect 24385 28053 26336 28067
rect 24385 28015 25307 28053
rect 24184 28001 25307 28015
rect 25359 28001 25385 28053
rect 25437 28001 25923 28053
rect 25975 28001 26001 28053
rect 26053 28015 26336 28053
rect 26388 28015 26410 28067
rect 26462 28015 26484 28067
rect 26536 28015 26537 28067
rect 26053 28001 26537 28015
rect 24184 27997 26537 28001
rect 24184 27945 24185 27997
rect 24237 27945 24259 27997
rect 24311 27945 24333 27997
rect 24385 27969 26336 27997
rect 24385 27945 25307 27969
rect 24184 27927 25307 27945
rect 24184 27875 24185 27927
rect 24237 27875 24259 27927
rect 24311 27875 24333 27927
rect 24385 27917 25307 27927
rect 25359 27917 25385 27969
rect 25437 27917 25923 27969
rect 25975 27917 26001 27969
rect 26053 27945 26336 27969
rect 26388 27945 26410 27997
rect 26462 27945 26484 27997
rect 26536 27945 26537 27997
rect 26053 27927 26537 27945
rect 26053 27917 26336 27927
rect 24385 27884 26336 27917
rect 24385 27875 25307 27884
rect 24184 27857 25307 27875
rect 24184 27805 24185 27857
rect 24237 27805 24259 27857
rect 24311 27805 24333 27857
rect 24385 27832 25307 27857
rect 25359 27832 25385 27884
rect 25437 27832 25923 27884
rect 25975 27832 26001 27884
rect 26053 27875 26336 27884
rect 26388 27875 26410 27927
rect 26462 27875 26484 27927
rect 26536 27875 26537 27927
rect 26053 27856 26537 27875
rect 26053 27832 26336 27856
rect 24385 27805 26336 27832
rect 24184 27804 26336 27805
rect 26388 27804 26410 27856
rect 26462 27804 26484 27856
rect 26536 27804 26537 27856
rect 24184 27799 26537 27804
rect 24184 27786 25307 27799
rect 24184 27734 24185 27786
rect 24237 27734 24259 27786
rect 24311 27734 24333 27786
rect 24385 27747 25307 27786
rect 25359 27747 25385 27799
rect 25437 27747 25923 27799
rect 25975 27747 26001 27799
rect 26053 27785 26537 27799
rect 26053 27747 26336 27785
rect 24385 27734 26336 27747
rect 24184 27733 26336 27734
rect 26388 27733 26410 27785
rect 26462 27733 26484 27785
rect 26536 27733 26537 27785
rect 24184 27715 26537 27733
rect 24184 27663 24185 27715
rect 24237 27663 24259 27715
rect 24311 27663 24333 27715
rect 24385 27714 26537 27715
rect 24385 27663 25307 27714
rect 24184 27662 25307 27663
rect 25359 27662 25385 27714
rect 25437 27662 25923 27714
rect 25975 27662 26001 27714
rect 26053 27662 26336 27714
rect 26388 27662 26410 27714
rect 26462 27662 26484 27714
rect 26536 27662 26537 27714
rect 24184 27656 26537 27662
rect 18906 26469 19032 27035
rect 24169 26791 26557 26797
rect 24169 26739 24185 26791
rect 24237 26739 24259 26791
rect 24311 26739 24333 26791
rect 24385 26739 25413 26791
rect 25465 26739 25491 26791
rect 25543 26739 25923 26791
rect 25975 26739 26001 26791
rect 26053 26739 26336 26791
rect 26388 26739 26410 26791
rect 26462 26739 26484 26791
rect 26536 26739 26557 26791
rect 24169 26721 26557 26739
rect 24169 26669 24185 26721
rect 24237 26669 24259 26721
rect 24311 26669 24333 26721
rect 24385 26707 26336 26721
rect 24385 26669 25413 26707
rect 24169 26655 25413 26669
rect 25465 26655 25491 26707
rect 25543 26655 25923 26707
rect 25975 26655 26001 26707
rect 26053 26669 26336 26707
rect 26388 26669 26410 26721
rect 26462 26669 26484 26721
rect 26536 26669 26557 26721
rect 26053 26655 26557 26669
rect 24169 26651 26557 26655
rect 24169 26599 24185 26651
rect 24237 26599 24259 26651
rect 24311 26599 24333 26651
rect 24385 26623 26336 26651
rect 24385 26599 25413 26623
rect 24169 26581 25413 26599
rect 24169 26529 24185 26581
rect 24237 26529 24259 26581
rect 24311 26529 24333 26581
rect 24385 26571 25413 26581
rect 25465 26571 25491 26623
rect 25543 26571 25923 26623
rect 25975 26571 26001 26623
rect 26053 26599 26336 26623
rect 26388 26599 26410 26651
rect 26462 26599 26484 26651
rect 26536 26599 26557 26651
rect 26053 26581 26557 26599
rect 26053 26571 26336 26581
rect 24385 26538 26336 26571
rect 24385 26529 25413 26538
rect 24169 26510 25413 26529
rect 24169 26458 24185 26510
rect 24237 26458 24259 26510
rect 24311 26458 24333 26510
rect 24385 26486 25413 26510
rect 25465 26486 25491 26538
rect 25543 26486 25923 26538
rect 25975 26486 26001 26538
rect 26053 26529 26336 26538
rect 26388 26529 26410 26581
rect 26462 26529 26484 26581
rect 26536 26529 26557 26581
rect 26053 26510 26557 26529
rect 26053 26486 26336 26510
rect 24385 26458 26336 26486
rect 26388 26458 26410 26510
rect 26462 26458 26484 26510
rect 26536 26458 26557 26510
rect 24169 26453 26557 26458
rect 24169 26439 25413 26453
rect 24169 26387 24185 26439
rect 24237 26387 24259 26439
rect 24311 26387 24333 26439
rect 24385 26401 25413 26439
rect 25465 26401 25491 26453
rect 25543 26401 25923 26453
rect 25975 26401 26001 26453
rect 26053 26439 26557 26453
rect 26053 26401 26336 26439
rect 24385 26387 26336 26401
rect 26388 26387 26410 26439
rect 26462 26387 26484 26439
rect 26536 26387 26557 26439
rect 24169 26368 26557 26387
rect 24169 26316 24185 26368
rect 24237 26316 24259 26368
rect 24311 26316 24333 26368
rect 24385 26316 25413 26368
rect 25465 26316 25491 26368
rect 25543 26316 25923 26368
rect 25975 26316 26001 26368
rect 26053 26316 26336 26368
rect 26388 26316 26410 26368
rect 26462 26316 26484 26368
rect 26536 26316 26557 26368
rect 24169 26310 26557 26316
rect 23264 25131 23316 25137
tri 23316 25100 23353 25137 sw
rect 23316 25079 25632 25100
rect 23264 25067 25632 25079
rect 23316 25048 25632 25067
rect 23264 25009 23316 25015
tri 23316 25011 23353 25048 nw
rect 23184 24637 23236 24643
rect 23236 24585 25509 24610
rect 23184 24573 25509 24585
rect 23236 24558 25509 24573
rect 23184 24515 23236 24521
rect 23445 24063 27223 24069
rect 23497 24011 27171 24063
rect 23445 23999 27223 24011
rect 23497 23947 27171 23999
rect 23445 23941 27223 23947
rect 24528 23560 24584 23569
tri 24512 23513 24528 23529 se
rect 23685 23507 23737 23513
tri 23737 23489 23761 23513 sw
tri 24488 23489 24512 23513 se
rect 24512 23504 24528 23513
rect 24512 23489 24584 23504
tri 24584 23489 24624 23529 sw
rect 23737 23462 25663 23489
rect 23737 23455 24528 23462
rect 23685 23443 24528 23455
rect 23737 23437 24528 23443
tri 23737 23397 23777 23437 nw
tri 24488 23397 24528 23437 ne
rect 24584 23437 25663 23462
rect 25715 23437 25727 23489
rect 25779 23437 25785 23489
rect 24528 23397 24584 23406
tri 24584 23397 24624 23437 nw
rect 23685 23385 23737 23391
rect 23361 23341 23737 23347
rect 23413 23289 23685 23341
rect 23361 23277 23737 23289
rect 23413 23225 23685 23277
rect 23361 23219 23737 23225
tri 26701 23136 26707 23142 se
rect 26707 23136 26759 23142
tri 26688 23123 26701 23136 se
rect 26701 23123 26707 23136
tri 26542 23084 26581 23123 se
rect 26581 23084 26707 23123
tri 26530 23072 26542 23084 se
rect 26542 23072 26759 23084
tri 26507 23049 26530 23072 se
rect 26530 23071 26707 23072
rect 26530 23049 26581 23071
tri 26581 23049 26603 23071 nw
tri 26669 23049 26691 23071 ne
rect 26691 23049 26707 23071
tri 26478 23020 26507 23049 se
rect 26507 23020 26552 23049
tri 26552 23020 26581 23049 nw
tri 26691 23033 26707 23049 ne
tri 26454 22996 26478 23020 se
rect 26478 22996 26507 23020
rect 23525 22990 23577 22996
tri 23577 22975 23598 22996 sw
tri 26433 22975 26454 22996 se
rect 26454 22975 26507 22996
tri 26507 22975 26552 23020 nw
rect 26707 23014 26759 23020
rect 23577 22974 23598 22975
tri 23598 22974 23599 22975 sw
tri 26432 22974 26433 22975 se
rect 26433 22974 26506 22975
tri 26506 22974 26507 22975 nw
rect 23577 22938 26454 22974
rect 23525 22926 26454 22938
rect 23577 22922 26454 22926
tri 26454 22922 26506 22974 nw
tri 23577 22896 23603 22922 nw
rect 23525 22868 23577 22874
rect 23525 22824 23577 22830
tri 27277 22813 27283 22819 se
rect 27283 22813 27335 22819
tri 27274 22810 27277 22813 se
rect 27277 22810 27283 22813
tri 23577 22784 23603 22810 sw
tri 27248 22784 27274 22810 se
rect 27274 22784 27283 22810
rect 23577 22772 27283 22784
rect 23525 22761 27283 22772
rect 23525 22760 27335 22761
tri 23499 22732 23525 22758 ne
rect 23577 22749 27335 22760
rect 23577 22732 27283 22749
rect 23525 22702 23577 22708
tri 23577 22706 23603 22732 nw
tri 27248 22706 27274 22732 ne
rect 27274 22706 27283 22732
tri 27274 22702 27278 22706 ne
rect 27278 22702 27283 22706
tri 27278 22697 27283 22702 ne
rect 27283 22691 27335 22697
rect 26633 22428 26685 22434
rect 23605 22417 23657 22423
tri 23657 22379 23683 22405 sw
tri 26607 22379 26633 22405 se
rect 23657 22376 26633 22379
rect 23657 22365 26685 22376
rect 23605 22364 26685 22365
rect 23605 22353 26633 22364
rect 23657 22327 26633 22353
rect 23657 22312 23668 22327
tri 23668 22312 23683 22327 nw
tri 26612 22312 26627 22327 ne
rect 26627 22312 26633 22327
rect 23657 22306 23662 22312
tri 23662 22306 23668 22312 nw
tri 26627 22306 26633 22312 ne
rect 26633 22306 26685 22312
tri 23657 22301 23662 22306 nw
rect 23605 22295 23657 22301
rect 24169 22263 26557 22269
rect 24169 22211 24185 22263
rect 24237 22211 24259 22263
rect 24311 22211 24333 22263
rect 24385 22211 25307 22263
rect 25359 22211 25385 22263
rect 25437 22211 25923 22263
rect 25975 22211 26001 22263
rect 26053 22211 26336 22263
rect 26388 22211 26410 22263
rect 26462 22211 26484 22263
rect 26536 22211 26557 22263
rect 24169 22198 26557 22211
rect 24169 22146 24185 22198
rect 24237 22146 24259 22198
rect 24311 22146 24333 22198
rect 24385 22165 26336 22198
rect 24385 22146 25307 22165
rect 24169 22133 25307 22146
rect 24169 22081 24185 22133
rect 24237 22081 24259 22133
rect 24311 22081 24333 22133
rect 24385 22113 25307 22133
rect 25359 22113 25385 22165
rect 25437 22113 25923 22165
rect 25975 22113 26001 22165
rect 26053 22146 26336 22165
rect 26388 22146 26410 22198
rect 26462 22146 26484 22198
rect 26536 22146 26557 22198
rect 26053 22133 26557 22146
rect 26053 22113 26336 22133
rect 24385 22081 26336 22113
rect 26388 22081 26410 22133
rect 26462 22081 26484 22133
rect 26536 22081 26557 22133
rect 24169 22067 26557 22081
rect 24169 22015 24185 22067
rect 24237 22015 24259 22067
rect 24311 22015 24333 22067
rect 24385 22015 25307 22067
rect 25359 22015 25385 22067
rect 25437 22015 25923 22067
rect 25975 22015 26001 22067
rect 26053 22015 26336 22067
rect 26388 22015 26410 22067
rect 26462 22015 26484 22067
rect 26536 22015 26557 22067
rect 24169 22009 26557 22015
rect 23445 21995 23497 22001
tri 23497 21984 23502 21989 sw
tri 27278 21984 27283 21989 se
rect 27283 21984 27335 21990
rect 23497 21955 23502 21984
tri 23502 21955 23531 21984 sw
tri 27249 21955 27278 21984 se
rect 27278 21955 27283 21984
rect 23497 21943 27283 21955
rect 23445 21932 27283 21943
rect 23445 21931 27335 21932
rect 23497 21920 27335 21931
rect 23497 21903 27283 21920
rect 23445 21873 23497 21879
tri 23497 21873 23527 21903 nw
tri 27249 21873 27279 21903 ne
rect 27279 21873 27283 21903
tri 27279 21869 27283 21873 ne
rect 27283 21862 27335 21868
tri 25019 21227 25032 21240 se
rect 25032 21227 25090 21240
tri 25090 21227 25103 21240 sw
tri 24998 21141 25032 21175 ne
rect 25032 21141 25088 21175
tri 25088 21141 25122 21175 nw
rect 27247 21042 27299 21048
tri 27238 21018 27247 21027 se
tri 25215 20992 25241 21018 nw
tri 27212 20992 27238 21018 se
rect 27238 20992 27247 21018
tri 27210 20990 27212 20992 se
rect 27212 20990 27247 20992
tri 27208 20988 27210 20990 se
rect 27210 20988 27299 20990
rect 23759 20982 23811 20988
tri 27206 20986 27208 20988 se
rect 27208 20986 27299 20988
tri 25735 20978 25743 20986 se
rect 25743 20978 27299 20986
tri 25730 20973 25735 20978 se
rect 25735 20973 27247 20978
tri 23811 20967 23817 20973 sw
tri 25724 20967 25730 20973 se
rect 25730 20967 27247 20973
rect 23811 20961 23817 20967
tri 23817 20961 23823 20967 sw
tri 25459 20961 25465 20967 se
rect 25465 20961 25517 20967
rect 23811 20939 23823 20961
tri 23823 20939 23845 20961 sw
tri 25437 20939 25459 20961 se
rect 25459 20939 25465 20961
rect 23811 20930 25465 20939
rect 23759 20918 25465 20930
rect 23811 20909 25465 20918
tri 25683 20926 25724 20967 se
rect 25724 20934 27247 20967
rect 25724 20926 25757 20934
tri 25757 20926 25765 20934 nw
tri 27233 20926 27241 20934 ne
rect 27241 20926 27247 20934
tri 25677 20920 25683 20926 se
rect 25683 20920 25751 20926
tri 25751 20920 25757 20926 nw
tri 27241 20920 27247 20926 ne
rect 27247 20920 27299 20926
tri 25669 20912 25677 20920 se
rect 25677 20912 25743 20920
tri 25743 20912 25751 20920 nw
rect 23811 20897 25517 20909
rect 23811 20887 25465 20897
rect 23759 20860 23811 20866
tri 23811 20860 23838 20887 nw
tri 25437 20860 25464 20887 ne
rect 25464 20860 25465 20887
tri 25464 20859 25465 20860 ne
rect 25465 20839 25517 20845
tri 25598 20841 25669 20912 se
rect 25669 20841 25672 20912
tri 25672 20841 25743 20912 nw
rect 25788 20864 25844 20873
tri 25596 20839 25598 20841 se
rect 25598 20839 25669 20841
tri 25595 20838 25596 20839 se
rect 25596 20838 25669 20839
tri 25669 20838 25672 20841 nw
tri 25588 20831 25595 20838 se
rect 25595 20831 25620 20838
tri 24777 20828 24780 20831 se
rect 24780 20828 24837 20831
tri 24837 20828 24840 20831 sw
tri 25585 20828 25588 20831 se
rect 25588 20828 25620 20831
rect 23363 20822 24414 20828
rect 23363 20770 23365 20822
rect 23417 20770 24414 20822
tri 25546 20789 25585 20828 se
rect 25585 20789 25620 20828
tri 25620 20789 25669 20838 nw
tri 25844 20847 25870 20873 sw
rect 25844 20841 27547 20847
rect 25844 20808 27495 20841
rect 25788 20789 27495 20808
tri 25534 20777 25546 20789 se
rect 25546 20777 25608 20789
tri 25608 20777 25620 20789 nw
rect 25788 20784 27547 20789
tri 25527 20770 25534 20777 se
rect 25534 20770 25601 20777
tri 25601 20770 25608 20777 nw
rect 23363 20758 24414 20770
rect 23363 20706 23365 20758
rect 23417 20706 24414 20758
tri 25383 20725 25428 20770 se
rect 25428 20725 25556 20770
tri 25556 20725 25601 20770 nw
rect 25844 20777 27547 20784
rect 25844 20728 27495 20777
rect 25788 20725 27495 20728
rect 23363 20700 24414 20706
tri 25358 20700 25383 20725 se
rect 25383 20718 25549 20725
tri 25549 20718 25556 20725 nw
rect 25788 20719 27547 20725
rect 25383 20700 25428 20718
tri 24757 20677 24780 20700 ne
rect 24780 20677 24836 20700
tri 24836 20677 24859 20700 nw
tri 25354 20696 25358 20700 se
rect 25358 20696 25428 20700
tri 25428 20696 25450 20718 nw
tri 25335 20677 25354 20696 se
tri 25323 20665 25335 20677 se
rect 25335 20665 25354 20677
rect 23125 20659 23177 20665
tri 25310 20652 25323 20665 se
rect 25323 20652 25354 20665
tri 23177 20622 23207 20652 sw
tri 25280 20622 25310 20652 se
rect 25310 20622 25354 20652
tri 25354 20622 25428 20696 nw
rect 23177 20618 23207 20622
tri 23207 20618 23211 20622 sw
tri 25276 20618 25280 20622 se
rect 25280 20618 25350 20622
tri 25350 20618 25354 20622 nw
rect 23177 20607 25298 20618
rect 23125 20595 25298 20607
rect 23177 20566 25298 20595
tri 25298 20566 25350 20618 nw
rect 23125 20537 23177 20543
tri 23177 20537 23206 20566 nw
rect 23282 20108 24906 20114
rect 23282 20056 23285 20108
rect 23337 20056 24906 20108
rect 23282 20018 24906 20056
rect 23282 19966 23285 20018
rect 23337 19966 24906 20018
rect 23282 19960 24906 19966
rect 25158 19923 25466 19932
rect 25214 19867 25410 19923
rect 25158 19843 25466 19867
rect 25214 19787 25410 19843
rect 25158 19778 25466 19787
rect 25284 19711 25718 19720
rect 25340 19655 25662 19711
rect 25284 19631 25718 19655
rect 25340 19575 25662 19631
rect 25284 19566 25718 19575
rect 25410 18583 25466 18592
rect 25410 18503 25466 18527
rect 25410 18438 25466 18447
rect 24169 18271 26557 18277
rect 24169 18219 24185 18271
rect 24237 18219 24259 18271
rect 24311 18219 24333 18271
rect 24385 18219 25307 18271
rect 25359 18219 25385 18271
rect 25437 18219 25923 18271
rect 25975 18219 26001 18271
rect 26053 18219 26336 18271
rect 26388 18219 26410 18271
rect 26462 18219 26484 18271
rect 26536 18219 26557 18271
rect 24169 18206 26557 18219
rect 24169 18154 24185 18206
rect 24237 18154 24259 18206
rect 24311 18154 24333 18206
rect 24385 18173 26336 18206
rect 24385 18154 25307 18173
rect 24169 18141 25307 18154
rect 24169 18089 24185 18141
rect 24237 18089 24259 18141
rect 24311 18089 24333 18141
rect 24385 18121 25307 18141
rect 25359 18121 25385 18173
rect 25437 18121 25923 18173
rect 25975 18121 26001 18173
rect 26053 18154 26336 18173
rect 26388 18154 26410 18206
rect 26462 18154 26484 18206
rect 26536 18154 26557 18206
rect 26053 18141 26557 18154
rect 26053 18121 26336 18141
rect 24385 18089 26336 18121
rect 26388 18089 26410 18141
rect 26462 18089 26484 18141
rect 26536 18089 26557 18141
rect 24169 18075 26557 18089
rect 24169 18023 24185 18075
rect 24237 18023 24259 18075
rect 24311 18023 24333 18075
rect 24385 18023 25307 18075
rect 25359 18023 25385 18075
rect 25437 18023 25923 18075
rect 25975 18023 26001 18075
rect 26053 18023 26336 18075
rect 26388 18023 26410 18075
rect 26462 18023 26484 18075
rect 26536 18023 26557 18075
rect 24169 18017 26557 18023
rect 23906 17846 24947 17855
rect 23906 17790 23917 17846
rect 23973 17790 24019 17846
rect 24075 17790 24121 17846
rect 24177 17790 24552 17846
rect 24608 17790 24634 17846
rect 24690 17790 24716 17846
rect 24772 17790 24798 17846
rect 24854 17790 24880 17846
rect 24936 17790 24947 17846
rect 23906 17753 24947 17790
rect 23906 17697 23917 17753
rect 23973 17697 24019 17753
rect 24075 17697 24121 17753
rect 24177 17697 24552 17753
rect 24608 17697 24634 17753
rect 24690 17697 24716 17753
rect 24772 17697 24798 17753
rect 24854 17697 24880 17753
rect 24936 17697 24947 17753
rect 23906 17660 24947 17697
rect 23906 17604 23917 17660
rect 23973 17604 24019 17660
rect 24075 17604 24121 17660
rect 24177 17604 24552 17660
rect 24608 17604 24634 17660
rect 24690 17604 24716 17660
rect 24772 17604 24798 17660
rect 24854 17604 24880 17660
rect 24936 17604 24947 17660
rect 23906 17567 24947 17604
rect 23906 17511 23917 17567
rect 23973 17511 24019 17567
rect 24075 17511 24121 17567
rect 24177 17511 24552 17567
rect 24608 17511 24634 17567
rect 24690 17511 24716 17567
rect 24772 17511 24798 17567
rect 24854 17511 24880 17567
rect 24936 17511 24947 17567
rect 23906 17473 24947 17511
rect 23906 17417 23917 17473
rect 23973 17417 24019 17473
rect 24075 17417 24121 17473
rect 24177 17417 24552 17473
rect 24608 17417 24634 17473
rect 24690 17417 24716 17473
rect 24772 17417 24798 17473
rect 24854 17417 24880 17473
rect 24936 17417 24947 17473
rect 23906 17379 24947 17417
rect 23906 17323 23917 17379
rect 23973 17323 24019 17379
rect 24075 17323 24121 17379
rect 24177 17323 24552 17379
rect 24608 17323 24634 17379
rect 24690 17323 24716 17379
rect 24772 17323 24798 17379
rect 24854 17323 24880 17379
rect 24936 17323 24947 17379
rect 23906 17314 24947 17323
rect 21049 8391 24947 8393
rect 21049 8342 24551 8391
rect 21049 8286 21060 8342
rect 21116 8286 21142 8342
rect 21198 8286 21224 8342
rect 21280 8286 21306 8342
rect 21362 8286 21388 8342
rect 21444 8286 21470 8342
rect 21526 8286 21551 8342
rect 21607 8286 21632 8342
rect 21688 8286 21713 8342
rect 21769 8286 21794 8342
rect 21850 8286 21875 8342
rect 21931 8335 24551 8342
rect 24607 8335 24634 8391
rect 24690 8335 24717 8391
rect 24773 8335 24800 8391
rect 24856 8335 24882 8391
rect 24938 8335 24947 8391
rect 21931 8305 24947 8335
rect 21931 8286 24551 8305
rect 21049 8262 24551 8286
rect 21049 8206 21060 8262
rect 21116 8206 21142 8262
rect 21198 8206 21224 8262
rect 21280 8206 21306 8262
rect 21362 8206 21388 8262
rect 21444 8206 21470 8262
rect 21526 8206 21551 8262
rect 21607 8206 21632 8262
rect 21688 8206 21713 8262
rect 21769 8206 21794 8262
rect 21850 8206 21875 8262
rect 21931 8249 24551 8262
rect 24607 8249 24634 8305
rect 24690 8249 24717 8305
rect 24773 8249 24800 8305
rect 24856 8249 24882 8305
rect 24938 8249 24947 8305
rect 21931 8219 24947 8249
rect 21931 8206 24551 8219
rect 21049 8182 24551 8206
rect 21049 8126 21060 8182
rect 21116 8126 21142 8182
rect 21198 8126 21224 8182
rect 21280 8126 21306 8182
rect 21362 8126 21388 8182
rect 21444 8126 21470 8182
rect 21526 8126 21551 8182
rect 21607 8126 21632 8182
rect 21688 8126 21713 8182
rect 21769 8126 21794 8182
rect 21850 8126 21875 8182
rect 21931 8163 24551 8182
rect 24607 8163 24634 8219
rect 24690 8163 24717 8219
rect 24773 8163 24800 8219
rect 24856 8163 24882 8219
rect 24938 8163 24947 8219
rect 21931 8133 24947 8163
rect 21931 8126 24551 8133
rect 21049 8077 24551 8126
rect 24607 8077 24634 8133
rect 24690 8077 24717 8133
rect 24773 8077 24800 8133
rect 24856 8077 24882 8133
rect 24938 8077 24947 8133
rect 21049 8075 24947 8077
rect 25284 4480 25340 4489
rect 25284 4400 25340 4424
rect 25284 4335 25340 4344
rect 25158 2793 25214 2802
rect 25158 2713 25214 2737
rect 25158 2648 25214 2657
rect 23269 2133 23385 2139
rect 23321 2081 23333 2133
rect 23269 2019 23385 2081
rect 23321 1967 23333 2019
rect 23269 1961 23385 1967
tri 23269 1949 23281 1961 ne
rect 23281 1956 23385 1961
tri 23279 1198 23281 1200 se
rect 23281 1198 23378 1956
tri 23378 1949 23385 1956 nw
rect 25764 1875 25770 1927
rect 25822 1875 25836 1927
rect 25888 1875 25894 1927
rect 25158 1723 25214 1732
tri 25138 1700 25158 1720 se
tri 25214 1700 25242 1728 sw
rect 25138 1648 25144 1700
rect 25196 1648 25208 1667
rect 25260 1648 25266 1700
tri 25138 1632 25154 1648 ne
rect 25154 1643 25214 1648
rect 25154 1632 25158 1643
tri 25214 1632 25230 1648 nw
rect 25158 1578 25214 1587
rect 25536 1212 25592 1221
tri 23248 1167 23279 1198 se
rect 23279 1167 23378 1198
rect 23248 1115 23254 1167
rect 23306 1115 23320 1167
rect 23372 1115 23378 1167
tri 25505 1167 25536 1198 se
tri 25592 1167 25633 1208 sw
rect 24139 1138 24195 1147
rect 23248 842 23378 1115
rect 24138 1125 24139 1131
rect 25505 1115 25511 1167
rect 25563 1132 25575 1156
rect 25627 1115 25633 1167
rect 25764 1167 25894 1875
rect 26857 1525 26863 1577
rect 26915 1525 26927 1577
rect 26979 1525 26985 1577
tri 26917 1497 26945 1525 ne
rect 25764 1115 25770 1167
rect 25822 1115 25836 1167
rect 25888 1115 25894 1167
rect 26945 1167 26985 1525
rect 27043 1420 27543 1421
rect 27043 1368 27049 1420
rect 27101 1416 27122 1420
rect 27174 1416 27195 1420
rect 27247 1416 27268 1420
rect 27320 1416 27341 1420
rect 27393 1416 27413 1420
rect 27465 1416 27485 1420
rect 27108 1368 27122 1416
rect 27194 1368 27195 1416
rect 27465 1368 27478 1416
rect 27537 1368 27543 1420
rect 27043 1360 27052 1368
rect 27108 1360 27138 1368
rect 27194 1360 27223 1368
rect 27279 1360 27308 1368
rect 27364 1360 27393 1368
rect 27449 1360 27478 1368
rect 27534 1360 27543 1368
rect 27043 1346 27543 1360
rect 27043 1294 27049 1346
rect 27101 1294 27122 1346
rect 27174 1294 27195 1346
rect 27247 1294 27268 1346
rect 27320 1294 27341 1346
rect 27393 1294 27413 1346
rect 27465 1294 27485 1346
rect 27537 1294 27543 1346
rect 27043 1280 27543 1294
rect 27043 1272 27052 1280
rect 27108 1272 27138 1280
rect 27194 1272 27223 1280
rect 27279 1272 27308 1280
rect 27364 1272 27393 1280
rect 27449 1272 27478 1280
rect 27534 1272 27543 1280
rect 27043 1220 27049 1272
rect 27108 1224 27122 1272
rect 27194 1224 27195 1272
rect 27465 1224 27478 1272
rect 27101 1220 27122 1224
rect 27174 1220 27195 1224
rect 27247 1220 27268 1224
rect 27320 1220 27341 1224
rect 27393 1220 27413 1224
rect 27465 1220 27485 1224
rect 27537 1220 27543 1272
rect 27043 1219 27543 1220
tri 26985 1167 26994 1176 sw
rect 26945 1158 26994 1167
tri 26945 1130 26973 1158 ne
rect 26973 1130 26994 1158
tri 26994 1130 27031 1167 sw
tri 26973 1118 26985 1130 ne
rect 26985 1118 27031 1130
tri 26985 1115 26988 1118 ne
rect 26988 1115 27031 1118
tri 27031 1115 27046 1130 sw
rect 27313 1115 27319 1167
rect 27371 1115 27383 1167
rect 27435 1115 27441 1167
tri 25505 1084 25536 1115 ne
rect 24190 1073 24195 1082
rect 24138 1061 24195 1073
tri 25592 1083 25624 1115 nw
rect 25536 1067 25592 1076
rect 24190 1058 24195 1061
rect 24138 1003 24139 1009
rect 24139 993 24195 1002
rect 24906 957 24962 966
rect 24716 919 24772 922
rect 23248 790 23254 842
rect 23306 790 23320 842
rect 23372 790 23378 842
rect 24681 913 24772 919
rect 24681 857 24716 861
rect 24681 849 24772 857
rect 24733 833 24772 849
rect 24906 877 24962 901
rect 24962 821 24977 848
rect 24906 807 24977 821
rect 24681 791 24716 797
rect 24716 768 24772 777
rect 25410 757 25466 766
tri 25374 684 25410 720 se
rect 25410 687 25466 701
tri 25466 687 25499 720 sw
rect 25410 684 25499 687
rect 23947 626 23953 678
rect 24005 626 24018 678
rect 24070 626 24076 678
rect 25371 632 25377 684
rect 25429 677 25441 684
rect 25493 632 25499 684
rect 25764 657 25894 1115
tri 26988 1072 27031 1115 ne
rect 27031 1072 27046 1115
tri 27046 1072 27089 1115 sw
tri 27031 1020 27083 1072 ne
rect 27083 1020 27092 1072
rect 27144 1020 27156 1072
rect 27208 1020 27214 1072
tri 25764 632 25789 657 ne
rect 25789 632 25894 657
tri 25894 632 25973 711 sw
rect 23947 614 24076 626
rect 23947 562 23953 614
rect 24005 562 24018 614
rect 24070 562 24076 614
tri 25390 612 25410 632 ne
rect 25410 612 25466 621
tri 25466 612 25486 632 nw
tri 25789 612 25809 632 ne
rect 25809 612 25973 632
tri 25973 612 25993 632 sw
tri 25809 598 25823 612 ne
rect 25823 598 25993 612
tri 25993 598 26007 612 sw
tri 25823 575 25846 598 ne
rect 25846 575 26007 598
rect 25662 566 25718 575
tri 25628 510 25662 544 se
tri 25846 547 25874 575 ne
rect 25874 547 26007 575
tri 25874 544 25877 547 ne
tri 25718 510 25726 518 sw
rect 25662 486 25726 510
tri 25628 430 25656 458 ne
rect 25656 430 25662 458
rect 25718 455 25726 486
tri 25718 447 25726 455 nw
tri 25656 424 25662 430 ne
rect 25662 421 25718 430
rect 25877 41 26007 547
rect 26160 518 26240 547
tri 26240 518 26269 547 nw
rect 26160 497 26219 518
tri 26219 497 26240 518 nw
rect 27043 439 27052 495
rect 27108 439 27138 495
rect 27194 439 27223 495
rect 27279 439 27308 495
rect 27364 439 27393 495
rect 27449 439 27478 495
rect 27534 439 27543 495
rect 27043 430 27543 439
rect 27043 378 27049 430
rect 27101 378 27158 430
rect 27210 378 27267 430
rect 27319 378 27376 430
rect 27428 378 27485 430
rect 27537 378 27543 430
rect 27043 359 27543 378
rect 27043 352 27052 359
rect 27043 300 27049 352
rect 27108 303 27138 359
rect 27194 352 27223 359
rect 27279 352 27308 359
rect 27364 352 27393 359
rect 27210 303 27223 352
rect 27364 303 27376 352
rect 27449 303 27478 359
rect 27534 352 27543 359
rect 27101 300 27158 303
rect 27210 300 27267 303
rect 27319 300 27376 303
rect 27428 300 27485 303
rect 27537 300 27543 352
rect 25877 -11 25883 41
rect 25935 -11 25949 41
rect 26001 -11 26007 41
rect 25158 -171 25214 -162
rect 25158 -256 25214 -227
tri 25154 -269 25158 -265 se
rect 25214 -269 25216 -265
tri 25216 -269 25220 -265 sw
rect 25158 -321 25214 -312
<< via2 >>
rect 13451 32067 13507 32123
rect 13531 32067 13587 32123
rect 3608 31904 3664 31960
rect 3608 31824 3664 31880
rect 2170 31674 2226 31730
rect 2250 31674 2306 31730
rect 3693 31666 3749 31722
rect 3773 31666 3829 31722
rect 3899 31599 3955 31655
rect 2174 31537 2230 31593
rect 2254 31537 2310 31593
rect 3899 31519 3955 31575
rect 19713 32564 19769 32620
rect 19811 32564 19867 32620
rect 19910 32564 19966 32620
rect 19359 32445 19415 32501
rect 19439 32445 19495 32501
rect 19713 32460 19769 32516
rect 19811 32460 19867 32516
rect 19910 32460 19966 32516
rect 18520 32193 18576 32249
rect 18600 32193 18656 32249
rect 14888 31517 14944 31573
rect 14970 31517 15026 31573
rect 15052 31517 15108 31573
rect 15134 31517 15190 31573
rect 15216 31517 15272 31573
rect 15298 31517 15354 31573
rect 15380 31517 15436 31573
rect 2176 31400 2232 31456
rect 2256 31400 2312 31456
rect 4025 31429 4081 31485
rect 1971 31310 2027 31366
rect 4025 31349 4081 31405
rect 14888 31436 14944 31492
rect 14970 31436 15026 31492
rect 15052 31436 15108 31492
rect 15134 31436 15190 31492
rect 15216 31436 15272 31492
rect 15298 31436 15354 31492
rect 15380 31436 15436 31492
rect 14888 31355 14944 31411
rect 14970 31355 15026 31411
rect 15052 31355 15108 31411
rect 15134 31355 15190 31411
rect 15216 31355 15272 31411
rect 15298 31355 15354 31411
rect 15380 31355 15436 31411
rect 1971 31230 2027 31286
rect 4151 31229 4207 31285
rect 4151 31149 4207 31205
rect 14888 31274 14944 31330
rect 14970 31274 15026 31330
rect 15052 31274 15108 31330
rect 15134 31274 15190 31330
rect 15216 31274 15272 31330
rect 15298 31274 15354 31330
rect 15380 31274 15436 31330
rect 14888 31193 14944 31249
rect 14970 31193 15026 31249
rect 15052 31193 15108 31249
rect 15134 31193 15190 31249
rect 15216 31193 15272 31249
rect 15298 31193 15354 31249
rect 15380 31193 15436 31249
rect 19360 31924 19416 31947
rect 19468 31924 19524 31947
rect 19575 31924 19631 31947
rect 19682 31924 19738 31947
rect 19789 31924 19845 31947
rect 19360 31891 19389 31924
rect 19389 31891 19402 31924
rect 19402 31891 19416 31924
rect 19468 31891 19519 31924
rect 19519 31891 19524 31924
rect 19575 31891 19584 31924
rect 19584 31891 19597 31924
rect 19597 31891 19631 31924
rect 19682 31891 19714 31924
rect 19714 31891 19726 31924
rect 19726 31891 19738 31924
rect 19789 31891 19790 31924
rect 19790 31891 19842 31924
rect 19842 31891 19845 31924
rect 19896 31891 19952 31947
rect 19360 31780 19416 31789
rect 19468 31780 19524 31789
rect 19575 31780 19631 31789
rect 19682 31780 19738 31789
rect 19789 31780 19845 31789
rect 19360 31733 19389 31780
rect 19389 31733 19402 31780
rect 19402 31733 19416 31780
rect 19468 31733 19519 31780
rect 19519 31733 19524 31780
rect 19575 31733 19584 31780
rect 19584 31733 19597 31780
rect 19597 31733 19631 31780
rect 19682 31733 19714 31780
rect 19714 31733 19726 31780
rect 19726 31733 19738 31780
rect 19789 31733 19790 31780
rect 19790 31733 19842 31780
rect 19842 31733 19845 31780
rect 19896 31733 19952 31789
rect 14888 31112 14944 31168
rect 14970 31112 15026 31168
rect 15052 31112 15108 31168
rect 15134 31112 15190 31168
rect 15216 31112 15272 31168
rect 15298 31112 15354 31168
rect 15380 31112 15436 31168
rect 14888 31031 14944 31087
rect 14970 31031 15026 31087
rect 15052 31031 15108 31087
rect 15134 31031 15190 31087
rect 15216 31031 15272 31087
rect 15298 31031 15354 31087
rect 15380 31031 15436 31087
rect 14888 30950 14944 31006
rect 14970 30950 15026 31006
rect 15052 30950 15108 31006
rect 15134 30950 15190 31006
rect 15216 30950 15272 31006
rect 15298 30950 15354 31006
rect 15380 30950 15436 31006
rect 14888 30868 14944 30924
rect 14970 30868 15026 30924
rect 15052 30868 15108 30924
rect 15134 30868 15190 30924
rect 15216 30868 15272 30924
rect 15298 30868 15354 30924
rect 15380 30868 15436 30924
rect 14888 30786 14944 30842
rect 14970 30786 15026 30842
rect 15052 30786 15108 30842
rect 15134 30786 15190 30842
rect 15216 30786 15272 30842
rect 15298 30786 15354 30842
rect 15380 30786 15436 30842
rect 14888 30704 14944 30760
rect 14970 30704 15026 30760
rect 15052 30704 15108 30760
rect 15134 30704 15190 30760
rect 15216 30704 15272 30760
rect 15298 30704 15354 30760
rect 15380 30704 15436 30760
rect 14888 30622 14944 30678
rect 14970 30622 15026 30678
rect 15052 30622 15108 30678
rect 15134 30622 15190 30678
rect 15216 30622 15272 30678
rect 15298 30622 15354 30678
rect 15380 30622 15436 30678
rect 20987 32594 21032 32620
rect 21032 32594 21043 32620
rect 21106 32594 21116 32620
rect 21116 32594 21148 32620
rect 21148 32594 21162 32620
rect 21225 32594 21232 32620
rect 21232 32594 21281 32620
rect 20987 32572 21043 32594
rect 21106 32572 21162 32594
rect 21225 32572 21281 32594
rect 20987 32564 21032 32572
rect 21032 32564 21043 32572
rect 21106 32564 21116 32572
rect 21116 32564 21148 32572
rect 21148 32564 21162 32572
rect 21225 32564 21232 32572
rect 21232 32564 21281 32572
rect 20987 32498 21043 32516
rect 21106 32498 21162 32516
rect 21225 32498 21281 32516
rect 20987 32460 21032 32498
rect 21032 32460 21043 32498
rect 21106 32460 21116 32498
rect 21116 32460 21148 32498
rect 21148 32460 21162 32498
rect 21225 32460 21232 32498
rect 21232 32460 21281 32498
rect 20978 31908 21034 31964
rect 21106 31908 21162 31964
rect 21234 31908 21290 31964
rect 20978 31798 21034 31854
rect 21106 31798 21162 31854
rect 21234 31798 21290 31854
rect 20978 31687 21034 31743
rect 21106 31687 21162 31743
rect 21234 31687 21290 31743
rect 20978 31576 21034 31632
rect 21106 31576 21162 31632
rect 21234 31576 21290 31632
rect 14888 30540 14944 30596
rect 14970 30540 15026 30596
rect 15052 30540 15108 30596
rect 15134 30540 15190 30596
rect 15216 30540 15272 30596
rect 15298 30540 15354 30596
rect 15380 30540 15436 30596
rect 26442 33433 26498 33489
rect 26522 33433 26578 33489
rect 26900 33433 26956 33489
rect 26980 33433 27036 33489
rect 14888 30493 14944 30514
rect 14970 30493 15026 30514
rect 15052 30493 15108 30514
rect 15134 30493 15190 30514
rect 15216 30493 15272 30514
rect 15298 30493 15354 30514
rect 15380 30493 15436 30514
rect 14888 30458 14895 30493
rect 14895 30458 14910 30493
rect 14910 30458 14944 30493
rect 14970 30458 14977 30493
rect 14977 30458 15026 30493
rect 15052 30458 15096 30493
rect 15096 30458 15108 30493
rect 15134 30458 15163 30493
rect 15163 30458 15178 30493
rect 15178 30458 15190 30493
rect 15216 30458 15230 30493
rect 15230 30458 15245 30493
rect 15245 30458 15272 30493
rect 15298 30458 15312 30493
rect 15312 30458 15354 30493
rect 15380 30458 15430 30493
rect 15430 30458 15436 30493
rect 14888 30409 14944 30432
rect 14970 30409 15026 30432
rect 15052 30409 15108 30432
rect 15134 30409 15190 30432
rect 15216 30409 15272 30432
rect 15298 30409 15354 30432
rect 15380 30409 15436 30432
rect 14888 30376 14895 30409
rect 14895 30376 14910 30409
rect 14910 30376 14944 30409
rect 14970 30376 14977 30409
rect 14977 30376 15026 30409
rect 15052 30376 15096 30409
rect 15096 30376 15108 30409
rect 15134 30376 15163 30409
rect 15163 30376 15178 30409
rect 15178 30376 15190 30409
rect 15216 30376 15230 30409
rect 15230 30376 15245 30409
rect 15245 30376 15272 30409
rect 15298 30376 15312 30409
rect 15312 30376 15354 30409
rect 15380 30376 15430 30409
rect 15430 30376 15436 30409
rect 14888 30325 14944 30350
rect 14970 30325 15026 30350
rect 15052 30325 15108 30350
rect 15134 30325 15190 30350
rect 15216 30325 15272 30350
rect 15298 30325 15354 30350
rect 15380 30325 15436 30350
rect 14888 30294 14895 30325
rect 14895 30294 14910 30325
rect 14910 30294 14944 30325
rect 14970 30294 14977 30325
rect 14977 30294 15026 30325
rect 15052 30294 15096 30325
rect 15096 30294 15108 30325
rect 15134 30294 15163 30325
rect 15163 30294 15178 30325
rect 15178 30294 15190 30325
rect 15216 30294 15230 30325
rect 15230 30294 15245 30325
rect 15245 30294 15272 30325
rect 15298 30294 15312 30325
rect 15312 30294 15354 30325
rect 15380 30294 15430 30325
rect 15430 30294 15436 30325
rect 14888 30212 14944 30268
rect 14970 30212 15026 30268
rect 15052 30212 15108 30268
rect 15134 30212 15190 30268
rect 15216 30212 15272 30268
rect 15298 30212 15354 30268
rect 15380 30212 15436 30268
rect 23275 32857 23276 32879
rect 23276 32857 23328 32879
rect 23328 32857 23331 32879
rect 23357 32857 23392 32879
rect 23392 32857 23413 32879
rect 23275 32823 23331 32857
rect 23357 32823 23413 32857
rect 25364 32749 25420 32805
rect 25506 32749 25562 32805
rect 25648 32804 25704 32805
rect 25648 32752 25663 32804
rect 25663 32752 25704 32804
rect 25648 32749 25704 32752
rect 25364 32630 25420 32686
rect 25506 32630 25562 32686
rect 25648 32674 25704 32686
rect 25648 32630 25663 32674
rect 25663 32630 25704 32674
rect 25364 32511 25420 32567
rect 25506 32511 25562 32567
rect 25648 32532 25703 32567
rect 25703 32532 25704 32567
rect 25648 32519 25704 32532
rect 25648 32511 25703 32519
rect 25703 32511 25704 32519
rect 25364 32391 25420 32447
rect 25506 32391 25562 32447
rect 25648 32402 25703 32447
rect 25703 32402 25704 32447
rect 25648 32391 25704 32402
rect 25364 32271 25420 32327
rect 25506 32271 25562 32327
rect 25648 32271 25704 32327
rect 25869 31951 25925 32007
rect 25869 31871 25925 31927
rect 27559 33241 27615 33297
rect 27559 33144 27615 33200
rect 27559 33047 27615 33103
rect 27559 32950 27615 33006
rect 26001 31951 26057 32007
rect 26001 31871 26057 31927
rect 26142 31951 26198 32007
rect 26142 31871 26198 31927
rect 27660 32038 27716 32068
rect 27773 32038 27829 32068
rect 27660 32012 27661 32038
rect 27661 32012 27689 32038
rect 27689 32012 27716 32038
rect 27773 32012 27821 32038
rect 27821 32012 27829 32038
rect 27885 32012 27941 32068
rect 27660 31962 27716 31964
rect 27773 31962 27829 31964
rect 27660 31910 27661 31962
rect 27661 31910 27689 31962
rect 27689 31910 27716 31962
rect 27773 31910 27821 31962
rect 27821 31910 27829 31962
rect 27660 31908 27716 31910
rect 27773 31908 27829 31910
rect 27885 31908 27941 31964
rect 26544 31438 26600 31454
rect 26544 31398 26546 31438
rect 26546 31398 26598 31438
rect 26598 31398 26600 31438
rect 26292 31346 26348 31362
rect 26292 31306 26294 31346
rect 26294 31306 26346 31346
rect 26346 31306 26348 31346
rect 26544 31322 26546 31374
rect 26546 31322 26598 31374
rect 26598 31322 26600 31374
rect 26544 31318 26600 31322
rect 26292 31230 26294 31282
rect 26294 31230 26346 31282
rect 26346 31230 26348 31282
rect 26292 31226 26348 31230
rect 26796 31240 26852 31256
rect 26796 31200 26798 31240
rect 26798 31200 26850 31240
rect 26850 31200 26852 31240
rect 26796 31124 26798 31176
rect 26798 31124 26850 31176
rect 26850 31124 26852 31176
rect 26796 31120 26852 31124
rect 26922 31096 26978 31112
rect 24402 30995 24458 31051
rect 26922 31056 26924 31096
rect 26924 31056 26976 31096
rect 26976 31056 26978 31096
rect 26922 30980 26924 31032
rect 26924 30980 26976 31032
rect 26976 30980 26978 31032
rect 24402 30915 24458 30971
rect 26670 30955 26726 30971
rect 26922 30976 26978 30980
rect 26670 30915 26672 30955
rect 26672 30915 26724 30955
rect 26724 30915 26726 30955
rect 26418 30868 26474 30884
rect 26418 30828 26420 30868
rect 26420 30828 26472 30868
rect 26472 30828 26474 30868
rect 26670 30839 26672 30891
rect 26672 30839 26724 30891
rect 26724 30839 26726 30891
rect 26670 30835 26726 30839
rect 26418 30752 26420 30804
rect 26420 30752 26472 30804
rect 26472 30752 26474 30804
rect 26418 30748 26474 30752
rect 24164 30639 24220 30695
rect 24268 30639 24324 30695
rect 24164 30587 24220 30600
rect 24268 30587 24324 30600
rect 24164 30544 24216 30587
rect 24216 30544 24220 30587
rect 24268 30544 24286 30587
rect 24286 30544 24304 30587
rect 24304 30544 24324 30587
rect 24164 30471 24216 30505
rect 24216 30471 24220 30505
rect 24268 30471 24286 30505
rect 24286 30471 24304 30505
rect 24304 30471 24324 30505
rect 24164 30459 24220 30471
rect 24268 30459 24324 30471
rect 24164 30449 24216 30459
rect 24216 30449 24220 30459
rect 24268 30449 24286 30459
rect 24286 30449 24304 30459
rect 24304 30449 24324 30459
rect 24164 30407 24216 30410
rect 24216 30407 24220 30410
rect 24268 30407 24286 30410
rect 24286 30407 24304 30410
rect 24304 30407 24324 30410
rect 24164 30395 24220 30407
rect 24268 30395 24324 30407
rect 24164 30354 24216 30395
rect 24216 30354 24220 30395
rect 24268 30354 24286 30395
rect 24286 30354 24304 30395
rect 24304 30354 24324 30395
rect 25732 30219 25788 30275
rect 25732 30139 25788 30195
rect 25410 29666 25466 29722
rect 25410 29586 25466 29642
rect 23765 28804 23821 28860
rect 24261 28804 24317 28860
rect 23765 28724 23821 28780
rect 24261 28724 24317 28780
rect 25536 28429 25592 28485
rect 25536 28349 25592 28405
rect 24528 23504 24584 23560
rect 24528 23406 24584 23462
rect 25788 20808 25844 20864
rect 25788 20728 25844 20784
rect 25158 19867 25214 19923
rect 25410 19867 25466 19923
rect 25158 19787 25214 19843
rect 25410 19787 25466 19843
rect 25284 19655 25340 19711
rect 25662 19655 25718 19711
rect 25284 19575 25340 19631
rect 25662 19575 25718 19631
rect 25410 18527 25466 18583
rect 25410 18447 25466 18503
rect 23917 17790 23973 17846
rect 24019 17790 24075 17846
rect 24121 17790 24177 17846
rect 24552 17790 24608 17846
rect 24634 17790 24690 17846
rect 24716 17790 24772 17846
rect 24798 17790 24854 17846
rect 24880 17790 24936 17846
rect 23917 17697 23973 17753
rect 24019 17697 24075 17753
rect 24121 17697 24177 17753
rect 24552 17697 24608 17753
rect 24634 17697 24690 17753
rect 24716 17697 24772 17753
rect 24798 17697 24854 17753
rect 24880 17697 24936 17753
rect 23917 17604 23973 17660
rect 24019 17604 24075 17660
rect 24121 17604 24177 17660
rect 24552 17604 24608 17660
rect 24634 17604 24690 17660
rect 24716 17604 24772 17660
rect 24798 17604 24854 17660
rect 24880 17604 24936 17660
rect 23917 17511 23973 17567
rect 24019 17511 24075 17567
rect 24121 17511 24177 17567
rect 24552 17511 24608 17567
rect 24634 17511 24690 17567
rect 24716 17511 24772 17567
rect 24798 17511 24854 17567
rect 24880 17511 24936 17567
rect 23917 17417 23973 17473
rect 24019 17417 24075 17473
rect 24121 17417 24177 17473
rect 24552 17417 24608 17473
rect 24634 17417 24690 17473
rect 24716 17417 24772 17473
rect 24798 17417 24854 17473
rect 24880 17417 24936 17473
rect 23917 17323 23973 17379
rect 24019 17323 24075 17379
rect 24121 17323 24177 17379
rect 24552 17323 24608 17379
rect 24634 17323 24690 17379
rect 24716 17323 24772 17379
rect 24798 17323 24854 17379
rect 24880 17323 24936 17379
rect 21060 8286 21116 8342
rect 21142 8286 21198 8342
rect 21224 8286 21280 8342
rect 21306 8286 21362 8342
rect 21388 8286 21444 8342
rect 21470 8286 21526 8342
rect 21551 8286 21607 8342
rect 21632 8286 21688 8342
rect 21713 8286 21769 8342
rect 21794 8286 21850 8342
rect 21875 8286 21931 8342
rect 24551 8335 24607 8391
rect 24634 8335 24690 8391
rect 24717 8335 24773 8391
rect 24800 8335 24856 8391
rect 24882 8335 24938 8391
rect 21060 8206 21116 8262
rect 21142 8206 21198 8262
rect 21224 8206 21280 8262
rect 21306 8206 21362 8262
rect 21388 8206 21444 8262
rect 21470 8206 21526 8262
rect 21551 8206 21607 8262
rect 21632 8206 21688 8262
rect 21713 8206 21769 8262
rect 21794 8206 21850 8262
rect 21875 8206 21931 8262
rect 24551 8249 24607 8305
rect 24634 8249 24690 8305
rect 24717 8249 24773 8305
rect 24800 8249 24856 8305
rect 24882 8249 24938 8305
rect 21060 8126 21116 8182
rect 21142 8126 21198 8182
rect 21224 8126 21280 8182
rect 21306 8126 21362 8182
rect 21388 8126 21444 8182
rect 21470 8126 21526 8182
rect 21551 8126 21607 8182
rect 21632 8126 21688 8182
rect 21713 8126 21769 8182
rect 21794 8126 21850 8182
rect 21875 8126 21931 8182
rect 24551 8163 24607 8219
rect 24634 8163 24690 8219
rect 24717 8163 24773 8219
rect 24800 8163 24856 8219
rect 24882 8163 24938 8219
rect 24551 8077 24607 8133
rect 24634 8077 24690 8133
rect 24717 8077 24773 8133
rect 24800 8077 24856 8133
rect 24882 8077 24938 8133
rect 25284 4424 25340 4480
rect 25284 4344 25340 4400
rect 25158 2737 25214 2793
rect 25158 2657 25214 2713
rect 25158 1700 25214 1723
rect 25158 1667 25196 1700
rect 25196 1667 25208 1700
rect 25208 1667 25214 1700
rect 25158 1587 25214 1643
rect 25536 1167 25592 1212
rect 24139 1125 24195 1138
rect 24139 1082 24190 1125
rect 24190 1082 24195 1125
rect 25536 1156 25563 1167
rect 25563 1156 25575 1167
rect 25575 1156 25592 1167
rect 25536 1115 25563 1132
rect 25563 1115 25575 1132
rect 25575 1115 25592 1132
rect 27052 1368 27101 1416
rect 27101 1368 27108 1416
rect 27138 1368 27174 1416
rect 27174 1368 27194 1416
rect 27223 1368 27247 1416
rect 27247 1368 27268 1416
rect 27268 1368 27279 1416
rect 27308 1368 27320 1416
rect 27320 1368 27341 1416
rect 27341 1368 27364 1416
rect 27393 1368 27413 1416
rect 27413 1368 27449 1416
rect 27478 1368 27485 1416
rect 27485 1368 27534 1416
rect 27052 1360 27108 1368
rect 27138 1360 27194 1368
rect 27223 1360 27279 1368
rect 27308 1360 27364 1368
rect 27393 1360 27449 1368
rect 27478 1360 27534 1368
rect 27052 1272 27108 1280
rect 27138 1272 27194 1280
rect 27223 1272 27279 1280
rect 27308 1272 27364 1280
rect 27393 1272 27449 1280
rect 27478 1272 27534 1280
rect 27052 1224 27101 1272
rect 27101 1224 27108 1272
rect 27138 1224 27174 1272
rect 27174 1224 27194 1272
rect 27223 1224 27247 1272
rect 27247 1224 27268 1272
rect 27268 1224 27279 1272
rect 27308 1224 27320 1272
rect 27320 1224 27341 1272
rect 27341 1224 27364 1272
rect 27393 1224 27413 1272
rect 27413 1224 27449 1272
rect 27478 1224 27485 1272
rect 27485 1224 27534 1272
rect 25536 1076 25592 1115
rect 24139 1009 24190 1058
rect 24190 1009 24195 1058
rect 24139 1002 24195 1009
rect 24716 861 24733 913
rect 24733 861 24772 913
rect 24716 857 24772 861
rect 24716 797 24733 833
rect 24733 797 24772 833
rect 24906 901 24962 957
rect 24906 821 24962 877
rect 24716 777 24772 797
rect 25410 701 25466 757
rect 25410 632 25429 677
rect 25429 632 25441 677
rect 25441 632 25466 677
rect 25410 621 25466 632
rect 25662 510 25718 566
rect 25662 430 25718 486
rect 27052 439 27108 495
rect 27138 439 27194 495
rect 27223 439 27279 495
rect 27308 439 27364 495
rect 27393 439 27449 495
rect 27478 439 27534 495
rect 27052 352 27108 359
rect 27052 303 27101 352
rect 27101 303 27108 352
rect 27138 352 27194 359
rect 27223 352 27279 359
rect 27308 352 27364 359
rect 27393 352 27449 359
rect 27138 303 27158 352
rect 27158 303 27194 352
rect 27223 303 27267 352
rect 27267 303 27279 352
rect 27308 303 27319 352
rect 27319 303 27364 352
rect 27393 303 27428 352
rect 27428 303 27449 352
rect 27478 352 27534 359
rect 27478 303 27485 352
rect 27485 303 27534 352
rect 25158 -227 25214 -171
rect 25158 -312 25214 -256
<< metal3 >>
rect 26437 33489 27041 33494
rect 26437 33433 26442 33489
rect 26498 33433 26522 33489
rect 26578 33433 26900 33489
rect 26956 33433 26980 33489
rect 27036 33433 27041 33489
rect 26437 33428 27041 33433
tri 4090 33384 4115 33409 se
rect 4115 33384 15530 33409
tri 15530 33384 15555 33409 sw
tri 4021 33315 4090 33384 se
rect 4090 33343 15555 33384
rect 4090 33315 4115 33343
tri 4115 33315 4143 33343 nw
tri 15502 33315 15530 33343 ne
rect 15530 33315 15555 33343
tri 4003 33297 4021 33315 se
rect 4021 33297 4097 33315
tri 4097 33297 4115 33315 nw
tri 15530 33297 15548 33315 ne
rect 15548 33312 15555 33315
tri 15555 33312 15627 33384 sw
rect 15548 33297 15627 33312
tri 15627 33297 15642 33312 sw
rect 27512 33297 27999 33312
tri 3996 33290 4003 33297 se
rect 4003 33290 4090 33297
tri 4090 33290 4097 33297 nw
tri 15548 33290 15555 33297 ne
rect 15555 33290 15642 33297
tri 15642 33290 15649 33297 sw
tri 3989 33283 3996 33290 se
rect 3996 33283 4083 33290
tri 4083 33283 4090 33290 nw
tri 15555 33283 15562 33290 ne
rect 15562 33283 15649 33290
tri 15649 33283 15656 33290 sw
tri 3964 33258 3989 33283 se
rect 3989 33258 4058 33283
tri 4058 33258 4083 33283 nw
tri 4144 33258 4169 33283 se
rect 4169 33258 15476 33283
tri 15476 33258 15501 33283 sw
tri 15562 33258 15587 33283 ne
rect 15587 33258 15656 33283
tri 15656 33258 15681 33283 sw
tri 3947 33241 3964 33258 se
rect 3964 33241 4041 33258
tri 4041 33241 4058 33258 nw
tri 4127 33241 4144 33258 se
rect 4144 33241 15501 33258
tri 15501 33241 15518 33258 sw
tri 15587 33241 15604 33258 ne
rect 15604 33241 15681 33258
tri 15681 33241 15698 33258 sw
rect 27512 33241 27559 33297
rect 27615 33241 27999 33297
tri 3927 33221 3947 33241 se
rect 3947 33229 4029 33241
tri 4029 33229 4041 33241 nw
tri 4115 33229 4127 33241 se
rect 4127 33229 15518 33241
rect 3947 33221 4021 33229
tri 4021 33221 4029 33229 nw
tri 4107 33221 4115 33229 se
rect 4115 33221 15518 33229
tri 3906 33200 3927 33221 se
rect 3927 33200 4000 33221
tri 4000 33200 4021 33221 nw
tri 4086 33200 4107 33221 se
rect 4107 33217 15518 33221
rect 4107 33200 4180 33217
tri 4180 33200 4197 33217 nw
tri 15448 33200 15465 33217 ne
rect 15465 33204 15518 33217
tri 15518 33204 15555 33241 sw
tri 15604 33204 15641 33241 ne
rect 15641 33204 15698 33241
rect 15465 33200 15555 33204
tri 15555 33200 15559 33204 sw
tri 15641 33200 15645 33204 ne
rect 15645 33200 15698 33204
tri 15698 33200 15739 33241 sw
rect 27512 33200 27999 33241
tri 3895 33189 3906 33200 se
rect 3906 33189 3989 33200
tri 3989 33189 4000 33200 nw
tri 4075 33189 4086 33200 se
rect 4086 33189 4169 33200
tri 4169 33189 4180 33200 nw
tri 15465 33189 15476 33200 ne
rect 15476 33196 15559 33200
tri 15559 33196 15563 33200 sw
tri 15645 33196 15649 33200 ne
rect 15649 33196 15739 33200
tri 15739 33196 15743 33200 sw
rect 15476 33189 15563 33196
tri 3870 33164 3895 33189 se
rect 3895 33164 3964 33189
tri 3964 33164 3989 33189 nw
tri 4050 33164 4075 33189 se
rect 4075 33164 4144 33189
tri 4144 33164 4169 33189 nw
tri 15476 33164 15501 33189 ne
rect 15501 33164 15563 33189
tri 15563 33164 15595 33196 sw
tri 15649 33164 15681 33196 ne
rect 15681 33164 15743 33196
tri 15743 33164 15775 33196 sw
tri 3863 33157 3870 33164 se
rect 3870 33157 3957 33164
tri 3957 33157 3964 33164 nw
tri 4043 33157 4050 33164 se
rect 4050 33157 4137 33164
tri 4137 33157 4144 33164 nw
tri 15501 33157 15508 33164 ne
rect 15508 33157 15595 33164
tri 15595 33157 15602 33164 sw
tri 15681 33157 15688 33164 ne
rect 15688 33157 15775 33164
tri 15775 33157 15782 33164 sw
tri 3850 33144 3863 33157 se
rect 3863 33144 3944 33157
tri 3944 33144 3957 33157 nw
tri 4030 33144 4043 33157 se
rect 4043 33144 4124 33157
tri 4124 33144 4137 33157 nw
tri 4210 33144 4223 33157 se
rect 4223 33144 15422 33157
tri 15422 33144 15435 33157 sw
tri 15508 33144 15521 33157 ne
rect 15521 33144 15602 33157
tri 15602 33144 15615 33157 sw
tri 15688 33144 15701 33157 ne
rect 15701 33144 15782 33157
tri 15782 33144 15795 33157 sw
rect 27512 33144 27559 33200
rect 27615 33144 27999 33200
tri 3838 33132 3850 33144 se
rect 3850 33135 3935 33144
tri 3935 33135 3944 33144 nw
tri 4021 33135 4030 33144 se
rect 4030 33135 4112 33144
rect 3850 33132 3932 33135
tri 3932 33132 3935 33135 nw
tri 4018 33132 4021 33135 se
rect 4021 33132 4112 33135
tri 4112 33132 4124 33144 nw
tri 4198 33132 4210 33144 se
rect 4210 33132 15435 33144
tri 15435 33132 15447 33144 sw
tri 15521 33132 15533 33144 ne
rect 15533 33132 15615 33144
tri 15615 33132 15627 33144 sw
tri 15701 33132 15713 33144 ne
rect 15713 33132 15795 33144
tri 15795 33132 15807 33144 sw
tri 3833 33127 3838 33132 se
rect 3838 33127 3927 33132
tri 3927 33127 3932 33132 nw
tri 4013 33127 4018 33132 se
rect 4018 33127 4083 33132
tri 3809 33103 3833 33127 se
rect 3833 33103 3903 33127
tri 3903 33103 3927 33127 nw
tri 3989 33103 4013 33127 se
rect 4013 33103 4083 33127
tri 4083 33103 4112 33132 nw
tri 4169 33103 4198 33132 se
rect 4198 33103 15447 33132
tri 15447 33103 15476 33132 sw
tri 15533 33103 15562 33132 ne
rect 15562 33110 15627 33132
tri 15627 33110 15649 33132 sw
tri 15713 33110 15735 33132 ne
rect 15735 33110 15807 33132
rect 15562 33103 15649 33110
tri 15649 33103 15656 33110 sw
tri 15735 33103 15742 33110 ne
rect 15742 33103 15807 33110
tri 15807 33103 15836 33132 sw
rect 27512 33103 27999 33144
tri 3801 33095 3809 33103 se
rect 3809 33095 3895 33103
tri 3895 33095 3903 33103 nw
tri 3981 33095 3989 33103 se
rect 3989 33095 4075 33103
tri 4075 33095 4083 33103 nw
tri 4161 33095 4169 33103 se
rect 4169 33095 15476 33103
tri 3772 33066 3801 33095 se
rect 3801 33066 3866 33095
tri 3866 33066 3895 33095 nw
tri 3952 33066 3981 33095 se
rect 3981 33066 4043 33095
rect 3772 33063 3863 33066
tri 3863 33063 3866 33066 nw
tri 3949 33063 3952 33066 se
rect 3952 33063 4043 33066
tri 4043 33063 4075 33095 nw
tri 4129 33063 4161 33095 se
rect 4161 33091 15476 33095
rect 4161 33063 4223 33091
tri 4223 33063 4251 33091 nw
tri 15394 33063 15422 33091 ne
rect 15422 33078 15476 33091
tri 15476 33078 15501 33103 sw
tri 15562 33078 15587 33103 ne
rect 15587 33102 15656 33103
tri 15656 33102 15657 33103 sw
tri 15742 33102 15743 33103 ne
rect 15743 33102 15836 33103
tri 15836 33102 15837 33103 sw
rect 15587 33078 15657 33102
rect 15422 33070 15501 33078
tri 15501 33070 15509 33078 sw
tri 15587 33070 15595 33078 ne
rect 15595 33070 15657 33078
tri 15657 33070 15689 33102 sw
tri 15743 33070 15775 33102 ne
rect 15775 33070 15837 33102
tri 15837 33070 15869 33102 sw
rect 15422 33063 15509 33070
rect 3772 33047 3847 33063
tri 3847 33047 3863 33063 nw
tri 3933 33047 3949 33063 se
rect 3949 33047 4027 33063
tri 4027 33047 4043 33063 nw
tri 4113 33047 4129 33063 se
rect 4129 33047 4207 33063
tri 4207 33047 4223 33063 nw
tri 15422 33047 15438 33063 ne
rect 15438 33047 15509 33063
tri 15509 33047 15532 33070 sw
tri 15595 33047 15618 33070 ne
rect 15618 33047 15689 33070
tri 15689 33047 15712 33070 sw
tri 15775 33047 15798 33070 ne
rect 15798 33047 15869 33070
tri 15869 33047 15892 33070 sw
rect 27512 33047 27559 33103
rect 27615 33047 27999 33103
rect 3772 33041 3841 33047
tri 3841 33041 3847 33047 nw
tri 3927 33041 3933 33047 se
rect 3933 33041 4018 33047
rect 3772 33038 3838 33041
tri 3838 33038 3841 33041 nw
tri 3924 33038 3927 33041 se
rect 3927 33038 4018 33041
tri 4018 33038 4027 33047 nw
tri 4104 33038 4113 33047 se
rect 4113 33038 4198 33047
tri 4198 33038 4207 33047 nw
tri 15438 33038 15447 33047 ne
rect 15447 33038 15532 33047
tri 15532 33038 15541 33047 sw
tri 15618 33038 15627 33047 ne
rect 15627 33038 15712 33047
tri 15712 33038 15721 33047 sw
tri 15798 33038 15807 33047 ne
rect 15807 33038 15892 33047
tri 15892 33038 15901 33047 sw
rect 3603 31960 3669 31965
rect 3603 31904 3608 31960
rect 3664 31904 3669 31960
rect 3603 31880 3669 31904
rect 3603 31824 3608 31880
rect 3664 31824 3669 31880
rect 3603 31819 3669 31824
tri 3759 31798 3772 31811 se
rect 3772 31798 3834 33038
tri 3834 33034 3838 33038 nw
tri 3920 33034 3924 33038 se
rect 3924 33034 4011 33038
tri 3917 33031 3920 33034 se
rect 3920 33031 4011 33034
tri 4011 33031 4018 33038 nw
tri 4097 33031 4104 33038 se
rect 4104 33031 4191 33038
tri 4191 33031 4198 33038 nw
tri 15447 33031 15454 33038 ne
rect 15454 33031 15541 33038
tri 15541 33031 15548 33038 sw
tri 15627 33031 15634 33038 ne
rect 15634 33031 15721 33038
tri 15721 33031 15728 33038 sw
tri 15807 33031 15814 33038 ne
rect 15814 33031 15901 33038
tri 15901 33031 15908 33038 sw
tri 3750 31789 3759 31798 se
rect 3759 31789 3834 31798
tri 3696 31735 3750 31789 se
rect 3750 31735 3834 31789
tri 1770 31733 1772 31735 se
rect 1772 31733 2311 31735
tri 3694 31733 3696 31735 se
rect 3696 31733 3834 31735
tri 1767 31730 1770 31733 se
rect 1770 31730 2311 31733
tri 1719 31682 1767 31730 se
rect 1767 31682 2170 31730
tri 1714 31677 1719 31682 se
rect 1719 31677 2170 31682
rect 1714 31674 2170 31677
rect 2226 31674 2250 31730
rect 2306 31674 2311 31730
rect 1714 31669 2311 31674
tri 3688 31727 3694 31733 se
rect 3694 31727 3834 31733
rect 3688 31722 3834 31727
rect 1714 31666 1848 31669
tri 1848 31666 1851 31669 nw
rect 3688 31666 3693 31722
rect 3749 31666 3773 31722
rect 3829 31666 3834 31722
rect 1714 31655 1837 31666
tri 1837 31655 1848 31666 nw
rect 3688 31661 3834 31666
tri 3898 33012 3917 33031 se
rect 3917 33012 3992 33031
tri 3992 33012 4011 33031 nw
tri 4078 33012 4097 33031 se
rect 4097 33012 4166 33031
rect 3898 33006 3986 33012
tri 3986 33006 3992 33012 nw
tri 4072 33006 4078 33012 se
rect 4078 33006 4166 33012
tri 4166 33006 4191 33031 nw
tri 4346 33006 4371 33031 se
rect 4371 33006 15368 33031
tri 15368 33006 15393 33031 sw
tri 15454 33006 15479 33031 ne
rect 15479 33006 15548 33031
tri 15548 33006 15573 33031 sw
tri 15634 33006 15659 33031 ne
rect 15659 33016 15728 33031
tri 15728 33016 15743 33031 sw
tri 15814 33016 15829 33031 ne
rect 15829 33016 15908 33031
rect 15659 33008 15743 33016
tri 15743 33008 15751 33016 sw
tri 15829 33008 15837 33016 ne
rect 15837 33008 15908 33016
tri 15908 33008 15931 33031 sw
rect 15659 33006 15751 33008
tri 15751 33006 15753 33008 sw
tri 15837 33006 15839 33008 ne
rect 15839 33006 15931 33008
tri 15931 33006 15933 33008 sw
rect 27512 33006 27999 33047
tri 3895 31661 3898 31664 se
rect 3898 31661 3960 33006
tri 3960 32980 3986 33006 nw
tri 4046 32980 4072 33006 se
rect 4072 32980 4129 33006
tri 4035 32969 4046 32980 se
rect 4046 32969 4129 32980
tri 4129 32969 4166 33006 nw
tri 4309 32969 4346 33006 se
rect 4346 32969 15393 33006
tri 3894 31660 3895 31661 se
rect 3895 31660 3960 31661
rect 3894 31655 3960 31660
rect 1714 31599 1781 31655
tri 1781 31599 1837 31655 nw
rect 3894 31599 3899 31655
rect 3955 31599 3960 31655
tri 1707 31230 1714 31237 se
rect 1714 31230 1780 31599
tri 1780 31598 1781 31599 nw
tri 1891 31593 1896 31598 se
rect 1896 31593 2315 31598
tri 1706 31229 1707 31230 se
rect 1707 31229 1780 31230
tri 1682 31205 1706 31229 se
rect 1706 31209 1780 31229
rect 1706 31205 1776 31209
tri 1776 31205 1780 31209 nw
tri 1840 31542 1891 31593 se
rect 1891 31542 2174 31593
rect 1840 31537 2174 31542
rect 2230 31537 2254 31593
rect 2310 31537 2315 31593
rect 1840 31532 2315 31537
rect 3894 31575 3960 31599
rect 1840 31519 1946 31532
tri 1946 31519 1959 31532 nw
rect 3894 31519 3899 31575
rect 3955 31519 3960 31575
rect 1840 31517 1944 31519
tri 1944 31517 1946 31519 nw
rect 1840 31514 1941 31517
tri 1941 31514 1944 31517 nw
rect 3894 31514 3960 31519
tri 4020 32954 4035 32969 se
rect 4035 32954 4114 32969
tri 4114 32954 4129 32969 nw
tri 4294 32954 4309 32969 se
rect 4309 32965 15393 32969
rect 4309 32954 4404 32965
rect 4020 32950 4110 32954
tri 4110 32950 4114 32954 nw
tri 4290 32950 4294 32954 se
rect 4294 32950 4404 32954
tri 4404 32950 4419 32965 nw
tri 15340 32950 15355 32965 ne
rect 15355 32952 15393 32965
tri 15393 32952 15447 33006 sw
tri 15479 32952 15533 33006 ne
rect 15533 32984 15573 33006
tri 15573 32984 15595 33006 sw
tri 15659 32984 15681 33006 ne
rect 15681 32984 15753 33006
rect 15533 32976 15595 32984
tri 15595 32976 15603 32984 sw
tri 15681 32976 15689 32984 ne
rect 15689 32976 15753 32984
tri 15753 32976 15783 33006 sw
tri 15839 32976 15869 33006 ne
rect 15869 32976 15933 33006
tri 15933 32976 15963 33006 sw
rect 15533 32952 15603 32976
rect 15355 32950 15447 32952
tri 15447 32950 15449 32952 sw
tri 15533 32950 15535 32952 ne
rect 15535 32950 15603 32952
tri 15603 32950 15629 32976 sw
tri 15689 32950 15715 32976 ne
rect 15715 32950 15783 32976
tri 15783 32950 15809 32976 sw
tri 15869 32950 15895 32976 ne
rect 15895 32950 15963 32976
tri 15963 32950 15989 32976 sw
rect 27512 32950 27559 33006
rect 27615 32950 27999 33006
rect 1840 31492 1919 31514
tri 1919 31492 1941 31514 nw
rect 1840 31485 1912 31492
tri 1912 31485 1919 31492 nw
rect 4020 31485 4086 32950
tri 4086 32926 4110 32950 nw
tri 4266 32926 4290 32950 se
rect 4290 32926 4371 32950
tri 4257 32917 4266 32926 se
rect 4266 32917 4371 32926
tri 4371 32917 4404 32950 nw
tri 15355 32917 15388 32950 ne
rect 15388 32944 15449 32950
tri 15449 32944 15455 32950 sw
tri 15535 32944 15541 32950 ne
rect 15541 32944 15629 32950
tri 15629 32944 15635 32950 sw
tri 15715 32944 15721 32950 ne
rect 15721 32944 15809 32950
tri 15809 32944 15815 32950 sw
tri 15895 32944 15901 32950 ne
rect 15901 32944 15989 32950
tri 15989 32944 15995 32950 sw
rect 15388 32917 15455 32944
tri 4252 32912 4257 32917 se
rect 4257 32912 4366 32917
tri 4366 32912 4371 32917 nw
tri 15388 32912 15393 32917 ne
rect 15393 32912 15455 32917
tri 15455 32912 15487 32944 sw
tri 15541 32912 15573 32944 ne
rect 15573 32912 15635 32944
tri 15635 32912 15667 32944 sw
tri 15721 32912 15753 32944 ne
rect 15753 32922 15815 32944
tri 15815 32922 15837 32944 sw
tri 15901 32922 15923 32944 ne
rect 15923 32922 15995 32944
rect 15753 32914 15837 32922
tri 15837 32914 15845 32922 sw
tri 15923 32914 15931 32922 ne
rect 15931 32914 15995 32922
tri 15995 32914 16025 32944 sw
rect 27512 32939 27999 32950
tri 27512 32914 27537 32939 ne
rect 27537 32914 27999 32939
rect 15753 32912 15845 32914
tri 15845 32912 15847 32914 sw
tri 15931 32912 15933 32914 ne
rect 15933 32912 16025 32914
tri 16025 32912 16027 32914 sw
tri 27537 32912 27539 32914 ne
rect 27539 32912 27999 32914
tri 4219 32879 4252 32912 se
rect 4252 32879 4333 32912
tri 4333 32879 4366 32912 nw
tri 15393 32879 15426 32912 ne
rect 15426 32884 15487 32912
tri 15487 32884 15515 32912 sw
tri 15573 32884 15601 32912 ne
rect 15601 32890 15667 32912
tri 15667 32890 15689 32912 sw
tri 15753 32890 15775 32912 ne
rect 15775 32890 15847 32912
rect 15601 32884 15689 32890
tri 15689 32884 15695 32890 sw
tri 15775 32884 15781 32890 ne
rect 15781 32884 15847 32890
tri 15847 32884 15875 32912 sw
tri 15933 32884 15961 32912 ne
rect 15961 32884 16027 32912
tri 16027 32884 16055 32912 sw
tri 27539 32884 27567 32912 ne
rect 27567 32884 27999 32912
rect 15426 32879 15515 32884
tri 15515 32879 15520 32884 sw
tri 15601 32879 15606 32884 ne
rect 15606 32882 15695 32884
tri 15695 32882 15697 32884 sw
tri 15781 32882 15783 32884 ne
rect 15783 32882 15875 32884
tri 15875 32882 15877 32884 sw
tri 15961 32882 15963 32884 ne
rect 15963 32882 16055 32884
tri 16055 32882 16057 32884 sw
rect 15606 32879 15697 32882
tri 15697 32879 15700 32882 sw
tri 15783 32879 15786 32882 ne
rect 15786 32879 15877 32882
tri 15877 32879 15880 32882 sw
tri 15963 32879 15966 32882 ne
rect 15966 32879 16057 32882
tri 16057 32879 16060 32882 sw
rect 23270 32879 23418 32884
tri 4163 32823 4219 32879 se
rect 4219 32823 4277 32879
tri 4277 32823 4333 32879 nw
tri 15426 32823 15482 32879 ne
rect 15482 32858 15520 32879
tri 15520 32858 15541 32879 sw
tri 15606 32858 15627 32879 ne
rect 15627 32858 15700 32879
rect 15482 32850 15541 32858
tri 15541 32850 15549 32858 sw
tri 15627 32850 15635 32858 ne
rect 15635 32850 15700 32858
tri 15700 32850 15729 32879 sw
tri 15786 32850 15815 32879 ne
rect 15815 32850 15880 32879
tri 15880 32850 15909 32879 sw
tri 15966 32850 15995 32879 ne
rect 15995 32850 16060 32879
tri 16060 32850 16089 32879 sw
rect 15482 32823 15549 32850
tri 15549 32823 15576 32850 sw
tri 15635 32823 15662 32850 ne
rect 15662 32823 15729 32850
tri 15729 32823 15756 32850 sw
tri 15815 32823 15842 32850 ne
rect 15842 32828 15909 32850
tri 15909 32828 15931 32850 sw
tri 15995 32828 16017 32850 ne
rect 16017 32828 16089 32850
rect 15842 32823 15931 32828
tri 15931 32823 15936 32828 sw
tri 16017 32823 16022 32828 ne
rect 16022 32823 16089 32828
tri 16089 32823 16116 32850 sw
rect 23270 32823 23275 32879
rect 23331 32823 23357 32879
rect 23413 32823 23418 32879
tri 4158 32818 4163 32823 se
rect 4163 32818 4272 32823
tri 4272 32818 4277 32823 nw
tri 15482 32818 15487 32823 ne
rect 15487 32818 15576 32823
tri 15576 32818 15581 32823 sw
tri 15662 32818 15667 32823 ne
rect 15667 32818 15756 32823
tri 15756 32818 15761 32823 sw
tri 15842 32818 15847 32823 ne
rect 15847 32820 15936 32823
tri 15936 32820 15939 32823 sw
tri 16022 32820 16025 32823 ne
rect 16025 32820 16116 32823
tri 16116 32820 16119 32823 sw
rect 15847 32818 15939 32820
tri 15939 32818 15941 32820 sw
tri 16025 32818 16027 32820 ne
rect 16027 32818 16119 32820
tri 16119 32818 16121 32820 sw
rect 23270 32818 23418 32823
tri 27567 32819 27632 32884 ne
rect 27632 32819 27999 32884
tri 1626 31149 1682 31205 se
rect 1682 31183 1754 31205
tri 1754 31183 1776 31205 nw
rect 1682 31175 1746 31183
tri 1746 31175 1754 31183 nw
tri 1832 31175 1840 31183 se
rect 1840 31175 1906 31485
tri 1906 31479 1912 31485 nw
rect 2171 31456 2317 31461
rect 2171 31400 2176 31456
rect 2232 31400 2256 31456
rect 2312 31400 2317 31456
rect 2171 31395 2317 31400
rect 4020 31429 4025 31485
rect 4081 31429 4086 31485
rect 4020 31405 4086 31429
rect 1682 31149 1720 31175
tri 1720 31149 1746 31175 nw
tri 1806 31149 1832 31175 se
rect 1832 31155 1906 31175
rect 1832 31149 1900 31155
tri 1900 31149 1906 31155 nw
rect 1966 31366 2032 31371
rect 1966 31310 1971 31366
rect 2027 31310 2032 31366
rect 1966 31286 2032 31310
rect 1966 31230 1971 31286
rect 2027 31230 2032 31286
tri 1620 31143 1626 31149 se
rect 1626 31143 1714 31149
tri 1714 31143 1720 31149 nw
tri 1800 31143 1806 31149 se
rect 1806 31143 1880 31149
tri 1589 31112 1620 31143 se
rect 1620 31112 1683 31143
tri 1683 31112 1714 31143 nw
tri 1786 31129 1800 31143 se
rect 1800 31129 1880 31143
tri 1880 31129 1900 31149 nw
tri 1769 31112 1786 31129 se
rect 1786 31112 1863 31129
tri 1863 31112 1880 31129 nw
tri 1949 31112 1966 31129 se
rect 1966 31112 2032 31230
tri 1564 31087 1589 31112 se
rect 1589 31089 1660 31112
tri 1660 31089 1683 31112 nw
tri 1746 31089 1769 31112 se
rect 1769 31089 1840 31112
tri 1840 31089 1863 31112 nw
tri 1926 31089 1949 31112 se
rect 1949 31101 2032 31112
rect 1949 31089 2018 31101
rect 1589 31087 1658 31089
tri 1658 31087 1660 31089 nw
tri 1744 31087 1746 31089 se
rect 1746 31087 1838 31089
tri 1838 31087 1840 31089 nw
tri 1924 31087 1926 31089 se
rect 1926 31087 2018 31089
tri 2018 31087 2032 31101 nw
tri 1526 31049 1564 31087 se
rect 1564 31081 1652 31087
tri 1652 31081 1658 31087 nw
tri 1738 31081 1744 31087 se
rect 1744 31081 1800 31087
rect 1564 31049 1620 31081
tri 1620 31049 1652 31081 nw
tri 1706 31049 1738 31081 se
rect 1738 31049 1800 31081
tri 1800 31049 1838 31087 nw
tri 1886 31049 1924 31087 se
rect 1924 31049 1966 31087
tri 1508 31031 1526 31049 se
rect 1526 31031 1602 31049
tri 1602 31031 1620 31049 nw
tri 1692 31035 1706 31049 se
rect 1706 31035 1786 31049
tri 1786 31035 1800 31049 nw
tri 1872 31035 1886 31049 se
rect 1886 31035 1966 31049
tri 1966 31035 2018 31087 nw
tri 1688 31031 1692 31035 se
rect 1692 31031 1782 31035
tri 1782 31031 1786 31035 nw
tri 1868 31031 1872 31035 se
rect 1872 31031 1962 31035
tri 1962 31031 1966 31035 nw
tri 1483 31006 1508 31031 se
rect 1508 31006 1577 31031
tri 1577 31006 1602 31031 nw
tri 1663 31006 1688 31031 se
rect 1688 31006 1757 31031
tri 1757 31006 1782 31031 nw
tri 1843 31006 1868 31031 se
rect 1868 31006 1937 31031
tri 1937 31006 1962 31031 nw
tri 1432 30955 1483 31006 se
rect 1483 30995 1566 31006
tri 1566 30995 1577 31006 nw
tri 1652 30995 1663 31006 se
rect 1663 31003 1754 31006
tri 1754 31003 1757 31006 nw
tri 1840 31003 1843 31006 se
rect 1843 31003 1881 31006
rect 1663 30995 1746 31003
tri 1746 30995 1754 31003 nw
tri 1832 30995 1840 31003 se
rect 1840 30995 1881 31003
rect 1483 30987 1558 30995
tri 1558 30987 1566 30995 nw
tri 1644 30987 1652 30995 se
rect 1652 30987 1706 30995
rect 1483 30955 1526 30987
tri 1526 30955 1558 30987 nw
tri 1612 30955 1644 30987 se
rect 1644 30955 1706 30987
tri 1706 30955 1746 30995 nw
tri 1792 30955 1832 30995 se
rect 1832 30955 1881 30995
tri 1427 30950 1432 30955 se
rect 1432 30950 1521 30955
tri 1521 30950 1526 30955 nw
tri 1607 30950 1612 30955 se
rect 1612 30950 1701 30955
tri 1701 30950 1706 30955 nw
tri 1787 30950 1792 30955 se
rect 1792 30950 1881 30955
tri 1881 30950 1937 31006 nw
tri 1401 30924 1427 30950 se
rect 1427 30924 1495 30950
tri 1495 30924 1521 30950 nw
tri 1598 30941 1607 30950 se
rect 1607 30941 1692 30950
tri 1692 30941 1701 30950 nw
tri 1778 30941 1787 30950 se
rect 1787 30941 1872 30950
tri 1872 30941 1881 30950 nw
tri 1581 30924 1598 30941 se
rect 1598 30924 1675 30941
tri 1675 30924 1692 30941 nw
tri 1761 30924 1778 30941 se
rect 1778 30924 1855 30941
tri 1855 30924 1872 30941 nw
tri 1345 30868 1401 30924 se
rect 1401 30901 1472 30924
tri 1472 30901 1495 30924 nw
tri 1558 30901 1581 30924 se
rect 1581 30909 1660 30924
tri 1660 30909 1675 30924 nw
tri 1746 30909 1761 30924 se
rect 1761 30909 1799 30924
rect 1581 30901 1652 30909
tri 1652 30901 1660 30909 nw
tri 1738 30901 1746 30909 se
rect 1746 30901 1799 30909
rect 1401 30893 1464 30901
tri 1464 30893 1472 30901 nw
tri 1550 30893 1558 30901 se
rect 1558 30893 1619 30901
rect 1401 30868 1439 30893
tri 1439 30868 1464 30893 nw
tri 1525 30868 1550 30893 se
rect 1550 30868 1619 30893
tri 1619 30868 1652 30901 nw
tri 1705 30868 1738 30901 se
rect 1738 30868 1799 30901
tri 1799 30868 1855 30924 nw
tri 1338 30861 1345 30868 se
rect 1345 30861 1432 30868
tri 1432 30861 1439 30868 nw
tri 1518 30861 1525 30868 se
rect 1525 30861 1612 30868
tri 1612 30861 1619 30868 nw
tri 1698 30861 1705 30868 se
rect 1705 30861 1778 30868
tri 1319 30842 1338 30861 se
rect 1338 30842 1413 30861
tri 1413 30842 1432 30861 nw
tri 1504 30847 1518 30861 se
rect 1518 30847 1598 30861
tri 1598 30847 1612 30861 nw
tri 1684 30847 1698 30861 se
rect 1698 30847 1778 30861
tri 1778 30847 1799 30868 nw
tri 1499 30842 1504 30847 se
rect 1504 30842 1593 30847
tri 1593 30842 1598 30847 nw
tri 1679 30842 1684 30847 se
rect 1684 30842 1773 30847
tri 1773 30842 1778 30847 nw
tri 1263 30786 1319 30842 se
rect 1319 30807 1378 30842
tri 1378 30807 1413 30842 nw
tri 1464 30807 1499 30842 se
rect 1499 30815 1566 30842
tri 1566 30815 1593 30842 nw
tri 1652 30815 1679 30842 se
rect 1679 30815 1717 30842
rect 1499 30807 1558 30815
tri 1558 30807 1566 30815 nw
tri 1644 30807 1652 30815 se
rect 1652 30807 1717 30815
rect 1319 30799 1370 30807
tri 1370 30799 1378 30807 nw
tri 1456 30799 1464 30807 se
rect 1464 30799 1537 30807
rect 1319 30786 1357 30799
tri 1357 30786 1370 30799 nw
tri 1443 30786 1456 30799 se
rect 1456 30786 1537 30799
tri 1537 30786 1558 30807 nw
tri 1623 30786 1644 30807 se
rect 1644 30786 1717 30807
tri 1717 30786 1773 30842 nw
tri 1244 30767 1263 30786 se
rect 1263 30767 1338 30786
tri 1338 30767 1357 30786 nw
tri 1424 30767 1443 30786 se
rect 1443 30767 1518 30786
tri 1518 30767 1537 30786 nw
tri 1604 30767 1623 30786 se
rect 1623 30767 1691 30786
tri 1237 30760 1244 30767 se
rect 1244 30760 1331 30767
tri 1331 30760 1338 30767 nw
tri 1417 30760 1424 30767 se
rect 1424 30760 1511 30767
tri 1511 30760 1518 30767 nw
tri 1597 30760 1604 30767 se
rect 1604 30760 1691 30767
tri 1691 30760 1717 30786 nw
tri 1189 30712 1237 30760 se
rect 1237 30713 1284 30760
tri 1284 30713 1331 30760 nw
tri 1410 30753 1417 30760 se
rect 1417 30753 1504 30760
tri 1504 30753 1511 30760 nw
tri 1590 30753 1597 30760 se
rect 1597 30753 1684 30760
tri 1684 30753 1691 30760 nw
tri 1370 30713 1410 30753 se
rect 1410 30721 1472 30753
tri 1472 30721 1504 30753 nw
tri 1558 30721 1590 30753 se
rect 1590 30721 1635 30753
rect 1410 30713 1464 30721
tri 1464 30713 1472 30721 nw
tri 1550 30713 1558 30721 se
rect 1558 30713 1635 30721
rect 1237 30712 1283 30713
tri 1283 30712 1284 30713 nw
tri 1369 30712 1370 30713 se
rect 1370 30712 1463 30713
tri 1463 30712 1464 30713 nw
tri 1549 30712 1550 30713 se
rect 1550 30712 1635 30713
rect 1189 30704 1275 30712
tri 1275 30704 1283 30712 nw
tri 1361 30704 1369 30712 se
rect 1369 30704 1455 30712
tri 1455 30704 1463 30712 nw
tri 1541 30704 1549 30712 se
rect 1549 30704 1635 30712
tri 1635 30704 1684 30753 nw
rect 1189 30695 1266 30704
tri 1266 30695 1275 30704 nw
tri 1352 30695 1361 30704 se
rect 1361 30695 1446 30704
tri 1446 30695 1455 30704 nw
tri 1532 30695 1541 30704 se
rect 1541 30695 1626 30704
tri 1626 30695 1635 30704 nw
rect 1189 27416 1249 30695
tri 1249 30678 1266 30695 nw
tri 1335 30678 1352 30695 se
rect 1352 30678 1429 30695
tri 1429 30678 1446 30695 nw
tri 1515 30678 1532 30695 se
rect 1532 30678 1609 30695
tri 1609 30678 1626 30695 nw
tri 1315 30658 1335 30678 se
rect 1335 30658 1409 30678
tri 1409 30658 1429 30678 nw
tri 1495 30658 1515 30678 se
rect 1515 30666 1598 30678
tri 1598 30667 1609 30678 nw
rect 1515 30658 1590 30666
tri 1590 30658 1598 30666 nw
tri 1309 30652 1315 30658 se
rect 1315 30652 1403 30658
tri 1403 30652 1409 30658 nw
tri 1489 30652 1495 30658 se
rect 1495 30652 1554 30658
rect 1309 30622 1373 30652
tri 1373 30622 1403 30652 nw
tri 1459 30622 1489 30652 se
rect 1489 30622 1554 30652
tri 1554 30622 1590 30658 nw
rect 1309 27417 1369 30622
tri 1369 30618 1373 30622 nw
tri 1455 30618 1459 30622 se
rect 1459 30618 1532 30622
tri 1437 30600 1455 30618 se
rect 1455 30600 1532 30618
tri 1532 30600 1554 30622 nw
tri 1433 30596 1437 30600 se
rect 1437 30596 1528 30600
tri 1528 30596 1532 30600 nw
tri 1429 30592 1433 30596 se
rect 1433 30592 1524 30596
tri 1524 30592 1528 30596 nw
rect 1429 27411 1489 30592
tri 1489 30557 1524 30592 nw
rect 2171 27669 2231 31395
tri 2231 31368 2258 31395 nw
rect 4020 31349 4025 31405
rect 4081 31349 4086 31405
rect 4020 31344 4086 31349
tri 4146 32806 4158 32818 se
rect 4158 32806 4260 32818
tri 4260 32806 4272 32818 nw
tri 15487 32806 15499 32818 ne
rect 15499 32806 15581 32818
rect 4146 32805 4259 32806
tri 4259 32805 4260 32806 nw
tri 15499 32805 15500 32806 ne
rect 15500 32805 15581 32806
tri 15581 32805 15594 32818 sw
tri 15667 32805 15680 32818 ne
rect 15680 32805 15761 32818
tri 15761 32805 15774 32818 sw
tri 15847 32805 15860 32818 ne
rect 15860 32805 15941 32818
tri 15941 32805 15954 32818 sw
tri 16027 32805 16040 32818 ne
rect 16040 32805 16121 32818
tri 16121 32805 16134 32818 sw
rect 25354 32805 27385 32819
rect 4146 31285 4212 32805
tri 4212 32758 4259 32805 nw
tri 15500 32758 15547 32805 ne
rect 15547 32764 15594 32805
tri 15594 32764 15635 32805 sw
tri 15680 32764 15721 32805 ne
rect 15721 32796 15774 32805
tri 15774 32796 15783 32805 sw
tri 15860 32796 15869 32805 ne
rect 15869 32796 15954 32805
rect 15721 32788 15783 32796
tri 15783 32788 15791 32796 sw
tri 15869 32788 15877 32796 ne
rect 15877 32788 15954 32796
tri 15954 32788 15971 32805 sw
tri 16040 32788 16057 32805 ne
rect 16057 32788 16134 32805
tri 16134 32788 16151 32805 sw
rect 15721 32764 15791 32788
rect 15547 32758 15635 32764
tri 15547 32749 15556 32758 ne
rect 15556 32756 15635 32758
tri 15635 32756 15643 32764 sw
tri 15721 32756 15729 32764 ne
rect 15729 32756 15791 32764
tri 15791 32756 15823 32788 sw
tri 15877 32756 15909 32788 ne
rect 15909 32756 15971 32788
tri 15971 32756 16003 32788 sw
tri 16057 32756 16089 32788 ne
rect 16089 32756 16151 32788
tri 16151 32756 16183 32788 sw
rect 15556 32749 15643 32756
tri 15643 32749 15650 32756 sw
tri 15729 32749 15736 32756 ne
rect 15736 32749 15823 32756
tri 15823 32749 15830 32756 sw
tri 15909 32749 15916 32756 ne
rect 15916 32749 16003 32756
tri 16003 32749 16010 32756 sw
tri 16089 32749 16096 32756 ne
rect 16096 32749 16183 32756
tri 16183 32749 16190 32756 sw
rect 25354 32749 25364 32805
rect 25420 32749 25506 32805
rect 25562 32749 25648 32805
rect 25704 32800 27385 32805
tri 27385 32800 27404 32819 sw
tri 27632 32800 27651 32819 ne
rect 25704 32749 27404 32800
tri 15556 32724 15581 32749 ne
rect 15581 32724 15650 32749
tri 15650 32724 15675 32749 sw
tri 15736 32724 15761 32749 ne
rect 15761 32724 15830 32749
tri 15830 32724 15855 32749 sw
tri 15916 32724 15941 32749 ne
rect 15941 32734 16010 32749
tri 16010 32734 16025 32749 sw
tri 16096 32734 16111 32749 ne
rect 16111 32734 16190 32749
rect 15941 32726 16025 32734
tri 16025 32726 16033 32734 sw
tri 16111 32726 16119 32734 ne
rect 16119 32726 16190 32734
tri 16190 32726 16213 32749 sw
rect 15941 32724 16033 32726
tri 16033 32724 16035 32726 sw
tri 16119 32724 16121 32726 ne
rect 16121 32724 16213 32726
tri 16213 32724 16215 32726 sw
tri 15581 32686 15619 32724 ne
rect 15619 32686 15675 32724
tri 15675 32686 15713 32724 sw
tri 15761 32686 15799 32724 ne
rect 15799 32702 15855 32724
tri 15855 32702 15877 32724 sw
tri 15941 32702 15963 32724 ne
rect 15963 32702 16035 32724
rect 15799 32694 15877 32702
tri 15877 32694 15885 32702 sw
tri 15963 32694 15971 32702 ne
rect 15971 32694 16035 32702
tri 16035 32694 16065 32724 sw
tri 16121 32694 16151 32724 ne
rect 16151 32694 16215 32724
tri 16215 32694 16245 32724 sw
rect 15799 32686 15885 32694
tri 15885 32686 15893 32694 sw
tri 15971 32686 15979 32694 ne
rect 15979 32686 16065 32694
tri 16065 32686 16073 32694 sw
tri 16151 32686 16159 32694 ne
rect 16159 32686 16245 32694
tri 16245 32686 16253 32694 sw
rect 25354 32686 27404 32749
tri 15619 32630 15675 32686 ne
rect 15675 32670 15713 32686
tri 15713 32670 15729 32686 sw
tri 15799 32670 15815 32686 ne
rect 15815 32670 15893 32686
rect 15675 32662 15729 32670
tri 15729 32662 15737 32670 sw
tri 15815 32662 15823 32670 ne
rect 15823 32662 15893 32670
tri 15893 32662 15917 32686 sw
tri 15979 32662 16003 32686 ne
rect 16003 32662 16073 32686
tri 16073 32662 16097 32686 sw
tri 16159 32662 16183 32686 ne
rect 16183 32662 16253 32686
tri 16253 32662 16277 32686 sw
rect 15675 32630 15737 32662
tri 15737 32630 15769 32662 sw
tri 15823 32630 15855 32662 ne
rect 15855 32630 15917 32662
tri 15917 32630 15949 32662 sw
tri 16003 32630 16035 32662 ne
rect 16035 32640 16097 32662
tri 16097 32640 16119 32662 sw
tri 16183 32640 16205 32662 ne
rect 16205 32640 16277 32662
rect 16035 32632 16119 32640
tri 16119 32632 16127 32640 sw
tri 16205 32632 16213 32640 ne
rect 16213 32632 16277 32640
tri 16277 32632 16307 32662 sw
rect 16035 32630 16127 32632
tri 16127 32630 16129 32632 sw
tri 16213 32630 16215 32632 ne
rect 16215 32630 19423 32632
tri 15675 32620 15685 32630 ne
rect 15685 32620 15769 32630
tri 15769 32620 15779 32630 sw
tri 15855 32620 15865 32630 ne
rect 15865 32620 15949 32630
tri 15949 32620 15959 32630 sw
tri 16035 32620 16045 32630 ne
rect 16045 32620 16129 32630
tri 16129 32620 16139 32630 sw
tri 16215 32620 16225 32630 ne
rect 16225 32620 19423 32630
rect 25354 32630 25364 32686
rect 25420 32630 25506 32686
rect 25562 32630 25648 32686
rect 25704 32661 27404 32686
tri 27404 32661 27543 32800 sw
rect 25704 32630 27543 32661
tri 15685 32564 15741 32620 ne
rect 15741 32576 15779 32620
tri 15779 32576 15823 32620 sw
tri 15865 32576 15909 32620 ne
rect 15909 32608 15959 32620
tri 15959 32608 15971 32620 sw
tri 16045 32608 16057 32620 ne
rect 16057 32608 16139 32620
rect 15909 32600 15971 32608
tri 15971 32600 15979 32608 sw
tri 16057 32600 16065 32608 ne
rect 16065 32600 16139 32608
tri 16139 32600 16159 32620 sw
tri 16225 32600 16245 32620 ne
rect 16245 32600 19423 32620
rect 15909 32576 15979 32600
rect 15741 32568 15823 32576
tri 15823 32568 15831 32576 sw
tri 15909 32568 15917 32576 ne
rect 15917 32568 15979 32576
tri 15979 32568 16011 32600 sw
tri 16065 32568 16097 32600 ne
rect 16097 32568 16159 32600
tri 16159 32568 16191 32600 sw
tri 16245 32568 16277 32600 ne
rect 16277 32568 19423 32600
rect 15741 32564 15831 32568
tri 15831 32564 15835 32568 sw
tri 15917 32564 15921 32568 ne
rect 15921 32564 16011 32568
tri 16011 32564 16015 32568 sw
tri 16097 32564 16101 32568 ne
rect 16101 32566 16191 32568
tri 16191 32566 16193 32568 sw
tri 16277 32566 16279 32568 ne
rect 16279 32566 19423 32568
rect 19704 32621 23313 32629
tri 23313 32621 23321 32629 sw
rect 19704 32620 23321 32621
rect 16101 32564 16193 32566
tri 16193 32564 16195 32566 sw
rect 19704 32564 19713 32620
rect 19769 32564 19811 32620
rect 19867 32564 19910 32620
rect 19966 32564 20987 32620
rect 21043 32564 21106 32620
rect 21162 32564 21225 32620
rect 21281 32567 23321 32620
tri 23321 32567 23375 32621 sw
rect 25354 32567 27543 32630
rect 21281 32566 23375 32567
tri 23375 32566 23376 32567 sw
rect 21281 32564 23376 32566
tri 15741 32536 15769 32564 ne
rect 15769 32536 15835 32564
tri 15835 32536 15863 32564 sw
tri 15921 32536 15949 32564 ne
rect 15949 32536 16015 32564
tri 16015 32536 16043 32564 sw
tri 16101 32536 16129 32564 ne
rect 16129 32536 16195 32564
tri 16195 32536 16223 32564 sw
rect 19704 32536 23376 32564
tri 23376 32536 23406 32566 sw
tri 15769 32516 15789 32536 ne
rect 15789 32516 15863 32536
tri 15863 32516 15883 32536 sw
tri 15949 32516 15969 32536 ne
rect 15969 32516 16043 32536
tri 16043 32516 16063 32536 sw
tri 16129 32516 16149 32536 ne
rect 16149 32516 16223 32536
tri 16223 32516 16243 32536 sw
rect 19704 32516 23406 32536
tri 15789 32501 15804 32516 ne
rect 15804 32506 15883 32516
tri 15883 32506 15893 32516 sw
tri 15969 32506 15979 32516 ne
rect 15979 32514 16063 32516
tri 16063 32514 16065 32516 sw
tri 16149 32514 16151 32516 ne
rect 16151 32514 16243 32516
rect 15979 32506 16065 32514
tri 16065 32506 16073 32514 sw
tri 16151 32506 16159 32514 ne
rect 16159 32506 16243 32514
tri 16243 32506 16253 32516 sw
rect 15804 32501 15893 32506
tri 15893 32501 15898 32506 sw
tri 15979 32501 15984 32506 ne
rect 15984 32501 16073 32506
tri 16073 32501 16078 32506 sw
tri 16159 32501 16164 32506 ne
rect 16164 32501 19500 32506
tri 15804 32445 15860 32501 ne
rect 15860 32482 15898 32501
tri 15898 32482 15917 32501 sw
tri 15984 32482 16003 32501 ne
rect 16003 32482 16078 32501
rect 15860 32474 15917 32482
tri 15917 32474 15925 32482 sw
tri 16003 32474 16011 32482 ne
rect 16011 32474 16078 32482
tri 16078 32474 16105 32501 sw
tri 16164 32474 16191 32501 ne
rect 16191 32474 19359 32501
rect 15860 32445 15925 32474
tri 15925 32445 15954 32474 sw
tri 16011 32445 16040 32474 ne
rect 16040 32445 16105 32474
tri 16105 32445 16134 32474 sw
tri 16191 32445 16220 32474 ne
rect 16220 32445 19359 32474
rect 19415 32445 19439 32501
rect 19495 32445 19500 32501
rect 19704 32460 19713 32516
rect 19769 32460 19811 32516
rect 19867 32460 19910 32516
rect 19966 32460 20987 32516
rect 21043 32460 21106 32516
rect 21162 32460 21225 32516
rect 21281 32511 23406 32516
tri 23406 32511 23431 32536 sw
rect 25354 32511 25364 32567
rect 25420 32511 25506 32567
rect 25562 32511 25648 32567
rect 25704 32511 27543 32567
rect 21281 32506 23431 32511
tri 23431 32506 23436 32511 sw
rect 21281 32460 23436 32506
rect 19704 32449 23436 32460
tri 23156 32447 23158 32449 ne
rect 23158 32447 23436 32449
tri 23436 32447 23495 32506 sw
rect 25354 32447 27543 32511
tri 15860 32442 15863 32445 ne
rect 15863 32442 15954 32445
tri 15954 32442 15957 32445 sw
tri 16040 32442 16043 32445 ne
rect 16043 32442 16134 32445
tri 16134 32442 16137 32445 sw
tri 16220 32442 16223 32445 ne
rect 16223 32442 19500 32445
tri 15863 32391 15914 32442 ne
rect 15914 32440 15957 32442
tri 15957 32440 15959 32442 sw
tri 16043 32440 16045 32442 ne
rect 16045 32440 16137 32442
tri 16137 32440 16139 32442 sw
tri 16223 32440 16225 32442 ne
rect 16225 32440 19500 32442
tri 23158 32440 23165 32447 ne
rect 23165 32440 23495 32447
tri 23495 32440 23502 32447 sw
rect 15914 32391 15959 32440
tri 15959 32391 16008 32440 sw
tri 16045 32391 16094 32440 ne
rect 16094 32391 16139 32440
tri 16139 32391 16188 32440 sw
tri 23165 32391 23214 32440 ne
rect 23214 32391 23502 32440
tri 23502 32391 23551 32440 sw
rect 25354 32391 25364 32447
rect 25420 32391 25506 32447
rect 25562 32391 25648 32447
rect 25704 32391 27543 32447
tri 15914 32348 15957 32391 ne
rect 15957 32388 16008 32391
tri 16008 32388 16011 32391 sw
tri 16094 32388 16097 32391 ne
rect 16097 32388 16188 32391
rect 15957 32380 16011 32388
tri 16011 32380 16019 32388 sw
tri 16097 32380 16105 32388 ne
rect 16105 32380 16188 32388
tri 16188 32380 16199 32391 sw
tri 23214 32380 23225 32391 ne
rect 23225 32380 23551 32391
tri 23551 32380 23562 32391 sw
rect 15957 32348 16019 32380
tri 16019 32348 16051 32380 sw
tri 16105 32348 16137 32380 ne
rect 16137 32348 18524 32380
tri 15957 32327 15978 32348 ne
rect 15978 32327 16051 32348
tri 16051 32327 16072 32348 sw
tri 16137 32327 16158 32348 ne
rect 16158 32327 18524 32348
tri 23225 32327 23278 32380 ne
rect 23278 32327 23562 32380
tri 23562 32327 23615 32380 sw
rect 25354 32327 27543 32391
tri 15978 32271 16034 32327 ne
rect 16034 32314 16072 32327
tri 16072 32314 16085 32327 sw
tri 16158 32314 16171 32327 ne
rect 16171 32314 18524 32327
tri 23278 32314 23291 32327 ne
rect 23291 32314 23615 32327
tri 23615 32314 23628 32327 sw
rect 16034 32271 16085 32314
tri 16085 32271 16128 32314 sw
tri 23291 32284 23321 32314 ne
rect 23321 32284 23628 32314
tri 23628 32284 23658 32314 sw
tri 23321 32271 23334 32284 ne
rect 23334 32271 23658 32284
tri 23658 32271 23671 32284 sw
rect 25354 32271 25364 32327
rect 25420 32271 25506 32327
rect 25562 32271 25648 32327
rect 25704 32271 27543 32327
tri 16034 32254 16051 32271 ne
rect 16051 32262 16128 32271
tri 16128 32262 16137 32271 sw
tri 23334 32262 23343 32271 ne
rect 23343 32262 23671 32271
tri 23671 32262 23680 32271 sw
rect 25354 32262 27543 32271
rect 16051 32254 16137 32262
tri 16137 32254 16145 32262 sw
tri 23343 32254 23351 32262 ne
rect 23351 32254 23680 32262
tri 23680 32254 23688 32262 sw
tri 26703 32254 26711 32262 ne
rect 26711 32254 27543 32262
tri 16051 32249 16056 32254 ne
rect 16056 32249 18334 32254
tri 16056 32193 16112 32249 ne
rect 16112 32193 18334 32249
tri 16112 32188 16117 32193 ne
rect 16117 32188 18334 32193
rect 18515 32249 18661 32254
rect 18515 32193 18520 32249
rect 18576 32193 18600 32249
rect 18656 32193 18661 32249
rect 18515 32188 18661 32193
tri 23351 32188 23417 32254 ne
rect 23417 32188 23688 32254
tri 23688 32188 23754 32254 sw
tri 26711 32188 26777 32254 ne
rect 26777 32188 27543 32254
tri 23417 32128 23477 32188 ne
rect 23477 32128 23754 32188
tri 23754 32128 23814 32188 sw
tri 26777 32128 26837 32188 ne
rect 26837 32128 27543 32188
rect 13446 32123 23004 32128
rect 13446 32067 13451 32123
rect 13507 32067 13531 32123
rect 13587 32068 23004 32123
tri 23004 32068 23064 32128 sw
tri 23477 32068 23537 32128 ne
rect 23537 32068 23814 32128
tri 23814 32068 23874 32128 sw
tri 26837 32068 26897 32128 ne
rect 26897 32068 27543 32128
rect 13587 32067 23064 32068
rect 13446 32062 23064 32067
tri 23064 32062 23070 32068 sw
tri 23537 32062 23543 32068 ne
rect 23543 32062 23874 32068
tri 23874 32062 23880 32068 sw
tri 26897 32062 26903 32068 ne
rect 26903 32062 27543 32068
tri 22976 32058 22980 32062 ne
rect 22980 32058 23070 32062
tri 23070 32058 23074 32062 sw
tri 23543 32058 23547 32062 ne
rect 23547 32058 23880 32062
tri 23880 32058 23884 32062 sw
tri 26903 32058 26907 32062 ne
rect 26907 32058 27543 32062
tri 22980 32034 23004 32058 ne
rect 23004 32034 23074 32058
tri 23004 32012 23026 32034 ne
rect 23026 32012 23074 32034
tri 23074 32012 23120 32058 sw
tri 23547 32012 23593 32058 ne
rect 23593 32012 23884 32058
tri 23884 32012 23930 32058 sw
tri 26907 32012 26953 32058 ne
rect 26953 32012 27543 32058
tri 23026 32007 23031 32012 ne
rect 23031 32007 23120 32012
tri 23120 32007 23125 32012 sw
tri 23593 32007 23598 32012 ne
rect 23598 32007 23930 32012
tri 23930 32007 23935 32012 sw
rect 25864 32007 25930 32012
tri 23031 31973 23065 32007 ne
rect 23065 31973 23125 32007
rect 19336 31964 21295 31973
tri 23065 31964 23074 31973 ne
rect 23074 31964 23125 31973
tri 23125 31964 23168 32007 sw
tri 23598 31964 23641 32007 ne
rect 23641 31964 23935 32007
tri 23935 31964 23978 32007 sw
rect 19336 31947 20978 31964
rect 19336 31891 19360 31947
rect 19416 31891 19468 31947
rect 19524 31891 19575 31947
rect 19631 31891 19682 31947
rect 19738 31891 19789 31947
rect 19845 31891 19896 31947
rect 19952 31908 20978 31947
rect 21034 31908 21106 31964
rect 21162 31908 21234 31964
rect 21290 31908 21295 31964
tri 23074 31951 23087 31964 ne
rect 23087 31951 23168 31964
tri 23168 31951 23181 31964 sw
tri 23641 31951 23654 31964 ne
rect 23654 31951 23978 31964
tri 23978 31951 23991 31964 sw
rect 25864 31951 25869 32007
rect 25925 31951 25930 32007
tri 23087 31927 23111 31951 ne
rect 23111 31927 23181 31951
tri 23181 31927 23205 31951 sw
tri 23654 31947 23658 31951 ne
rect 23658 31947 23991 31951
tri 23991 31947 23995 31951 sw
tri 23658 31927 23678 31947 ne
rect 23678 31927 23995 31947
tri 23995 31927 24015 31947 sw
rect 25864 31927 25930 31951
rect 19952 31891 21295 31908
rect 19336 31854 21295 31891
tri 23111 31871 23167 31927 ne
rect 23167 31871 23205 31927
tri 23205 31871 23261 31927 sw
tri 23678 31871 23734 31927 ne
rect 23734 31871 24015 31927
tri 24015 31871 24071 31927 sw
rect 25864 31871 25869 31927
rect 25925 31871 25930 31927
tri 23167 31870 23168 31871 ne
rect 23168 31870 23261 31871
tri 23261 31870 23262 31871 sw
tri 23734 31870 23735 31871 ne
rect 23735 31870 24071 31871
tri 24071 31870 24072 31871 sw
rect 19336 31798 20978 31854
rect 21034 31798 21106 31854
rect 21162 31798 21234 31854
rect 21290 31798 21295 31854
rect 19336 31789 21295 31798
rect 19336 31733 19360 31789
rect 19416 31733 19468 31789
rect 19524 31733 19575 31789
rect 19631 31733 19682 31789
rect 19738 31733 19789 31789
rect 19845 31733 19896 31789
rect 19952 31743 21295 31789
tri 23168 31776 23262 31870 ne
tri 23262 31776 23356 31870 sw
tri 23735 31776 23829 31870 ne
rect 23829 31776 24072 31870
tri 24072 31776 24166 31870 sw
rect 19952 31733 20978 31743
rect 19336 31687 20978 31733
rect 21034 31687 21106 31743
rect 21162 31687 21234 31743
rect 21290 31687 21295 31743
rect 19336 31632 21295 31687
tri 23262 31682 23356 31776 ne
tri 23356 31682 23450 31776 sw
tri 23829 31682 23923 31776 ne
rect 23923 31682 24166 31776
tri 24166 31682 24260 31776 sw
rect 4146 31229 4151 31285
rect 4207 31229 4212 31285
rect 4146 31205 4212 31229
rect 4146 31149 4151 31205
rect 4207 31149 4212 31205
rect 4146 31144 4212 31149
rect 14879 31573 15445 31578
rect 14879 31517 14888 31573
rect 14944 31517 14970 31573
rect 15026 31517 15052 31573
rect 15108 31517 15134 31573
rect 15190 31517 15216 31573
rect 15272 31517 15298 31573
rect 15354 31517 15380 31573
rect 15436 31517 15445 31573
rect 19336 31576 20978 31632
rect 21034 31576 21106 31632
rect 21162 31576 21234 31632
rect 21290 31576 21295 31632
tri 23356 31588 23450 31682 ne
tri 23450 31588 23544 31682 sw
tri 23923 31610 23995 31682 ne
rect 23995 31610 24260 31682
tri 24260 31610 24332 31682 sw
tri 23995 31588 24017 31610 ne
rect 24017 31588 24332 31610
rect 19336 31567 21295 31576
tri 23450 31567 23471 31588 ne
rect 23471 31567 23544 31588
rect 14879 31492 15445 31517
tri 23471 31494 23544 31567 ne
tri 23544 31494 23638 31588 sw
tri 24017 31494 24111 31588 ne
rect 24111 31494 24332 31588
rect 14879 31436 14888 31492
rect 14944 31436 14970 31492
rect 15026 31436 15052 31492
rect 15108 31436 15134 31492
rect 15190 31436 15216 31492
rect 15272 31436 15298 31492
rect 15354 31436 15380 31492
rect 15436 31436 15445 31492
tri 23544 31454 23584 31494 ne
rect 23584 31454 23638 31494
tri 23638 31454 23678 31494 sw
tri 24111 31454 24151 31494 ne
rect 24151 31454 24332 31494
rect 14879 31411 15445 31436
rect 14879 31355 14888 31411
rect 14944 31355 14970 31411
rect 15026 31355 15052 31411
rect 15108 31355 15134 31411
rect 15190 31355 15216 31411
rect 15272 31355 15298 31411
rect 15354 31355 15380 31411
rect 15436 31355 15445 31411
tri 23584 31400 23638 31454 ne
rect 23638 31400 23678 31454
tri 23678 31400 23732 31454 sw
tri 24151 31453 24152 31454 ne
tri 23638 31398 23640 31400 ne
rect 23640 31398 23732 31400
tri 23732 31398 23734 31400 sw
tri 23640 31374 23664 31398 ne
rect 23664 31374 23734 31398
tri 23734 31374 23758 31398 sw
tri 23664 31362 23676 31374 ne
rect 23676 31362 23758 31374
tri 23758 31362 23770 31374 sw
rect 14879 31330 15445 31355
rect 14879 31274 14888 31330
rect 14944 31274 14970 31330
rect 15026 31274 15052 31330
rect 15108 31274 15134 31330
rect 15190 31274 15216 31330
rect 15272 31274 15298 31330
rect 15354 31274 15380 31330
rect 15436 31274 15445 31330
tri 23676 31306 23732 31362 ne
rect 23732 31306 23770 31362
tri 23770 31306 23826 31362 sw
tri 23732 31282 23756 31306 ne
rect 23756 31282 23826 31306
tri 23756 31278 23760 31282 ne
rect 14879 31249 15445 31274
rect 14879 31193 14888 31249
rect 14944 31193 14970 31249
rect 15026 31193 15052 31249
rect 15108 31193 15134 31249
rect 15190 31193 15216 31249
rect 15272 31193 15298 31249
rect 15354 31193 15380 31249
rect 15436 31193 15445 31249
rect 14879 31168 15445 31193
rect 14879 31112 14888 31168
rect 14944 31112 14970 31168
rect 15026 31112 15052 31168
rect 15108 31112 15134 31168
rect 15190 31112 15216 31168
rect 15272 31112 15298 31168
rect 15354 31112 15380 31168
rect 15436 31112 15445 31168
rect 14879 31087 15445 31112
rect 14879 31031 14888 31087
rect 14944 31031 14970 31087
rect 15026 31031 15052 31087
rect 15108 31031 15134 31087
rect 15190 31031 15216 31087
rect 15272 31031 15298 31087
rect 15354 31031 15380 31087
rect 15436 31031 15445 31087
rect 14879 31006 15445 31031
rect 14879 30950 14888 31006
rect 14944 30950 14970 31006
rect 15026 30950 15052 31006
rect 15108 30950 15134 31006
rect 15190 30950 15216 31006
rect 15272 30950 15298 31006
rect 15354 30950 15380 31006
rect 15436 30950 15445 31006
rect 14879 30924 15445 30950
rect 14879 30868 14888 30924
rect 14944 30868 14970 30924
rect 15026 30868 15052 30924
rect 15108 30868 15134 30924
rect 15190 30868 15216 30924
rect 15272 30868 15298 30924
rect 15354 30868 15380 30924
rect 15436 30868 15445 30924
rect 14879 30842 15445 30868
rect 14879 30786 14888 30842
rect 14944 30786 14970 30842
rect 15026 30786 15052 30842
rect 15108 30786 15134 30842
rect 15190 30786 15216 30842
rect 15272 30786 15298 30842
rect 15354 30786 15380 30842
rect 15436 30786 15445 30842
rect 14879 30760 15445 30786
rect 14879 30704 14888 30760
rect 14944 30704 14970 30760
rect 15026 30704 15052 30760
rect 15108 30704 15134 30760
rect 15190 30704 15216 30760
rect 15272 30704 15298 30760
rect 15354 30704 15380 30760
rect 15436 30704 15445 30760
rect 14879 30678 15445 30704
rect 14879 30622 14888 30678
rect 14944 30622 14970 30678
rect 15026 30622 15052 30678
rect 15108 30622 15134 30678
rect 15190 30622 15216 30678
rect 15272 30622 15298 30678
rect 15354 30622 15380 30678
rect 15436 30622 15445 30678
rect 14879 30596 15445 30622
rect 14879 30540 14888 30596
rect 14944 30540 14970 30596
rect 15026 30540 15052 30596
rect 15108 30540 15134 30596
rect 15190 30540 15216 30596
rect 15272 30540 15298 30596
rect 15354 30540 15380 30596
rect 15436 30540 15445 30596
rect 14879 30514 15445 30540
rect 14879 30458 14888 30514
rect 14944 30458 14970 30514
rect 15026 30458 15052 30514
rect 15108 30458 15134 30514
rect 15190 30458 15216 30514
rect 15272 30458 15298 30514
rect 15354 30458 15380 30514
rect 15436 30458 15445 30514
rect 14879 30432 15445 30458
rect 14879 30376 14888 30432
rect 14944 30376 14970 30432
rect 15026 30376 15052 30432
rect 15108 30376 15134 30432
rect 15190 30376 15216 30432
rect 15272 30376 15298 30432
rect 15354 30376 15380 30432
rect 15436 30376 15445 30432
rect 14879 30350 15445 30376
rect 14879 30294 14888 30350
rect 14944 30294 14970 30350
rect 15026 30294 15052 30350
rect 15108 30294 15134 30350
rect 15190 30294 15216 30350
rect 15272 30294 15298 30350
rect 15354 30294 15380 30350
rect 15436 30294 15445 30350
rect 14879 30268 15445 30294
rect 14879 30212 14888 30268
rect 14944 30212 14970 30268
rect 15026 30212 15052 30268
rect 15108 30212 15134 30268
rect 15190 30212 15216 30268
rect 15272 30212 15298 30268
rect 15354 30212 15380 30268
rect 15436 30212 15445 30268
rect 14879 30207 15445 30212
rect 23760 28860 23826 31282
rect 24152 30695 24332 31454
rect 24397 31051 24463 31056
rect 24397 30995 24402 31051
rect 24458 30995 24463 31051
rect 24397 30971 24463 30995
rect 24397 30915 24402 30971
rect 24458 30915 24463 30971
rect 24397 30910 24463 30915
rect 24152 30639 24164 30695
rect 24220 30639 24268 30695
rect 24324 30639 24332 30695
rect 24152 30600 24332 30639
rect 24152 30544 24164 30600
rect 24220 30544 24268 30600
rect 24324 30544 24332 30600
rect 24152 30505 24332 30544
tri 25771 30529 25864 30622 se
rect 25864 30595 25930 31871
tri 25864 30529 25930 30595 nw
rect 25996 32007 26062 32012
rect 25996 31951 26001 32007
rect 26057 31951 26062 32007
rect 25996 31927 26062 31951
rect 25996 31871 26001 31927
rect 26057 31871 26062 31927
rect 24152 30449 24164 30505
rect 24220 30449 24268 30505
rect 24324 30449 24332 30505
rect 24152 30410 24332 30449
tri 25678 30436 25771 30529 se
tri 25771 30436 25864 30529 nw
tri 25906 30436 25996 30526 se
rect 25996 30498 26062 31871
rect 24152 30354 24164 30410
rect 24220 30354 24268 30410
rect 24324 30354 24332 30410
tri 24098 29586 24152 29640 se
rect 24152 29586 24332 30354
tri 25585 30343 25678 30436 se
tri 25678 30343 25771 30436 nw
tri 25902 30432 25906 30436 se
rect 25906 30432 25996 30436
tri 25996 30432 26062 30498 nw
rect 26137 32007 26203 32012
rect 26137 31951 26142 32007
rect 26198 31951 26203 32007
tri 26953 31964 27001 32012 ne
rect 27001 31964 27543 32012
rect 26137 31927 26203 31951
rect 26137 31871 26142 31927
rect 26198 31871 26203 31927
tri 27001 31922 27043 31964 ne
tri 25813 30343 25902 30432 se
tri 25527 30285 25585 30343 se
rect 25585 30285 25620 30343
tri 25620 30285 25678 30343 nw
tri 25808 30338 25813 30343 se
rect 25813 30338 25902 30343
tri 25902 30338 25996 30432 nw
tri 25755 30285 25808 30338 se
rect 25808 30285 25849 30338
tri 25849 30285 25902 30338 nw
tri 25517 30275 25527 30285 se
rect 25527 30275 25610 30285
tri 25610 30275 25620 30285 nw
tri 25750 30280 25755 30285 se
rect 25755 30280 25826 30285
rect 25727 30275 25826 30280
tri 25492 30250 25517 30275 se
rect 25517 30250 25585 30275
tri 25585 30250 25610 30275 nw
tri 25461 30219 25492 30250 se
rect 25492 30219 25554 30250
tri 25554 30219 25585 30250 nw
rect 25727 30219 25732 30275
rect 25788 30262 25826 30275
tri 25826 30262 25849 30285 nw
tri 26114 30262 26137 30285 se
rect 26137 30262 26203 31871
rect 26539 31454 26605 31459
rect 26539 31398 26544 31454
rect 26600 31398 26605 31454
rect 26539 31374 26605 31398
rect 25788 30250 25814 30262
tri 25814 30250 25826 30262 nw
tri 26102 30250 26114 30262 se
rect 26114 30257 26203 30262
rect 26114 30250 26137 30257
rect 25788 30219 25793 30250
tri 25793 30229 25814 30250 nw
tri 26081 30229 26102 30250 se
rect 26102 30229 26137 30250
tri 25437 30195 25461 30219 se
rect 25461 30195 25530 30219
tri 25530 30195 25554 30219 nw
rect 25727 30195 25793 30219
tri 25433 30191 25437 30195 se
rect 25437 30191 25526 30195
tri 25526 30191 25530 30195 nw
tri 25399 30157 25433 30191 se
rect 25433 30157 25492 30191
tri 25492 30157 25526 30191 nw
tri 25381 30139 25399 30157 se
rect 25399 30139 25474 30157
tri 25474 30139 25492 30157 nw
rect 25727 30139 25732 30195
rect 25788 30139 25793 30195
tri 26043 30191 26081 30229 se
rect 26081 30191 26137 30229
tri 26137 30191 26203 30257 nw
rect 26287 31362 26353 31367
rect 26287 31306 26292 31362
rect 26348 31306 26353 31362
rect 26287 31282 26353 31306
rect 26287 31226 26292 31282
rect 26348 31226 26353 31282
tri 25339 30097 25381 30139 se
rect 25381 30097 25432 30139
tri 25432 30097 25474 30139 nw
rect 25727 30134 25793 30139
tri 25986 30134 26043 30191 se
tri 25949 30097 25986 30134 se
rect 25986 30097 26043 30134
tri 26043 30097 26137 30191 nw
tri 25306 30064 25339 30097 se
rect 25339 30064 25399 30097
tri 25399 30064 25432 30097 nw
tri 25916 30064 25949 30097 se
tri 25280 30038 25306 30064 se
rect 25306 30038 25373 30064
tri 25373 30038 25399 30064 nw
tri 25890 30038 25916 30064 se
rect 25916 30038 25949 30064
rect 23760 28804 23765 28860
rect 23821 28804 23826 28860
rect 23760 28780 23826 28804
rect 23760 28724 23765 28780
rect 23821 28724 23826 28780
rect 23760 28715 23826 28724
tri 23906 29394 24098 29586 se
rect 24098 29394 24332 29586
rect 23906 29377 24332 29394
tri 2171 27614 2226 27669 ne
rect 2226 27614 2231 27669
tri 2231 27614 2312 27695 sw
tri 2226 27609 2231 27614 ne
rect 2231 27609 2312 27614
tri 2231 27589 2251 27609 ne
rect 2251 27471 2312 27609
rect 20566 27158 20743 27455
rect 2646 18462 2686 18491
rect 23906 17846 24187 29377
tri 24187 29232 24332 29377 nw
rect 23906 17790 23917 17846
rect 23973 17790 24019 17846
rect 24075 17790 24121 17846
rect 24177 17790 24187 17846
rect 23906 17753 24187 17790
rect 23906 17697 23917 17753
rect 23973 17697 24019 17753
rect 24075 17697 24121 17753
rect 24177 17697 24187 17753
rect 23906 17660 24187 17697
rect 23906 17604 23917 17660
rect 23973 17604 24019 17660
rect 24075 17604 24121 17660
rect 24177 17604 24187 17660
rect 23906 17567 24187 17604
rect 23906 17511 23917 17567
rect 23973 17511 24019 17567
rect 24075 17511 24121 17567
rect 24177 17511 24187 17567
rect 23906 17473 24187 17511
rect 23906 17417 23917 17473
rect 23973 17417 24019 17473
rect 24075 17417 24121 17473
rect 24177 17417 24187 17473
rect 23906 17379 24187 17417
rect 23906 17323 23917 17379
rect 23973 17323 24019 17379
rect 24075 17323 24121 17379
rect 24177 17323 24187 17379
rect 23906 17314 24187 17323
rect 24256 28860 24322 28881
rect 24256 28804 24261 28860
rect 24317 28804 24322 28860
rect 24256 28780 24322 28804
rect 24256 28724 24261 28780
rect 24317 28724 24322 28780
rect 21051 8342 21940 8347
rect 21051 8286 21060 8342
rect 21116 8286 21142 8342
rect 21198 8286 21224 8342
rect 21280 8286 21306 8342
rect 21362 8286 21388 8342
rect 21444 8286 21470 8342
rect 21526 8286 21551 8342
rect 21607 8286 21632 8342
rect 21688 8286 21713 8342
rect 21769 8286 21794 8342
rect 21850 8286 21875 8342
rect 21931 8286 21940 8342
rect 21051 8262 21940 8286
rect 21051 8206 21060 8262
rect 21116 8206 21142 8262
rect 21198 8206 21224 8262
rect 21280 8206 21306 8262
rect 21362 8206 21388 8262
rect 21444 8206 21470 8262
rect 21526 8206 21551 8262
rect 21607 8206 21632 8262
rect 21688 8206 21713 8262
rect 21769 8206 21794 8262
rect 21850 8206 21875 8262
rect 21931 8206 21940 8262
rect 21051 8182 21940 8206
rect 21051 8126 21060 8182
rect 21116 8126 21142 8182
rect 21198 8126 21224 8182
rect 21280 8126 21306 8182
rect 21362 8126 21388 8182
rect 21444 8126 21470 8182
rect 21526 8126 21551 8182
rect 21607 8126 21632 8182
rect 21688 8126 21713 8182
rect 21769 8126 21794 8182
rect 21850 8126 21875 8182
rect 21931 8126 21940 8182
rect 21051 8121 21940 8126
tri 24222 1156 24256 1190 se
rect 24256 1156 24322 28724
tri 24209 1143 24222 1156 se
rect 24222 1143 24322 1156
rect 24134 1138 24322 1143
rect 24134 1082 24139 1138
rect 24195 1082 24322 1138
rect 24134 1058 24322 1082
rect 24134 1002 24139 1058
rect 24195 1002 24322 1058
rect 24134 997 24322 1002
rect 24397 329 24463 29767
rect 24523 23560 24589 23565
rect 24523 23504 24528 23560
rect 24584 23504 24589 23560
rect 24523 23462 24589 23504
rect 24523 23406 24528 23462
rect 24584 23406 24589 23462
rect 24523 23401 24589 23406
tri 25241 20066 25280 20105 se
rect 25280 20066 25345 30038
tri 25345 30010 25373 30038 nw
tri 25862 30010 25890 30038 se
rect 25890 30010 25949 30038
tri 25855 30003 25862 30010 se
rect 25862 30003 25949 30010
tri 25949 30003 26043 30097 nw
tri 25761 29909 25855 30003 se
tri 25855 29909 25949 30003 nw
tri 25667 29815 25761 29909 se
tri 25761 29815 25855 29909 nw
tri 25657 29805 25667 29815 se
rect 25667 29805 25751 29815
tri 25751 29805 25761 29815 nw
rect 25027 20000 25345 20066
rect 25405 29722 25471 29734
rect 25405 29666 25410 29722
rect 25466 29666 25471 29722
rect 25405 29642 25471 29666
rect 25405 29586 25410 29642
rect 25466 29586 25471 29642
rect 24542 17846 24947 17855
rect 24542 17790 24552 17846
rect 24608 17790 24634 17846
rect 24690 17790 24716 17846
rect 24772 17790 24798 17846
rect 24854 17790 24880 17846
rect 24936 17790 24947 17846
rect 24542 17753 24947 17790
rect 24542 17697 24552 17753
rect 24608 17697 24634 17753
rect 24690 17697 24716 17753
rect 24772 17697 24798 17753
rect 24854 17697 24880 17753
rect 24936 17697 24947 17753
rect 24542 17660 24947 17697
rect 24542 17604 24552 17660
rect 24608 17604 24634 17660
rect 24690 17604 24716 17660
rect 24772 17604 24798 17660
rect 24854 17604 24880 17660
rect 24936 17604 24947 17660
rect 24542 17567 24947 17604
rect 24542 17511 24552 17567
rect 24608 17511 24634 17567
rect 24690 17511 24716 17567
rect 24772 17511 24798 17567
rect 24854 17511 24880 17567
rect 24936 17511 24947 17567
rect 24542 17473 24947 17511
rect 24542 17417 24552 17473
rect 24608 17417 24634 17473
rect 24690 17417 24716 17473
rect 24772 17417 24798 17473
rect 24854 17417 24880 17473
rect 24936 17417 24947 17473
rect 24542 17379 24947 17417
rect 24542 17323 24552 17379
rect 24608 17323 24634 17379
rect 24690 17323 24716 17379
rect 24772 17323 24798 17379
rect 24854 17323 24880 17379
rect 24936 17323 24947 17379
rect 24542 8391 24947 17323
rect 24542 8335 24551 8391
rect 24607 8335 24634 8391
rect 24690 8335 24717 8391
rect 24773 8335 24800 8391
rect 24856 8335 24882 8391
rect 24938 8335 24947 8391
rect 24542 8305 24947 8335
rect 24542 8249 24551 8305
rect 24607 8249 24634 8305
rect 24690 8249 24717 8305
rect 24773 8249 24800 8305
rect 24856 8249 24882 8305
rect 24938 8249 24947 8305
rect 24542 8219 24947 8249
rect 24542 8163 24551 8219
rect 24607 8163 24634 8219
rect 24690 8163 24717 8219
rect 24773 8163 24800 8219
rect 24856 8163 24882 8219
rect 24938 8163 24947 8219
rect 24542 8133 24947 8163
rect 24542 8077 24551 8133
rect 24607 8077 24634 8133
rect 24690 8077 24717 8133
rect 24773 8077 24800 8133
rect 24856 8077 24882 8133
rect 24938 8077 24947 8133
rect 24542 8070 24947 8077
rect 24901 957 24967 962
rect 24711 913 24841 918
rect 24711 857 24716 913
rect 24772 857 24841 913
rect 24711 833 24841 857
rect 24711 777 24716 833
rect 24772 777 24841 833
rect 24711 772 24841 777
tri 24744 757 24759 772 ne
rect 24759 757 24841 772
tri 24759 741 24775 757 ne
rect 24775 49 24841 757
rect 24901 901 24906 957
rect 24962 901 24967 957
rect 24901 877 24967 901
rect 24901 821 24906 877
rect 24962 821 24967 877
rect 24901 49 24967 821
rect 25027 43 25093 20000
tri 25093 19961 25132 20000 nw
rect 25153 19923 25219 19932
rect 25153 19867 25158 19923
rect 25214 19867 25219 19923
rect 25153 19843 25219 19867
rect 25153 19787 25158 19843
rect 25214 19787 25219 19843
rect 25153 2793 25219 19787
rect 25405 19923 25471 29586
rect 25405 19867 25410 19923
rect 25466 19867 25471 19923
rect 25405 19843 25471 19867
rect 25405 19787 25410 19843
rect 25466 19787 25471 19843
rect 25405 19782 25471 19787
rect 25531 28485 25597 28504
rect 25531 28429 25536 28485
rect 25592 28429 25597 28485
rect 25531 28405 25597 28429
rect 25531 28349 25536 28405
rect 25592 28349 25597 28405
rect 25153 2737 25158 2793
rect 25214 2737 25219 2793
rect 25153 2713 25219 2737
rect 25153 2657 25158 2713
rect 25214 2657 25219 2713
rect 25153 1723 25219 2657
rect 25153 1667 25158 1723
rect 25214 1667 25219 1723
rect 25153 1643 25219 1667
rect 25153 1587 25158 1643
rect 25214 1587 25219 1643
rect 25153 1571 25219 1587
rect 25279 19711 25345 19720
rect 25279 19655 25284 19711
rect 25340 19655 25345 19711
rect 25279 19631 25345 19655
rect 25279 19575 25284 19631
rect 25340 19575 25345 19631
rect 25279 4480 25345 19575
rect 25279 4424 25284 4480
rect 25340 4424 25345 4480
rect 25279 4400 25345 4424
rect 25279 4344 25284 4400
rect 25340 4344 25345 4400
rect 25153 -171 25219 1506
rect 25279 26 25345 4344
rect 25405 18583 25471 18607
rect 25405 18527 25410 18583
rect 25466 18527 25471 18583
rect 25405 18503 25471 18527
rect 25405 18447 25410 18503
rect 25466 18447 25471 18503
rect 25405 757 25471 18447
rect 25531 1212 25597 28349
rect 25657 19711 25723 29805
tri 25723 29777 25751 29805 nw
rect 25657 19655 25662 19711
rect 25718 19655 25723 19711
rect 25657 19631 25723 19655
rect 25657 19575 25662 19631
rect 25718 19575 25723 19631
rect 25657 19570 25723 19575
rect 25783 20864 25849 20869
rect 25783 20808 25788 20864
rect 25844 20808 25849 20864
rect 25783 20784 25849 20808
rect 25783 20728 25788 20784
rect 25844 20728 25849 20784
rect 25783 20723 25849 20728
tri 25678 19425 25783 19530 se
rect 25783 19485 25843 20723
tri 25843 20717 25849 20723 nw
tri 25783 19425 25843 19485 nw
rect 25531 1156 25536 1212
rect 25592 1156 25597 1212
rect 25531 1132 25597 1156
rect 25531 1076 25536 1132
rect 25592 1076 25597 1132
rect 25531 1043 25597 1076
tri 25657 19404 25678 19425 se
rect 25678 19404 25762 19425
tri 25762 19404 25783 19425 nw
rect 25405 701 25410 757
rect 25466 701 25471 757
rect 25405 677 25471 701
rect 25405 621 25410 677
rect 25466 621 25471 677
rect 25405 615 25471 621
rect 25657 566 25723 19404
tri 25723 19365 25762 19404 nw
rect 25657 510 25662 566
rect 25718 510 25723 566
rect 25657 486 25723 510
rect 25657 430 25662 486
rect 25718 430 25723 486
rect 25657 425 25723 430
rect 26287 -19 26353 31226
rect 26539 31318 26544 31374
rect 26600 31318 26605 31374
rect 26413 30884 26479 30889
rect 26413 30828 26418 30884
rect 26474 30828 26479 30884
rect 26413 30804 26479 30828
rect 26413 30748 26418 30804
rect 26474 30748 26479 30804
rect 26413 -19 26479 30748
rect 26539 -19 26605 31318
rect 26791 31256 26857 31261
rect 26791 31200 26796 31256
rect 26852 31200 26857 31256
rect 26791 31176 26857 31200
rect 26791 31120 26796 31176
rect 26852 31120 26857 31176
rect 26665 30971 26731 30976
rect 26665 30915 26670 30971
rect 26726 30915 26731 30971
rect 26665 30891 26731 30915
rect 26665 30835 26670 30891
rect 26726 30835 26731 30891
rect 26665 -19 26731 30835
rect 26791 -19 26857 31120
rect 26917 31112 26983 31128
rect 26917 31056 26922 31112
rect 26978 31056 26983 31112
rect 26917 31032 26983 31056
rect 26917 30976 26922 31032
rect 26978 30976 26983 31032
rect 26917 -19 26983 30976
rect 27043 1416 27543 31964
rect 27043 1360 27052 1416
rect 27108 1360 27138 1416
rect 27194 1360 27223 1416
rect 27279 1360 27308 1416
rect 27364 1360 27393 1416
rect 27449 1360 27478 1416
rect 27534 1360 27543 1416
rect 27043 1280 27543 1360
rect 27043 1224 27052 1280
rect 27108 1224 27138 1280
rect 27194 1224 27223 1280
rect 27279 1224 27308 1280
rect 27364 1224 27393 1280
rect 27449 1224 27478 1280
rect 27534 1224 27543 1280
rect 27043 495 27543 1224
rect 27043 439 27052 495
rect 27108 439 27138 495
rect 27194 439 27223 495
rect 27279 439 27308 495
rect 27364 439 27393 495
rect 27449 439 27478 495
rect 27534 439 27543 495
rect 27043 359 27543 439
rect 27043 303 27052 359
rect 27108 303 27138 359
rect 27194 303 27223 359
rect 27279 303 27308 359
rect 27364 303 27393 359
rect 27449 303 27478 359
rect 27534 303 27543 359
rect 25153 -227 25158 -171
rect 25214 -227 25219 -171
rect 25153 -256 25219 -227
rect 25153 -312 25158 -256
rect 25214 -312 25219 -256
rect 25153 -317 25219 -312
rect 27043 -5849 27543 303
rect 27651 32068 27999 32819
rect 27651 32012 27660 32068
rect 27716 32012 27773 32068
rect 27829 32012 27885 32068
rect 27941 32012 27999 32068
rect 27651 31964 27999 32012
rect 27651 31908 27660 31964
rect 27716 31908 27773 31964
rect 27829 31908 27885 31964
rect 27941 31908 27999 31964
rect 27651 -5849 27999 31908
use sky130_fd_io__gpio_ovtv2_hvsbt_inv_x2_1  sky130_fd_io__gpio_ovtv2_hvsbt_inv_x2_1_0
timestamp 1694700623
transform 1 0 21872 0 1 29860
box -107 21 459 1369
use sky130_fd_io__gpio_ovtv2_hvsbt_inv_x2_1  sky130_fd_io__gpio_ovtv2_hvsbt_inv_x2_1_1
timestamp 1694700623
transform 1 0 20336 0 1 29860
box -107 21 459 1369
use sky130_fd_io__gpio_ovtv2_obpredrvr_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_obpredrvr_i2c_fix_leak_fix_0
timestamp 1694700623
transform 1 0 0 0 1 0
box 206 9097 28083 33907
use sky130_fd_io__gpio_ovtv2_octl_i2c_fix  sky130_fd_io__gpio_ovtv2_octl_i2c_fix_0
timestamp 1694700623
transform 1 0 20322 0 -1 33684
box -251 12 7522 3737
use sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix  sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix_0
timestamp 1694700623
transform -1 0 27820 0 -1 2305
box -349 -581 12658 2367
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1694700623
transform -1 0 21872 0 1 29860
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1694700623
transform -1 0 21192 0 1 29860
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_1
timestamp 1694700623
transform 1 0 21192 0 1 29860
box -107 21 487 1369
<< labels >>
flabel metal3 s 2646 18462 2686 18491 0 FreeSans 200 0 0 0 NGHS_H
port 21 nsew
flabel metal3 s 27651 32483 27999 32585 3 FreeSans 520 0 0 0 VCCD
port 1 nsew
flabel metal3 s 27043 31221 27543 31379 3 FreeSans 520 0 0 0 VSSD
port 2 nsew
flabel metal3 s 25027 43 25093 149 3 FreeSans 520 90 0 0 SLOW
port 3 nsew
flabel metal3 s 24901 49 24967 184 3 FreeSans 520 90 0 0 OE_N
port 4 nsew
flabel metal3 s 24775 49 24841 118 3 FreeSans 520 90 0 0 OUT
port 5 nsew
flabel metal3 s 26287 -17 26353 124 3 FreeSans 520 90 0 0 DM_H_N[2]
port 19 nsew
flabel metal3 s 2171 27784 2231 27925 3 FreeSans 520 90 0 0 SLEW_CTL_H[0]
port 6 nsew
flabel metal3 s 1429 27807 1489 27948 3 FreeSans 520 90 0 0 SLEW_CTL_H[1]
port 7 nsew
flabel metal3 s 1309 27806 1369 27947 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[0]
port 8 nsew
flabel metal3 s 1189 27807 1249 27948 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[1]
port 9 nsew
flabel metal3 s 25657 438 25723 579 3 FreeSans 520 90 0 0 DRVHI_H
port 10 nsew
flabel metal3 s 24397 329 24463 427 3 FreeSans 520 90 0 0 SLOW_H_N
port 11 nsew
flabel metal3 s 25279 26 25345 152 3 FreeSans 520 90 0 0 HLD_I_H_N
port 12 nsew
flabel metal3 s 25153 26 25219 152 3 FreeSans 520 90 0 0 OD_H
port 13 nsew
flabel metal3 s 26917 -17 26983 124 3 FreeSans 520 90 0 0 DM_H[0]
port 14 nsew
flabel metal3 s 26791 -17 26857 124 3 FreeSans 520 90 0 0 DM_H[1]
port 15 nsew
flabel metal3 s 26665 -17 26731 124 3 FreeSans 520 90 0 0 DM_H[2]
port 16 nsew
flabel metal3 s 26539 -17 26605 124 3 FreeSans 520 90 0 0 DM_H_N[0]
port 17 nsew
flabel metal3 s 26413 -17 26479 124 3 FreeSans 520 90 0 0 DM_H_N[1]
port 18 nsew
flabel metal3 s 20566 27158 20743 27455 3 FreeSans 520 0 0 0 VSSIO
port 20 nsew
flabel metal2 s 18906 26469 19032 27035 3 FreeSans 520 0 0 0 PAD
port 23 nsew
flabel metal2 s 8162 28590 8339 28887 3 FreeSans 520 0 0 0 VSSIO
port 20 nsew
flabel metal2 s 24403 27765 24580 28062 3 FreeSans 520 0 0 0 VSSIO
port 20 nsew
flabel metal1 s 23626 15958 23678 16046 3 FreeSans 520 90 0 0 OE_HS_H
port 25 nsew
flabel metal1 s 18821 33497 19162 33656 3 FreeSans 520 0 0 0 VDDIO
port 26 nsew
flabel metal1 s 23525 16019 23577 16108 3 FreeSans 520 90 0 0 PD_H[0]
port 27 nsew
flabel metal1 s 23445 16019 23497 16108 3 FreeSans 520 90 0 0 PD_H[1]
port 28 nsew
flabel metal1 s 23365 16019 23417 16108 3 FreeSans 520 90 0 0 PD_H[2]
port 29 nsew
flabel metal1 s 23285 16019 23337 16108 3 FreeSans 520 90 0 0 PD_H[3]
port 30 nsew
flabel metal1 s 23205 15957 23257 16046 3 FreeSans 520 90 0 0 PU_H_N[0]
port 31 nsew
flabel metal1 s 23125 15957 23177 16046 3 FreeSans 520 90 0 0 PU_H_N[1]
port 32 nsew
flabel metal1 s 23045 15957 23097 16046 3 FreeSans 520 90 0 0 PU_H_N[2]
port 33 nsew
flabel metal1 s 22965 15957 23017 16046 3 FreeSans 520 90 0 0 PU_H_N[3]
port 34 nsew
flabel metal1 s 23083 1691 23153 1780 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 35 nsew
flabel metal1 s 19389 31740 19686 31917 3 FreeSans 520 90 0 0 VDDIO
port 26 nsew
flabel metal1 s 22370 1898 22620 2182 3 FreeSans 520 0 0 0 VPWR_KA
port 36 nsew
flabel metal1 s 18821 86 19162 245 3 FreeSans 520 0 0 0 VDDIO
port 26 nsew
flabel comment s 26939 2789 26939 2789 0 FreeSans 600 90 0 0 DM_H[0]
flabel comment s 26826 2782 26826 2782 0 FreeSans 600 90 0 0 DM_H[1]
flabel comment s 26699 2772 26699 2772 0 FreeSans 600 90 0 0 DM_H[2]
flabel comment s 25581 1637 25581 1637 0 FreeSans 440 90 0 0 OE_H
flabel comment s 25432 1602 25432 1602 0 FreeSans 440 90 0 0 DRVLO_H_N
flabel comment s 25705 2758 25705 2758 0 FreeSans 440 90 0 0 DRVHI_H
flabel comment s 428 28951 428 28951 0 FreeSans 440 90 0 0 LV_NET
flabel comment s 26084 2682 26084 2682 0 FreeSans 440 90 0 0 SLEW_CTL_H_N[0]
flabel comment s 25831 2757 25831 2757 0 FreeSans 440 90 0 0 SLEW_CTL_H[1]
flabel comment s 25950 2747 25950 2747 0 FreeSans 440 90 0 0 SLEW_CTL_H[0]
flabel comment s 26214 2803 26214 2803 0 FreeSans 440 90 0 0 SLEW_CTL_H_N<>
flabel comment s 20136 32612 20136 32612 0 FreeSans 440 0 0 0 SLEW_CTL_H_N<>
flabel comment s 20015 32482 20015 32482 0 FreeSans 440 0 0 0 SLEW_CTL_H_N[0]
flabel comment s 20080 32348 20080 32348 0 FreeSans 440 0 0 0 SLEW_CTL_H[0]
flabel comment s 20090 32229 20090 32229 0 FreeSans 440 0 0 0 SLEW_CTL_H[1]
flabel comment s 22041 30395 22041 30395 0 FreeSans 440 90 0 0 OE_HS_H
flabel comment s 20904 29914 20904 29914 0 FreeSans 440 0 0 0 OE_H
flabel comment s 22041 30784 22041 30784 0 FreeSans 440 90 0 0 OE_HS_H
flabel comment s 24420 16590 24420 16590 0 FreeSans 440 90 0 0 SLOW_H_N
flabel comment s 26939 30876 26939 30876 0 FreeSans 200 90 0 0 DM_H[0]
flabel comment s 26826 30869 26826 30869 0 FreeSans 200 90 0 0 DM_H[1]
flabel comment s 26699 30859 26699 30859 0 FreeSans 200 90 0 0 DM_H[2]
flabel comment s 26575 30853 26575 30853 0 FreeSans 200 90 0 0 DM_H_N[0]
flabel comment s 26440 30841 26440 30841 0 FreeSans 200 90 0 0 DM_H_N[1]
flabel comment s 26317 30832 26317 30832 0 FreeSans 200 90 0 0 DM_H_N[2]
flabel comment s 26575 2766 26575 2766 0 FreeSans 600 90 0 0 DM_H_N[0]
flabel comment s 26440 2754 26440 2754 0 FreeSans 600 90 0 0 DM_H_N[1]
flabel comment s 26317 2745 26317 2745 0 FreeSans 600 90 0 0 DM_H_N[2]
<< properties >>
string GDS_END 38326494
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 38188572
<< end >>
