magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 4577 -193 5282 539
rect 5775 333 6109 605
rect 4727 -1281 5065 -650
<< pwell >>
rect 4830 3207 4916 3237
rect 4830 2357 5202 3207
rect 4802 2271 5395 2357
rect 4802 2242 5157 2271
rect 4799 1915 5157 2242
rect 4799 1713 5971 1915
rect 5165 1524 5971 1713
rect 4674 1263 5971 1524
rect 4674 942 5720 1263
rect 4674 612 5484 942
rect 5373 290 5625 442
rect 5373 104 6096 290
rect 5782 38 6096 104
<< nmos >>
rect 5861 64 5911 264
rect 5967 64 6017 264
<< mvnmos >>
rect 4878 2066 5078 2216
rect 4878 1739 5078 1889
rect 4753 1298 4873 1498
rect 4929 1298 5049 1498
rect 5244 1289 5364 1889
rect 5420 1289 5540 1889
rect 5596 1289 5716 1889
rect 5772 1289 5892 1889
<< mvpmos >>
rect 4867 -127 4987 473
rect 5043 -127 5163 473
rect 4846 -866 4946 -716
rect 4846 -1215 4946 -1065
<< mvnnmos >>
rect 4753 968 4933 1168
rect 4989 968 5169 1168
rect 5225 968 5405 1168
rect 5461 968 5641 1168
rect 4753 638 4933 838
rect 4989 638 5169 838
rect 5225 638 5405 838
rect 5399 183 5599 363
<< pmoshvt >>
rect 5864 369 5914 569
rect 5970 369 6020 569
<< nmoslvt >>
rect 4976 3098 5176 3128
rect 4976 3012 5176 3042
rect 4976 2926 5176 2956
rect 4976 2840 5176 2870
rect 4976 2754 5176 2784
rect 4976 2668 5176 2698
rect 4976 2582 5176 2612
rect 4976 2496 5176 2526
<< ndiff >>
rect 4976 3173 5176 3181
rect 4976 3139 4988 3173
rect 5022 3139 5056 3173
rect 5090 3139 5124 3173
rect 5158 3139 5176 3173
rect 4976 3128 5176 3139
rect 4976 3087 5176 3098
rect 4976 3053 4988 3087
rect 5022 3053 5056 3087
rect 5090 3053 5124 3087
rect 5158 3053 5176 3087
rect 4976 3042 5176 3053
rect 4976 3001 5176 3012
rect 4976 2967 4988 3001
rect 5022 2967 5056 3001
rect 5090 2967 5124 3001
rect 5158 2967 5176 3001
rect 4976 2956 5176 2967
rect 4976 2915 5176 2926
rect 4976 2881 4988 2915
rect 5022 2881 5056 2915
rect 5090 2881 5124 2915
rect 5158 2881 5176 2915
rect 4976 2870 5176 2881
rect 4976 2829 5176 2840
rect 4976 2795 4988 2829
rect 5022 2795 5056 2829
rect 5090 2795 5124 2829
rect 5158 2795 5176 2829
rect 4976 2784 5176 2795
rect 4976 2743 5176 2754
rect 4976 2709 4988 2743
rect 5022 2709 5056 2743
rect 5090 2709 5124 2743
rect 5158 2709 5176 2743
rect 4976 2698 5176 2709
rect 4976 2657 5176 2668
rect 4976 2623 4988 2657
rect 5022 2623 5056 2657
rect 5090 2623 5124 2657
rect 5158 2623 5176 2657
rect 4976 2612 5176 2623
rect 4976 2571 5176 2582
rect 4976 2537 4988 2571
rect 5022 2537 5056 2571
rect 5090 2537 5124 2571
rect 5158 2537 5176 2571
rect 4976 2526 5176 2537
rect 4976 2485 5176 2496
rect 4976 2451 4988 2485
rect 5022 2451 5056 2485
rect 5090 2451 5124 2485
rect 5158 2451 5176 2485
rect 4976 2443 5176 2451
rect 5808 246 5861 264
rect 5808 212 5816 246
rect 5850 212 5861 246
rect 5808 178 5861 212
rect 5808 144 5816 178
rect 5850 144 5861 178
rect 5808 110 5861 144
rect 5808 76 5816 110
rect 5850 76 5861 110
rect 5808 64 5861 76
rect 5911 246 5967 264
rect 5911 212 5922 246
rect 5956 212 5967 246
rect 5911 178 5967 212
rect 5911 144 5922 178
rect 5956 144 5967 178
rect 5911 110 5967 144
rect 5911 76 5922 110
rect 5956 76 5967 110
rect 5911 64 5967 76
rect 6017 246 6070 264
rect 6017 212 6028 246
rect 6062 212 6070 246
rect 6017 178 6070 212
rect 6017 144 6028 178
rect 6062 144 6070 178
rect 6017 110 6070 144
rect 6017 76 6028 110
rect 6062 76 6070 110
rect 6017 64 6070 76
<< pdiff >>
rect 5811 551 5864 569
rect 5811 517 5819 551
rect 5853 517 5864 551
rect 5811 483 5864 517
rect 5811 449 5819 483
rect 5853 449 5864 483
rect 5811 415 5864 449
rect 5811 381 5819 415
rect 5853 381 5864 415
rect 5811 369 5864 381
rect 5914 551 5970 569
rect 5914 517 5925 551
rect 5959 517 5970 551
rect 5914 483 5970 517
rect 5914 449 5925 483
rect 5959 449 5970 483
rect 5914 415 5970 449
rect 5914 381 5925 415
rect 5959 381 5970 415
rect 5914 369 5970 381
rect 6020 551 6073 569
rect 6020 517 6031 551
rect 6065 517 6073 551
rect 6020 483 6073 517
rect 6020 449 6031 483
rect 6065 449 6073 483
rect 6020 415 6073 449
rect 6020 381 6031 415
rect 6065 381 6073 415
rect 6020 369 6073 381
<< mvndiff >>
rect 4825 2204 4878 2216
rect 4825 2170 4833 2204
rect 4867 2170 4878 2204
rect 4825 2136 4878 2170
rect 4825 2102 4833 2136
rect 4867 2102 4878 2136
rect 4825 2066 4878 2102
rect 5078 2204 5131 2216
rect 5078 2170 5089 2204
rect 5123 2170 5131 2204
rect 5078 2136 5131 2170
rect 5078 2102 5089 2136
rect 5123 2102 5131 2136
rect 5078 2066 5131 2102
rect 4825 1853 4878 1889
rect 4825 1819 4833 1853
rect 4867 1819 4878 1853
rect 4825 1785 4878 1819
rect 4825 1751 4833 1785
rect 4867 1751 4878 1785
rect 4825 1739 4878 1751
rect 5078 1853 5131 1889
rect 5078 1819 5089 1853
rect 5123 1819 5131 1853
rect 5078 1785 5131 1819
rect 5078 1751 5089 1785
rect 5123 1751 5131 1785
rect 5078 1739 5131 1751
rect 5191 1811 5244 1889
rect 5191 1777 5199 1811
rect 5233 1777 5244 1811
rect 5191 1743 5244 1777
rect 5191 1709 5199 1743
rect 5233 1709 5244 1743
rect 5191 1675 5244 1709
rect 5191 1641 5199 1675
rect 5233 1641 5244 1675
rect 5191 1607 5244 1641
rect 5191 1573 5199 1607
rect 5233 1573 5244 1607
rect 5191 1539 5244 1573
rect 5191 1505 5199 1539
rect 5233 1505 5244 1539
rect 4700 1480 4753 1498
rect 4700 1446 4708 1480
rect 4742 1446 4753 1480
rect 4700 1412 4753 1446
rect 4700 1378 4708 1412
rect 4742 1378 4753 1412
rect 4700 1344 4753 1378
rect 4700 1310 4708 1344
rect 4742 1310 4753 1344
rect 4700 1298 4753 1310
rect 4873 1480 4929 1498
rect 4873 1446 4884 1480
rect 4918 1446 4929 1480
rect 4873 1412 4929 1446
rect 4873 1378 4884 1412
rect 4918 1378 4929 1412
rect 4873 1344 4929 1378
rect 4873 1310 4884 1344
rect 4918 1310 4929 1344
rect 4873 1298 4929 1310
rect 5049 1480 5102 1498
rect 5049 1446 5060 1480
rect 5094 1446 5102 1480
rect 5049 1412 5102 1446
rect 5049 1378 5060 1412
rect 5094 1378 5102 1412
rect 5049 1344 5102 1378
rect 5049 1310 5060 1344
rect 5094 1310 5102 1344
rect 5049 1298 5102 1310
rect 5191 1471 5244 1505
rect 5191 1437 5199 1471
rect 5233 1437 5244 1471
rect 5191 1403 5244 1437
rect 5191 1369 5199 1403
rect 5233 1369 5244 1403
rect 5191 1335 5244 1369
rect 5191 1301 5199 1335
rect 5233 1301 5244 1335
rect 5191 1289 5244 1301
rect 5364 1811 5420 1889
rect 5364 1777 5375 1811
rect 5409 1777 5420 1811
rect 5364 1743 5420 1777
rect 5364 1709 5375 1743
rect 5409 1709 5420 1743
rect 5364 1675 5420 1709
rect 5364 1641 5375 1675
rect 5409 1641 5420 1675
rect 5364 1607 5420 1641
rect 5364 1573 5375 1607
rect 5409 1573 5420 1607
rect 5364 1539 5420 1573
rect 5364 1505 5375 1539
rect 5409 1505 5420 1539
rect 5364 1471 5420 1505
rect 5364 1437 5375 1471
rect 5409 1437 5420 1471
rect 5364 1403 5420 1437
rect 5364 1369 5375 1403
rect 5409 1369 5420 1403
rect 5364 1335 5420 1369
rect 5364 1301 5375 1335
rect 5409 1301 5420 1335
rect 5364 1289 5420 1301
rect 5540 1811 5596 1889
rect 5540 1777 5551 1811
rect 5585 1777 5596 1811
rect 5540 1743 5596 1777
rect 5540 1709 5551 1743
rect 5585 1709 5596 1743
rect 5540 1675 5596 1709
rect 5540 1641 5551 1675
rect 5585 1641 5596 1675
rect 5540 1607 5596 1641
rect 5540 1573 5551 1607
rect 5585 1573 5596 1607
rect 5540 1539 5596 1573
rect 5540 1505 5551 1539
rect 5585 1505 5596 1539
rect 5540 1471 5596 1505
rect 5540 1437 5551 1471
rect 5585 1437 5596 1471
rect 5540 1403 5596 1437
rect 5540 1369 5551 1403
rect 5585 1369 5596 1403
rect 5540 1335 5596 1369
rect 5540 1301 5551 1335
rect 5585 1301 5596 1335
rect 5540 1289 5596 1301
rect 5716 1811 5772 1889
rect 5716 1777 5727 1811
rect 5761 1777 5772 1811
rect 5716 1743 5772 1777
rect 5716 1709 5727 1743
rect 5761 1709 5772 1743
rect 5716 1675 5772 1709
rect 5716 1641 5727 1675
rect 5761 1641 5772 1675
rect 5716 1607 5772 1641
rect 5716 1573 5727 1607
rect 5761 1573 5772 1607
rect 5716 1539 5772 1573
rect 5716 1505 5727 1539
rect 5761 1505 5772 1539
rect 5716 1471 5772 1505
rect 5716 1437 5727 1471
rect 5761 1437 5772 1471
rect 5716 1403 5772 1437
rect 5716 1369 5727 1403
rect 5761 1369 5772 1403
rect 5716 1335 5772 1369
rect 5716 1301 5727 1335
rect 5761 1301 5772 1335
rect 5716 1289 5772 1301
rect 5892 1811 5945 1889
rect 5892 1777 5903 1811
rect 5937 1777 5945 1811
rect 5892 1743 5945 1777
rect 5892 1709 5903 1743
rect 5937 1709 5945 1743
rect 5892 1675 5945 1709
rect 5892 1641 5903 1675
rect 5937 1641 5945 1675
rect 5892 1607 5945 1641
rect 5892 1573 5903 1607
rect 5937 1573 5945 1607
rect 5892 1539 5945 1573
rect 5892 1505 5903 1539
rect 5937 1505 5945 1539
rect 5892 1471 5945 1505
rect 5892 1437 5903 1471
rect 5937 1437 5945 1471
rect 5892 1403 5945 1437
rect 5892 1369 5903 1403
rect 5937 1369 5945 1403
rect 5892 1335 5945 1369
rect 5892 1301 5903 1335
rect 5937 1301 5945 1335
rect 5892 1289 5945 1301
rect 4700 1150 4753 1168
rect 4700 1116 4708 1150
rect 4742 1116 4753 1150
rect 4700 1082 4753 1116
rect 4700 1048 4708 1082
rect 4742 1048 4753 1082
rect 4700 1014 4753 1048
rect 4700 980 4708 1014
rect 4742 980 4753 1014
rect 4700 968 4753 980
rect 4933 1150 4989 1168
rect 4933 1116 4944 1150
rect 4978 1116 4989 1150
rect 4933 1082 4989 1116
rect 4933 1048 4944 1082
rect 4978 1048 4989 1082
rect 4933 1014 4989 1048
rect 4933 980 4944 1014
rect 4978 980 4989 1014
rect 4933 968 4989 980
rect 5169 1150 5225 1168
rect 5169 1116 5180 1150
rect 5214 1116 5225 1150
rect 5169 1082 5225 1116
rect 5169 1048 5180 1082
rect 5214 1048 5225 1082
rect 5169 1014 5225 1048
rect 5169 980 5180 1014
rect 5214 980 5225 1014
rect 5169 968 5225 980
rect 5405 1150 5461 1168
rect 5405 1116 5416 1150
rect 5450 1116 5461 1150
rect 5405 1082 5461 1116
rect 5405 1048 5416 1082
rect 5450 1048 5461 1082
rect 5405 1014 5461 1048
rect 5405 980 5416 1014
rect 5450 980 5461 1014
rect 5405 968 5461 980
rect 5641 1150 5694 1168
rect 5641 1116 5652 1150
rect 5686 1116 5694 1150
rect 5641 1082 5694 1116
rect 5641 1048 5652 1082
rect 5686 1048 5694 1082
rect 5641 1014 5694 1048
rect 5641 980 5652 1014
rect 5686 980 5694 1014
rect 5641 968 5694 980
rect 4700 820 4753 838
rect 4700 786 4708 820
rect 4742 786 4753 820
rect 4700 752 4753 786
rect 4700 718 4708 752
rect 4742 718 4753 752
rect 4700 684 4753 718
rect 4700 650 4708 684
rect 4742 650 4753 684
rect 4700 638 4753 650
rect 4933 820 4989 838
rect 4933 786 4944 820
rect 4978 786 4989 820
rect 4933 752 4989 786
rect 4933 718 4944 752
rect 4978 718 4989 752
rect 4933 684 4989 718
rect 4933 650 4944 684
rect 4978 650 4989 684
rect 4933 638 4989 650
rect 5169 820 5225 838
rect 5169 786 5180 820
rect 5214 786 5225 820
rect 5169 752 5225 786
rect 5169 718 5180 752
rect 5214 718 5225 752
rect 5169 684 5225 718
rect 5169 650 5180 684
rect 5214 650 5225 684
rect 5169 638 5225 650
rect 5405 820 5458 838
rect 5405 786 5416 820
rect 5450 786 5458 820
rect 5405 752 5458 786
rect 5405 718 5416 752
rect 5450 718 5458 752
rect 5405 684 5458 718
rect 5405 650 5416 684
rect 5450 650 5458 684
rect 5405 638 5458 650
rect 5399 408 5599 416
rect 5399 374 5417 408
rect 5451 374 5485 408
rect 5519 374 5553 408
rect 5587 374 5599 408
rect 5399 363 5599 374
rect 5399 172 5599 183
rect 5399 138 5417 172
rect 5451 138 5485 172
rect 5519 138 5553 172
rect 5587 138 5599 172
rect 5399 130 5599 138
<< mvpdiff >>
rect 4814 461 4867 473
rect 4814 427 4822 461
rect 4856 427 4867 461
rect 4814 393 4867 427
rect 4814 359 4822 393
rect 4856 359 4867 393
rect 4814 325 4867 359
rect 4814 291 4822 325
rect 4856 291 4867 325
rect 4814 257 4867 291
rect 4814 223 4822 257
rect 4856 223 4867 257
rect 4814 189 4867 223
rect 4814 155 4822 189
rect 4856 155 4867 189
rect 4814 121 4867 155
rect 4814 87 4822 121
rect 4856 87 4867 121
rect 4814 53 4867 87
rect 4814 19 4822 53
rect 4856 19 4867 53
rect 4814 -15 4867 19
rect 4814 -49 4822 -15
rect 4856 -49 4867 -15
rect 4814 -127 4867 -49
rect 4987 461 5043 473
rect 4987 427 4998 461
rect 5032 427 5043 461
rect 4987 393 5043 427
rect 4987 359 4998 393
rect 5032 359 5043 393
rect 4987 325 5043 359
rect 4987 291 4998 325
rect 5032 291 5043 325
rect 4987 257 5043 291
rect 4987 223 4998 257
rect 5032 223 5043 257
rect 4987 189 5043 223
rect 4987 155 4998 189
rect 5032 155 5043 189
rect 4987 121 5043 155
rect 4987 87 4998 121
rect 5032 87 5043 121
rect 4987 53 5043 87
rect 4987 19 4998 53
rect 5032 19 5043 53
rect 4987 -15 5043 19
rect 4987 -49 4998 -15
rect 5032 -49 5043 -15
rect 4987 -127 5043 -49
rect 5163 461 5216 473
rect 5163 427 5174 461
rect 5208 427 5216 461
rect 5163 393 5216 427
rect 5163 359 5174 393
rect 5208 359 5216 393
rect 5163 325 5216 359
rect 5163 291 5174 325
rect 5208 291 5216 325
rect 5163 257 5216 291
rect 5163 223 5174 257
rect 5208 223 5216 257
rect 5163 189 5216 223
rect 5163 155 5174 189
rect 5208 155 5216 189
rect 5163 121 5216 155
rect 5163 87 5174 121
rect 5208 87 5216 121
rect 5163 53 5216 87
rect 5163 19 5174 53
rect 5208 19 5216 53
rect 5163 -15 5216 19
rect 5163 -49 5174 -15
rect 5208 -49 5216 -15
rect 5163 -127 5216 -49
rect 4793 -752 4846 -716
rect 4793 -786 4801 -752
rect 4835 -786 4846 -752
rect 4793 -820 4846 -786
rect 4793 -854 4801 -820
rect 4835 -854 4846 -820
rect 4793 -866 4846 -854
rect 4946 -752 4999 -716
rect 4946 -786 4957 -752
rect 4991 -786 4999 -752
rect 4946 -820 4999 -786
rect 4946 -854 4957 -820
rect 4991 -854 4999 -820
rect 4946 -866 4999 -854
rect 4793 -1101 4846 -1065
rect 4793 -1135 4801 -1101
rect 4835 -1135 4846 -1101
rect 4793 -1169 4846 -1135
rect 4793 -1203 4801 -1169
rect 4835 -1203 4846 -1169
rect 4793 -1215 4846 -1203
rect 4946 -1101 4999 -1065
rect 4946 -1135 4957 -1101
rect 4991 -1135 4999 -1101
rect 4946 -1169 4999 -1135
rect 4946 -1203 4957 -1169
rect 4991 -1203 4999 -1169
rect 4946 -1215 4999 -1203
<< ndiffc >>
rect 4988 3139 5022 3173
rect 5056 3139 5090 3173
rect 5124 3139 5158 3173
rect 4988 3053 5022 3087
rect 5056 3053 5090 3087
rect 5124 3053 5158 3087
rect 4988 2967 5022 3001
rect 5056 2967 5090 3001
rect 5124 2967 5158 3001
rect 4988 2881 5022 2915
rect 5056 2881 5090 2915
rect 5124 2881 5158 2915
rect 4988 2795 5022 2829
rect 5056 2795 5090 2829
rect 5124 2795 5158 2829
rect 4988 2709 5022 2743
rect 5056 2709 5090 2743
rect 5124 2709 5158 2743
rect 4988 2623 5022 2657
rect 5056 2623 5090 2657
rect 5124 2623 5158 2657
rect 4988 2537 5022 2571
rect 5056 2537 5090 2571
rect 5124 2537 5158 2571
rect 4988 2451 5022 2485
rect 5056 2451 5090 2485
rect 5124 2451 5158 2485
rect 5816 212 5850 246
rect 5816 144 5850 178
rect 5816 76 5850 110
rect 5922 212 5956 246
rect 5922 144 5956 178
rect 5922 76 5956 110
rect 6028 212 6062 246
rect 6028 144 6062 178
rect 6028 76 6062 110
<< pdiffc >>
rect 5819 517 5853 551
rect 5819 449 5853 483
rect 5819 381 5853 415
rect 5925 517 5959 551
rect 5925 449 5959 483
rect 5925 381 5959 415
rect 6031 517 6065 551
rect 6031 449 6065 483
rect 6031 381 6065 415
<< mvndiffc >>
rect 4833 2170 4867 2204
rect 4833 2102 4867 2136
rect 5089 2170 5123 2204
rect 5089 2102 5123 2136
rect 4833 1819 4867 1853
rect 4833 1751 4867 1785
rect 5089 1819 5123 1853
rect 5089 1751 5123 1785
rect 5199 1777 5233 1811
rect 5199 1709 5233 1743
rect 5199 1641 5233 1675
rect 5199 1573 5233 1607
rect 5199 1505 5233 1539
rect 4708 1446 4742 1480
rect 4708 1378 4742 1412
rect 4708 1310 4742 1344
rect 4884 1446 4918 1480
rect 4884 1378 4918 1412
rect 4884 1310 4918 1344
rect 5060 1446 5094 1480
rect 5060 1378 5094 1412
rect 5060 1310 5094 1344
rect 5199 1437 5233 1471
rect 5199 1369 5233 1403
rect 5199 1301 5233 1335
rect 5375 1777 5409 1811
rect 5375 1709 5409 1743
rect 5375 1641 5409 1675
rect 5375 1573 5409 1607
rect 5375 1505 5409 1539
rect 5375 1437 5409 1471
rect 5375 1369 5409 1403
rect 5375 1301 5409 1335
rect 5551 1777 5585 1811
rect 5551 1709 5585 1743
rect 5551 1641 5585 1675
rect 5551 1573 5585 1607
rect 5551 1505 5585 1539
rect 5551 1437 5585 1471
rect 5551 1369 5585 1403
rect 5551 1301 5585 1335
rect 5727 1777 5761 1811
rect 5727 1709 5761 1743
rect 5727 1641 5761 1675
rect 5727 1573 5761 1607
rect 5727 1505 5761 1539
rect 5727 1437 5761 1471
rect 5727 1369 5761 1403
rect 5727 1301 5761 1335
rect 5903 1777 5937 1811
rect 5903 1709 5937 1743
rect 5903 1641 5937 1675
rect 5903 1573 5937 1607
rect 5903 1505 5937 1539
rect 5903 1437 5937 1471
rect 5903 1369 5937 1403
rect 5903 1301 5937 1335
rect 4708 1116 4742 1150
rect 4708 1048 4742 1082
rect 4708 980 4742 1014
rect 4944 1116 4978 1150
rect 4944 1048 4978 1082
rect 4944 980 4978 1014
rect 5180 1116 5214 1150
rect 5180 1048 5214 1082
rect 5180 980 5214 1014
rect 5416 1116 5450 1150
rect 5416 1048 5450 1082
rect 5416 980 5450 1014
rect 5652 1116 5686 1150
rect 5652 1048 5686 1082
rect 5652 980 5686 1014
rect 4708 786 4742 820
rect 4708 718 4742 752
rect 4708 650 4742 684
rect 4944 786 4978 820
rect 4944 718 4978 752
rect 4944 650 4978 684
rect 5180 786 5214 820
rect 5180 718 5214 752
rect 5180 650 5214 684
rect 5416 786 5450 820
rect 5416 718 5450 752
rect 5416 650 5450 684
rect 5417 374 5451 408
rect 5485 374 5519 408
rect 5553 374 5587 408
rect 5417 138 5451 172
rect 5485 138 5519 172
rect 5553 138 5587 172
<< mvpdiffc >>
rect 4822 427 4856 461
rect 4822 359 4856 393
rect 4822 291 4856 325
rect 4822 223 4856 257
rect 4822 155 4856 189
rect 4822 87 4856 121
rect 4822 19 4856 53
rect 4822 -49 4856 -15
rect 4998 427 5032 461
rect 4998 359 5032 393
rect 4998 291 5032 325
rect 4998 223 5032 257
rect 4998 155 5032 189
rect 4998 87 5032 121
rect 4998 19 5032 53
rect 4998 -49 5032 -15
rect 5174 427 5208 461
rect 5174 359 5208 393
rect 5174 291 5208 325
rect 5174 223 5208 257
rect 5174 155 5208 189
rect 5174 87 5208 121
rect 5174 19 5208 53
rect 5174 -49 5208 -15
rect 4801 -786 4835 -752
rect 4801 -854 4835 -820
rect 4957 -786 4991 -752
rect 4957 -854 4991 -820
rect 4801 -1135 4835 -1101
rect 4801 -1203 4835 -1169
rect 4957 -1135 4991 -1101
rect 4957 -1203 4991 -1169
<< psubdiff >>
rect 4856 3177 4890 3211
rect 4856 3071 4890 3143
rect 4856 2965 4890 3037
rect 4856 2859 4890 2931
rect 4856 2753 4890 2825
rect 4856 2647 4890 2719
rect 4856 2541 4890 2613
rect 4856 2473 4890 2507
<< mvpsubdiff >>
rect 4828 2297 4852 2331
rect 4886 2297 4929 2331
rect 4963 2297 5006 2331
rect 5040 2297 5083 2331
rect 5117 2297 5159 2331
rect 5193 2297 5235 2331
rect 5269 2297 5311 2331
rect 5345 2297 5369 2331
<< mvnsubdiff >>
rect 4643 449 4677 473
rect 4643 375 4677 415
rect 4643 301 4677 341
rect 4643 227 4677 267
rect 4643 153 4677 193
rect 4643 79 4677 119
rect 4643 5 4677 45
rect 4643 -69 4677 -29
rect 4643 -127 4677 -103
<< psubdiffcont >>
rect 4856 3143 4890 3177
rect 4856 3037 4890 3071
rect 4856 2931 4890 2965
rect 4856 2825 4890 2859
rect 4856 2719 4890 2753
rect 4856 2613 4890 2647
rect 4856 2507 4890 2541
<< mvpsubdiffcont >>
rect 4852 2297 4886 2331
rect 4929 2297 4963 2331
rect 5006 2297 5040 2331
rect 5083 2297 5117 2331
rect 5159 2297 5193 2331
rect 5235 2297 5269 2331
rect 5311 2297 5345 2331
<< mvnsubdiffcont >>
rect 4643 415 4677 449
rect 4643 341 4677 375
rect 4643 267 4677 301
rect 4643 193 4677 227
rect 4643 119 4677 153
rect 4643 45 4677 79
rect 4643 -29 4677 5
rect 4643 -103 4677 -69
<< poly >>
rect 4944 3098 4976 3128
rect 5176 3112 5274 3128
rect 5176 3098 5224 3112
rect 5208 3078 5224 3098
rect 5258 3078 5274 3112
rect 5208 3042 5274 3078
rect 4944 3012 4976 3042
rect 5176 3038 5274 3042
rect 5176 3012 5224 3038
rect 5208 3004 5224 3012
rect 5258 3004 5274 3038
rect 5208 2964 5274 3004
rect 5208 2956 5224 2964
rect 4944 2926 4976 2956
rect 5176 2930 5224 2956
rect 5258 2930 5274 2964
rect 5176 2926 5274 2930
rect 5208 2890 5274 2926
rect 5208 2870 5224 2890
rect 4944 2840 4976 2870
rect 5176 2856 5224 2870
rect 5258 2856 5274 2890
rect 5176 2840 5274 2856
rect 4944 2754 4976 2784
rect 5176 2768 5274 2784
rect 5176 2754 5224 2768
rect 5208 2734 5224 2754
rect 5258 2734 5274 2768
rect 5208 2698 5274 2734
rect 4944 2668 4976 2698
rect 5176 2694 5274 2698
rect 5176 2668 5224 2694
rect 5208 2660 5224 2668
rect 5258 2660 5274 2694
rect 5208 2620 5274 2660
rect 5208 2612 5224 2620
rect 4944 2582 4976 2612
rect 5176 2586 5224 2612
rect 5258 2586 5274 2620
rect 5176 2582 5274 2586
rect 5208 2546 5274 2582
rect 5208 2526 5224 2546
rect 4944 2496 4976 2526
rect 5176 2512 5224 2526
rect 5258 2512 5274 2546
rect 5176 2496 5274 2512
rect 4878 2216 5078 2248
rect 4878 2018 5078 2066
rect 4878 1984 4894 2018
rect 4928 1984 5028 2018
rect 5062 1984 5078 2018
rect 4878 1968 5078 1984
rect 5244 2048 5364 2064
rect 5244 2014 5289 2048
rect 5323 2014 5364 2048
rect 5244 1980 5364 2014
rect 5244 1946 5289 1980
rect 5323 1946 5364 1980
rect 4878 1889 5078 1921
rect 5244 1889 5364 1946
rect 5420 2048 5540 2064
rect 5420 2014 5464 2048
rect 5498 2014 5540 2048
rect 5420 1980 5540 2014
rect 5420 1946 5464 1980
rect 5498 1946 5540 1980
rect 5420 1889 5540 1946
rect 5596 2048 5716 2085
rect 5596 2014 5629 2048
rect 5663 2014 5716 2048
rect 5596 1980 5716 2014
rect 5596 1946 5629 1980
rect 5663 1946 5716 1980
rect 5596 1889 5716 1946
rect 5772 2048 5892 2064
rect 5772 2014 5814 2048
rect 5848 2014 5892 2048
rect 5772 1980 5892 2014
rect 5772 1946 5814 1980
rect 5848 1946 5892 1980
rect 5772 1889 5892 1946
rect 4878 1691 5078 1739
rect 4878 1657 4894 1691
rect 4928 1657 5008 1691
rect 5042 1657 5078 1691
rect 4878 1641 5078 1657
rect 4739 1580 4873 1596
rect 4739 1546 4755 1580
rect 4789 1546 4823 1580
rect 4857 1546 4873 1580
rect 4739 1530 4873 1546
rect 4753 1498 4873 1530
rect 4929 1580 5063 1596
rect 4929 1546 4945 1580
rect 4979 1546 5013 1580
rect 5047 1546 5063 1580
rect 4929 1530 5063 1546
rect 4929 1498 5049 1530
rect 4753 1266 4873 1298
rect 4929 1266 5049 1298
rect 5244 1257 5364 1289
rect 5420 1257 5540 1289
rect 5596 1257 5716 1289
rect 5772 1257 5892 1289
rect 4753 1168 4933 1200
rect 4989 1168 5169 1200
rect 5225 1168 5405 1200
rect 5461 1168 5641 1200
rect 4753 936 4933 968
rect 4989 936 5169 968
rect 5225 936 5405 968
rect 5461 936 5641 968
rect 4753 920 5641 936
rect 4753 886 4769 920
rect 4803 886 4837 920
rect 4871 886 4905 920
rect 4939 886 4973 920
rect 5007 886 5041 920
rect 5075 886 5109 920
rect 5143 886 5177 920
rect 5211 886 5246 920
rect 5280 886 5315 920
rect 5349 886 5384 920
rect 5418 886 5453 920
rect 5487 886 5522 920
rect 5556 886 5591 920
rect 5625 886 5641 920
rect 4753 870 5641 886
rect 4753 838 4933 870
rect 4989 838 5169 870
rect 5225 838 5405 870
rect 5895 700 6029 716
rect 5895 666 5911 700
rect 5945 666 5979 700
rect 6013 666 6029 700
rect 5895 650 6029 666
rect 4753 606 4933 638
rect 4989 606 5169 638
rect 5225 606 5405 638
rect 5864 569 5914 595
rect 5970 569 6020 650
rect 4867 473 4987 505
rect 5043 473 5163 505
rect 5367 183 5399 363
rect 5599 347 5697 363
rect 5599 313 5647 347
rect 5681 313 5697 347
rect 5864 343 5914 369
rect 5970 343 6020 369
rect 5599 233 5697 313
rect 5861 290 5914 343
rect 5967 290 6020 343
rect 5861 264 5911 290
rect 5967 264 6017 290
rect 5599 199 5647 233
rect 5681 199 5697 233
rect 5599 183 5697 199
rect 5861 -4 5911 64
rect 5967 38 6017 64
rect 5848 -20 5914 -4
rect 5848 -54 5864 -20
rect 5898 -54 5914 -20
rect 5848 -88 5914 -54
rect 5848 -122 5864 -88
rect 5898 -122 5914 -88
rect 4867 -159 4987 -127
rect 4853 -175 4987 -159
rect 4853 -209 4869 -175
rect 4903 -209 4937 -175
rect 4971 -209 4987 -175
rect 4853 -225 4987 -209
rect 5043 -159 5163 -127
rect 5848 -138 5914 -122
rect 5043 -175 5177 -159
rect 5043 -209 5059 -175
rect 5093 -209 5127 -175
rect 5161 -209 5177 -175
rect 5043 -225 5177 -209
rect 4846 -634 4980 -618
rect 4846 -668 4862 -634
rect 4896 -668 4930 -634
rect 4964 -668 4980 -634
rect 4846 -684 4980 -668
rect 4846 -716 4946 -684
rect 4846 -898 4946 -866
rect 4846 -983 4980 -967
rect 4846 -1017 4862 -983
rect 4896 -1017 4930 -983
rect 4964 -1017 4980 -983
rect 4846 -1033 4980 -1017
rect 4846 -1065 4946 -1033
rect 4846 -1247 4946 -1215
<< polycont >>
rect 5224 3078 5258 3112
rect 5224 3004 5258 3038
rect 5224 2930 5258 2964
rect 5224 2856 5258 2890
rect 5224 2734 5258 2768
rect 5224 2660 5258 2694
rect 5224 2586 5258 2620
rect 5224 2512 5258 2546
rect 4894 1984 4928 2018
rect 5028 1984 5062 2018
rect 5289 2014 5323 2048
rect 5289 1946 5323 1980
rect 5464 2014 5498 2048
rect 5464 1946 5498 1980
rect 5629 2014 5663 2048
rect 5629 1946 5663 1980
rect 5814 2014 5848 2048
rect 5814 1946 5848 1980
rect 4894 1657 4928 1691
rect 5008 1657 5042 1691
rect 4755 1546 4789 1580
rect 4823 1546 4857 1580
rect 4945 1546 4979 1580
rect 5013 1546 5047 1580
rect 4769 886 4803 920
rect 4837 886 4871 920
rect 4905 886 4939 920
rect 4973 886 5007 920
rect 5041 886 5075 920
rect 5109 886 5143 920
rect 5177 886 5211 920
rect 5246 886 5280 920
rect 5315 886 5349 920
rect 5384 886 5418 920
rect 5453 886 5487 920
rect 5522 886 5556 920
rect 5591 886 5625 920
rect 5911 666 5945 700
rect 5979 666 6013 700
rect 5647 313 5681 347
rect 5647 199 5681 233
rect 5864 -54 5898 -20
rect 5864 -122 5898 -88
rect 4869 -209 4903 -175
rect 4937 -209 4971 -175
rect 5059 -209 5093 -175
rect 5127 -209 5161 -175
rect 4862 -668 4896 -634
rect 4930 -668 4964 -634
rect 4862 -1017 4896 -983
rect 4930 -1017 4964 -983
<< locali >>
rect 4856 3177 4890 3211
rect 4884 3138 4890 3143
rect 4956 3139 4988 3173
rect 5028 3139 5056 3173
rect 5090 3139 5124 3173
rect 5158 3139 5174 3173
rect 4850 3097 4890 3138
rect 4884 3071 4890 3097
rect 5224 3112 5232 3128
rect 4850 3037 4856 3063
rect 4972 3053 4988 3087
rect 5022 3053 5056 3087
rect 5114 3053 5124 3087
rect 5258 3078 5266 3094
rect 4850 3022 4890 3037
rect 4884 2988 4890 3022
rect 5224 3044 5266 3078
rect 5224 3038 5232 3044
rect 5258 3004 5266 3010
rect 4850 2965 4890 2988
rect 4956 2967 4988 3001
rect 5028 2967 5056 3001
rect 5090 2967 5124 3001
rect 5158 2967 5174 3001
rect 4850 2947 4856 2965
rect 4884 2913 4890 2931
rect 5224 2964 5266 3004
rect 5258 2959 5266 2964
rect 5224 2925 5232 2930
rect 4850 2871 4890 2913
rect 4972 2881 4988 2915
rect 5022 2881 5056 2915
rect 5114 2881 5124 2915
rect 5224 2890 5266 2925
rect 4884 2859 4890 2871
rect 5258 2874 5266 2890
rect 5224 2840 5232 2856
rect 4850 2825 4856 2837
rect 4850 2795 4890 2825
rect 4956 2795 4988 2829
rect 5028 2795 5056 2829
rect 5090 2795 5124 2829
rect 5158 2795 5174 2829
rect 4884 2761 4890 2795
rect 4850 2753 4890 2761
rect 4850 2719 4856 2753
rect 5224 2768 5258 2784
rect 4884 2685 4890 2719
rect 4972 2709 4988 2743
rect 5022 2709 5056 2743
rect 5114 2709 5124 2743
rect 5224 2726 5258 2734
rect 4850 2647 4890 2685
rect 5224 2694 5232 2726
rect 5258 2660 5266 2692
rect 4850 2643 4856 2647
rect 4956 2623 4988 2657
rect 5028 2623 5056 2657
rect 5090 2623 5124 2657
rect 5158 2623 5174 2657
rect 5224 2628 5266 2660
rect 4884 2609 4890 2613
rect 4850 2567 4890 2609
rect 5224 2620 5232 2628
rect 5258 2586 5266 2594
rect 4884 2541 4890 2567
rect 4972 2537 4988 2571
rect 5022 2537 5056 2571
rect 5114 2537 5124 2571
rect 5224 2546 5266 2586
rect 4850 2507 4856 2533
rect 4850 2491 4890 2507
rect 5258 2530 5266 2546
rect 5224 2496 5232 2512
rect 4884 2473 4890 2491
rect 4956 2451 4988 2485
rect 5028 2451 5056 2485
rect 5090 2451 5124 2485
rect 5158 2451 5174 2485
rect 4828 2297 4839 2331
rect 4886 2297 4920 2331
rect 4963 2297 5001 2331
rect 5040 2297 5082 2331
rect 5117 2297 5159 2331
rect 5196 2297 5235 2331
rect 5276 2297 5311 2331
rect 5356 2297 5369 2331
rect 5088 2236 5425 2263
rect 4833 2204 4867 2220
rect 4833 2136 4867 2169
rect 5088 2204 5383 2236
rect 5088 2170 5089 2204
rect 5123 2202 5383 2204
rect 5417 2202 5425 2236
rect 5123 2170 5425 2202
rect 5088 2164 5425 2170
rect 5088 2136 5383 2164
rect 5088 2102 5089 2136
rect 5123 2130 5383 2136
rect 5417 2130 5425 2164
rect 5123 2102 5425 2130
rect 5088 2098 5425 2102
rect 4833 2086 4867 2097
rect 5089 2086 5123 2098
rect 5289 2048 5323 2064
rect 4878 1984 4894 2018
rect 4928 1984 5028 2018
rect 5062 1984 5123 2018
rect 4878 1923 5123 1984
rect 4833 1853 4867 1869
rect 4833 1788 4867 1819
rect 5089 1853 5123 1923
rect 5289 1980 5323 2008
rect 5289 1896 5323 1936
rect 5464 2048 5498 2064
rect 5464 1980 5498 2008
rect 5464 1930 5498 1936
rect 5629 2048 5663 2064
rect 5629 1980 5663 2008
rect 5629 1930 5663 1936
rect 5802 2048 5851 2064
rect 5802 2014 5814 2048
rect 5848 2014 5851 2048
rect 5802 2012 5851 2014
rect 5802 1946 5814 2012
rect 5848 1946 5851 2012
rect 5802 1940 5851 1946
rect 5802 1906 5814 1940
rect 5848 1906 5851 1940
rect 5802 1896 5851 1906
rect 5288 1861 5851 1896
rect 4858 1785 4896 1788
rect 4867 1754 4896 1785
rect 5089 1785 5123 1787
rect 4833 1735 4867 1751
rect 5089 1749 5123 1751
rect 5184 1811 5233 1844
rect 5184 1777 5199 1811
rect 5184 1743 5233 1777
rect 5184 1709 5199 1743
rect 4878 1657 4894 1691
rect 4928 1657 5008 1691
rect 5042 1657 5063 1691
rect 4929 1587 5063 1657
rect 4929 1580 4957 1587
rect 4991 1580 5029 1587
rect 4739 1546 4755 1580
rect 4789 1569 4796 1580
rect 4789 1546 4823 1569
rect 4857 1546 4873 1580
rect 4929 1546 4945 1580
rect 4991 1553 5013 1580
rect 4979 1546 5013 1553
rect 5047 1546 5063 1553
rect 5184 1675 5233 1709
rect 5184 1641 5199 1675
rect 5184 1607 5233 1641
rect 5184 1573 5199 1607
rect 4796 1531 4830 1546
rect 5184 1539 5233 1573
rect 5184 1505 5199 1539
rect 4708 1425 4742 1446
rect 4708 1344 4742 1378
rect 4708 1294 4742 1310
rect 4884 1480 4918 1496
rect 5062 1480 5100 1502
rect 5094 1468 5100 1480
rect 5184 1471 5233 1505
rect 4884 1412 4918 1446
rect 4884 1344 4918 1377
rect 4884 1294 4918 1305
rect 5060 1412 5094 1446
rect 5060 1344 5094 1378
rect 5060 1294 5094 1310
rect 5184 1437 5199 1471
rect 5184 1403 5233 1437
rect 5184 1369 5199 1403
rect 5184 1335 5233 1369
rect 5184 1301 5199 1335
rect 5184 1166 5233 1301
rect 5349 1821 5409 1827
rect 5383 1811 5409 1821
rect 5349 1777 5375 1787
rect 5349 1749 5409 1777
rect 5383 1743 5409 1749
rect 5349 1709 5375 1715
rect 5349 1675 5409 1709
rect 5349 1641 5375 1675
rect 5349 1607 5409 1641
rect 5349 1573 5375 1607
rect 5349 1539 5409 1573
rect 5349 1505 5375 1539
rect 5349 1471 5409 1505
rect 5349 1437 5375 1471
rect 5349 1403 5409 1437
rect 5551 1811 5585 1827
rect 5551 1743 5585 1777
rect 5551 1675 5585 1709
rect 5551 1607 5585 1641
rect 5551 1539 5585 1573
rect 5551 1471 5585 1505
rect 5551 1411 5585 1437
rect 5349 1369 5375 1403
rect 5349 1335 5409 1369
rect 5349 1301 5375 1335
rect 5583 1403 5585 1411
rect 5549 1369 5551 1377
rect 5549 1339 5585 1369
rect 5583 1335 5585 1339
rect 5349 1285 5409 1301
rect 5551 1285 5585 1301
rect 5727 1811 5761 1827
rect 5727 1743 5761 1770
rect 5727 1702 5761 1709
rect 5727 1607 5761 1641
rect 5727 1539 5761 1573
rect 5727 1471 5761 1505
rect 5727 1403 5761 1437
rect 5727 1335 5761 1369
rect 5727 1285 5761 1301
rect 5903 1811 5937 1827
rect 5903 1743 5937 1777
rect 5903 1675 5937 1709
rect 5903 1607 5937 1641
rect 5903 1539 5937 1573
rect 5903 1471 5937 1475
rect 5903 1426 5937 1437
rect 5903 1335 5937 1369
rect 5903 1285 5937 1301
rect 5349 1284 5383 1285
rect 4708 1150 4742 1166
rect 4944 1150 4978 1166
rect 4708 1082 4742 1116
rect 5180 1150 5233 1166
rect 4978 1116 4982 1145
rect 4944 1111 4982 1116
rect 5214 1116 5233 1150
rect 5416 1150 5450 1166
rect 4944 1082 4978 1111
rect 4742 1035 4780 1069
rect 5180 1082 5233 1116
rect 5415 1116 5416 1145
rect 5652 1150 5686 1166
rect 5450 1116 5453 1145
rect 5415 1111 5453 1116
rect 4708 1014 4742 1035
rect 4708 964 4742 980
rect 4944 1014 4978 1048
rect 5178 1048 5180 1069
rect 5214 1069 5233 1082
rect 5416 1082 5450 1111
rect 5214 1048 5216 1069
rect 5178 1035 5216 1048
rect 5652 1082 5686 1116
rect 4944 964 4978 980
rect 5180 1014 5233 1035
rect 5214 980 5233 1014
rect 5180 964 5233 980
rect 5416 1014 5450 1048
rect 5614 1035 5652 1069
rect 5416 964 5450 980
rect 5652 1014 5686 1035
rect 5652 964 5686 980
rect 5184 961 5233 964
rect 4753 886 4769 920
rect 4803 886 4821 920
rect 4871 886 4894 920
rect 4939 886 4967 920
rect 5007 886 5040 920
rect 5075 886 5109 920
rect 5147 886 5177 920
rect 5220 886 5246 920
rect 5293 886 5315 920
rect 5367 886 5384 920
rect 5441 886 5453 920
rect 5515 886 5522 920
rect 5589 886 5591 920
rect 5625 886 5641 920
rect 5417 836 5604 840
rect 4708 820 4742 836
rect 4708 752 4742 786
rect 4944 820 4978 836
rect 4944 752 4978 786
rect 4708 684 4742 718
rect 4942 718 4944 732
rect 5180 820 5214 836
rect 5180 752 5214 786
rect 4978 718 4980 732
rect 4942 698 4980 718
rect 5416 820 5604 836
rect 5450 786 5604 820
rect 5416 752 5604 786
rect 4944 684 4978 698
rect 4742 622 4780 656
rect 5180 684 5214 718
rect 5413 718 5416 732
rect 5450 732 5604 752
rect 5450 718 5451 732
rect 5413 698 5451 718
rect 5485 698 5604 732
rect 4944 634 4978 650
rect 5179 650 5180 656
rect 5416 684 5604 698
rect 5214 650 5217 656
rect 5179 622 5217 650
rect 5450 650 5604 684
rect 5416 634 5604 650
rect 5417 493 5604 634
rect 4643 449 4677 473
rect 4643 387 4677 415
rect 4822 472 4856 477
rect 4822 393 4856 427
rect 4643 375 4718 387
rect 4677 353 4718 375
rect 4677 341 4752 353
rect 4643 309 4752 341
rect 4643 301 4718 309
rect 4677 275 4718 301
rect 4677 267 4752 275
rect 4643 231 4752 267
rect 4643 227 4718 231
rect 4677 197 4718 227
rect 4677 193 4752 197
rect 4643 153 4752 193
rect 4677 152 4752 153
rect 4677 119 4718 152
rect 4643 118 4718 119
rect 4643 79 4752 118
rect 4677 73 4752 79
rect 4677 45 4718 73
rect 4643 39 4718 45
rect 4643 5 4752 39
rect 4677 -6 4752 5
rect 4677 -29 4718 -6
rect 4643 -40 4718 -29
rect 4643 -69 4752 -40
rect 4822 325 4856 353
rect 4822 257 4856 268
rect 4822 217 4856 223
rect 4822 121 4856 155
rect 4822 53 4856 87
rect 4822 -15 4856 19
rect 4822 -65 4856 -49
rect 4998 461 5032 477
rect 4998 393 5032 427
rect 4998 329 5032 359
rect 4998 257 5032 291
rect 4998 189 5032 219
rect 4998 121 5032 143
rect 4998 53 5032 66
rect 4998 -15 5032 -11
rect 4998 -65 5032 -49
rect 5174 461 5208 477
rect 5174 399 5208 427
rect 5417 459 5561 493
rect 5595 459 5604 493
rect 5417 421 5604 459
rect 5417 408 5561 421
rect 5401 374 5417 408
rect 5451 374 5485 408
rect 5519 374 5553 408
rect 5595 387 5604 421
rect 5587 374 5604 387
rect 5782 700 6029 746
rect 5782 666 5911 700
rect 5945 666 5979 700
rect 6013 666 6029 700
rect 5782 615 5853 666
rect 5816 581 5853 615
rect 5782 551 5853 581
rect 5782 543 5819 551
rect 5816 517 5819 543
rect 5816 509 5853 517
rect 5782 483 5853 509
rect 5782 449 5819 483
rect 5782 415 5853 449
rect 5782 381 5819 415
rect 5174 327 5208 359
rect 5174 257 5208 291
rect 5174 189 5208 223
rect 5647 360 5681 363
rect 5647 241 5681 313
rect 5647 183 5681 199
rect 5782 246 5853 381
rect 5925 560 5959 598
rect 5925 483 5959 517
rect 5925 415 5959 449
rect 5925 365 5959 381
rect 6028 551 6065 567
rect 6028 517 6031 551
rect 6028 483 6065 517
rect 6028 449 6031 483
rect 6028 415 6065 449
rect 6028 381 6031 415
rect 6028 365 6065 381
rect 5782 212 5816 246
rect 5850 212 5853 246
rect 5782 178 5853 212
rect 5174 121 5208 155
rect 5401 138 5417 172
rect 5451 138 5471 172
rect 5519 138 5553 172
rect 5782 144 5816 178
rect 5850 144 5853 178
rect 5174 53 5208 87
rect 5782 110 5853 144
rect 5782 76 5816 110
rect 5850 76 5853 110
rect 5922 246 5956 262
rect 5922 178 5956 212
rect 5922 110 5956 144
rect 5782 58 5853 76
rect 5921 76 5922 89
rect 6028 246 6062 365
rect 6028 178 6062 212
rect 6028 110 6062 144
rect 5956 76 5959 89
rect 5921 55 5959 76
rect 5174 -15 5208 19
rect 5869 -20 5907 1
rect 5898 -33 5907 -20
rect 5174 -65 5208 -49
rect 4677 -85 4752 -69
rect 4677 -103 4718 -85
rect 4643 -119 4718 -103
rect 5864 -88 5898 -54
rect 6028 -76 6062 76
rect 4643 -127 4677 -119
rect 6037 -110 6075 -76
rect 6028 -111 6062 -110
rect 5864 -138 5898 -122
rect 5083 -175 5121 -163
rect 4853 -208 4856 -175
rect 4853 -209 4869 -208
rect 4903 -209 4937 -175
rect 4971 -209 4987 -175
rect 5043 -197 5049 -175
rect 5093 -197 5121 -175
rect 5043 -209 5059 -197
rect 5093 -209 5127 -197
rect 5161 -209 5177 -175
rect 4856 -246 4890 -209
rect 4846 -668 4862 -634
rect 4896 -645 4930 -634
rect 4909 -668 4930 -645
rect 4964 -668 4980 -634
rect 4875 -717 4909 -679
rect 4801 -791 4835 -786
rect 4801 -939 4835 -854
rect 4957 -752 4991 -736
rect 4957 -789 4958 -786
rect 4957 -820 4992 -789
rect 4991 -827 4992 -820
rect 4957 -861 4958 -854
rect 4957 -870 4991 -861
rect 4801 -983 4985 -939
rect 4801 -1017 4862 -983
rect 4896 -1017 4930 -983
rect 4964 -1017 4985 -983
rect 4801 -1023 4985 -1017
rect 4801 -1094 4835 -1085
rect 4801 -1166 4835 -1135
rect 4801 -1219 4835 -1203
rect 4957 -1091 4991 -1085
rect 4957 -1101 4958 -1091
rect 4991 -1135 4992 -1125
rect 4957 -1163 4992 -1135
rect 4957 -1169 4958 -1163
rect 4957 -1219 4991 -1203
<< viali >>
rect 4850 3143 4856 3172
rect 4856 3143 4884 3172
rect 4850 3138 4884 3143
rect 4922 3139 4956 3173
rect 4994 3139 5022 3173
rect 5022 3139 5028 3173
rect 4850 3071 4884 3097
rect 5232 3112 5266 3128
rect 5232 3094 5258 3112
rect 5258 3094 5266 3112
rect 4850 3063 4856 3071
rect 4856 3063 4884 3071
rect 5080 3053 5090 3087
rect 5090 3053 5114 3087
rect 5152 3053 5158 3087
rect 5158 3053 5186 3087
rect 4850 2988 4884 3022
rect 5232 3038 5266 3044
rect 5232 3010 5258 3038
rect 5258 3010 5266 3038
rect 4922 2967 4956 3001
rect 4994 2967 5022 3001
rect 5022 2967 5028 3001
rect 4850 2931 4856 2947
rect 4856 2931 4884 2947
rect 4850 2913 4884 2931
rect 5232 2930 5258 2959
rect 5258 2930 5266 2959
rect 5232 2925 5266 2930
rect 5080 2881 5090 2915
rect 5090 2881 5114 2915
rect 5152 2881 5158 2915
rect 5158 2881 5186 2915
rect 4850 2859 4884 2871
rect 4850 2837 4856 2859
rect 4856 2837 4884 2859
rect 5232 2856 5258 2874
rect 5258 2856 5266 2874
rect 5232 2840 5266 2856
rect 4922 2795 4956 2829
rect 4994 2795 5022 2829
rect 5022 2795 5028 2829
rect 4850 2761 4884 2795
rect 4850 2685 4884 2719
rect 5080 2709 5090 2743
rect 5090 2709 5114 2743
rect 5152 2709 5158 2743
rect 5158 2709 5186 2743
rect 5232 2694 5266 2726
rect 5232 2692 5258 2694
rect 5258 2692 5266 2694
rect 4850 2613 4856 2643
rect 4856 2613 4884 2643
rect 4922 2623 4956 2657
rect 4994 2623 5022 2657
rect 5022 2623 5028 2657
rect 4850 2609 4884 2613
rect 5232 2620 5266 2628
rect 5232 2594 5258 2620
rect 5258 2594 5266 2620
rect 4850 2541 4884 2567
rect 4850 2533 4856 2541
rect 4856 2533 4884 2541
rect 5080 2537 5090 2571
rect 5090 2537 5114 2571
rect 5152 2537 5158 2571
rect 5158 2537 5186 2571
rect 5232 2512 5258 2530
rect 5258 2512 5266 2530
rect 5232 2496 5266 2512
rect 4850 2457 4884 2491
rect 4922 2451 4956 2485
rect 4994 2451 5022 2485
rect 5022 2451 5028 2485
rect 4839 2297 4852 2331
rect 4852 2297 4873 2331
rect 4920 2297 4929 2331
rect 4929 2297 4954 2331
rect 5001 2297 5006 2331
rect 5006 2297 5035 2331
rect 5082 2297 5083 2331
rect 5083 2297 5116 2331
rect 5162 2297 5193 2331
rect 5193 2297 5196 2331
rect 5242 2297 5269 2331
rect 5269 2297 5276 2331
rect 5322 2297 5345 2331
rect 5345 2297 5356 2331
rect 4833 2170 4867 2203
rect 4833 2169 4867 2170
rect 4833 2102 4867 2131
rect 4833 2097 4867 2102
rect 5383 2202 5417 2236
rect 5383 2130 5417 2164
rect 5289 2014 5323 2042
rect 5289 2008 5323 2014
rect 5289 1946 5323 1970
rect 5289 1936 5323 1946
rect 5464 2014 5498 2042
rect 5464 2008 5498 2014
rect 5464 1946 5498 1970
rect 5464 1936 5498 1946
rect 5629 2014 5663 2042
rect 5629 2008 5663 2014
rect 5629 1946 5663 1970
rect 5629 1936 5663 1946
rect 5814 1980 5848 2012
rect 5814 1978 5848 1980
rect 5814 1906 5848 1940
rect 5089 1819 5123 1821
rect 4824 1785 4858 1788
rect 4824 1754 4833 1785
rect 4833 1754 4858 1785
rect 4896 1754 4930 1788
rect 5089 1787 5123 1819
rect 5089 1715 5123 1749
rect 4796 1580 4830 1603
rect 4957 1580 4991 1587
rect 5029 1580 5063 1587
rect 4796 1569 4823 1580
rect 4823 1569 4830 1580
rect 4957 1553 4979 1580
rect 4979 1553 4991 1580
rect 5029 1553 5047 1580
rect 5047 1553 5063 1580
rect 4796 1497 4830 1531
rect 4708 1480 4742 1497
rect 4708 1463 4742 1480
rect 4708 1412 4742 1425
rect 4708 1391 4742 1412
rect 5028 1480 5062 1502
rect 5028 1468 5060 1480
rect 5060 1468 5062 1480
rect 5100 1468 5134 1502
rect 4884 1378 4918 1411
rect 4884 1377 4918 1378
rect 4884 1310 4918 1339
rect 4884 1305 4918 1310
rect 5349 1811 5383 1821
rect 5349 1787 5375 1811
rect 5375 1787 5383 1811
rect 5349 1743 5383 1749
rect 5349 1715 5375 1743
rect 5375 1715 5383 1743
rect 5549 1403 5583 1411
rect 5549 1377 5551 1403
rect 5551 1377 5583 1403
rect 5549 1335 5583 1339
rect 5549 1305 5551 1335
rect 5551 1305 5583 1335
rect 5727 1777 5761 1804
rect 5727 1770 5761 1777
rect 5727 1675 5761 1702
rect 5727 1668 5761 1675
rect 5903 1505 5937 1509
rect 5903 1475 5937 1505
rect 5903 1403 5937 1426
rect 5903 1392 5937 1403
rect 4910 1111 4944 1145
rect 4982 1111 5016 1145
rect 4708 1048 4742 1069
rect 4708 1035 4742 1048
rect 4780 1035 4814 1069
rect 5381 1111 5415 1145
rect 5453 1111 5487 1145
rect 5144 1035 5178 1069
rect 5216 1035 5250 1069
rect 5580 1035 5614 1069
rect 5652 1048 5686 1069
rect 5652 1035 5686 1048
rect 4821 886 4837 920
rect 4837 886 4855 920
rect 4894 886 4905 920
rect 4905 886 4928 920
rect 4967 886 4973 920
rect 4973 886 5001 920
rect 5040 886 5041 920
rect 5041 886 5074 920
rect 5113 886 5143 920
rect 5143 886 5147 920
rect 5186 886 5211 920
rect 5211 886 5220 920
rect 5259 886 5280 920
rect 5280 886 5293 920
rect 5333 886 5349 920
rect 5349 886 5367 920
rect 5407 886 5418 920
rect 5418 886 5441 920
rect 5481 886 5487 920
rect 5487 886 5515 920
rect 5555 886 5556 920
rect 5556 886 5589 920
rect 4908 698 4942 732
rect 4980 698 5014 732
rect 4708 650 4742 656
rect 4708 622 4742 650
rect 4780 622 4814 656
rect 5379 698 5413 732
rect 5451 698 5485 732
rect 5145 622 5179 656
rect 5217 622 5251 656
rect 4822 461 4856 472
rect 4822 438 4856 461
rect 4718 353 4752 387
rect 4718 275 4752 309
rect 4718 197 4752 231
rect 4718 118 4752 152
rect 4718 39 4752 73
rect 4718 -40 4752 -6
rect 4822 359 4856 387
rect 4822 353 4856 359
rect 4822 291 4856 302
rect 4822 268 4856 291
rect 4822 189 4856 217
rect 4822 183 4856 189
rect 4998 325 5032 329
rect 4998 295 5032 325
rect 4998 223 5032 253
rect 4998 219 5032 223
rect 4998 155 5032 177
rect 4998 143 5032 155
rect 4998 87 5032 100
rect 4998 66 5032 87
rect 4998 19 5032 23
rect 4998 -11 5032 19
rect 5561 459 5595 493
rect 5561 408 5595 421
rect 5174 393 5208 399
rect 5174 365 5208 393
rect 5561 387 5587 408
rect 5587 387 5595 408
rect 5782 581 5816 615
rect 5782 509 5816 543
rect 5174 325 5208 327
rect 5174 293 5208 325
rect 5647 347 5681 360
rect 5647 326 5681 347
rect 5647 233 5681 241
rect 5647 207 5681 233
rect 5925 598 5959 632
rect 5925 551 5959 560
rect 5925 526 5959 551
rect 5471 138 5485 172
rect 5485 138 5505 172
rect 5571 138 5587 172
rect 5587 138 5605 172
rect 5887 55 5921 89
rect 5959 55 5993 89
rect 5835 -20 5869 1
rect 5835 -33 5864 -20
rect 5864 -33 5869 -20
rect 5907 -33 5941 1
rect 4718 -119 4752 -85
rect 6003 -110 6037 -76
rect 6075 -110 6109 -76
rect 4856 -175 4890 -174
rect 5049 -175 5083 -163
rect 5121 -175 5155 -163
rect 4856 -208 4869 -175
rect 4869 -208 4890 -175
rect 5049 -197 5059 -175
rect 5059 -197 5083 -175
rect 5121 -197 5127 -175
rect 5127 -197 5155 -175
rect 4856 -280 4890 -246
rect 4875 -668 4896 -645
rect 4896 -668 4909 -645
rect 4875 -679 4909 -668
rect 4801 -752 4835 -719
rect 4875 -751 4909 -717
rect 4801 -753 4835 -752
rect 4801 -820 4835 -791
rect 4801 -825 4835 -820
rect 4958 -786 4991 -755
rect 4991 -786 4992 -755
rect 4958 -789 4992 -786
rect 4958 -854 4991 -827
rect 4991 -854 4992 -827
rect 4958 -861 4992 -854
rect 4801 -1101 4835 -1094
rect 4801 -1128 4835 -1101
rect 4801 -1169 4835 -1166
rect 4801 -1200 4835 -1169
rect 4958 -1101 4992 -1091
rect 4958 -1125 4991 -1101
rect 4991 -1125 4992 -1101
rect 4958 -1169 4992 -1163
rect 4958 -1197 4991 -1169
rect 4991 -1197 4992 -1169
<< metal1 >>
tri 5068 3240 5163 3335 se
rect 5163 3329 5397 3335
rect 5163 3277 5345 3329
rect 5163 3265 5397 3277
rect 5163 3240 5345 3265
rect 5068 3213 5345 3240
rect 5068 3205 5397 3213
rect 5068 3184 5230 3205
tri 5230 3184 5251 3205 nw
rect 4809 3178 5040 3184
rect 4861 3172 4891 3178
rect 4943 3173 5040 3178
rect 4884 3138 4891 3172
rect 4956 3139 4994 3173
rect 5028 3139 5040 3173
rect 4861 3126 4891 3138
rect 4943 3126 5040 3139
rect 4809 3111 5040 3126
rect 4861 3097 4891 3111
rect 4884 3063 4891 3097
rect 4861 3059 4891 3063
rect 4943 3059 5040 3111
rect 4809 3044 5040 3059
rect 4861 3022 4891 3044
rect 4884 2992 4891 3022
rect 4943 3001 5040 3044
rect 4809 2988 4850 2992
rect 4884 2988 4922 2992
rect 4809 2977 4922 2988
rect 4861 2947 4891 2977
rect 4956 2967 4994 3001
rect 5028 2967 5040 3001
rect 4884 2925 4891 2947
rect 4943 2925 5040 2967
rect 4809 2913 4850 2925
rect 4884 2913 5040 2925
rect 4809 2910 5040 2913
rect 4861 2871 4891 2910
rect 4884 2858 4891 2871
rect 4943 2858 5040 2910
rect 5068 3087 5198 3184
tri 5198 3152 5230 3184 nw
rect 5068 3053 5080 3087
rect 5114 3053 5152 3087
rect 5186 3053 5198 3087
rect 5068 2915 5198 3053
rect 5068 2881 5080 2915
rect 5114 2881 5152 2915
rect 5186 2881 5198 2915
rect 5068 2875 5198 2881
rect 5226 3128 5272 3140
rect 5226 3094 5232 3128
rect 5266 3094 5272 3128
rect 5226 3074 5272 3094
tri 5272 3074 5338 3140 sw
rect 5226 3068 5434 3074
rect 5226 3044 5382 3068
rect 5226 3010 5232 3044
rect 5266 3016 5382 3044
rect 5266 3010 5434 3016
rect 5226 3004 5434 3010
rect 5226 2959 5382 3004
rect 5226 2925 5232 2959
rect 5266 2952 5382 2959
rect 5266 2946 5434 2952
rect 5266 2925 5272 2946
rect 4809 2843 4850 2858
rect 4884 2843 5040 2858
rect 4884 2837 4891 2843
rect 4861 2795 4891 2837
rect 4943 2829 5040 2843
rect 4956 2795 4994 2829
rect 5028 2795 5040 2829
rect 5226 2874 5272 2925
rect 5226 2840 5232 2874
rect 5266 2840 5272 2874
rect 5226 2828 5272 2840
tri 5272 2828 5390 2946 nw
rect 4884 2791 4891 2795
rect 4943 2791 5040 2795
rect 4809 2775 4850 2791
rect 4884 2775 5040 2791
rect 4884 2761 4891 2775
rect 4861 2723 4891 2761
rect 4943 2723 5040 2775
rect 4809 2719 5040 2723
rect 4809 2707 4850 2719
rect 4884 2707 5040 2719
rect 4884 2685 4891 2707
rect 4861 2655 4891 2685
rect 4943 2657 5040 2707
rect 4809 2643 4922 2655
rect 4809 2639 4850 2643
rect 4884 2639 4922 2643
rect 4884 2609 4891 2639
rect 4956 2623 4994 2657
rect 5028 2623 5040 2657
rect 4861 2587 4891 2609
rect 4943 2587 5040 2623
rect 4809 2571 5040 2587
rect 4861 2567 4891 2571
rect 4884 2533 4891 2567
rect 4861 2519 4891 2533
rect 4943 2519 5040 2571
rect 4809 2503 5040 2519
rect 4861 2491 4891 2503
rect 4884 2457 4891 2491
rect 4943 2485 5040 2503
rect 4861 2451 4891 2457
rect 4956 2451 4994 2485
rect 5028 2451 5040 2485
rect 4809 2445 5040 2451
rect 5068 2743 5198 2749
rect 5068 2709 5080 2743
rect 5114 2709 5152 2743
rect 5186 2709 5198 2743
rect 5068 2571 5198 2709
rect 5068 2537 5080 2571
rect 5114 2537 5152 2571
rect 5186 2537 5198 2571
rect 5068 2445 5198 2537
rect 5226 2726 5272 2738
rect 5226 2692 5232 2726
rect 5266 2692 5272 2726
rect 5226 2678 5272 2692
tri 5272 2678 5332 2738 sw
rect 5226 2672 5587 2678
rect 5226 2628 5535 2672
rect 5226 2594 5232 2628
rect 5266 2620 5535 2628
rect 5266 2608 5587 2620
rect 5266 2594 5535 2608
rect 5226 2556 5535 2594
rect 5226 2550 5587 2556
rect 5226 2530 5272 2550
rect 5226 2496 5232 2530
rect 5266 2496 5272 2530
rect 5226 2484 5272 2496
tri 5272 2484 5338 2550 nw
tri 5198 2445 5223 2470 sw
rect 5068 2443 5223 2445
tri 5223 2443 5225 2445 sw
rect 5068 2391 5507 2443
tri 5402 2379 5414 2391 ne
rect 5414 2379 5507 2391
tri 5414 2340 5453 2379 ne
rect 5453 2373 5507 2379
rect 5453 2340 5455 2373
rect 4809 2288 4815 2340
rect 4867 2331 4885 2340
rect 4937 2338 4943 2340
tri 4943 2338 4945 2340 sw
tri 5453 2338 5455 2340 ne
rect 4937 2337 4945 2338
tri 4945 2337 4946 2338 sw
rect 4937 2331 5368 2337
rect 4873 2297 4885 2331
rect 4954 2297 5001 2331
rect 5035 2297 5082 2331
rect 5116 2297 5162 2331
rect 5196 2297 5242 2331
rect 5276 2297 5322 2331
rect 5356 2297 5368 2331
rect 4867 2288 4885 2297
rect 4937 2291 5368 2297
rect 5455 2309 5507 2321
rect 4937 2288 4943 2291
tri 4943 2288 4946 2291 nw
rect 5455 2251 5507 2257
rect 5377 2236 5423 2248
rect 4809 2163 4815 2215
rect 4867 2163 4879 2215
rect 4931 2163 4937 2215
rect 4809 2135 4937 2163
rect 4809 2083 4815 2135
rect 4867 2083 4879 2135
rect 4931 2083 4937 2135
rect 5377 2202 5383 2236
rect 5417 2202 5423 2236
rect 5377 2164 5423 2202
rect 5377 2130 5383 2164
rect 5417 2130 5423 2164
rect 5283 2052 5329 2054
rect 5280 2046 5332 2052
rect 5280 1982 5332 1994
rect 5280 1924 5332 1930
rect 5377 1885 5423 2130
rect 5452 2048 5504 2054
rect 5452 1984 5504 1996
rect 5452 1926 5504 1932
rect 5458 1924 5504 1926
rect 5623 2042 5669 2054
rect 5623 2008 5629 2042
rect 5663 2008 5669 2042
rect 5623 1970 5669 2008
rect 5765 1974 5771 2026
rect 5823 2012 5835 2026
rect 5823 1974 5835 1978
rect 5887 1974 5893 2026
rect 5623 1936 5629 1970
rect 5663 1936 5669 1970
tri 5769 1940 5803 1974 ne
rect 5803 1940 5854 1974
rect 5623 1924 5669 1936
tri 5803 1935 5808 1940 ne
rect 5808 1906 5814 1940
rect 5848 1906 5854 1940
tri 5854 1939 5889 1974 nw
tri 5377 1883 5379 1885 ne
rect 5379 1883 5423 1885
tri 5423 1883 5445 1905 sw
rect 5808 1894 5854 1906
tri 5379 1839 5423 1883 ne
rect 5423 1839 5445 1883
tri 5423 1833 5429 1839 ne
rect 5429 1833 5445 1839
tri 5445 1833 5495 1883 sw
tri 5070 1821 5082 1833 se
rect 5082 1821 5389 1833
tri 5049 1800 5070 1821 se
rect 5070 1800 5089 1821
rect 4809 1748 4815 1800
rect 4867 1748 4884 1800
rect 4936 1748 4942 1800
tri 5043 1794 5049 1800 se
rect 5049 1794 5089 1800
tri 5036 1787 5043 1794 se
rect 5043 1787 5089 1794
rect 5123 1787 5349 1821
rect 5383 1787 5389 1821
tri 5429 1817 5445 1833 ne
rect 5445 1817 5495 1833
tri 5495 1817 5511 1833 sw
tri 5445 1804 5458 1817 ne
rect 5458 1804 5511 1817
tri 5511 1804 5524 1817 sw
rect 5718 1810 5770 1816
tri 5019 1770 5036 1787 se
rect 5036 1770 5389 1787
tri 5458 1770 5492 1804 ne
rect 5492 1770 5524 1804
tri 5524 1770 5558 1804 sw
tri 4998 1749 5019 1770 se
rect 5019 1749 5389 1770
tri 5492 1751 5511 1770 ne
rect 5511 1764 5558 1770
tri 5558 1764 5564 1770 sw
rect 5511 1758 5577 1764
rect 5511 1751 5525 1758
tri 4997 1748 4998 1749 se
rect 4998 1748 5089 1749
tri 4965 1716 4997 1748 se
rect 4997 1716 5089 1748
rect 4786 1715 5089 1716
rect 5123 1715 5349 1749
rect 5383 1715 5389 1749
tri 5511 1737 5525 1751 ne
rect 4786 1703 5389 1715
rect 4786 1702 5027 1703
tri 5027 1702 5028 1703 nw
rect 4786 1670 4995 1702
tri 4995 1670 5027 1702 nw
rect 5525 1694 5577 1706
rect 4786 1668 4889 1670
tri 4889 1668 4891 1670 nw
rect 4786 1643 4864 1668
tri 4864 1643 4889 1668 nw
rect 4786 1603 4838 1643
tri 4838 1617 4864 1643 nw
tri 5499 1617 5525 1643 se
rect 5718 1746 5770 1758
rect 5718 1668 5727 1694
rect 5761 1668 5770 1694
rect 5718 1656 5770 1668
rect 5525 1629 5577 1642
rect 5525 1617 5546 1629
rect 4786 1569 4796 1603
rect 4830 1569 4838 1603
tri 5480 1598 5499 1617 se
rect 5499 1598 5546 1617
tri 5546 1598 5577 1629 nw
rect 4786 1531 4838 1569
rect 4945 1587 5142 1598
rect 4945 1553 4957 1587
rect 4991 1553 5029 1587
rect 5063 1553 5142 1587
rect 4945 1546 5142 1553
rect 5194 1546 5206 1598
rect 5258 1546 5494 1598
tri 5494 1546 5546 1598 nw
rect 4702 1497 4754 1509
rect 4702 1476 4708 1497
rect 4742 1476 4754 1497
rect 4702 1412 4708 1424
rect 4742 1412 4754 1424
rect 4702 1354 4754 1360
rect 4786 1497 4796 1531
rect 4830 1497 4838 1531
rect 5894 1515 5946 1521
rect 4786 1245 4838 1497
rect 5016 1502 5057 1514
rect 5109 1502 5121 1514
rect 5016 1468 5028 1502
rect 5016 1462 5057 1468
rect 5109 1462 5121 1468
rect 5173 1462 5179 1514
tri 5619 1462 5623 1466 se
tri 5613 1456 5619 1462 se
rect 5619 1456 5623 1462
tri 5585 1428 5613 1456 se
rect 5613 1428 5623 1456
tri 5675 1428 5703 1456 sw
rect 5894 1438 5946 1463
rect 4878 1423 5022 1428
rect 4878 1422 5589 1423
rect 4930 1370 4970 1422
rect 5022 1411 5589 1422
rect 5022 1377 5549 1411
rect 5583 1377 5589 1411
rect 5894 1380 5946 1386
rect 5022 1370 5589 1377
rect 4878 1355 5589 1370
rect 4930 1303 4970 1355
rect 5022 1339 5589 1355
rect 5022 1305 5549 1339
rect 5583 1305 5589 1339
rect 5022 1303 5589 1305
rect 4878 1293 5589 1303
rect 4878 1288 5022 1293
rect 4930 1236 4970 1288
rect 4878 1230 5022 1236
rect 4786 1181 4838 1193
rect 4786 1123 4838 1129
rect 4886 1105 4892 1157
rect 4944 1105 4956 1157
rect 5008 1145 5499 1157
rect 5016 1111 5381 1145
rect 5415 1111 5453 1145
rect 5487 1111 5499 1145
rect 5008 1105 5499 1111
rect 4696 1069 5698 1075
rect 4696 1035 4708 1069
rect 4742 1035 4780 1069
rect 4814 1035 5144 1069
rect 5178 1035 5216 1069
rect 5250 1035 5580 1069
rect 5614 1035 5652 1069
rect 5686 1035 5698 1069
rect 4696 1029 5698 1035
rect 4809 920 5856 926
rect 4809 886 4821 920
rect 4855 886 4894 920
rect 4928 886 4967 920
rect 5001 886 5040 920
rect 5074 886 5113 920
rect 5147 886 5186 920
rect 5220 886 5259 920
rect 5293 886 5333 920
rect 5367 886 5407 920
rect 5441 886 5481 920
rect 5515 886 5555 920
rect 5589 919 5856 920
tri 5856 919 5863 926 sw
rect 5589 886 5863 919
rect 4809 880 5863 886
tri 5863 880 5902 919 sw
tri 5836 853 5863 880 ne
rect 5863 852 5902 880
tri 5902 852 5930 880 sw
rect 5772 814 5824 820
tri 5717 738 5772 793 se
rect 5772 750 5824 762
rect 4896 732 5772 738
rect 4896 698 4908 732
rect 4942 698 4980 732
rect 5014 698 5379 732
rect 5413 698 5451 732
rect 5485 698 5772 732
rect 4896 692 5824 698
tri 5523 662 5553 692 ne
rect 5553 662 5601 692
tri 5601 664 5629 692 nw
rect 4696 656 5511 662
tri 5553 660 5555 662 ne
rect 4696 622 4708 656
rect 4742 622 4780 656
rect 4814 622 5145 656
rect 5179 622 5217 656
rect 5251 622 5459 656
rect 4696 616 5459 622
tri 5401 615 5402 616 ne
rect 5402 615 5459 616
tri 5402 581 5436 615 ne
rect 5436 604 5459 615
rect 5436 592 5511 604
rect 5436 581 5459 592
tri 5436 571 5446 581 ne
rect 5446 571 5459 581
rect 4702 565 5108 571
rect 4754 560 5108 565
tri 5108 560 5119 571 sw
tri 5446 560 5457 571 ne
rect 5457 560 5459 571
rect 4754 558 5119 560
tri 5119 558 5121 560 sw
tri 5457 558 5459 560 ne
rect 4754 543 5121 558
tri 5121 543 5136 558 sw
rect 4754 539 5136 543
tri 5136 539 5140 543 sw
rect 4754 519 5140 539
rect 4754 513 4785 519
rect 4702 509 4785 513
tri 4785 509 4795 519 nw
tri 5086 509 5096 519 ne
rect 5096 509 5140 519
tri 5140 509 5170 539 sw
rect 5305 529 5357 535
rect 4702 501 4769 509
rect 4754 493 4769 501
tri 4769 493 4785 509 nw
tri 5096 493 5112 509 ne
rect 5112 497 5170 509
tri 5170 497 5182 509 sw
rect 5112 493 5182 497
tri 5182 493 5186 497 sw
rect 4754 484 4760 493
tri 4760 484 4769 493 nw
tri 5112 484 5121 493 ne
rect 5121 484 5186 493
tri 5186 484 5195 493 sw
tri 4754 478 4760 484 nw
rect 4816 478 4952 484
rect 4702 443 4754 449
rect 4816 472 4900 478
rect 4816 438 4822 472
rect 4856 438 4900 472
rect 4816 426 4900 438
tri 5121 465 5140 484 ne
rect 5140 465 5195 484
tri 5195 465 5214 484 sw
tri 5140 459 5146 465 ne
rect 5146 459 5214 465
tri 5146 437 5168 459 ne
rect 4816 414 4952 426
rect 4712 387 4758 399
rect 4712 353 4718 387
rect 4752 353 4758 387
rect 4712 309 4758 353
rect 4712 275 4718 309
rect 4752 275 4758 309
rect 4712 231 4758 275
rect 4712 197 4718 231
rect 4752 197 4758 231
rect 4712 152 4758 197
rect 4816 387 4900 414
rect 4816 353 4822 387
rect 4856 362 4900 387
rect 4856 356 4952 362
rect 5168 399 5214 459
rect 5168 365 5174 399
rect 5208 365 5214 399
rect 4856 353 4895 356
rect 4816 329 4895 353
tri 4895 329 4922 356 nw
rect 4992 329 5038 341
rect 4816 302 4862 329
rect 4816 268 4822 302
rect 4856 268 4862 302
tri 4862 296 4895 329 nw
rect 4816 217 4862 268
rect 4992 295 4998 329
rect 5032 295 5038 329
rect 4992 281 5038 295
rect 5168 327 5214 365
rect 5168 293 5174 327
rect 5208 293 5214 327
tri 5038 281 5046 289 sw
rect 5168 281 5214 293
rect 5305 465 5357 477
rect 4992 255 5046 281
tri 5046 255 5072 281 sw
rect 4816 183 4822 217
rect 4856 183 4862 217
rect 4816 171 4862 183
rect 4894 249 4946 255
rect 4894 185 4946 197
rect 4712 118 4718 152
rect 4752 118 4758 152
rect 4712 73 4758 118
rect 4712 39 4718 73
rect 4752 39 4758 73
rect 4712 -6 4758 39
rect 4712 -40 4718 -6
rect 4752 -40 4758 -6
rect 4712 -85 4758 -40
tri 4893 -76 4894 -75 se
rect 4894 -76 4946 133
rect 4992 253 5072 255
rect 4992 219 4998 253
rect 5032 241 5072 253
tri 5072 241 5086 255 sw
rect 5032 219 5086 241
rect 4992 207 5086 219
tri 5086 207 5120 241 sw
rect 4992 66 4998 207
rect 5114 91 5120 207
rect 5305 151 5357 413
rect 5459 235 5511 540
rect 5555 493 5601 662
rect 5863 662 5930 852
tri 5930 662 5943 675 sw
rect 5863 644 5943 662
tri 5943 644 5961 662 sw
rect 5863 632 6166 644
rect 5774 621 5826 627
rect 5774 555 5826 569
rect 5774 497 5826 503
rect 5863 598 5925 632
rect 5959 598 6166 632
rect 5863 560 6166 598
rect 5863 526 5925 560
rect 5959 526 6166 560
rect 5863 514 6166 526
rect 5863 497 5937 514
tri 5937 497 5954 514 nw
rect 5555 459 5561 493
rect 5595 459 5601 493
rect 5555 421 5601 459
rect 5555 387 5561 421
rect 5595 387 5601 421
rect 5555 375 5601 387
tri 5797 381 5863 447 se
rect 5863 427 5909 497
tri 5909 469 5937 497 nw
tri 5863 381 5909 427 nw
tri 5791 375 5797 381 se
rect 5797 375 5854 381
tri 5788 372 5791 375 se
rect 5791 372 5854 375
tri 5854 372 5863 381 nw
rect 5641 360 5752 372
rect 5641 326 5647 360
rect 5681 326 5752 360
rect 5641 270 5752 326
tri 5752 270 5854 372 nw
rect 5641 241 5687 270
tri 5511 235 5515 239 sw
rect 5459 207 5515 235
tri 5515 207 5543 235 sw
rect 5641 207 5647 241
rect 5681 207 5687 241
tri 5687 235 5722 270 nw
rect 5459 178 5543 207
tri 5543 178 5572 207 sw
rect 5641 195 5687 207
rect 5459 172 5617 178
tri 5305 141 5315 151 ne
rect 5315 141 5357 151
tri 5357 141 5381 165 sw
tri 5315 138 5318 141 ne
rect 5318 138 5381 141
tri 5381 138 5384 141 sw
rect 5459 138 5471 172
rect 5505 138 5571 172
rect 5605 138 5617 172
tri 5318 99 5357 138 ne
rect 5357 99 5384 138
rect 5032 89 5118 91
tri 5118 89 5120 91 nw
tri 5357 89 5367 99 ne
rect 5367 95 5384 99
tri 5384 95 5427 138 sw
rect 5459 132 5617 138
rect 5367 89 5427 95
tri 5427 89 5433 95 sw
rect 5874 89 6052 95
rect 5032 75 5104 89
tri 5104 75 5118 89 nw
tri 5367 75 5381 89 ne
rect 5381 75 5433 89
tri 5433 75 5447 89 sw
rect 5032 66 5091 75
rect 4992 62 5091 66
tri 5091 62 5104 75 nw
tri 5381 62 5394 75 ne
rect 5394 62 5658 75
tri 5658 62 5671 75 sw
rect 4992 55 5084 62
tri 5084 55 5091 62 nw
tri 5394 55 5401 62 ne
rect 5401 55 5671 62
tri 5671 55 5678 62 sw
rect 5874 55 5887 89
rect 5921 55 5959 89
rect 5993 55 6052 89
rect 4992 29 5058 55
tri 5058 29 5084 55 nw
tri 5401 29 5427 55 ne
rect 5427 43 5678 55
tri 5678 43 5690 55 sw
rect 5874 43 6052 55
rect 5427 29 5690 43
rect 4992 23 5038 29
rect 4992 -11 4998 23
rect 5032 -11 5038 23
tri 5038 9 5058 29 nw
tri 5638 9 5658 29 ne
rect 5658 9 5690 29
tri 5658 1 5666 9 ne
rect 5666 7 5690 9
tri 5690 7 5726 43 sw
rect 5666 1 5726 7
tri 5726 1 5732 7 sw
rect 5823 1 5953 7
tri 5666 -4 5671 1 ne
rect 5671 -4 5732 1
tri 5732 -4 5737 1 sw
rect 4992 -23 5038 -11
tri 5671 -23 5690 -4 ne
rect 5690 -23 5737 -4
tri 5690 -33 5700 -23 ne
rect 5700 -33 5737 -23
tri 5737 -33 5766 -4 sw
rect 5823 -33 5835 1
rect 5869 -33 5907 1
rect 5941 -33 5953 1
tri 5700 -70 5737 -33 ne
rect 5737 -39 5766 -33
tri 5766 -39 5772 -33 sw
rect 5823 -39 5953 -33
rect 5737 -70 5772 -39
tri 5772 -70 5803 -39 sw
tri 5737 -76 5743 -70 ne
rect 5743 -76 6121 -70
rect 4712 -119 4718 -85
rect 4752 -119 4758 -85
tri 4880 -89 4893 -76 se
rect 4893 -89 4946 -76
tri 4859 -110 4880 -89 se
rect 4880 -110 4925 -89
tri 4925 -110 4946 -89 nw
tri 5743 -110 5777 -76 ne
rect 5777 -110 6003 -76
rect 6037 -110 6075 -76
rect 6109 -110 6121 -76
rect 4712 -817 4758 -119
tri 4850 -119 4859 -110 se
rect 4859 -119 4896 -110
rect 4850 -174 4896 -119
tri 4896 -139 4925 -110 nw
tri 5777 -116 5783 -110 ne
rect 5783 -116 6121 -110
rect 4978 -122 5030 -116
rect 4850 -208 4856 -174
rect 4890 -208 4896 -174
rect 4850 -246 4896 -208
tri 5030 -157 5071 -116 sw
rect 5030 -163 5167 -157
rect 5030 -174 5049 -163
rect 4978 -186 5049 -174
tri 4943 -244 4978 -209 se
rect 5030 -197 5049 -186
rect 5083 -197 5121 -163
rect 5155 -197 5167 -163
rect 5030 -203 5167 -197
rect 5030 -238 5037 -203
rect 4978 -244 5037 -238
tri 5037 -244 5078 -203 nw
rect 4850 -280 4856 -246
rect 4890 -280 4896 -246
tri 4830 -463 4850 -443 se
rect 4850 -463 4896 -280
tri 4795 -498 4830 -463 se
rect 4830 -498 4854 -463
rect 4795 -505 4854 -498
tri 4854 -505 4896 -463 nw
tri 4938 -249 4943 -244 se
rect 4943 -249 4989 -244
rect 4938 -292 4989 -249
tri 4989 -292 5037 -244 nw
rect 4795 -719 4841 -505
tri 4841 -518 4854 -505 nw
tri 4925 -518 4938 -505 se
rect 4938 -518 4984 -292
tri 4984 -297 4989 -292 nw
tri 4922 -521 4925 -518 se
rect 4925 -521 4984 -518
tri 4915 -528 4922 -521 se
rect 4922 -528 4977 -521
tri 4977 -528 4984 -521 nw
tri 4892 -551 4915 -528 se
rect 4915 -551 4954 -528
tri 4954 -551 4977 -528 nw
rect 4795 -753 4801 -719
rect 4835 -753 4841 -719
rect 4795 -791 4841 -753
tri 4758 -817 4764 -811 sw
rect 4712 -823 4764 -817
rect 4795 -825 4801 -791
rect 4835 -825 4841 -791
rect 4795 -837 4841 -825
tri 4869 -574 4892 -551 se
rect 4892 -574 4915 -551
rect 4869 -645 4915 -574
tri 4915 -590 4954 -551 nw
rect 4869 -679 4875 -645
rect 4909 -679 4915 -645
rect 4869 -717 4915 -679
rect 4869 -751 4875 -717
rect 4909 -751 4915 -717
rect 4712 -887 4764 -875
rect 4712 -945 4764 -939
tri 4863 -945 4869 -939 se
rect 4869 -945 4915 -751
tri 4849 -959 4863 -945 se
rect 4863 -959 4915 -945
tri 4841 -967 4849 -959 se
rect 4849 -967 4907 -959
tri 4907 -967 4915 -959 nw
rect 4952 -755 4998 -743
rect 4952 -789 4958 -755
rect 4992 -789 4998 -755
rect 4952 -827 4998 -789
rect 4952 -861 4958 -827
rect 4992 -861 4998 -827
rect 4952 -967 4998 -861
tri 4998 -967 4999 -966 sw
tri 4795 -1013 4841 -967 se
rect 4795 -1094 4841 -1013
tri 4841 -1033 4907 -967 nw
rect 4952 -1033 4999 -967
tri 4999 -1033 5065 -967 sw
rect 4795 -1128 4801 -1094
rect 4835 -1128 4841 -1094
rect 4795 -1166 4841 -1128
rect 4795 -1200 4801 -1166
rect 4835 -1200 4841 -1166
rect 4795 -1212 4841 -1200
rect 4952 -1069 5065 -1033
tri 5065 -1069 5101 -1033 sw
rect 4952 -1070 5191 -1069
rect 4952 -1076 5260 -1070
rect 4952 -1091 5134 -1076
rect 4952 -1125 4958 -1091
rect 4992 -1125 5134 -1091
rect 4952 -1128 5134 -1125
rect 5186 -1128 5208 -1076
rect 4952 -1142 5260 -1128
rect 4952 -1163 5134 -1142
rect 4952 -1197 4958 -1163
rect 4992 -1194 5134 -1163
rect 5186 -1194 5208 -1142
rect 4992 -1197 5260 -1194
rect 4952 -1208 5260 -1197
rect 4952 -1214 5134 -1208
rect 4952 -1266 4970 -1214
rect 5022 -1266 5034 -1214
rect 5086 -1260 5134 -1214
rect 5186 -1260 5208 -1208
rect 5086 -1266 5260 -1260
rect 4952 -1272 5158 -1266
<< via1 >>
rect 5345 3277 5397 3329
rect 5345 3213 5397 3265
rect 4809 3172 4861 3178
rect 4891 3173 4943 3178
rect 4809 3138 4850 3172
rect 4850 3138 4861 3172
rect 4891 3139 4922 3173
rect 4922 3139 4943 3173
rect 4809 3126 4861 3138
rect 4891 3126 4943 3139
rect 4809 3097 4861 3111
rect 4809 3063 4850 3097
rect 4850 3063 4861 3097
rect 4809 3059 4861 3063
rect 4891 3059 4943 3111
rect 4809 3022 4861 3044
rect 4809 2992 4850 3022
rect 4850 2992 4861 3022
rect 4891 3001 4943 3044
rect 4891 2992 4922 3001
rect 4922 2992 4943 3001
rect 4809 2947 4861 2977
rect 4891 2967 4922 2977
rect 4922 2967 4943 2977
rect 4809 2925 4850 2947
rect 4850 2925 4861 2947
rect 4891 2925 4943 2967
rect 4809 2871 4861 2910
rect 4809 2858 4850 2871
rect 4850 2858 4861 2871
rect 4891 2858 4943 2910
rect 5382 3016 5434 3068
rect 5382 2952 5434 3004
rect 4809 2837 4850 2843
rect 4850 2837 4861 2843
rect 4809 2795 4861 2837
rect 4891 2829 4943 2843
rect 4891 2795 4922 2829
rect 4922 2795 4943 2829
rect 4809 2791 4850 2795
rect 4850 2791 4861 2795
rect 4891 2791 4943 2795
rect 4809 2761 4850 2775
rect 4850 2761 4861 2775
rect 4809 2723 4861 2761
rect 4891 2723 4943 2775
rect 4809 2685 4850 2707
rect 4850 2685 4861 2707
rect 4809 2655 4861 2685
rect 4891 2657 4943 2707
rect 4891 2655 4922 2657
rect 4922 2655 4943 2657
rect 4809 2609 4850 2639
rect 4850 2609 4861 2639
rect 4891 2623 4922 2639
rect 4922 2623 4943 2639
rect 4809 2587 4861 2609
rect 4891 2587 4943 2623
rect 4809 2567 4861 2571
rect 4809 2533 4850 2567
rect 4850 2533 4861 2567
rect 4809 2519 4861 2533
rect 4891 2519 4943 2571
rect 4809 2491 4861 2503
rect 4809 2457 4850 2491
rect 4850 2457 4861 2491
rect 4891 2485 4943 2503
rect 4809 2451 4861 2457
rect 4891 2451 4922 2485
rect 4922 2451 4943 2485
rect 5535 2620 5587 2672
rect 5535 2556 5587 2608
rect 4815 2331 4867 2340
rect 4885 2331 4937 2340
rect 4815 2297 4839 2331
rect 4839 2297 4867 2331
rect 4885 2297 4920 2331
rect 4920 2297 4937 2331
rect 4815 2288 4867 2297
rect 4885 2288 4937 2297
rect 5455 2321 5507 2373
rect 5455 2257 5507 2309
rect 4815 2203 4867 2215
rect 4815 2169 4833 2203
rect 4833 2169 4867 2203
rect 4815 2163 4867 2169
rect 4879 2163 4931 2215
rect 4815 2131 4867 2135
rect 4815 2097 4833 2131
rect 4833 2097 4867 2131
rect 4815 2083 4867 2097
rect 4879 2083 4931 2135
rect 5280 2042 5332 2046
rect 5280 2008 5289 2042
rect 5289 2008 5323 2042
rect 5323 2008 5332 2042
rect 5280 1994 5332 2008
rect 5280 1970 5332 1982
rect 5280 1936 5289 1970
rect 5289 1936 5323 1970
rect 5323 1936 5332 1970
rect 5280 1930 5332 1936
rect 5452 2042 5504 2048
rect 5452 2008 5464 2042
rect 5464 2008 5498 2042
rect 5498 2008 5504 2042
rect 5452 1996 5504 2008
rect 5452 1970 5504 1984
rect 5452 1936 5464 1970
rect 5464 1936 5498 1970
rect 5498 1936 5504 1970
rect 5452 1932 5504 1936
rect 5771 2012 5823 2026
rect 5835 2012 5887 2026
rect 5771 1978 5814 2012
rect 5814 1978 5823 2012
rect 5835 1978 5848 2012
rect 5848 1978 5887 2012
rect 5771 1974 5823 1978
rect 5835 1974 5887 1978
rect 4815 1788 4867 1800
rect 4815 1754 4824 1788
rect 4824 1754 4858 1788
rect 4858 1754 4867 1788
rect 4815 1748 4867 1754
rect 4884 1788 4936 1800
rect 4884 1754 4896 1788
rect 4896 1754 4930 1788
rect 4930 1754 4936 1788
rect 4884 1748 4936 1754
rect 5718 1804 5770 1810
rect 5718 1770 5727 1804
rect 5727 1770 5761 1804
rect 5761 1770 5770 1804
rect 5525 1706 5577 1758
rect 5525 1642 5577 1694
rect 5718 1758 5770 1770
rect 5718 1702 5770 1746
rect 5718 1694 5727 1702
rect 5727 1694 5761 1702
rect 5761 1694 5770 1702
rect 5142 1546 5194 1598
rect 5206 1546 5258 1598
rect 4702 1463 4708 1476
rect 4708 1463 4742 1476
rect 4742 1463 4754 1476
rect 4702 1425 4754 1463
rect 4702 1424 4708 1425
rect 4708 1424 4742 1425
rect 4742 1424 4754 1425
rect 4702 1391 4708 1412
rect 4708 1391 4742 1412
rect 4742 1391 4754 1412
rect 4702 1360 4754 1391
rect 5057 1502 5109 1514
rect 5121 1502 5173 1514
rect 5057 1468 5062 1502
rect 5062 1468 5100 1502
rect 5100 1468 5109 1502
rect 5121 1468 5134 1502
rect 5134 1468 5173 1502
rect 5057 1462 5109 1468
rect 5121 1462 5173 1468
rect 5894 1509 5946 1515
rect 5894 1475 5903 1509
rect 5903 1475 5937 1509
rect 5937 1475 5946 1509
rect 5894 1463 5946 1475
rect 4786 1193 4838 1245
rect 5894 1426 5946 1438
rect 4878 1411 4930 1422
rect 4878 1377 4884 1411
rect 4884 1377 4918 1411
rect 4918 1377 4930 1411
rect 4878 1370 4930 1377
rect 4970 1370 5022 1422
rect 5894 1392 5903 1426
rect 5903 1392 5937 1426
rect 5937 1392 5946 1426
rect 5894 1386 5946 1392
rect 4878 1339 4930 1355
rect 4878 1305 4884 1339
rect 4884 1305 4918 1339
rect 4918 1305 4930 1339
rect 4878 1303 4930 1305
rect 4970 1303 5022 1355
rect 4878 1236 4930 1288
rect 4970 1236 5022 1288
rect 4786 1129 4838 1181
rect 4892 1145 4944 1157
rect 4892 1111 4910 1145
rect 4910 1111 4944 1145
rect 4892 1105 4944 1111
rect 4956 1145 5008 1157
rect 4956 1111 4982 1145
rect 4982 1111 5008 1145
rect 4956 1105 5008 1111
rect 5772 762 5824 814
rect 5772 698 5824 750
rect 5459 604 5511 656
rect 4702 513 4754 565
rect 5459 540 5511 592
rect 4702 449 4754 501
rect 4900 426 4952 478
rect 4900 362 4952 414
rect 5305 477 5357 529
rect 5305 413 5357 465
rect 4894 197 4946 249
rect 4894 133 4946 185
rect 4998 177 5114 207
rect 4998 143 5032 177
rect 5032 143 5114 177
rect 4998 100 5114 143
rect 4998 91 5032 100
rect 5032 91 5114 100
rect 5774 615 5826 621
rect 5774 581 5782 615
rect 5782 581 5816 615
rect 5816 581 5826 615
rect 5774 569 5826 581
rect 5774 543 5826 555
rect 5774 509 5782 543
rect 5782 509 5816 543
rect 5816 509 5826 543
rect 5774 503 5826 509
rect 4978 -174 5030 -122
rect 4978 -238 5030 -186
rect 4712 -875 4764 -823
rect 4712 -939 4764 -887
rect 5134 -1128 5186 -1076
rect 5208 -1128 5260 -1076
rect 5134 -1194 5186 -1142
rect 5208 -1194 5260 -1142
rect 4970 -1266 5022 -1214
rect 5034 -1266 5086 -1214
rect 5134 -1260 5186 -1208
rect 5208 -1260 5260 -1208
<< metal2 >>
rect 5341 3344 5397 3353
rect 5341 3277 5345 3288
rect 5341 3265 5397 3277
rect 5341 3264 5345 3265
rect 5341 3199 5397 3208
rect 4809 3178 4943 3184
rect 4861 3126 4891 3178
rect 4809 3111 4943 3126
rect 4861 3059 4891 3111
rect 4809 3044 4943 3059
rect 4861 2992 4891 3044
rect 4809 2977 4943 2992
rect 4861 2925 4891 2977
rect 5378 3083 5434 3092
rect 5378 3016 5382 3027
rect 5378 3004 5434 3016
rect 5378 3003 5382 3004
rect 5378 2938 5434 2947
rect 4809 2910 4943 2925
rect 4861 2858 4891 2910
rect 4809 2843 4943 2858
rect 4861 2791 4891 2843
rect 4809 2775 4943 2791
rect 4861 2723 4891 2775
rect 4809 2707 4943 2723
rect 4861 2655 4891 2707
rect 4809 2639 4943 2655
rect 4861 2587 4891 2639
rect 4809 2571 4943 2587
rect 4861 2519 4891 2571
rect 5535 2672 5721 2678
rect 5587 2669 5721 2672
rect 5587 2620 5665 2669
rect 5535 2613 5665 2620
rect 5535 2608 5721 2613
rect 5587 2589 5721 2608
rect 5587 2556 5665 2589
rect 5535 2533 5665 2556
rect 5535 2524 5721 2533
rect 4809 2503 4943 2519
rect 4861 2451 4891 2503
rect 4809 2340 4943 2451
rect 4809 2288 4815 2340
rect 4867 2288 4885 2340
rect 4937 2288 4943 2340
rect 4809 2215 4943 2288
rect 5455 2383 5511 2392
rect 5507 2321 5511 2327
rect 5455 2309 5511 2321
rect 5507 2303 5511 2309
rect 5455 2238 5511 2247
rect 4809 2163 4815 2215
rect 4867 2163 4879 2215
rect 4931 2163 4943 2215
rect 4809 2135 4943 2163
rect 4809 2083 4815 2135
rect 4867 2083 4879 2135
rect 4931 2083 4943 2135
rect 4809 1800 4943 2083
rect 5280 2046 5332 2052
rect 5280 1982 5332 1994
rect 5280 1924 5332 1930
rect 5452 2048 5504 2054
rect 5452 1984 5504 1996
rect 5765 1974 5771 2026
rect 5823 1974 5835 2026
rect 5887 1974 5893 2026
rect 5452 1926 5504 1932
tri 5712 1810 5718 1816 se
rect 5718 1810 5770 1816
rect 4809 1748 4815 1800
rect 4867 1748 4884 1800
rect 4936 1748 4943 1800
tri 5676 1774 5712 1810 se
rect 5712 1774 5718 1810
rect 4809 1694 4943 1748
rect 5525 1758 5718 1774
rect 5577 1746 5770 1758
rect 5577 1722 5718 1746
rect 5577 1706 5587 1722
tri 4943 1694 4949 1700 sw
rect 5525 1694 5587 1706
tri 5587 1694 5615 1722 nw
tri 5684 1694 5712 1722 ne
rect 5712 1694 5718 1722
rect 4809 1644 4949 1694
tri 4809 1642 4811 1644 ne
rect 4811 1642 4949 1644
tri 4949 1642 5001 1694 sw
rect 5577 1688 5581 1694
tri 5581 1688 5587 1694 nw
tri 5712 1688 5718 1694 ne
rect 5718 1688 5770 1694
tri 5577 1684 5581 1688 nw
tri 4811 1621 4832 1642 ne
rect 4832 1621 5001 1642
tri 5001 1621 5022 1642 sw
rect 5525 1636 5577 1642
tri 4832 1598 4855 1621 ne
rect 4855 1598 5022 1621
tri 4855 1575 4878 1598 ne
rect 4702 1476 4754 1482
rect 4702 1412 4754 1424
rect 4702 565 4754 1360
rect 4878 1422 5022 1598
rect 5136 1546 5142 1598
rect 5194 1546 5206 1598
rect 5258 1546 5264 1598
tri 5187 1521 5212 1546 ne
rect 5051 1462 5057 1514
rect 5109 1462 5121 1514
rect 5173 1462 5179 1514
tri 5051 1453 5060 1462 ne
rect 5060 1453 5131 1462
tri 5131 1453 5140 1462 nw
rect 4930 1370 4970 1422
rect 4878 1355 5022 1370
rect 4930 1303 4970 1355
rect 4878 1288 5022 1303
rect 4786 1245 4838 1251
rect 4930 1236 4970 1288
rect 4878 1230 5022 1236
rect 5060 1438 5116 1453
tri 5116 1438 5131 1453 nw
rect 4786 1181 4838 1193
tri 4917 1157 4929 1169 se
rect 4929 1160 4985 1169
tri 4985 1157 4997 1169 sw
tri 4838 1141 4851 1154 sw
rect 4838 1129 4851 1141
rect 4786 1123 4851 1129
tri 4786 1110 4799 1123 ne
rect 4702 501 4754 513
rect 4702 24 4754 449
rect 4799 91 4851 1123
rect 4886 1105 4892 1157
rect 5008 1105 5014 1157
tri 4886 1062 4929 1105 ne
rect 4929 1080 4985 1104
tri 4985 1076 5014 1105 nw
rect 4929 1015 4985 1024
tri 4984 849 5060 925 se
rect 5060 849 5112 1438
tri 5112 1434 5116 1438 nw
rect 4984 808 5112 849
tri 5187 814 5212 839 se
rect 5212 817 5264 1546
rect 5894 1515 5946 1521
rect 5894 1438 5946 1463
tri 5820 1199 5894 1273 se
rect 5894 1251 5946 1386
tri 5894 1199 5946 1251 nw
rect 5212 814 5261 817
tri 5261 814 5264 817 nw
tri 5772 1151 5820 1199 se
rect 5820 1151 5846 1199
tri 5846 1151 5894 1199 nw
rect 5772 814 5824 1151
tri 5824 1129 5846 1151 nw
rect 4984 765 5069 808
tri 5069 765 5112 808 nw
tri 5138 765 5187 814 se
rect 5187 765 5212 814
tri 5212 765 5261 814 nw
rect 4984 762 5066 765
tri 5066 762 5069 765 nw
tri 5135 762 5138 765 se
rect 5138 762 5209 765
tri 5209 762 5212 765 nw
rect 4984 754 5058 762
tri 5058 754 5066 762 nw
tri 5127 754 5135 762 se
rect 5135 754 5197 762
tri 4980 750 4984 754 se
rect 4984 750 5054 754
tri 5054 750 5058 754 nw
tri 5123 750 5127 754 se
rect 5127 750 5197 754
tri 5197 750 5209 762 nw
rect 5772 750 5824 762
tri 4928 698 4980 750 se
rect 4980 739 5043 750
tri 5043 739 5054 750 nw
tri 5112 739 5123 750 se
rect 5123 739 5145 750
rect 4980 698 5002 739
tri 5002 698 5043 739 nw
tri 5071 698 5112 739 se
rect 5112 698 5145 739
tri 5145 698 5197 750 nw
tri 4921 691 4928 698 se
rect 4928 691 4995 698
tri 4995 691 5002 698 nw
tri 5064 691 5071 698 se
rect 5071 691 5138 698
tri 5138 691 5145 698 nw
rect 5772 692 5824 698
tri 4910 680 4921 691 se
rect 4921 680 4984 691
tri 4984 680 4995 691 nw
tri 5055 682 5064 691 se
rect 5064 682 5129 691
tri 5129 682 5138 691 nw
rect 5055 680 5127 682
tri 5127 680 5129 682 nw
tri 4900 670 4910 680 se
rect 4910 670 4974 680
tri 4974 670 4984 680 nw
rect 4900 656 4960 670
tri 4960 656 4974 670 nw
rect 4900 478 4952 656
tri 4952 648 4960 656 nw
rect 4900 414 4952 426
rect 4900 356 4952 362
tri 5018 356 5055 393 se
rect 5055 371 5107 680
tri 5107 660 5127 680 nw
rect 5455 672 5511 681
rect 5455 604 5459 616
rect 5455 592 5511 604
rect 5303 549 5359 558
rect 5455 527 5511 536
rect 5770 638 5826 647
rect 5770 569 5774 582
rect 5770 558 5826 569
rect 5770 493 5826 502
rect 5303 477 5305 493
rect 5357 477 5359 493
rect 5303 469 5359 477
rect 5303 404 5359 413
tri 4981 319 5018 356 se
rect 5018 319 5055 356
tri 5055 319 5107 371 nw
tri 4917 255 4981 319 se
rect 4981 255 4986 319
rect 4894 250 4986 255
tri 4986 250 5055 319 nw
rect 4894 249 4946 250
tri 4946 210 4986 250 nw
rect 4894 185 4946 197
rect 4894 127 4946 133
tri 4851 91 4858 98 sw
rect 4992 91 4998 207
rect 5114 91 5120 207
tri 5120 91 5125 96 sw
rect 4799 84 4858 91
tri 4799 51 4832 84 ne
rect 4832 51 4858 84
tri 4858 51 4898 91 sw
rect 4992 83 5125 91
tri 5125 83 5133 91 sw
rect 4992 51 5133 83
tri 5133 51 5165 83 sw
tri 4832 46 4837 51 ne
rect 4837 46 4898 51
tri 4898 46 4903 51 sw
rect 4992 46 5165 51
tri 5165 46 5170 51 sw
tri 4702 20 4706 24 ne
rect 4706 20 4754 24
tri 4754 20 4780 46 sw
tri 4837 32 4851 46 ne
rect 4851 32 4903 46
tri 4851 20 4863 32 ne
rect 4863 20 4903 32
tri 4903 20 4929 46 sw
rect 4992 42 5170 46
tri 5170 42 5174 46 sw
tri 4992 20 5014 42 ne
rect 5014 20 5174 42
tri 4706 -28 4754 20 ne
rect 4754 -15 4780 20
tri 4780 -15 4815 20 sw
tri 4863 -15 4898 20 ne
rect 4898 -15 4929 20
tri 4929 -15 4964 20 sw
tri 5014 -15 5049 20 ne
rect 5049 -15 5174 20
rect 4754 -28 4815 -15
tri 4754 -54 4780 -28 ne
rect 4780 -54 4815 -28
tri 4815 -54 4854 -15 sw
tri 4898 -54 4937 -15 ne
rect 4937 -43 4964 -15
tri 4964 -43 4992 -15 sw
tri 5049 -43 5077 -15 ne
rect 5077 -43 5174 -15
rect 4937 -54 4992 -43
tri 4992 -54 5003 -43 sw
tri 5077 -54 5088 -43 ne
rect 5088 -45 5174 -43
tri 5174 -45 5261 42 sw
rect 5088 -54 5261 -45
tri 4780 -122 4848 -54 ne
rect 4848 -81 4854 -54
tri 4854 -81 4881 -54 sw
tri 4937 -81 4964 -54 ne
rect 4964 -81 5003 -54
tri 5003 -81 5030 -54 sw
rect 4848 -122 4881 -81
tri 4881 -122 4922 -81 sw
tri 4964 -95 4978 -81 ne
rect 4978 -122 5030 -81
tri 5088 -99 5133 -54 ne
tri 4848 -128 4854 -122 ne
rect 4854 -128 4922 -122
tri 4922 -128 4928 -122 sw
tri 4854 -150 4876 -128 ne
rect 4712 -823 4764 -817
rect 4712 -887 4764 -875
rect 4712 -1128 4764 -939
rect 4876 -987 4928 -128
rect 4978 -186 5030 -174
rect 4978 -244 5030 -238
tri 4928 -987 5004 -911 sw
tri 4764 -1128 4782 -1110 sw
rect 4712 -1132 4782 -1128
tri 4712 -1140 4720 -1132 ne
rect 4720 -1140 4782 -1132
tri 4782 -1140 4794 -1128 sw
tri 4720 -1142 4722 -1140 ne
rect 4722 -1141 4794 -1140
tri 4794 -1141 4795 -1140 sw
rect 4876 -1141 4948 -987
rect 5133 -1076 5261 -54
rect 5133 -1128 5134 -1076
rect 5186 -1128 5208 -1076
rect 5260 -1128 5261 -1076
rect 4722 -1142 4795 -1141
tri 4795 -1142 4796 -1141 sw
rect 5133 -1142 5261 -1128
tri 4722 -1184 4764 -1142 ne
rect 4764 -1184 4796 -1142
tri 4764 -1194 4774 -1184 ne
rect 4774 -1194 4796 -1184
tri 4796 -1194 4848 -1142 sw
rect 5133 -1194 5134 -1142
rect 5186 -1194 5208 -1142
rect 5260 -1194 5261 -1142
tri 4774 -1208 4788 -1194 ne
rect 4788 -1208 4848 -1194
tri 4848 -1208 4862 -1194 sw
rect 5133 -1208 5261 -1194
tri 4788 -1214 4794 -1208 ne
rect 4794 -1214 4862 -1208
tri 4862 -1214 4868 -1208 sw
tri 4794 -1266 4846 -1214 ne
rect 4846 -1266 4970 -1214
rect 5022 -1266 5034 -1214
rect 5086 -1266 5092 -1214
rect 5133 -1260 5134 -1208
rect 5186 -1260 5208 -1208
rect 5260 -1260 5261 -1208
rect 5133 -1266 5261 -1260
<< via2 >>
rect 5341 3329 5397 3344
rect 5341 3288 5345 3329
rect 5345 3288 5397 3329
rect 5341 3213 5345 3264
rect 5345 3213 5397 3264
rect 5341 3208 5397 3213
rect 5378 3068 5434 3083
rect 5378 3027 5382 3068
rect 5382 3027 5434 3068
rect 5378 2952 5382 3003
rect 5382 2952 5434 3003
rect 5378 2947 5434 2952
rect 5665 2613 5721 2669
rect 5665 2533 5721 2589
rect 5455 2373 5511 2383
rect 5455 2327 5507 2373
rect 5507 2327 5511 2373
rect 5455 2257 5507 2303
rect 5507 2257 5511 2303
rect 5455 2247 5511 2257
rect 4929 1157 4985 1160
rect 4929 1105 4944 1157
rect 4944 1105 4956 1157
rect 4956 1105 4985 1157
rect 4929 1104 4985 1105
rect 4929 1024 4985 1080
rect 5455 656 5511 672
rect 5455 616 5459 656
rect 5459 616 5511 656
rect 5303 529 5359 549
rect 5303 493 5305 529
rect 5305 493 5357 529
rect 5357 493 5359 529
rect 5455 540 5459 592
rect 5459 540 5511 592
rect 5455 536 5511 540
rect 5770 621 5826 638
rect 5770 582 5774 621
rect 5774 582 5826 621
rect 5770 555 5826 558
rect 5770 503 5774 555
rect 5774 503 5826 555
rect 5770 502 5826 503
rect 5303 465 5359 469
rect 5303 413 5305 465
rect 5305 413 5357 465
rect 5357 413 5359 465
<< metal3 >>
tri 5278 3344 5283 3349 se
rect 5283 3344 5402 3349
tri 5222 3288 5278 3344 se
rect 5278 3288 5341 3344
rect 5397 3288 5402 3344
tri 5198 3264 5222 3288 se
rect 5222 3264 5402 3288
rect 5198 3208 5341 3264
rect 5397 3208 5402 3264
rect 5198 3203 5402 3208
tri 5104 1387 5198 1481 se
rect 5198 1453 5264 3203
tri 5264 3108 5359 3203 nw
rect 5373 3083 5439 3088
rect 5373 3027 5378 3083
rect 5434 3027 5439 3083
rect 5373 3003 5439 3027
rect 5373 2947 5378 3003
rect 5434 2947 5439 3003
tri 5198 1387 5264 1453 nw
tri 5324 2765 5373 2814 se
rect 5373 2786 5439 2947
rect 5373 2765 5418 2786
tri 5418 2765 5439 2786 nw
tri 5010 1293 5104 1387 se
tri 5104 1293 5198 1387 nw
tri 4924 1207 5010 1293 se
rect 5010 1207 5018 1293
tri 5018 1207 5104 1293 nw
rect 4924 1160 4990 1207
tri 4990 1179 5018 1207 nw
rect 4924 1104 4929 1160
rect 4985 1104 4990 1160
rect 4924 1080 4990 1104
rect 4924 1024 4929 1080
rect 4985 1024 4990 1080
rect 4924 1019 4990 1024
tri 5298 1073 5324 1099 se
rect 5324 1073 5390 2765
tri 5390 2737 5418 2765 nw
rect 5660 2669 5726 2674
rect 5660 2613 5665 2669
rect 5721 2613 5726 2669
rect 5660 2610 5726 2613
tri 5726 2610 5737 2621 sw
rect 5660 2589 5737 2610
rect 5660 2533 5665 2589
rect 5721 2533 5737 2589
rect 5660 2528 5737 2533
tri 5725 2516 5737 2528 ne
tri 5737 2516 5831 2610 sw
tri 5737 2488 5765 2516 ne
rect 5298 1071 5390 1073
rect 5298 549 5364 1071
tri 5364 1045 5390 1071 nw
rect 5450 2383 5516 2388
rect 5450 2327 5455 2383
rect 5511 2327 5516 2383
rect 5450 2303 5516 2327
rect 5450 2247 5455 2303
rect 5511 2247 5516 2303
rect 5298 493 5303 549
rect 5359 493 5364 549
rect 5450 672 5516 2247
rect 5450 616 5455 672
rect 5511 616 5516 672
rect 5450 592 5516 616
rect 5450 536 5455 592
rect 5511 536 5516 592
rect 5450 531 5516 536
rect 5765 638 5831 2516
rect 5765 582 5770 638
rect 5826 582 5831 638
rect 5765 558 5831 582
rect 5765 502 5770 558
rect 5826 502 5831 558
rect 5765 497 5831 502
rect 5298 469 5364 493
rect 5298 413 5303 469
rect 5359 413 5364 469
rect 5298 408 5364 413
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_0
timestamp 1694700623
transform 1 0 5244 0 1 1289
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_1
timestamp 1694700623
transform -1 0 5540 0 1 1289
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_2
timestamp 1694700623
transform 1 0 5596 0 1 1289
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_3
timestamp 1694700623
transform -1 0 5892 0 1 1289
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808618  sky130_fd_pr__nfet_01v8__example_55959141808618_0
timestamp 1694700623
transform 0 -1 5599 -1 0 363
box -1 0 181 1
use sky130_fd_pr__nfet_01v8__example_55959141808619  sky130_fd_pr__nfet_01v8__example_55959141808619_0
timestamp 1694700623
transform -1 0 5405 0 1 638
box -1 0 653 1
use sky130_fd_pr__nfet_01v8__example_55959141808620  sky130_fd_pr__nfet_01v8__example_55959141808620_0
timestamp 1694700623
transform -1 0 5911 0 1 64
box -1 0 51 1
use sky130_fd_pr__nfet_01v8__example_55959141808620  sky130_fd_pr__nfet_01v8__example_55959141808620_1
timestamp 1694700623
transform 1 0 5967 0 1 64
box -1 0 51 1
use sky130_fd_pr__nfet_01v8__example_55959141808621  sky130_fd_pr__nfet_01v8__example_55959141808621_0
timestamp 1694700623
transform -1 0 5641 0 1 968
box -1 0 889 1
use sky130_fd_pr__nfet_01v8__example_55959141808622  sky130_fd_pr__nfet_01v8__example_55959141808622_0
timestamp 1694700623
transform 0 1 4976 1 0 2496
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808622  sky130_fd_pr__nfet_01v8__example_55959141808622_1
timestamp 1694700623
transform 0 1 4976 1 0 2840
box -1 0 289 1
use sky130_fd_pr__nfet_01v8__example_55959141808623  sky130_fd_pr__nfet_01v8__example_55959141808623_0
timestamp 1694700623
transform 1 0 4878 0 1 1739
box -1 0 201 1
use sky130_fd_pr__nfet_01v8__example_55959141808623  sky130_fd_pr__nfet_01v8__example_55959141808623_1
timestamp 1694700623
transform 1 0 4878 0 -1 2216
box -1 0 201 1
use sky130_fd_pr__nfet_01v8__example_55959141808624  sky130_fd_pr__nfet_01v8__example_55959141808624_0
timestamp 1694700623
transform -1 0 4873 0 1 1298
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808624  sky130_fd_pr__nfet_01v8__example_55959141808624_1
timestamp 1694700623
transform 1 0 4929 0 1 1298
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180813  sky130_fd_pr__pfet_01v8__example_5595914180813_0
timestamp 1694700623
transform 1 0 5043 0 -1 473
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180813  sky130_fd_pr__pfet_01v8__example_5595914180813_1
timestamp 1694700623
transform -1 0 4987 0 -1 473
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_5595914180822  sky130_fd_pr__pfet_01v8__example_5595914180822_0
timestamp 1694700623
transform -1 0 4946 0 1 -1215
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_5595914180822  sky130_fd_pr__pfet_01v8__example_5595914180822_1
timestamp 1694700623
transform -1 0 4946 0 1 -866
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808430  sky130_fd_pr__pfet_01v8__example_55959141808430_0
timestamp 1694700623
transform 1 0 5864 0 1 369
box -1 0 157 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1694700623
transform 0 -1 5959 1 0 526
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1694700623
transform -1 0 5993 0 -1 89
box 0 0 1 1
<< labels >>
flabel metal1 s 5452 1974 5504 2026 3 FreeSans 200 0 0 0 SET_H
port 2 nsew
flabel metal1 s 5811 1973 5852 2025 3 FreeSans 200 0 0 0 HLD_H_N
port 3 nsew
flabel metal1 s 5286 1976 5327 2028 3 FreeSans 200 0 0 0 HLD_H_N
port 3 nsew
flabel metal1 s 4838 2127 4890 2179 3 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 4707 1421 4743 1473 3 FreeSans 200 0 0 0 OUT_H
port 5 nsew
flabel metal1 s 4817 372 4858 424 3 FreeSans 200 0 0 0 OUT_H_N
port 6 nsew
flabel metal1 s 5623 1970 5669 2022 3 FreeSans 200 0 0 0 RST_H
port 7 nsew
flabel metal1 s 4856 2547 4908 2599 3 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 5905 -18 5905 -18 3 FreeSans 520 0 0 0 IN
flabel metal1 s 5931 555 5983 595 3 FreeSans 200 0 0 0 VPWR
port 8 nsew
flabel metal1 s 5875 43 5927 95 3 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 5137 -1259 5184 -1234 3 FreeSans 520 0 0 0 VCC_IO
port 9 nsew
<< properties >>
string GDS_END 7910480
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7861298
<< end >>
