magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 2 21 1064 203
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 177
rect 164 47 194 177
rect 352 47 382 177
rect 436 47 466 177
rect 520 47 550 177
rect 604 47 634 177
rect 704 47 734 177
rect 788 47 818 177
rect 872 47 902 177
rect 956 47 986 177
<< scpmoshvt >>
rect 80 297 110 497
rect 164 297 194 497
rect 352 297 382 497
rect 436 297 466 497
rect 520 297 550 497
rect 604 297 634 497
rect 704 297 734 497
rect 788 297 818 497
rect 872 297 902 497
rect 956 297 986 497
<< ndiff >>
rect 28 163 80 177
rect 28 129 36 163
rect 70 129 80 163
rect 28 95 80 129
rect 28 61 36 95
rect 70 61 80 95
rect 28 47 80 61
rect 110 163 164 177
rect 110 129 120 163
rect 154 129 164 163
rect 110 47 164 129
rect 194 163 246 177
rect 194 129 204 163
rect 238 129 246 163
rect 194 95 246 129
rect 194 61 204 95
rect 238 61 246 95
rect 194 47 246 61
rect 300 95 352 177
rect 300 61 308 95
rect 342 61 352 95
rect 300 47 352 61
rect 382 163 436 177
rect 382 129 392 163
rect 426 129 436 163
rect 382 47 436 129
rect 466 95 520 177
rect 466 61 476 95
rect 510 61 520 95
rect 466 47 520 61
rect 550 163 604 177
rect 550 129 560 163
rect 594 129 604 163
rect 550 47 604 129
rect 634 163 704 177
rect 634 129 653 163
rect 687 129 704 163
rect 634 95 704 129
rect 634 61 653 95
rect 687 61 704 95
rect 634 47 704 61
rect 734 95 788 177
rect 734 61 744 95
rect 778 61 788 95
rect 734 47 788 61
rect 818 163 872 177
rect 818 129 828 163
rect 862 129 872 163
rect 818 95 872 129
rect 818 61 828 95
rect 862 61 872 95
rect 818 47 872 61
rect 902 95 956 177
rect 902 61 912 95
rect 946 61 956 95
rect 902 47 956 61
rect 986 163 1038 177
rect 986 129 996 163
rect 1030 129 1038 163
rect 986 95 1038 129
rect 986 61 996 95
rect 1030 61 1038 95
rect 986 47 1038 61
<< pdiff >>
rect 28 483 80 497
rect 28 449 36 483
rect 70 449 80 483
rect 28 415 80 449
rect 28 381 36 415
rect 70 381 80 415
rect 28 347 80 381
rect 28 313 36 347
rect 70 313 80 347
rect 28 297 80 313
rect 110 477 164 497
rect 110 443 120 477
rect 154 443 164 477
rect 110 409 164 443
rect 110 375 120 409
rect 154 375 164 409
rect 110 341 164 375
rect 110 307 120 341
rect 154 307 164 341
rect 110 297 164 307
rect 194 477 352 497
rect 194 443 204 477
rect 238 443 308 477
rect 342 443 352 477
rect 194 297 352 443
rect 382 477 436 497
rect 382 443 392 477
rect 426 443 436 477
rect 382 297 436 443
rect 466 409 520 497
rect 466 375 476 409
rect 510 375 520 409
rect 466 297 520 375
rect 550 477 604 497
rect 550 443 560 477
rect 594 443 604 477
rect 550 297 604 443
rect 634 477 704 497
rect 634 443 644 477
rect 678 443 704 477
rect 634 297 704 443
rect 734 477 788 497
rect 734 443 744 477
rect 778 443 788 477
rect 734 297 788 443
rect 818 409 872 497
rect 818 375 828 409
rect 862 375 872 409
rect 818 297 872 375
rect 902 477 956 497
rect 902 443 912 477
rect 946 443 956 477
rect 902 409 956 443
rect 902 375 912 409
rect 946 375 956 409
rect 902 297 956 375
rect 986 477 1043 497
rect 986 443 997 477
rect 1031 443 1043 477
rect 986 409 1043 443
rect 986 375 997 409
rect 1031 375 1043 409
rect 986 341 1043 375
rect 986 307 997 341
rect 1031 307 1043 341
rect 986 297 1043 307
<< ndiffc >>
rect 36 129 70 163
rect 36 61 70 95
rect 120 129 154 163
rect 204 129 238 163
rect 204 61 238 95
rect 308 61 342 95
rect 392 129 426 163
rect 476 61 510 95
rect 560 129 594 163
rect 653 129 687 163
rect 653 61 687 95
rect 744 61 778 95
rect 828 129 862 163
rect 828 61 862 95
rect 912 61 946 95
rect 996 129 1030 163
rect 996 61 1030 95
<< pdiffc >>
rect 36 449 70 483
rect 36 381 70 415
rect 36 313 70 347
rect 120 443 154 477
rect 120 375 154 409
rect 120 307 154 341
rect 204 443 238 477
rect 308 443 342 477
rect 392 443 426 477
rect 476 375 510 409
rect 560 443 594 477
rect 644 443 678 477
rect 744 443 778 477
rect 828 375 862 409
rect 912 443 946 477
rect 912 375 946 409
rect 997 443 1031 477
rect 997 375 1031 409
rect 997 307 1031 341
<< poly >>
rect 80 497 110 523
rect 164 497 194 523
rect 352 497 382 523
rect 436 497 466 523
rect 520 497 550 523
rect 604 497 634 523
rect 704 497 734 523
rect 788 497 818 523
rect 872 497 902 523
rect 956 497 986 523
rect 80 265 110 297
rect 164 265 194 297
rect 352 265 382 297
rect 436 265 466 297
rect 520 265 550 297
rect 604 265 634 297
rect 704 265 734 297
rect 788 265 818 297
rect 872 265 902 297
rect 956 265 986 297
rect 21 249 194 265
rect 21 215 37 249
rect 71 215 194 249
rect 21 199 194 215
rect 340 249 394 265
rect 340 215 350 249
rect 384 215 394 249
rect 340 199 394 215
rect 436 249 550 265
rect 436 215 476 249
rect 510 215 550 249
rect 436 199 550 215
rect 592 249 646 265
rect 592 215 602 249
rect 636 215 646 249
rect 592 199 646 215
rect 692 249 746 265
rect 692 215 702 249
rect 736 215 746 249
rect 692 199 746 215
rect 788 249 902 265
rect 788 215 828 249
rect 862 215 902 249
rect 788 199 902 215
rect 944 249 998 265
rect 944 215 954 249
rect 988 215 998 249
rect 944 199 998 215
rect 80 177 110 199
rect 164 177 194 199
rect 352 177 382 199
rect 436 177 466 199
rect 520 177 550 199
rect 604 177 634 199
rect 704 177 734 199
rect 788 177 818 199
rect 872 177 902 199
rect 956 177 986 199
rect 80 21 110 47
rect 164 21 194 47
rect 352 21 382 47
rect 436 21 466 47
rect 520 21 550 47
rect 604 21 634 47
rect 704 21 734 47
rect 788 21 818 47
rect 872 21 902 47
rect 956 21 986 47
<< polycont >>
rect 37 215 71 249
rect 350 215 384 249
rect 476 215 510 249
rect 602 215 636 249
rect 702 215 736 249
rect 828 215 862 249
rect 954 215 988 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 28 483 78 527
rect 28 449 36 483
rect 70 449 78 483
rect 28 415 78 449
rect 28 381 36 415
rect 70 381 78 415
rect 28 347 78 381
rect 28 313 36 347
rect 70 313 78 347
rect 28 291 78 313
rect 112 477 162 493
rect 112 443 120 477
rect 154 443 162 477
rect 112 409 162 443
rect 196 477 350 527
rect 196 443 204 477
rect 238 443 308 477
rect 342 443 350 477
rect 196 425 350 443
rect 384 477 602 493
rect 384 443 392 477
rect 426 459 560 477
rect 426 443 434 459
rect 384 425 434 443
rect 552 443 560 459
rect 594 443 602 477
rect 552 425 602 443
rect 636 477 702 527
rect 636 443 644 477
rect 678 443 702 477
rect 636 425 702 443
rect 736 477 954 493
rect 736 443 744 477
rect 778 459 912 477
rect 778 443 786 459
rect 736 425 786 443
rect 904 443 912 459
rect 946 443 954 477
rect 112 375 120 409
rect 154 391 162 409
rect 468 409 518 425
rect 468 391 476 409
rect 154 375 476 391
rect 510 391 518 409
rect 820 409 870 425
rect 820 391 828 409
rect 510 375 828 391
rect 862 375 870 409
rect 112 357 870 375
rect 904 409 954 443
rect 904 375 912 409
rect 946 375 954 409
rect 904 357 954 375
rect 997 477 1038 527
rect 1031 443 1038 477
rect 997 409 1038 443
rect 1031 375 1038 409
rect 112 341 170 357
rect 112 307 120 341
rect 154 307 170 341
rect 997 341 1038 375
rect 112 289 170 307
rect 17 249 87 255
rect 17 215 37 249
rect 71 215 87 249
rect 20 163 70 179
rect 121 173 170 289
rect 204 289 652 323
rect 204 249 407 289
rect 204 215 350 249
rect 384 215 407 249
rect 441 249 552 255
rect 441 215 476 249
rect 510 215 552 249
rect 586 249 652 289
rect 586 215 602 249
rect 636 215 652 249
rect 686 289 963 323
rect 1031 307 1038 341
rect 997 291 1038 307
rect 686 249 752 289
rect 929 255 963 289
rect 686 215 702 249
rect 736 215 752 249
rect 796 249 895 255
rect 796 215 828 249
rect 862 215 895 249
rect 929 249 1087 255
rect 929 215 954 249
rect 988 215 1087 249
rect 20 129 36 163
rect 104 163 170 173
rect 104 129 120 163
rect 154 129 170 163
rect 204 163 610 181
rect 238 129 392 163
rect 426 129 560 163
rect 594 129 610 163
rect 644 163 1046 181
rect 644 129 653 163
rect 687 147 828 163
rect 687 129 710 147
rect 20 95 70 129
rect 204 95 254 129
rect 644 95 710 129
rect 812 129 828 147
rect 862 145 996 163
rect 862 129 878 145
rect 20 61 36 95
rect 70 61 204 95
rect 238 61 254 95
rect 20 51 254 61
rect 292 61 308 95
rect 342 61 476 95
rect 510 61 653 95
rect 687 61 710 95
rect 292 51 710 61
rect 744 95 778 111
rect 744 17 778 61
rect 812 95 878 129
rect 980 129 996 145
rect 1030 129 1046 163
rect 812 61 828 95
rect 862 61 878 95
rect 812 51 878 61
rect 912 95 946 111
rect 912 17 946 61
rect 980 95 1046 129
rect 980 61 996 95
rect 1030 61 1046 95
rect 980 51 1046 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 493 221 527 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 309 357 343 391 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 861 221 895 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 1045 221 1079 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o221ai_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 834742
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 826076
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.520 0.000 
<< end >>
