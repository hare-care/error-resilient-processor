magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 614 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 234 47 264 177
rect 318 47 348 177
rect 402 47 432 177
rect 502 47 532 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 318 297 348 497
rect 402 297 432 497
rect 502 297 532 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 234 177
rect 109 127 190 161
rect 224 127 234 161
rect 109 93 234 127
rect 109 59 174 93
rect 208 59 234 93
rect 109 47 234 59
rect 264 93 318 177
rect 264 59 274 93
rect 308 59 318 93
rect 264 47 318 59
rect 348 161 402 177
rect 348 127 358 161
rect 392 127 402 161
rect 348 93 402 127
rect 348 59 358 93
rect 392 59 402 93
rect 348 47 402 59
rect 432 93 502 177
rect 432 59 458 93
rect 492 59 502 93
rect 432 47 502 59
rect 532 161 588 177
rect 532 127 542 161
rect 576 127 588 161
rect 532 93 588 127
rect 532 59 542 93
rect 576 59 588 93
rect 532 47 588 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 297 318 497
rect 348 297 402 497
rect 432 297 502 497
rect 532 485 588 497
rect 532 451 542 485
rect 576 451 588 485
rect 532 417 588 451
rect 532 383 542 417
rect 576 383 588 417
rect 532 349 588 383
rect 532 315 542 349
rect 576 315 588 349
rect 532 297 588 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 190 127 224 161
rect 174 59 208 93
rect 274 59 308 93
rect 358 127 392 161
rect 358 59 392 93
rect 458 59 492 93
rect 542 127 576 161
rect 542 59 576 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 542 451 576 485
rect 542 383 576 417
rect 542 315 576 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 318 497 348 523
rect 402 497 432 523
rect 502 497 532 523
rect 79 261 109 297
rect 21 249 109 261
rect 21 215 38 249
rect 72 215 109 249
rect 21 203 109 215
rect 163 259 193 297
rect 318 265 348 297
rect 402 265 432 297
rect 502 265 532 297
rect 163 249 264 259
rect 163 215 214 249
rect 248 215 264 249
rect 163 205 264 215
rect 79 177 109 203
rect 234 177 264 205
rect 306 249 360 265
rect 306 215 316 249
rect 350 215 360 249
rect 306 199 360 215
rect 402 249 460 265
rect 402 215 416 249
rect 450 215 460 249
rect 402 199 460 215
rect 502 249 560 265
rect 502 215 516 249
rect 550 215 560 249
rect 502 199 560 215
rect 318 177 348 199
rect 402 177 432 199
rect 502 177 532 199
rect 79 21 109 47
rect 234 21 264 47
rect 318 21 348 47
rect 402 21 432 47
rect 502 21 532 47
<< polycont >>
rect 38 215 72 249
rect 214 215 248 249
rect 316 215 350 249
rect 416 215 450 249
rect 516 215 550 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 289 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 526 485 592 527
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 103 315 119 349
rect 153 315 169 349
rect 103 297 169 315
rect 21 249 88 255
rect 21 215 38 249
rect 72 215 88 249
rect 122 181 156 297
rect 203 249 264 471
rect 198 215 214 249
rect 248 215 264 249
rect 300 249 364 471
rect 398 283 466 471
rect 526 451 542 485
rect 576 451 592 485
rect 526 417 592 451
rect 526 383 542 417
rect 576 383 592 417
rect 526 349 592 383
rect 526 315 542 349
rect 576 315 592 349
rect 526 299 592 315
rect 400 249 466 283
rect 300 215 316 249
rect 350 215 366 249
rect 400 215 416 249
rect 450 215 466 249
rect 500 249 616 265
rect 500 215 516 249
rect 550 215 616 249
rect 17 161 156 181
rect 17 127 35 161
rect 69 147 156 161
rect 190 161 592 181
rect 69 127 85 147
rect 17 93 85 127
rect 224 147 358 161
rect 190 113 224 127
rect 342 127 358 147
rect 392 147 542 161
rect 392 127 408 147
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 158 93 224 113
rect 158 59 174 93
rect 208 59 224 93
rect 158 51 224 59
rect 258 93 308 113
rect 258 59 274 93
rect 258 17 308 59
rect 342 93 408 127
rect 526 127 542 147
rect 576 127 592 161
rect 342 59 358 93
rect 392 59 408 93
rect 342 51 408 59
rect 442 93 492 113
rect 442 59 458 93
rect 442 17 492 59
rect 526 93 592 127
rect 526 59 542 93
rect 576 59 592 93
rect 526 51 592 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 398 425 432 459 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 357 432 391 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 425 340 459 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 306 357 340 391 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 306 289 340 323 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 214 425 248 459 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 214 357 248 391 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 214 289 248 323 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 85 64 119 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B1
port 5 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o41ai_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 719410
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 712164
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
