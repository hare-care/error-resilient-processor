magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 3350 582
<< pwell >>
rect 79 21 3273 203
rect 29 -17 63 17
<< locali >>
rect 17 199 133 265
rect 1937 325 1987 425
rect 2105 325 2155 425
rect 2273 325 2323 425
rect 2441 325 2491 425
rect 2609 325 2659 425
rect 2777 325 2827 425
rect 2945 325 2995 425
rect 3113 325 3163 425
rect 1937 291 3295 325
rect 1890 215 3130 257
rect 17 51 63 199
rect 3164 181 3295 291
rect 585 145 3295 181
rect 585 51 651 145
rect 753 51 819 145
rect 921 51 987 145
rect 1089 51 1155 145
rect 1257 51 1323 145
rect 1425 51 1491 145
rect 1593 51 1659 145
rect 1761 51 1827 145
rect 1929 51 1995 145
rect 2097 51 2163 145
rect 2265 51 2331 145
rect 2433 51 2499 145
rect 2601 51 2667 145
rect 2769 51 2835 145
rect 2937 51 3003 145
rect 3105 51 3171 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 60 299 103 527
rect 137 299 203 493
rect 167 257 203 299
rect 237 291 271 527
rect 305 257 371 493
rect 405 291 454 527
rect 495 333 559 493
rect 593 367 643 527
rect 677 333 727 493
rect 761 367 811 527
rect 845 333 895 493
rect 929 367 979 527
rect 1013 333 1063 493
rect 1097 367 1147 527
rect 1181 333 1231 493
rect 1265 367 1315 527
rect 1349 333 1399 493
rect 1433 367 1483 527
rect 1517 333 1567 493
rect 1601 367 1651 527
rect 1685 333 1735 493
rect 1769 367 1819 527
rect 1853 459 3247 493
rect 1853 333 1903 459
rect 495 291 1903 333
rect 2021 359 2071 459
rect 2189 359 2239 459
rect 2357 359 2407 459
rect 2525 359 2575 459
rect 2693 359 2743 459
rect 2861 359 2911 459
rect 3029 359 3079 459
rect 3197 359 3247 459
rect 167 215 1856 257
rect 167 213 407 215
rect 97 17 163 165
rect 197 51 239 213
rect 273 17 323 179
rect 357 51 407 213
rect 441 17 551 181
rect 685 17 719 111
rect 853 17 887 111
rect 1021 17 1055 111
rect 1189 17 1223 111
rect 1357 17 1391 111
rect 1525 17 1559 111
rect 1693 17 1727 111
rect 1861 17 1895 111
rect 2029 17 2063 111
rect 2197 17 2231 111
rect 2365 17 2399 111
rect 2533 17 2567 111
rect 2701 17 2735 111
rect 2869 17 2903 111
rect 3037 17 3071 111
rect 3205 17 3259 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 3157 527 3191 561
rect 3249 527 3283 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
rect 3157 -17 3191 17
rect 3249 -17 3283 17
<< metal1 >>
rect 0 561 3312 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3312 561
rect 0 496 3312 527
rect 0 17 3312 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3312 17
rect 0 -48 3312 -17
<< labels >>
rlabel locali s 17 51 63 199 6 A
port 1 nsew signal input
rlabel locali s 17 199 133 265 6 A
port 1 nsew signal input
rlabel locali s 1890 215 3130 257 6 SLEEP
port 2 nsew signal input
rlabel metal1 s 0 -48 3312 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 3350 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 3312 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 3105 51 3171 145 6 X
port 7 nsew signal output
rlabel locali s 2937 51 3003 145 6 X
port 7 nsew signal output
rlabel locali s 2769 51 2835 145 6 X
port 7 nsew signal output
rlabel locali s 2601 51 2667 145 6 X
port 7 nsew signal output
rlabel locali s 2433 51 2499 145 6 X
port 7 nsew signal output
rlabel locali s 2265 51 2331 145 6 X
port 7 nsew signal output
rlabel locali s 2097 51 2163 145 6 X
port 7 nsew signal output
rlabel locali s 1929 51 1995 145 6 X
port 7 nsew signal output
rlabel locali s 1761 51 1827 145 6 X
port 7 nsew signal output
rlabel locali s 1593 51 1659 145 6 X
port 7 nsew signal output
rlabel locali s 1425 51 1491 145 6 X
port 7 nsew signal output
rlabel locali s 1257 51 1323 145 6 X
port 7 nsew signal output
rlabel locali s 1089 51 1155 145 6 X
port 7 nsew signal output
rlabel locali s 921 51 987 145 6 X
port 7 nsew signal output
rlabel locali s 753 51 819 145 6 X
port 7 nsew signal output
rlabel locali s 585 51 651 145 6 X
port 7 nsew signal output
rlabel locali s 585 145 3295 181 6 X
port 7 nsew signal output
rlabel locali s 3164 181 3295 291 6 X
port 7 nsew signal output
rlabel locali s 1937 291 3295 325 6 X
port 7 nsew signal output
rlabel locali s 3113 325 3163 425 6 X
port 7 nsew signal output
rlabel locali s 2945 325 2995 425 6 X
port 7 nsew signal output
rlabel locali s 2777 325 2827 425 6 X
port 7 nsew signal output
rlabel locali s 2609 325 2659 425 6 X
port 7 nsew signal output
rlabel locali s 2441 325 2491 425 6 X
port 7 nsew signal output
rlabel locali s 2273 325 2323 425 6 X
port 7 nsew signal output
rlabel locali s 2105 325 2155 425 6 X
port 7 nsew signal output
rlabel locali s 1937 325 1987 425 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3312 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2422542
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2398934
<< end >>
