// input external delay: 4 ns
// in delay: 0.011365 ns
// input delay: 0.010861 ns
// output delay: 0.175128 ns
// out delay: 0.000627 ns
// total extra delay: 4.197981 ns
// critical path time: 11.947532  ns
// total inverter delay needed: 11.947532 - 4.197981 = 7.647751 ns
// average one inverter delay: 0.03012 ns
// inverters needed: 256

module inverter(input wire a, output wire y);
     not (y, a);
endmodule

module multiplier_replica(input wire in, output wire out);
    wire [253:0] interconnections; // Wires to connect inverters

    // Instantiate inverters individually with connections from 1 to 318
    inverter inv1(in, interconnections[0]);
    inverter inv2(interconnections[0], interconnections[1]);
    inverter inv3(interconnections[1], interconnections[2]);
    inverter inv4(interconnections[2], interconnections[3]);
    inverter inv5(interconnections[3], interconnections[4]);
    inverter inv6(interconnections[4], interconnections[5]);
    inverter inv7(interconnections[5], interconnections[6]);
    inverter inv8(interconnections[6], interconnections[7]);
    inverter inv9(interconnections[7], interconnections[8]);
    inverter inv10(interconnections[8], interconnections[9]);
    inverter inv11(interconnections[9], interconnections[10]);
    inverter inv12(interconnections[10], interconnections[11]);
    inverter inv13(interconnections[11], interconnections[12]);
    inverter inv14(interconnections[12], interconnections[13]);
    inverter inv15(interconnections[13], interconnections[14]);
    inverter inv16(interconnections[14], interconnections[15]);
    inverter inv17(interconnections[15], interconnections[16]);
    inverter inv18(interconnections[16], interconnections[17]);
    inverter inv19(interconnections[17], interconnections[18]);
    inverter inv20(interconnections[18], interconnections[19]);
    inverter inv21(interconnections[19], interconnections[20]);
    inverter inv22(interconnections[20], interconnections[21]);
    inverter inv23(interconnections[21], interconnections[22]);
    inverter inv24(interconnections[22], interconnections[23]);
    inverter inv25(interconnections[23], interconnections[24]);
    inverter inv26(interconnections[24], interconnections[25]);
    inverter inv27(interconnections[25], interconnections[26]);
    inverter inv28(interconnections[26], interconnections[27]);
    inverter inv29(interconnections[27], interconnections[28]);
    inverter inv30(interconnections[28], interconnections[29]);
    inverter inv31(interconnections[29], interconnections[30]);
    inverter inv32(interconnections[30], interconnections[31]);
    inverter inv33(interconnections[31], interconnections[32]);
    inverter inv34(interconnections[32], interconnections[33]);
    inverter inv35(interconnections[33], interconnections[34]);
    inverter inv36(interconnections[34], interconnections[35]);
    inverter inv37(interconnections[35], interconnections[36]);
    inverter inv38(interconnections[36], interconnections[37]);
    inverter inv39(interconnections[37], interconnections[38]);
    inverter inv40(interconnections[38], interconnections[39]);
    inverter inv41(interconnections[39], interconnections[40]);
    inverter inv42(interconnections[40], interconnections[41]);
    inverter inv43(interconnections[41], interconnections[42]);
    inverter inv44(interconnections[42], interconnections[43]);
    inverter inv45(interconnections[43], interconnections[44]);
    inverter inv46(interconnections[44], interconnections[45]);
    inverter inv47(interconnections[45], interconnections[46]);
    inverter inv48(interconnections[46], interconnections[47]);
    inverter inv49(interconnections[47], interconnections[48]);
    inverter inv50(interconnections[48], interconnections[49]);
    inverter inv51(interconnections[49], interconnections[50]);
    inverter inv52(interconnections[50], interconnections[51]);
    inverter inv53(interconnections[51], interconnections[52]);
    inverter inv54(interconnections[52], interconnections[53]);
    inverter inv55(interconnections[53], interconnections[54]);
    inverter inv56(interconnections[54], interconnections[55]);
    inverter inv57(interconnections[55], interconnections[56]);
    inverter inv58(interconnections[56], interconnections[57]);
    inverter inv59(interconnections[57], interconnections[58]);
    inverter inv60(interconnections[58], interconnections[59]);
    inverter inv61(interconnections[59], interconnections[60]);
    inverter inv62(interconnections[60], interconnections[61]);
    inverter inv63(interconnections[61], interconnections[62]);
    inverter inv64(interconnections[62], interconnections[63]);
    inverter inv65(interconnections[63], interconnections[64]);
    inverter inv66(interconnections[64], interconnections[65]);
    inverter inv67(interconnections[65], interconnections[66]);
    inverter inv68(interconnections[66], interconnections[67]);
    inverter inv69(interconnections[67], interconnections[68]);
    inverter inv70(interconnections[68], interconnections[69]);
    inverter inv71(interconnections[69], interconnections[70]);
    inverter inv72(interconnections[70], interconnections[71]);
    inverter inv73(interconnections[71], interconnections[72]);
    inverter inv74(interconnections[72], interconnections[73]);
    inverter inv75(interconnections[73], interconnections[74]);
    inverter inv76(interconnections[74], interconnections[75]);
    inverter inv77(interconnections[75], interconnections[76]);
    inverter inv78(interconnections[76], interconnections[77]);
    inverter inv79(interconnections[77], interconnections[78]);
    inverter inv80(interconnections[78], interconnections[79]);
    inverter inv81(interconnections[79], interconnections[80]);
    inverter inv82(interconnections[80], interconnections[81]);
    inverter inv83(interconnections[81], interconnections[82]);
    inverter inv84(interconnections[82], interconnections[83]);
    inverter inv85(interconnections[83], interconnections[84]);
    inverter inv86(interconnections[84], interconnections[85]);
    inverter inv87(interconnections[85], interconnections[86]);
    inverter inv88(interconnections[86], interconnections[87]);
    inverter inv89(interconnections[87], interconnections[88]);
    inverter inv90(interconnections[88], interconnections[89]);
    inverter inv91(interconnections[89], interconnections[90]);
    inverter inv92(interconnections[90], interconnections[91]);
    inverter inv93(interconnections[91], interconnections[92]);
    inverter inv94(interconnections[92], interconnections[93]);
    inverter inv95(interconnections[93], interconnections[94]);
    inverter inv96(interconnections[94], interconnections[95]);
    inverter inv97(interconnections[95], interconnections[96]);
    inverter inv98(interconnections[96], interconnections[97]);
    inverter inv99(interconnections[97], interconnections[98]);
    inverter inv100(interconnections[98], interconnections[99]);
    inverter inv101(interconnections[99], interconnections[100]);
    inverter inv102(interconnections[100], interconnections[101]);
    inverter inv103(interconnections[101], interconnections[102]);
    inverter inv104(interconnections[102], interconnections[103]);
    inverter inv105(interconnections[103], interconnections[104]);
    inverter inv106(interconnections[104], interconnections[105]);
    inverter inv107(interconnections[105], interconnections[106]);
    inverter inv108(interconnections[106], interconnections[107]);
    inverter inv109(interconnections[107], interconnections[108]);
    inverter inv110(interconnections[108], interconnections[109]);
    inverter inv111(interconnections[109], interconnections[110]);
    inverter inv112(interconnections[110], interconnections[111]);
    inverter inv113(interconnections[111], interconnections[112]);
    inverter inv114(interconnections[112], interconnections[113]);
    inverter inv115(interconnections[113], interconnections[114]);
    inverter inv116(interconnections[114], interconnections[115]);
    inverter inv117(interconnections[115], interconnections[116]);
    inverter inv118(interconnections[116], interconnections[117]);
    inverter inv119(interconnections[117], interconnections[118]);
    inverter inv120(interconnections[118], interconnections[119]);
    inverter inv121(interconnections[119], interconnections[120]);
    inverter inv122(interconnections[120], interconnections[121]);
    inverter inv123(interconnections[121], interconnections[122]);
    inverter inv124(interconnections[122], interconnections[123]);
    inverter inv125(interconnections[123], interconnections[124]);
    inverter inv126(interconnections[124], interconnections[125]);
    inverter inv127(interconnections[125], interconnections[126]);
    inverter inv128(interconnections[126], interconnections[127]);
    inverter inv129(interconnections[127], interconnections[128]);
    inverter inv130(interconnections[128], interconnections[129]);
    inverter inv131(interconnections[129], interconnections[130]);
    inverter inv132(interconnections[130], interconnections[131]);
    inverter inv133(interconnections[131], interconnections[132]);
    inverter inv134(interconnections[132], interconnections[133]);
    inverter inv135(interconnections[133], interconnections[134]);
    inverter inv136(interconnections[134], interconnections[135]);
    inverter inv137(interconnections[135], interconnections[136]);
    inverter inv138(interconnections[136], interconnections[137]);
    inverter inv139(interconnections[137], interconnections[138]);
    inverter inv140(interconnections[138], interconnections[139]);
    inverter inv141(interconnections[139], interconnections[140]);
    inverter inv142(interconnections[140], interconnections[141]);
    inverter inv143(interconnections[141], interconnections[142]);
    inverter inv144(interconnections[142], interconnections[143]);
    inverter inv145(interconnections[143], interconnections[144]);
    inverter inv146(interconnections[144], interconnections[145]);
    inverter inv147(interconnections[145], interconnections[146]);
    inverter inv148(interconnections[146], interconnections[147]);
    inverter inv149(interconnections[147], interconnections[148]);
    inverter inv150(interconnections[148], interconnections[149]);
    inverter inv151(interconnections[149], interconnections[150]);
    inverter inv152(interconnections[150], interconnections[151]);
    inverter inv153(interconnections[151], interconnections[152]);
    inverter inv154(interconnections[152], interconnections[153]);
    inverter inv155(interconnections[153], interconnections[154]);
    inverter inv156(interconnections[154], interconnections[155]);
    inverter inv157(interconnections[155], interconnections[156]);
    inverter inv158(interconnections[156], interconnections[157]);
    inverter inv159(interconnections[157], interconnections[158]);
    inverter inv160(interconnections[158], interconnections[159]);
    inverter inv161(interconnections[159], interconnections[160]);
    inverter inv162(interconnections[160], interconnections[161]);
    inverter inv163(interconnections[161], interconnections[162]);
    inverter inv164(interconnections[162], interconnections[163]);
    inverter inv165(interconnections[163], interconnections[164]);
    inverter inv166(interconnections[164], interconnections[165]);
    inverter inv167(interconnections[165], interconnections[166]);
    inverter inv168(interconnections[166], interconnections[167]);
    inverter inv169(interconnections[167], interconnections[168]);
    inverter inv170(interconnections[168], interconnections[169]);
    inverter inv171(interconnections[169], interconnections[170]);
    inverter inv172(interconnections[170], interconnections[171]);
    inverter inv173(interconnections[171], interconnections[172]);
    inverter inv174(interconnections[172], interconnections[173]);
    inverter inv175(interconnections[173], interconnections[174]);
    inverter inv176(interconnections[174], interconnections[175]);
    inverter inv177(interconnections[175], interconnections[176]);
    inverter inv178(interconnections[176], interconnections[177]);
    inverter inv179(interconnections[177], interconnections[178]);
    inverter inv180(interconnections[178], interconnections[179]);
    inverter inv181(interconnections[179], interconnections[180]);
    inverter inv182(interconnections[180], interconnections[181]);
    inverter inv183(interconnections[181], interconnections[182]);
    inverter inv184(interconnections[182], interconnections[183]);
    inverter inv185(interconnections[183], interconnections[184]);
    inverter inv186(interconnections[184], interconnections[185]);
    inverter inv187(interconnections[185], interconnections[186]);
    inverter inv188(interconnections[186], interconnections[187]);
    inverter inv189(interconnections[187], interconnections[188]);
    inverter inv190(interconnections[188], interconnections[189]);
    inverter inv191(interconnections[189], interconnections[190]);
    inverter inv192(interconnections[190], interconnections[191]);
    inverter inv193(interconnections[191], interconnections[192]);
    inverter inv194(interconnections[192], interconnections[193]);
    inverter inv195(interconnections[193], interconnections[194]);
    inverter inv196(interconnections[194], interconnections[195]);
    inverter inv197(interconnections[195], interconnections[196]);
    inverter inv198(interconnections[196], interconnections[197]);
    inverter inv199(interconnections[197], interconnections[198]);
    inverter inv200(interconnections[198], interconnections[199]);
    inverter inv201(interconnections[199], interconnections[200]);
    inverter inv202(interconnections[200], interconnections[201]);
    inverter inv203(interconnections[201], interconnections[202]);
    inverter inv204(interconnections[202], interconnections[203]);
    inverter inv205(interconnections[203], interconnections[204]);
    inverter inv206(interconnections[204], interconnections[205]);
    inverter inv207(interconnections[205], interconnections[206]);
    inverter inv208(interconnections[206], interconnections[207]);
    inverter inv209(interconnections[207], interconnections[208]);
    inverter inv210(interconnections[208], interconnections[209]);
    inverter inv211(interconnections[209], interconnections[210]);
    inverter inv212(interconnections[210], interconnections[211]);
    inverter inv213(interconnections[211], interconnections[212]);
    inverter inv214(interconnections[212], interconnections[213]);
    inverter inv215(interconnections[213], interconnections[214]);
    inverter inv216(interconnections[214], interconnections[215]);
    inverter inv217(interconnections[215], interconnections[216]);
    inverter inv218(interconnections[216], interconnections[217]);
    inverter inv219(interconnections[217], interconnections[218]);
    inverter inv220(interconnections[218], interconnections[219]);
    inverter inv221(interconnections[219], interconnections[220]);
    inverter inv222(interconnections[220], interconnections[221]);
    inverter inv223(interconnections[221], interconnections[222]);
    inverter inv224(interconnections[222], interconnections[223]);
    inverter inv225(interconnections[223], interconnections[224]);
    inverter inv226(interconnections[224], interconnections[225]);
    inverter inv227(interconnections[225], interconnections[226]);
    inverter inv228(interconnections[226], interconnections[227]);
    inverter inv229(interconnections[227], interconnections[228]);
    inverter inv230(interconnections[228], interconnections[229]);
    inverter inv231(interconnections[229], interconnections[230]);
    inverter inv232(interconnections[230], interconnections[231]);
    inverter inv233(interconnections[231], interconnections[232]);
    inverter inv234(interconnections[232], interconnections[233]);
    inverter inv235(interconnections[233], interconnections[234]);
    inverter inv236(interconnections[234], interconnections[235]);
    inverter inv237(interconnections[235], interconnections[236]);
    inverter inv238(interconnections[236], interconnections[237]);
    inverter inv239(interconnections[237], interconnections[238]);
    inverter inv240(interconnections[238], interconnections[239]);
    inverter inv241(interconnections[239], interconnections[240]);
    inverter inv242(interconnections[240], interconnections[241]);
    inverter inv243(interconnections[241], interconnections[242]);
    inverter inv244(interconnections[242], interconnections[243]);
    inverter inv245(interconnections[243], interconnections[244]);
    inverter inv246(interconnections[244], interconnections[245]);
    inverter inv247(interconnections[245], interconnections[246]);
    inverter inv248(interconnections[246], interconnections[247]);
    inverter inv249(interconnections[247], interconnections[248]);
    inverter inv250(interconnections[248], interconnections[249]);
    inverter inv251(interconnections[249], interconnections[250]);
    inverter inv252(interconnections[250], interconnections[251]);
    inverter inv253(interconnections[251], interconnections[252]);
    inverter inv254(interconnections[252], interconnections[253]);
    inverter inv255(interconnections[253], out);

endmodule