magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 269 203
rect 1 21 827 157
rect 30 -17 64 21
<< locali >>
rect 103 319 165 493
rect 103 150 137 319
rect 455 263 618 325
rect 455 256 489 263
rect 103 51 153 150
rect 363 153 489 256
rect 525 147 618 205
rect 672 151 710 325
rect 580 84 618 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 299 69 527
rect 205 435 263 527
rect 297 451 559 485
rect 297 401 331 451
rect 665 435 709 527
rect 743 401 810 493
rect 199 367 331 401
rect 365 367 810 401
rect 18 17 69 177
rect 199 265 233 367
rect 365 333 399 367
rect 171 199 233 265
rect 267 299 399 333
rect 267 199 301 299
rect 199 161 233 199
rect 199 127 321 161
rect 287 93 321 127
rect 187 17 253 93
rect 287 59 546 93
rect 670 17 710 117
rect 744 51 810 367
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 363 153 489 256 6 A0
port 1 nsew signal input
rlabel locali s 455 256 489 263 6 A0
port 1 nsew signal input
rlabel locali s 455 263 618 325 6 A0
port 1 nsew signal input
rlabel locali s 580 84 618 147 6 A1
port 2 nsew signal input
rlabel locali s 525 147 618 205 6 A1
port 2 nsew signal input
rlabel locali s 672 151 710 325 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 827 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 157 269 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 51 153 150 6 X
port 8 nsew signal output
rlabel locali s 103 150 137 319 6 X
port 8 nsew signal output
rlabel locali s 103 319 165 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1682210
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1675020
<< end >>
