magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 4 43 662 283
rect -26 -43 698 43
<< mvnmos >>
rect 83 173 183 257
rect 337 107 437 257
rect 479 107 579 257
<< mvpmos >>
rect 102 447 202 597
rect 313 443 413 743
rect 479 443 579 743
<< mvndiff >>
rect 30 232 83 257
rect 30 198 38 232
rect 72 198 83 232
rect 30 173 83 198
rect 183 249 337 257
rect 183 215 194 249
rect 228 215 292 249
rect 326 215 337 249
rect 183 173 337 215
rect 212 149 337 173
rect 212 115 224 149
rect 258 115 292 149
rect 326 115 337 149
rect 212 107 337 115
rect 437 107 479 257
rect 579 249 636 257
rect 579 215 590 249
rect 624 215 636 249
rect 579 149 636 215
rect 579 115 590 149
rect 624 115 636 149
rect 579 107 636 115
<< mvpdiff >>
rect 246 735 313 743
rect 246 701 258 735
rect 292 701 313 735
rect 246 655 313 701
rect 246 621 258 655
rect 292 621 313 655
rect 246 597 313 621
rect 45 589 102 597
rect 45 555 57 589
rect 91 555 102 589
rect 45 489 102 555
rect 45 455 57 489
rect 91 455 102 489
rect 45 447 102 455
rect 202 574 313 597
rect 202 540 258 574
rect 292 540 313 574
rect 202 494 313 540
rect 202 460 258 494
rect 292 460 313 494
rect 202 447 313 460
rect 263 443 313 447
rect 413 443 479 743
rect 579 735 636 743
rect 579 701 590 735
rect 624 701 636 735
rect 579 652 636 701
rect 579 618 590 652
rect 624 618 636 652
rect 579 568 636 618
rect 579 534 590 568
rect 624 534 636 568
rect 579 485 636 534
rect 579 451 590 485
rect 624 451 636 485
rect 579 443 636 451
<< mvndiffc >>
rect 38 198 72 232
rect 194 215 228 249
rect 292 215 326 249
rect 224 115 258 149
rect 292 115 326 149
rect 590 215 624 249
rect 590 115 624 149
<< mvpdiffc >>
rect 258 701 292 735
rect 258 621 292 655
rect 57 555 91 589
rect 57 455 91 489
rect 258 540 292 574
rect 258 460 292 494
rect 590 701 624 735
rect 590 618 624 652
rect 590 534 624 568
rect 590 451 624 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
<< poly >>
rect 313 743 413 769
rect 479 743 579 769
rect 102 597 202 623
rect 102 421 202 447
rect 313 421 413 443
rect 83 399 413 421
rect 479 411 579 443
rect 83 365 119 399
rect 153 365 187 399
rect 221 388 413 399
rect 455 395 579 411
rect 221 365 237 388
rect 83 321 237 365
rect 455 361 471 395
rect 505 361 579 395
rect 279 329 413 346
rect 455 345 579 361
rect 83 257 183 321
rect 279 295 295 329
rect 329 295 363 329
rect 397 303 413 329
rect 479 329 579 345
rect 397 295 437 303
rect 279 279 437 295
rect 337 257 437 279
rect 479 295 522 329
rect 556 295 579 329
rect 479 257 579 295
rect 83 147 183 173
rect 337 81 437 107
rect 479 81 579 107
<< polycont >>
rect 119 365 153 399
rect 187 365 221 399
rect 471 361 505 395
rect 295 295 329 329
rect 363 295 397 329
rect 522 295 556 329
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 148 735 554 751
rect 148 701 154 735
rect 188 701 226 735
rect 292 701 298 735
rect 332 701 370 735
rect 404 701 442 735
rect 476 701 514 735
rect 548 701 554 735
rect 148 655 554 701
rect 148 621 258 655
rect 292 621 554 655
rect 18 589 107 605
rect 18 555 57 589
rect 91 555 107 589
rect 18 489 107 555
rect 18 455 57 489
rect 91 460 107 489
rect 148 574 554 621
rect 148 540 258 574
rect 292 542 554 574
rect 590 735 647 751
rect 624 701 647 735
rect 590 652 647 701
rect 624 618 647 652
rect 590 568 647 618
rect 292 540 421 542
rect 148 494 421 540
rect 624 534 647 568
rect 148 460 258 494
rect 292 460 421 494
rect 18 439 91 455
rect 18 329 69 439
rect 127 405 359 424
rect 103 399 359 405
rect 103 365 119 399
rect 153 365 187 399
rect 221 365 359 399
rect 455 395 556 508
rect 455 361 471 395
rect 505 361 556 395
rect 455 345 556 361
rect 501 329 556 345
rect 18 295 295 329
rect 329 295 363 329
rect 397 295 413 329
rect 18 285 413 295
rect 501 295 522 329
rect 18 232 88 285
rect 18 198 38 232
rect 72 198 88 232
rect 18 182 88 198
rect 122 215 194 249
rect 228 215 292 249
rect 326 215 467 249
rect 501 232 556 295
rect 590 485 647 534
rect 624 451 647 485
rect 590 249 647 451
rect 122 180 467 215
rect 624 215 647 249
rect 122 149 554 180
rect 122 148 224 149
rect 88 115 224 148
rect 258 115 292 149
rect 326 115 554 149
rect 88 113 554 115
rect 122 79 160 113
rect 194 79 232 113
rect 266 79 304 113
rect 338 79 376 113
rect 410 79 448 113
rect 482 79 520 113
rect 590 149 647 215
rect 624 115 647 149
rect 590 99 647 115
rect 88 73 554 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 154 701 188 735
rect 226 701 258 735
rect 258 701 260 735
rect 298 701 332 735
rect 370 701 404 735
rect 442 701 476 735
rect 514 701 548 735
rect 88 79 122 113
rect 160 79 194 113
rect 232 79 266 113
rect 304 79 338 113
rect 376 79 410 113
rect 448 79 482 113
rect 520 79 554 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 154 735
rect 188 701 226 735
rect 260 701 298 735
rect 332 701 370 735
rect 404 701 442 735
rect 476 701 514 735
rect 548 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 88 113
rect 122 79 160 113
rect 194 79 232 113
rect 266 79 304 113
rect 338 79 376 113
rect 410 79 448 113
rect 482 79 520 113
rect 554 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvn_1
flabel metal1 s 0 51 672 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 672 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 672 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 672 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 612 641 646 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string GDS_END 1229982
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1220214
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
