magic
tech sky130A
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_0
timestamp 1694700623
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_1
timestamp 1694700623
transform 1 0 416 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_1
timestamp 1694700623
transform 1 0 652 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 7857454
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7855440
<< end >>
