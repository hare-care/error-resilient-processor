magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1924 201 2391 203
rect 780 157 1235 201
rect 1557 157 2391 201
rect 1 21 2391 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 446 47 476 119
rect 551 47 581 119
rect 647 47 677 131
rect 761 47 791 131
rect 857 47 887 175
rect 941 47 971 175
rect 1129 47 1159 175
rect 1249 47 1279 119
rect 1333 47 1363 119
rect 1428 47 1458 131
rect 1525 47 1555 131
rect 1633 47 1663 175
rect 1717 47 1747 175
rect 1905 47 1935 131
rect 2000 47 2030 177
rect 2188 47 2218 131
rect 2283 47 2313 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 413 381 497
rect 443 413 473 497
rect 527 413 557 497
rect 647 413 677 497
rect 753 413 783 497
rect 861 329 891 497
rect 945 329 975 497
rect 1082 329 1112 497
rect 1226 413 1256 497
rect 1310 413 1340 497
rect 1415 413 1445 497
rect 1536 413 1566 497
rect 1642 329 1672 497
rect 1714 329 1744 497
rect 1903 301 1933 429
rect 2000 297 2030 497
rect 2188 353 2218 481
rect 2283 297 2313 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 806 131 857 175
rect 596 119 647 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 551 119
rect 476 59 496 93
rect 530 59 551 93
rect 476 47 551 59
rect 581 47 647 119
rect 677 89 761 131
rect 677 55 717 89
rect 751 55 761 89
rect 677 47 761 55
rect 791 95 857 131
rect 791 61 801 95
rect 835 61 857 95
rect 791 47 857 61
rect 887 153 941 175
rect 887 119 897 153
rect 931 119 941 153
rect 887 47 941 119
rect 971 127 1023 175
rect 971 93 981 127
rect 1015 93 1023 127
rect 971 47 1023 93
rect 1077 93 1129 175
rect 1077 59 1085 93
rect 1119 59 1129 93
rect 1077 47 1129 59
rect 1159 119 1209 175
rect 1583 131 1633 175
rect 1378 119 1428 131
rect 1159 47 1249 119
rect 1279 93 1333 119
rect 1279 59 1289 93
rect 1323 59 1333 93
rect 1279 47 1333 59
rect 1363 47 1428 119
rect 1458 89 1525 131
rect 1458 55 1481 89
rect 1515 55 1525 89
rect 1458 47 1525 55
rect 1555 109 1633 131
rect 1555 75 1565 109
rect 1599 75 1633 109
rect 1555 47 1633 75
rect 1663 167 1717 175
rect 1663 133 1673 167
rect 1707 133 1717 167
rect 1663 47 1717 133
rect 1747 101 1799 175
rect 1950 131 2000 177
rect 1747 67 1757 101
rect 1791 67 1799 101
rect 1747 47 1799 67
rect 1853 103 1905 131
rect 1853 69 1861 103
rect 1895 69 1905 103
rect 1853 47 1905 69
rect 1935 93 2000 131
rect 1935 59 1956 93
rect 1990 59 2000 93
rect 1935 47 2000 59
rect 2030 127 2082 177
rect 2233 131 2283 177
rect 2030 93 2040 127
rect 2074 93 2082 127
rect 2030 47 2082 93
rect 2136 119 2188 131
rect 2136 85 2144 119
rect 2178 85 2188 119
rect 2136 47 2188 85
rect 2218 93 2283 131
rect 2218 59 2239 93
rect 2273 59 2283 93
rect 2218 47 2283 59
rect 2313 129 2365 177
rect 2313 95 2323 129
rect 2357 95 2365 129
rect 2313 47 2365 95
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 413 351 427
rect 381 477 443 497
rect 381 443 391 477
rect 425 443 443 477
rect 381 413 443 443
rect 473 484 527 497
rect 473 450 483 484
rect 517 450 527 484
rect 473 413 527 450
rect 557 413 647 497
rect 677 475 753 497
rect 677 441 697 475
rect 731 441 753 475
rect 677 413 753 441
rect 783 459 861 497
rect 783 425 817 459
rect 851 425 861 459
rect 783 413 861 425
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 799 391 861 413
rect 799 357 817 391
rect 851 357 861 391
rect 799 329 861 357
rect 891 329 945 497
rect 975 485 1082 497
rect 975 451 991 485
rect 1025 451 1082 485
rect 975 417 1082 451
rect 975 383 991 417
rect 1025 383 1082 417
rect 975 329 1082 383
rect 1112 413 1226 497
rect 1256 484 1310 497
rect 1256 450 1266 484
rect 1300 450 1310 484
rect 1256 413 1310 450
rect 1340 413 1415 497
rect 1445 485 1536 497
rect 1445 451 1480 485
rect 1514 451 1536 485
rect 1445 413 1536 451
rect 1566 459 1642 497
rect 1566 425 1588 459
rect 1622 425 1642 459
rect 1566 413 1642 425
rect 1112 329 1164 413
rect 1592 329 1642 413
rect 1672 329 1714 497
rect 1744 485 1796 497
rect 1744 451 1754 485
rect 1788 451 1796 485
rect 1948 485 2000 497
rect 1744 329 1796 451
rect 1948 451 1956 485
rect 1990 451 2000 485
rect 1948 429 2000 451
rect 1850 349 1903 429
rect 1850 315 1858 349
rect 1892 315 1903 349
rect 1850 301 1903 315
rect 1933 301 2000 429
rect 1950 297 2000 301
rect 2030 448 2082 497
rect 2233 481 2283 497
rect 2030 414 2040 448
rect 2074 414 2082 448
rect 2030 380 2082 414
rect 2030 346 2040 380
rect 2074 346 2082 380
rect 2136 467 2188 481
rect 2136 433 2144 467
rect 2178 433 2188 467
rect 2136 399 2188 433
rect 2136 365 2144 399
rect 2178 365 2188 399
rect 2136 353 2188 365
rect 2218 473 2283 481
rect 2218 439 2239 473
rect 2273 439 2283 473
rect 2218 405 2283 439
rect 2218 371 2239 405
rect 2273 371 2283 405
rect 2218 353 2283 371
rect 2030 297 2082 346
rect 2233 297 2283 353
rect 2313 449 2365 497
rect 2313 415 2323 449
rect 2357 415 2365 449
rect 2313 381 2365 415
rect 2313 347 2323 381
rect 2357 347 2365 381
rect 2313 297 2365 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 496 59 530 93
rect 717 55 751 89
rect 801 61 835 95
rect 897 119 931 153
rect 981 93 1015 127
rect 1085 59 1119 93
rect 1289 59 1323 93
rect 1481 55 1515 89
rect 1565 75 1599 109
rect 1673 133 1707 167
rect 1757 67 1791 101
rect 1861 69 1895 103
rect 1956 59 1990 93
rect 2040 93 2074 127
rect 2144 85 2178 119
rect 2239 59 2273 93
rect 2323 95 2357 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 307 427 341 461
rect 391 443 425 477
rect 483 450 517 484
rect 697 441 731 475
rect 817 425 851 459
rect 203 375 237 409
rect 817 357 851 391
rect 991 451 1025 485
rect 991 383 1025 417
rect 1266 450 1300 484
rect 1480 451 1514 485
rect 1588 425 1622 459
rect 1754 451 1788 485
rect 1956 451 1990 485
rect 1858 315 1892 349
rect 2040 414 2074 448
rect 2040 346 2074 380
rect 2144 433 2178 467
rect 2144 365 2178 399
rect 2239 439 2273 473
rect 2239 371 2273 405
rect 2323 415 2357 449
rect 2323 347 2357 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 443 497 473 523
rect 527 497 557 523
rect 647 497 677 523
rect 753 497 783 523
rect 861 497 891 523
rect 945 497 975 523
rect 1082 497 1112 523
rect 1226 497 1256 523
rect 1310 497 1340 523
rect 1415 497 1445 523
rect 1536 497 1566 523
rect 1642 497 1672 523
rect 1714 497 1744 523
rect 2000 497 2030 523
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 117 264 193 274
rect 351 267 381 413
rect 443 279 473 413
rect 527 375 557 413
rect 647 381 677 413
rect 515 365 581 375
rect 515 331 531 365
rect 565 331 581 365
rect 515 321 581 331
rect 647 365 711 381
rect 647 331 667 365
rect 701 331 711 365
rect 647 315 711 331
rect 117 230 133 264
rect 167 230 193 264
rect 117 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 339 251 393 267
rect 339 217 349 251
rect 383 217 393 251
rect 443 249 581 279
rect 339 201 393 217
rect 551 219 581 249
rect 351 131 381 201
rect 446 191 509 207
rect 446 157 465 191
rect 499 157 509 191
rect 446 141 509 157
rect 551 203 605 219
rect 551 169 561 203
rect 595 169 605 203
rect 551 153 605 169
rect 446 119 476 141
rect 551 119 581 153
rect 647 131 677 315
rect 753 229 783 413
rect 1226 381 1256 413
rect 1202 365 1256 381
rect 1310 375 1340 413
rect 1415 381 1445 413
rect 1202 331 1212 365
rect 1246 331 1256 365
rect 861 297 891 329
rect 945 297 975 329
rect 825 281 891 297
rect 825 247 835 281
rect 869 247 891 281
rect 825 231 891 247
rect 941 281 1031 297
rect 941 247 987 281
rect 1021 247 1031 281
rect 941 231 1031 247
rect 1082 263 1112 329
rect 1202 315 1256 331
rect 1298 365 1364 375
rect 1298 331 1314 365
rect 1348 331 1364 365
rect 1298 321 1364 331
rect 1415 365 1494 381
rect 1415 331 1450 365
rect 1484 331 1494 365
rect 1415 315 1494 331
rect 1226 279 1256 315
rect 1082 247 1159 263
rect 1226 249 1363 279
rect 1082 233 1115 247
rect 723 213 783 229
rect 723 179 733 213
rect 767 193 783 213
rect 767 179 791 193
rect 723 163 791 179
rect 857 175 887 231
rect 941 175 971 231
rect 1105 213 1115 233
rect 1149 213 1159 247
rect 1105 197 1159 213
rect 1129 175 1159 197
rect 1237 191 1291 207
rect 761 131 791 163
rect 1237 157 1247 191
rect 1281 157 1291 191
rect 1237 141 1291 157
rect 1249 119 1279 141
rect 1333 119 1363 249
rect 1428 131 1458 315
rect 1536 236 1566 413
rect 1903 429 1933 455
rect 1642 281 1672 329
rect 1501 213 1566 236
rect 1608 265 1672 281
rect 1608 231 1618 265
rect 1652 231 1672 265
rect 1714 297 1744 329
rect 1714 281 1798 297
rect 1714 247 1754 281
rect 1788 247 1798 281
rect 1903 269 1933 301
rect 2188 481 2218 507
rect 2283 497 2313 523
rect 2188 337 2218 353
rect 2163 307 2218 337
rect 1714 231 1798 247
rect 1853 253 1935 269
rect 2000 265 2030 297
rect 1608 215 1672 231
rect 1501 179 1511 213
rect 1545 206 1566 213
rect 1545 179 1555 206
rect 1501 163 1555 179
rect 1633 175 1663 215
rect 1717 175 1747 231
rect 1853 219 1863 253
rect 1897 219 1935 253
rect 1853 203 1935 219
rect 1525 131 1555 163
rect 1905 131 1935 203
rect 1981 259 2035 265
rect 2163 259 2193 307
rect 2283 265 2313 297
rect 1981 249 2193 259
rect 1981 215 1991 249
rect 2025 215 2193 249
rect 1981 205 2193 215
rect 1981 199 2030 205
rect 2000 177 2030 199
rect 2163 176 2193 205
rect 2255 249 2314 265
rect 2255 215 2265 249
rect 2299 215 2314 249
rect 2255 199 2314 215
rect 2283 177 2313 199
rect 2163 146 2218 176
rect 2188 131 2218 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 551 21 581 47
rect 647 21 677 47
rect 761 21 791 47
rect 857 21 887 47
rect 941 21 971 47
rect 1129 21 1159 47
rect 1249 21 1279 47
rect 1333 21 1363 47
rect 1428 21 1458 47
rect 1525 21 1555 47
rect 1633 21 1663 47
rect 1717 21 1747 47
rect 1905 21 1935 47
rect 2000 21 2030 47
rect 2188 21 2218 47
rect 2283 21 2313 47
<< polycont >>
rect 31 230 65 264
rect 531 331 565 365
rect 667 331 701 365
rect 133 230 167 264
rect 349 217 383 251
rect 465 157 499 191
rect 561 169 595 203
rect 1212 331 1246 365
rect 835 247 869 281
rect 987 247 1021 281
rect 1314 331 1348 365
rect 1450 331 1484 365
rect 733 179 767 213
rect 1115 213 1149 247
rect 1247 157 1281 191
rect 1618 231 1652 265
rect 1754 247 1788 281
rect 1511 179 1545 213
rect 1863 219 1897 253
rect 1991 215 2025 249
rect 2265 215 2299 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 247 493
rect 237 443 247 477
rect 203 409 247 443
rect 286 461 357 527
rect 286 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 467 450 483 484
rect 517 450 633 484
rect 69 375 168 393
rect 35 359 168 375
rect 17 264 87 325
rect 17 230 31 264
rect 65 230 87 264
rect 17 195 87 230
rect 122 264 168 359
rect 122 230 133 264
rect 167 230 168 264
rect 122 187 168 230
rect 35 153 122 161
rect 156 153 168 187
rect 35 127 168 153
rect 237 391 247 409
rect 391 393 425 443
rect 203 357 213 375
rect 35 119 69 127
rect 203 119 247 357
rect 281 359 425 393
rect 281 165 315 359
rect 465 357 489 391
rect 523 365 565 391
rect 523 357 531 365
rect 465 331 531 357
rect 349 251 431 325
rect 383 217 431 251
rect 349 201 431 217
rect 465 315 565 331
rect 465 191 509 315
rect 599 281 633 450
rect 681 475 757 527
rect 975 485 1041 527
rect 681 441 697 475
rect 731 441 757 475
rect 817 459 851 475
rect 817 407 851 425
rect 975 451 991 485
rect 1025 451 1041 485
rect 1464 485 1540 527
rect 975 417 1041 451
rect 1250 450 1266 484
rect 1300 450 1416 484
rect 1464 451 1480 485
rect 1514 451 1540 485
rect 1728 485 2006 527
rect 1588 459 1622 475
rect 667 391 937 407
rect 667 365 817 391
rect 701 357 817 365
rect 851 357 937 391
rect 975 383 991 417
rect 1025 383 1041 417
rect 1212 391 1259 397
rect 701 331 717 357
rect 667 315 717 331
rect 819 281 869 297
rect 599 247 835 281
rect 599 239 683 247
rect 281 127 425 165
rect 499 157 509 191
rect 465 141 509 157
rect 545 169 561 203
rect 595 187 615 203
rect 545 153 581 169
rect 545 129 615 153
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 247 119
rect 391 111 425 127
rect 203 69 247 85
rect 103 17 169 59
rect 286 59 307 93
rect 341 59 357 93
rect 649 93 683 239
rect 825 231 869 247
rect 903 213 937 357
rect 1212 365 1225 391
rect 1246 331 1259 357
rect 971 323 1172 331
rect 971 289 1133 323
rect 1167 289 1172 323
rect 1212 315 1259 331
rect 1307 365 1348 381
rect 1307 331 1314 365
rect 971 283 1172 289
rect 971 281 1037 283
rect 971 247 987 281
rect 1021 247 1037 281
rect 1307 261 1348 331
rect 1213 255 1348 261
rect 1099 213 1115 247
rect 1149 213 1165 247
rect 717 179 733 213
rect 767 193 783 213
rect 767 187 799 193
rect 717 153 765 179
rect 903 179 1165 213
rect 1213 221 1225 255
rect 1259 225 1348 255
rect 1382 281 1416 450
rect 1728 451 1754 485
rect 1788 451 1956 485
rect 1990 451 2006 485
rect 1588 417 1622 425
rect 2040 448 2097 493
rect 1450 383 2006 417
rect 1450 365 1500 383
rect 1484 331 1500 365
rect 1450 315 1500 331
rect 1382 265 1652 281
rect 1382 247 1618 265
rect 1259 221 1281 225
rect 1213 212 1281 221
rect 1237 191 1281 212
rect 903 153 947 179
rect 717 147 799 153
rect 881 119 897 153
rect 931 119 947 153
rect 1237 157 1247 191
rect 981 127 1015 143
rect 1237 141 1281 157
rect 391 61 425 77
rect 286 17 357 59
rect 480 59 496 93
rect 530 59 683 93
rect 480 53 683 59
rect 717 89 751 105
rect 717 17 751 55
rect 785 95 851 101
rect 785 61 801 95
rect 835 85 851 95
rect 1382 93 1416 247
rect 1608 231 1618 247
rect 1608 215 1652 231
rect 1456 179 1511 213
rect 1545 187 1565 213
rect 1456 153 1515 179
rect 1549 153 1565 187
rect 1686 168 1720 383
rect 1754 323 1858 349
rect 1754 289 1771 323
rect 1805 315 1858 323
rect 1892 315 1911 349
rect 1805 289 1811 315
rect 1754 281 1811 289
rect 1788 247 1811 281
rect 1972 265 2006 383
rect 2074 414 2097 448
rect 2040 380 2097 414
rect 2074 346 2097 380
rect 2040 326 2097 346
rect 1754 222 1811 247
rect 1767 185 1811 222
rect 1847 253 1938 265
rect 1847 219 1863 253
rect 1897 219 1938 253
rect 1972 249 2025 265
rect 1972 215 1991 249
rect 1972 199 2025 215
rect 1686 167 1723 168
rect 1456 147 1565 153
rect 1643 133 1673 167
rect 1707 133 1723 167
rect 1767 151 1895 185
rect 981 85 1015 93
rect 835 61 1015 85
rect 785 51 1015 61
rect 1065 59 1085 93
rect 1119 59 1135 93
rect 1065 17 1135 59
rect 1260 59 1289 93
rect 1323 59 1416 93
rect 1260 53 1416 59
rect 1450 89 1515 105
rect 1450 55 1481 89
rect 1450 17 1515 55
rect 1549 75 1565 109
rect 1599 85 1615 109
rect 1757 101 1791 117
rect 1599 75 1757 85
rect 1549 67 1757 75
rect 1549 51 1791 67
rect 1853 103 1895 151
rect 1853 69 1861 103
rect 1853 53 1895 69
rect 1945 93 2006 161
rect 2061 143 2097 326
rect 1945 59 1956 93
rect 1990 59 2006 93
rect 1945 17 2006 59
rect 2040 127 2097 143
rect 2074 93 2097 127
rect 2040 51 2097 93
rect 2132 467 2195 483
rect 2132 433 2144 467
rect 2178 433 2195 467
rect 2132 399 2195 433
rect 2132 365 2144 399
rect 2178 365 2195 399
rect 2132 265 2195 365
rect 2231 473 2289 527
rect 2231 439 2239 473
rect 2273 439 2289 473
rect 2231 405 2289 439
rect 2231 371 2239 405
rect 2273 371 2289 405
rect 2231 353 2289 371
rect 2323 449 2375 493
rect 2357 415 2375 449
rect 2323 381 2375 415
rect 2357 347 2375 381
rect 2323 291 2375 347
rect 2132 249 2299 265
rect 2132 215 2265 249
rect 2132 199 2299 215
rect 2132 119 2195 199
rect 2333 165 2375 291
rect 2132 85 2144 119
rect 2178 85 2195 119
rect 2323 129 2375 165
rect 2132 51 2195 85
rect 2230 93 2289 109
rect 2230 59 2239 93
rect 2273 59 2289 93
rect 2230 17 2289 59
rect 2357 95 2375 129
rect 2323 51 2375 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 122 153 156 187
rect 213 375 237 391
rect 237 375 247 391
rect 213 357 247 375
rect 489 357 523 391
rect 581 169 595 187
rect 595 169 615 187
rect 581 153 615 169
rect 1225 365 1259 391
rect 1225 357 1246 365
rect 1246 357 1259 365
rect 1133 289 1167 323
rect 765 179 767 187
rect 767 179 799 187
rect 765 153 799 179
rect 1225 221 1259 255
rect 1515 179 1545 187
rect 1545 179 1549 187
rect 1515 153 1549 179
rect 1771 289 1805 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 477 391 535 397
rect 477 388 489 391
rect 247 360 489 388
rect 247 357 259 360
rect 201 351 259 357
rect 477 357 489 360
rect 523 388 535 391
rect 1213 391 1271 397
rect 1213 388 1225 391
rect 523 360 1225 388
rect 523 357 535 360
rect 477 351 535 357
rect 1213 357 1225 360
rect 1259 357 1271 391
rect 1213 351 1271 357
rect 1121 323 1179 329
rect 1121 289 1133 323
rect 1167 320 1179 323
rect 1759 323 1817 329
rect 1759 320 1771 323
rect 1167 292 1771 320
rect 1167 289 1179 292
rect 1121 283 1179 289
rect 1759 289 1771 292
rect 1805 289 1817 323
rect 1759 283 1817 289
rect 1213 255 1271 261
rect 1213 252 1225 255
rect 584 224 1225 252
rect 584 193 627 224
rect 1213 221 1225 224
rect 1259 221 1271 255
rect 1213 215 1271 221
rect 110 187 168 193
rect 110 153 122 187
rect 156 184 168 187
rect 569 187 627 193
rect 569 184 581 187
rect 156 156 581 184
rect 156 153 168 156
rect 110 147 168 153
rect 569 153 581 156
rect 615 153 627 187
rect 569 147 627 153
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1503 187 1561 193
rect 1503 184 1515 187
rect 799 156 1515 184
rect 799 153 811 156
rect 753 147 811 153
rect 1503 153 1515 156
rect 1549 153 1561 187
rect 1503 147 1561 153
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel locali s 1869 221 1903 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 765 153 799 187 0 FreeSans 400 0 0 0 SET_B
port 4 nsew signal input
flabel locali s 2329 85 2363 119 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2329 357 2363 391 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2329 425 2363 459 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 397 289 431 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2053 425 2087 459 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2053 357 2087 391 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2053 85 2087 119 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 3 FreeSans 400 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 3 FreeSans 400 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dfbbn_1
rlabel locali s 1456 147 1565 213 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1503 184 1561 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1503 147 1561 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 753 184 811 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 753 156 1561 184 1 SET_B
port 4 nsew signal input
rlabel metal1 s 753 147 811 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2392 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_END 3384708
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3365158
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
