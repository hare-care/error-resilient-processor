magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 11 21 643 203
rect 29 -17 63 21
<< locali >>
rect 137 333 203 493
rect 305 333 371 493
rect 473 337 539 493
rect 473 333 627 337
rect 137 299 627 333
rect 21 215 523 265
rect 557 181 627 299
rect 153 145 627 181
rect 153 51 187 145
rect 321 51 355 145
rect 489 51 523 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 26 299 85 527
rect 237 367 271 527
rect 405 367 439 527
rect 573 435 607 527
rect 26 17 79 109
rect 237 17 271 109
rect 405 17 439 109
rect 557 17 607 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 21 215 523 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 11 21 643 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 489 51 523 145 6 Y
port 6 nsew signal output
rlabel locali s 321 51 355 145 6 Y
port 6 nsew signal output
rlabel locali s 153 51 187 145 6 Y
port 6 nsew signal output
rlabel locali s 153 145 627 181 6 Y
port 6 nsew signal output
rlabel locali s 557 181 627 299 6 Y
port 6 nsew signal output
rlabel locali s 137 299 627 333 6 Y
port 6 nsew signal output
rlabel locali s 473 333 627 337 6 Y
port 6 nsew signal output
rlabel locali s 473 337 539 493 6 Y
port 6 nsew signal output
rlabel locali s 305 333 371 493 6 Y
port 6 nsew signal output
rlabel locali s 137 333 203 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2214768
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2208818
<< end >>
