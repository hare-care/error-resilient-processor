VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO dcache_tag_ram
   CLASS BLOCK ;
   SIZE 403.42 BY 378.58 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.7 0.0 76.08 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.54 0.0 81.92 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.38 0.0 87.76 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.22 0.0 93.6 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.06 0.0 99.44 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.9 0.0 105.28 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.74 0.0 111.12 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.58 0.0 116.96 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.42 0.0 122.8 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.26 0.0 128.64 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.1 0.0 134.48 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.94 0.0 140.32 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.78 0.0 146.16 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.62 0.0 152.0 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.46 0.0 157.84 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.3 0.0 163.68 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.14 0.0 169.52 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.98 0.0 175.36 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.82 0.0 181.2 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.66 0.0 187.04 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.5 0.0 192.88 0.38 ;
      END
   END din0[20]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  69.86 0.0 70.24 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 108.68 0.38 109.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 117.18 0.38 117.56 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 122.82 0.38 123.2 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 131.32 0.38 131.7 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.96 0.38 137.34 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 145.46 0.38 145.84 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.1 0.38 151.48 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.34 378.2 327.72 378.58 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  403.04 63.54 403.42 63.92 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  347.09 0.0 347.47 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  342.735 0.0 343.115 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  346.4 0.0 346.78 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  343.425 0.0 343.805 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.115 0.0 344.495 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.86 0.0 345.24 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  403.04 363.33 403.42 363.71 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.26 0.0 30.64 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  372.78 378.2 373.16 378.58 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.425 378.2 136.805 378.58 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.665 378.2 143.045 378.58 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.905 378.2 149.285 378.58 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.145 378.2 155.525 378.58 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.385 378.2 161.765 378.58 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.625 378.2 168.005 378.58 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.865 378.2 174.245 378.58 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.105 378.2 180.485 378.58 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.345 378.2 186.725 378.58 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.585 378.2 192.965 378.58 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.825 378.2 199.205 378.58 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.065 378.2 205.445 378.58 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.305 378.2 211.685 378.58 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.545 378.2 217.925 378.58 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.785 378.2 224.165 378.58 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.025 378.2 230.405 378.58 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.265 378.2 236.645 378.58 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.505 378.2 242.885 378.58 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.745 378.2 249.125 378.58 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  254.985 378.2 255.365 378.58 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  261.225 378.2 261.605 378.58 ;
      END
   END dout1[20]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 378.58 ;
         LAYER met3 ;
         RECT  0.0 0.0 403.42 1.74 ;
         LAYER met4 ;
         RECT  401.68 0.0 403.42 378.58 ;
         LAYER met3 ;
         RECT  0.0 376.84 403.42 378.58 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 375.1 ;
         LAYER met3 ;
         RECT  3.48 3.48 399.94 5.22 ;
         LAYER met3 ;
         RECT  3.48 373.36 399.94 375.1 ;
         LAYER met4 ;
         RECT  398.2 3.48 399.94 375.1 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 402.8 377.96 ;
   LAYER  met2 ;
      RECT  0.62 0.62 402.8 377.96 ;
   LAYER  met3 ;
      RECT  0.98 108.08 402.8 109.66 ;
      RECT  0.62 109.66 0.98 116.58 ;
      RECT  0.62 118.16 0.98 122.22 ;
      RECT  0.62 123.8 0.98 130.72 ;
      RECT  0.62 132.3 0.98 136.36 ;
      RECT  0.62 137.94 0.98 144.86 ;
      RECT  0.62 146.44 0.98 150.5 ;
      RECT  0.98 62.94 402.44 64.52 ;
      RECT  0.98 64.52 402.44 108.08 ;
      RECT  402.44 64.52 402.8 108.08 ;
      RECT  0.62 15.85 0.98 108.08 ;
      RECT  0.98 109.66 402.44 362.73 ;
      RECT  0.98 362.73 402.44 364.31 ;
      RECT  402.44 109.66 402.8 362.73 ;
      RECT  402.44 2.34 402.8 62.94 ;
      RECT  0.62 2.34 0.98 14.27 ;
      RECT  0.62 152.08 0.98 376.24 ;
      RECT  402.44 364.31 402.8 376.24 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 62.94 ;
      RECT  2.88 2.34 400.54 2.88 ;
      RECT  2.88 5.82 400.54 62.94 ;
      RECT  400.54 2.34 402.44 2.88 ;
      RECT  400.54 2.88 402.44 5.82 ;
      RECT  400.54 5.82 402.44 62.94 ;
      RECT  0.98 364.31 2.88 372.76 ;
      RECT  0.98 372.76 2.88 375.7 ;
      RECT  0.98 375.7 2.88 376.24 ;
      RECT  2.88 364.31 400.54 372.76 ;
      RECT  2.88 375.7 400.54 376.24 ;
      RECT  400.54 364.31 402.44 372.76 ;
      RECT  400.54 372.76 402.44 375.7 ;
      RECT  400.54 375.7 402.44 376.24 ;
   LAYER  met4 ;
      RECT  75.1 0.98 76.68 377.96 ;
      RECT  76.68 0.62 80.94 0.98 ;
      RECT  82.52 0.62 86.78 0.98 ;
      RECT  88.36 0.62 92.62 0.98 ;
      RECT  94.2 0.62 98.46 0.98 ;
      RECT  100.04 0.62 104.3 0.98 ;
      RECT  105.88 0.62 110.14 0.98 ;
      RECT  111.72 0.62 115.98 0.98 ;
      RECT  117.56 0.62 121.82 0.98 ;
      RECT  123.4 0.62 127.66 0.98 ;
      RECT  129.24 0.62 133.5 0.98 ;
      RECT  135.08 0.62 139.34 0.98 ;
      RECT  140.92 0.62 145.18 0.98 ;
      RECT  146.76 0.62 151.02 0.98 ;
      RECT  152.6 0.62 156.86 0.98 ;
      RECT  158.44 0.62 162.7 0.98 ;
      RECT  164.28 0.62 168.54 0.98 ;
      RECT  170.12 0.62 174.38 0.98 ;
      RECT  175.96 0.62 180.22 0.98 ;
      RECT  181.8 0.62 186.06 0.98 ;
      RECT  187.64 0.62 191.9 0.98 ;
      RECT  70.84 0.62 75.1 0.98 ;
      RECT  76.68 0.98 326.74 377.6 ;
      RECT  326.74 0.98 328.32 377.6 ;
      RECT  193.48 0.62 342.135 0.98 ;
      RECT  31.24 0.62 69.26 0.98 ;
      RECT  328.32 377.6 372.18 377.96 ;
      RECT  76.68 377.6 135.825 377.96 ;
      RECT  137.405 377.6 142.065 377.96 ;
      RECT  143.645 377.6 148.305 377.96 ;
      RECT  149.885 377.6 154.545 377.96 ;
      RECT  156.125 377.6 160.785 377.96 ;
      RECT  162.365 377.6 167.025 377.96 ;
      RECT  168.605 377.6 173.265 377.96 ;
      RECT  174.845 377.6 179.505 377.96 ;
      RECT  181.085 377.6 185.745 377.96 ;
      RECT  187.325 377.6 191.985 377.96 ;
      RECT  193.565 377.6 198.225 377.96 ;
      RECT  199.805 377.6 204.465 377.96 ;
      RECT  206.045 377.6 210.705 377.96 ;
      RECT  212.285 377.6 216.945 377.96 ;
      RECT  218.525 377.6 223.185 377.96 ;
      RECT  224.765 377.6 229.425 377.96 ;
      RECT  231.005 377.6 235.665 377.96 ;
      RECT  237.245 377.6 241.905 377.96 ;
      RECT  243.485 377.6 248.145 377.96 ;
      RECT  249.725 377.6 254.385 377.96 ;
      RECT  255.965 377.6 260.625 377.96 ;
      RECT  262.205 377.6 326.74 377.96 ;
      RECT  2.34 0.62 29.66 0.98 ;
      RECT  348.07 0.62 401.08 0.98 ;
      RECT  373.76 377.6 401.08 377.96 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 375.7 ;
      RECT  2.34 375.7 2.88 377.96 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 375.7 5.82 377.96 ;
      RECT  5.82 0.98 75.1 2.88 ;
      RECT  5.82 2.88 75.1 375.7 ;
      RECT  5.82 375.7 75.1 377.96 ;
      RECT  328.32 0.98 397.6 2.88 ;
      RECT  328.32 2.88 397.6 375.7 ;
      RECT  328.32 375.7 397.6 377.6 ;
      RECT  397.6 0.98 400.54 2.88 ;
      RECT  397.6 375.7 400.54 377.6 ;
      RECT  400.54 0.98 401.08 2.88 ;
      RECT  400.54 2.88 401.08 375.7 ;
      RECT  400.54 375.7 401.08 377.6 ;
   END
END    dcache_tag_ram
END    LIBRARY
