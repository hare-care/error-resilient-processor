magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 0 0 536 806
<< pmos >>
rect 204 102 240 704
rect 296 102 332 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 692 296 704
rect 240 658 251 692
rect 285 658 296 692
rect 240 624 296 658
rect 240 590 251 624
rect 285 590 296 624
rect 240 556 296 590
rect 240 522 251 556
rect 285 522 296 556
rect 240 488 296 522
rect 240 454 251 488
rect 285 454 296 488
rect 240 420 296 454
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 692 388 704
rect 332 658 343 692
rect 377 658 388 692
rect 332 624 388 658
rect 332 590 343 624
rect 377 590 388 624
rect 332 556 388 590
rect 332 522 343 556
rect 377 522 388 556
rect 332 488 388 522
rect 332 454 343 488
rect 377 454 388 488
rect 332 420 388 454
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 658 285 692
rect 251 590 285 624
rect 251 522 285 556
rect 251 454 285 488
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 658 377 692
rect 343 590 377 624
rect 343 522 377 556
rect 343 454 377 488
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 442 658 500 704
rect 442 624 454 658
rect 488 624 500 658
rect 442 590 500 624
rect 442 556 454 590
rect 488 556 500 590
rect 442 522 500 556
rect 442 488 454 522
rect 488 488 500 522
rect 442 454 500 488
rect 442 420 454 454
rect 488 420 500 454
rect 442 386 500 420
rect 442 352 454 386
rect 488 352 500 386
rect 442 318 500 352
rect 442 284 454 318
rect 488 284 500 318
rect 442 250 500 284
rect 442 216 454 250
rect 488 216 500 250
rect 442 182 500 216
rect 442 148 454 182
rect 488 148 500 182
rect 442 102 500 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 454 624 488 658
rect 454 556 488 590
rect 454 488 488 522
rect 454 420 488 454
rect 454 352 488 386
rect 454 284 488 318
rect 454 216 488 250
rect 454 148 488 182
<< poly >>
rect 167 786 369 806
rect 167 752 183 786
rect 217 752 251 786
rect 285 752 319 786
rect 353 752 369 786
rect 167 736 369 752
rect 204 704 240 736
rect 296 704 332 736
rect 204 70 240 102
rect 296 70 332 102
rect 167 54 369 70
rect 167 20 183 54
rect 217 20 251 54
rect 285 20 319 54
rect 353 20 369 54
rect 167 0 369 20
<< polycont >>
rect 183 752 217 786
rect 251 752 285 786
rect 319 752 353 786
rect 183 20 217 54
rect 251 20 285 54
rect 319 20 353 54
<< locali >>
rect 167 752 179 786
rect 217 752 251 786
rect 285 752 319 786
rect 357 752 369 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 251 692 285 708
rect 251 624 285 638
rect 251 556 285 566
rect 251 488 285 494
rect 251 420 285 422
rect 251 384 285 386
rect 251 312 285 318
rect 251 240 285 250
rect 251 168 285 182
rect 251 98 285 114
rect 343 692 377 708
rect 343 624 377 638
rect 343 556 377 566
rect 343 488 377 494
rect 343 420 377 422
rect 343 384 377 386
rect 343 312 377 318
rect 343 240 377 250
rect 343 168 377 182
rect 454 672 488 674
rect 454 600 488 624
rect 454 528 488 556
rect 454 456 488 488
rect 454 386 488 420
rect 454 318 488 350
rect 454 250 488 278
rect 454 182 488 206
rect 454 132 488 134
rect 343 98 377 114
rect 167 20 179 54
rect 217 20 251 54
rect 285 20 319 54
rect 357 20 369 54
<< viali >>
rect 179 752 183 786
rect 183 752 213 786
rect 251 752 285 786
rect 323 752 353 786
rect 353 752 357 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 251 658 285 672
rect 251 638 285 658
rect 251 590 285 600
rect 251 566 285 590
rect 251 522 285 528
rect 251 494 285 522
rect 251 454 285 456
rect 251 422 285 454
rect 251 352 285 384
rect 251 350 285 352
rect 251 284 285 312
rect 251 278 285 284
rect 251 216 285 240
rect 251 206 285 216
rect 251 148 285 168
rect 251 134 285 148
rect 343 658 377 672
rect 343 638 377 658
rect 343 590 377 600
rect 343 566 377 590
rect 343 522 377 528
rect 343 494 377 522
rect 343 454 377 456
rect 343 422 377 454
rect 343 352 377 384
rect 343 350 377 352
rect 343 284 377 312
rect 343 278 377 284
rect 343 216 377 240
rect 343 206 377 216
rect 343 148 377 168
rect 343 134 377 148
rect 454 658 488 672
rect 454 638 488 658
rect 454 590 488 600
rect 454 566 488 590
rect 454 522 488 528
rect 454 494 488 522
rect 454 454 488 456
rect 454 422 488 454
rect 454 352 488 384
rect 454 350 488 352
rect 454 284 488 312
rect 454 278 488 284
rect 454 216 488 240
rect 454 206 488 216
rect 454 148 488 168
rect 454 134 488 148
rect 179 20 183 54
rect 183 20 213 54
rect 251 20 285 54
rect 323 20 353 54
rect 353 20 357 54
<< metal1 >>
rect 167 786 369 806
rect 167 752 179 786
rect 213 752 251 786
rect 285 752 323 786
rect 357 752 369 786
rect 167 740 369 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 242 678 294 684
rect 242 614 294 626
rect 242 550 294 562
rect 242 494 251 498
rect 285 494 294 498
rect 242 486 294 494
rect 242 422 251 434
rect 285 422 294 434
rect 242 384 294 422
rect 242 350 251 384
rect 285 350 294 384
rect 242 312 294 350
rect 242 278 251 312
rect 285 278 294 312
rect 242 240 294 278
rect 242 206 251 240
rect 285 206 294 240
rect 242 168 294 206
rect 242 134 251 168
rect 285 134 294 168
rect 242 122 294 134
rect 334 672 386 684
rect 334 638 343 672
rect 377 638 386 672
rect 334 600 386 638
rect 334 566 343 600
rect 377 566 386 600
rect 334 528 386 566
rect 334 494 343 528
rect 377 494 386 528
rect 334 456 386 494
rect 334 422 343 456
rect 377 422 386 456
rect 334 384 386 422
rect 334 372 343 384
rect 377 372 386 384
rect 334 312 386 320
rect 334 308 343 312
rect 377 308 386 312
rect 334 244 386 256
rect 334 180 386 192
rect 334 122 386 128
rect 442 672 500 684
rect 442 638 454 672
rect 488 638 500 672
rect 442 600 500 638
rect 442 566 454 600
rect 488 566 500 600
rect 442 528 500 566
rect 442 494 454 528
rect 488 494 500 528
rect 442 456 500 494
rect 442 422 454 456
rect 488 422 500 456
rect 442 384 500 422
rect 442 350 454 384
rect 488 350 500 384
rect 442 312 500 350
rect 442 278 454 312
rect 488 278 500 312
rect 442 240 500 278
rect 442 206 454 240
rect 488 206 500 240
rect 442 168 500 206
rect 442 134 454 168
rect 488 134 500 168
rect 442 122 500 134
rect 167 54 369 66
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
rect 167 0 369 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 242 672 294 678
rect 242 638 251 672
rect 251 638 285 672
rect 285 638 294 672
rect 242 626 294 638
rect 242 600 294 614
rect 242 566 251 600
rect 251 566 285 600
rect 285 566 294 600
rect 242 562 294 566
rect 242 528 294 550
rect 242 498 251 528
rect 251 498 285 528
rect 285 498 294 528
rect 242 456 294 486
rect 242 434 251 456
rect 251 434 285 456
rect 285 434 294 456
rect 334 350 343 372
rect 343 350 377 372
rect 377 350 386 372
rect 334 320 386 350
rect 334 278 343 308
rect 343 278 377 308
rect 377 278 386 308
rect 334 256 386 278
rect 334 240 386 244
rect 334 206 343 240
rect 343 206 377 240
rect 377 206 386 240
rect 334 192 386 206
rect 334 168 386 180
rect 334 134 343 168
rect 343 134 377 168
rect 377 134 386 168
rect 334 128 386 134
<< metal2 >>
rect 10 678 526 684
rect 10 626 242 678
rect 294 626 526 678
rect 10 614 526 626
rect 10 562 242 614
rect 294 562 526 614
rect 10 550 526 562
rect 10 498 242 550
rect 294 498 526 550
rect 10 486 526 498
rect 10 434 242 486
rect 294 434 526 486
rect 10 428 526 434
rect 10 372 526 378
rect 10 320 150 372
rect 202 320 334 372
rect 386 320 526 372
rect 10 308 526 320
rect 10 256 150 308
rect 202 256 334 308
rect 386 256 526 308
rect 10 244 526 256
rect 10 192 150 244
rect 202 192 334 244
rect 386 192 526 244
rect 10 180 526 192
rect 10 128 150 180
rect 202 128 334 180
rect 386 128 526 180
rect 10 122 526 128
<< labels >>
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
port 2 nsew
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
port 3 nsew
flabel metal1 s 167 740 369 806 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 167 0 369 66 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 442 122 500 138 3 FreeSans 300 90 0 0 BULK
port 5 nsew
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 9273642
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9262726
<< end >>
