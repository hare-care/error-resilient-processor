magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 1986 897
<< pwell >>
rect 23 43 1901 317
rect -26 -43 1946 43
<< mvnmos >>
rect 106 141 206 291
rect 314 141 414 291
rect 470 141 570 291
rect 626 141 726 291
rect 782 141 882 291
rect 938 141 1038 291
rect 1094 141 1194 291
rect 1250 141 1350 291
rect 1406 141 1506 291
rect 1562 141 1662 291
rect 1718 141 1818 291
<< mvpmos >>
rect 102 443 202 743
rect 314 443 414 743
rect 470 443 570 743
rect 626 443 726 743
rect 782 443 882 743
rect 938 443 1038 743
rect 1094 443 1194 743
rect 1250 443 1350 743
rect 1406 443 1506 743
rect 1562 443 1662 743
rect 1718 443 1818 743
<< mvndiff >>
rect 49 279 106 291
rect 49 245 57 279
rect 91 245 106 279
rect 49 211 106 245
rect 49 177 57 211
rect 91 177 106 211
rect 49 141 106 177
rect 206 273 314 291
rect 206 239 225 273
rect 259 239 314 273
rect 206 205 314 239
rect 206 171 225 205
rect 259 171 314 205
rect 206 141 314 171
rect 414 264 470 291
rect 414 230 425 264
rect 459 230 470 264
rect 414 196 470 230
rect 414 162 425 196
rect 459 162 470 196
rect 414 141 470 162
rect 570 273 626 291
rect 570 239 581 273
rect 615 239 626 273
rect 570 205 626 239
rect 570 171 581 205
rect 615 171 626 205
rect 570 141 626 171
rect 726 279 782 291
rect 726 245 737 279
rect 771 245 782 279
rect 726 211 782 245
rect 726 177 737 211
rect 771 177 782 211
rect 726 141 782 177
rect 882 273 938 291
rect 882 239 893 273
rect 927 239 938 273
rect 882 205 938 239
rect 882 171 893 205
rect 927 171 938 205
rect 882 141 938 171
rect 1038 279 1094 291
rect 1038 245 1049 279
rect 1083 245 1094 279
rect 1038 211 1094 245
rect 1038 177 1049 211
rect 1083 177 1094 211
rect 1038 141 1094 177
rect 1194 273 1250 291
rect 1194 239 1205 273
rect 1239 239 1250 273
rect 1194 205 1250 239
rect 1194 171 1205 205
rect 1239 171 1250 205
rect 1194 141 1250 171
rect 1350 279 1406 291
rect 1350 245 1361 279
rect 1395 245 1406 279
rect 1350 211 1406 245
rect 1350 177 1361 211
rect 1395 177 1406 211
rect 1350 141 1406 177
rect 1506 273 1562 291
rect 1506 239 1517 273
rect 1551 239 1562 273
rect 1506 205 1562 239
rect 1506 171 1517 205
rect 1551 171 1562 205
rect 1506 141 1562 171
rect 1662 279 1718 291
rect 1662 245 1673 279
rect 1707 245 1718 279
rect 1662 211 1718 245
rect 1662 177 1673 211
rect 1707 177 1718 211
rect 1662 141 1718 177
rect 1818 273 1875 291
rect 1818 239 1833 273
rect 1867 239 1875 273
rect 1818 205 1875 239
rect 1818 171 1833 205
rect 1867 171 1875 205
rect 1818 141 1875 171
<< mvpdiff >>
rect 45 693 102 743
rect 45 659 53 693
rect 87 659 102 693
rect 45 625 102 659
rect 45 591 53 625
rect 87 591 102 625
rect 45 557 102 591
rect 45 523 53 557
rect 87 523 102 557
rect 45 489 102 523
rect 45 455 53 489
rect 87 455 102 489
rect 45 443 102 455
rect 202 731 314 743
rect 202 697 213 731
rect 247 697 314 731
rect 202 663 314 697
rect 202 629 213 663
rect 247 629 314 663
rect 202 595 314 629
rect 202 561 213 595
rect 247 561 314 595
rect 202 527 314 561
rect 202 493 213 527
rect 247 493 314 527
rect 202 443 314 493
rect 414 689 470 743
rect 414 655 425 689
rect 459 655 470 689
rect 414 621 470 655
rect 414 587 425 621
rect 459 587 470 621
rect 414 553 470 587
rect 414 519 425 553
rect 459 519 470 553
rect 414 485 470 519
rect 414 451 425 485
rect 459 451 470 485
rect 414 443 470 451
rect 570 731 626 743
rect 570 697 581 731
rect 615 697 626 731
rect 570 663 626 697
rect 570 629 581 663
rect 615 629 626 663
rect 570 595 626 629
rect 570 561 581 595
rect 615 561 626 595
rect 570 527 626 561
rect 570 493 581 527
rect 615 493 626 527
rect 570 443 626 493
rect 726 689 782 743
rect 726 655 737 689
rect 771 655 782 689
rect 726 621 782 655
rect 726 587 737 621
rect 771 587 782 621
rect 726 553 782 587
rect 726 519 737 553
rect 771 519 782 553
rect 726 485 782 519
rect 726 451 737 485
rect 771 451 782 485
rect 726 443 782 451
rect 882 731 938 743
rect 882 697 893 731
rect 927 697 938 731
rect 882 663 938 697
rect 882 629 893 663
rect 927 629 938 663
rect 882 595 938 629
rect 882 561 893 595
rect 927 561 938 595
rect 882 527 938 561
rect 882 493 893 527
rect 927 493 938 527
rect 882 443 938 493
rect 1038 689 1094 743
rect 1038 655 1049 689
rect 1083 655 1094 689
rect 1038 621 1094 655
rect 1038 587 1049 621
rect 1083 587 1094 621
rect 1038 553 1094 587
rect 1038 519 1049 553
rect 1083 519 1094 553
rect 1038 485 1094 519
rect 1038 451 1049 485
rect 1083 451 1094 485
rect 1038 443 1094 451
rect 1194 731 1250 743
rect 1194 697 1205 731
rect 1239 697 1250 731
rect 1194 663 1250 697
rect 1194 629 1205 663
rect 1239 629 1250 663
rect 1194 595 1250 629
rect 1194 561 1205 595
rect 1239 561 1250 595
rect 1194 527 1250 561
rect 1194 493 1205 527
rect 1239 493 1250 527
rect 1194 443 1250 493
rect 1350 689 1406 743
rect 1350 655 1361 689
rect 1395 655 1406 689
rect 1350 621 1406 655
rect 1350 587 1361 621
rect 1395 587 1406 621
rect 1350 553 1406 587
rect 1350 519 1361 553
rect 1395 519 1406 553
rect 1350 485 1406 519
rect 1350 451 1361 485
rect 1395 451 1406 485
rect 1350 443 1406 451
rect 1506 731 1562 743
rect 1506 697 1517 731
rect 1551 697 1562 731
rect 1506 663 1562 697
rect 1506 629 1517 663
rect 1551 629 1562 663
rect 1506 595 1562 629
rect 1506 561 1517 595
rect 1551 561 1562 595
rect 1506 527 1562 561
rect 1506 493 1517 527
rect 1551 493 1562 527
rect 1506 443 1562 493
rect 1662 689 1718 743
rect 1662 655 1673 689
rect 1707 655 1718 689
rect 1662 621 1718 655
rect 1662 587 1673 621
rect 1707 587 1718 621
rect 1662 553 1718 587
rect 1662 519 1673 553
rect 1707 519 1718 553
rect 1662 485 1718 519
rect 1662 451 1673 485
rect 1707 451 1718 485
rect 1662 443 1718 451
rect 1818 731 1871 743
rect 1818 697 1829 731
rect 1863 697 1871 731
rect 1818 663 1871 697
rect 1818 629 1829 663
rect 1863 629 1871 663
rect 1818 595 1871 629
rect 1818 561 1829 595
rect 1863 561 1871 595
rect 1818 527 1871 561
rect 1818 493 1829 527
rect 1863 493 1871 527
rect 1818 443 1871 493
<< mvndiffc >>
rect 57 245 91 279
rect 57 177 91 211
rect 225 239 259 273
rect 225 171 259 205
rect 425 230 459 264
rect 425 162 459 196
rect 581 239 615 273
rect 581 171 615 205
rect 737 245 771 279
rect 737 177 771 211
rect 893 239 927 273
rect 893 171 927 205
rect 1049 245 1083 279
rect 1049 177 1083 211
rect 1205 239 1239 273
rect 1205 171 1239 205
rect 1361 245 1395 279
rect 1361 177 1395 211
rect 1517 239 1551 273
rect 1517 171 1551 205
rect 1673 245 1707 279
rect 1673 177 1707 211
rect 1833 239 1867 273
rect 1833 171 1867 205
<< mvpdiffc >>
rect 53 659 87 693
rect 53 591 87 625
rect 53 523 87 557
rect 53 455 87 489
rect 213 697 247 731
rect 213 629 247 663
rect 213 561 247 595
rect 213 493 247 527
rect 425 655 459 689
rect 425 587 459 621
rect 425 519 459 553
rect 425 451 459 485
rect 581 697 615 731
rect 581 629 615 663
rect 581 561 615 595
rect 581 493 615 527
rect 737 655 771 689
rect 737 587 771 621
rect 737 519 771 553
rect 737 451 771 485
rect 893 697 927 731
rect 893 629 927 663
rect 893 561 927 595
rect 893 493 927 527
rect 1049 655 1083 689
rect 1049 587 1083 621
rect 1049 519 1083 553
rect 1049 451 1083 485
rect 1205 697 1239 731
rect 1205 629 1239 663
rect 1205 561 1239 595
rect 1205 493 1239 527
rect 1361 655 1395 689
rect 1361 587 1395 621
rect 1361 519 1395 553
rect 1361 451 1395 485
rect 1517 697 1551 731
rect 1517 629 1551 663
rect 1517 561 1551 595
rect 1517 493 1551 527
rect 1673 655 1707 689
rect 1673 587 1707 621
rect 1673 519 1707 553
rect 1673 451 1707 485
rect 1829 697 1863 731
rect 1829 629 1863 663
rect 1829 561 1863 595
rect 1829 493 1863 527
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
<< poly >>
rect 102 743 202 769
rect 314 743 414 769
rect 470 743 570 769
rect 626 743 726 769
rect 782 743 882 769
rect 938 743 1038 769
rect 1094 743 1194 769
rect 1250 743 1350 769
rect 1406 743 1506 769
rect 1562 743 1662 769
rect 1718 743 1818 769
rect 102 413 202 443
rect 314 413 414 443
rect 470 413 570 443
rect 102 363 570 413
rect 102 329 330 363
rect 364 329 570 363
rect 102 313 570 329
rect 106 291 206 313
rect 314 291 414 313
rect 470 291 570 313
rect 626 421 726 443
rect 782 421 882 443
rect 938 421 1038 443
rect 1094 421 1194 443
rect 1250 421 1350 443
rect 1406 421 1506 443
rect 1562 421 1662 443
rect 1718 421 1818 443
rect 626 375 1818 421
rect 626 341 642 375
rect 676 341 1818 375
rect 626 321 1818 341
rect 626 291 726 321
rect 782 291 882 321
rect 938 291 1038 321
rect 1094 291 1194 321
rect 1250 291 1350 321
rect 1406 291 1506 321
rect 1562 291 1662 321
rect 1718 291 1818 321
rect 106 115 206 141
rect 314 115 414 141
rect 470 115 570 141
rect 626 115 726 141
rect 782 115 882 141
rect 938 115 1038 141
rect 1094 115 1194 141
rect 1250 115 1350 141
rect 1406 115 1506 141
rect 1562 115 1662 141
rect 1718 115 1818 141
<< polycont >>
rect 330 329 364 363
rect 642 341 676 375
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 123 731 1901 759
rect 123 729 213 731
rect 247 729 581 731
rect 615 729 893 731
rect 927 729 1205 731
rect 1239 729 1517 731
rect 49 693 87 709
rect 49 659 53 693
rect 49 625 87 659
rect 49 591 53 625
rect 49 557 87 591
rect 49 523 53 557
rect 49 489 87 523
rect 157 695 195 729
rect 247 697 267 729
rect 229 695 267 697
rect 301 695 339 729
rect 373 725 554 729
rect 123 663 373 695
rect 553 695 554 725
rect 615 697 626 729
rect 588 695 626 697
rect 660 725 821 729
rect 660 695 687 725
rect 123 629 213 663
rect 247 629 373 663
rect 123 595 373 629
rect 123 561 213 595
rect 247 561 373 595
rect 123 527 373 561
rect 123 493 213 527
rect 247 493 373 527
rect 123 489 373 493
rect 409 655 425 689
rect 459 655 519 689
rect 409 621 519 655
rect 409 587 425 621
rect 459 587 519 621
rect 409 553 519 587
rect 409 519 425 553
rect 459 519 519 553
rect 49 455 53 489
rect 49 453 87 455
rect 409 485 519 519
rect 409 453 425 485
rect 49 451 425 453
rect 459 451 519 485
rect 553 663 687 695
rect 855 695 893 729
rect 927 695 965 729
rect 999 725 1133 729
rect 553 629 581 663
rect 615 629 687 663
rect 553 595 687 629
rect 553 561 581 595
rect 615 561 687 595
rect 553 527 687 561
rect 553 493 581 527
rect 615 493 687 527
rect 553 477 687 493
rect 721 655 737 689
rect 771 655 787 689
rect 721 621 787 655
rect 721 587 737 621
rect 771 587 787 621
rect 721 553 787 587
rect 721 519 737 553
rect 771 519 787 553
rect 721 485 787 519
rect 49 419 519 451
rect 49 295 87 419
rect 485 391 519 419
rect 721 451 737 485
rect 771 451 787 485
rect 821 663 999 695
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 725 1446 729
rect 821 629 893 663
rect 927 629 999 663
rect 821 595 999 629
rect 821 561 893 595
rect 927 561 999 595
rect 821 527 999 561
rect 821 493 893 527
rect 927 493 999 527
rect 821 477 999 493
rect 1033 655 1049 689
rect 1083 655 1099 689
rect 1033 621 1099 655
rect 1033 587 1049 621
rect 1083 587 1099 621
rect 1033 553 1099 587
rect 1033 519 1049 553
rect 1083 519 1099 553
rect 1033 485 1099 519
rect 721 441 787 451
rect 1033 451 1049 485
rect 1083 451 1099 485
rect 1133 663 1311 695
rect 1445 695 1446 725
rect 1480 697 1517 729
rect 1551 729 1829 731
rect 1863 729 1901 731
rect 1551 697 1589 729
rect 1480 695 1589 697
rect 1623 725 1781 729
rect 1815 697 1829 729
rect 1815 695 1853 697
rect 1887 695 1901 729
rect 1133 629 1205 663
rect 1239 629 1311 663
rect 1133 595 1311 629
rect 1133 561 1205 595
rect 1239 561 1311 595
rect 1133 527 1311 561
rect 1133 493 1205 527
rect 1239 493 1311 527
rect 1133 477 1311 493
rect 1345 655 1361 689
rect 1395 655 1411 689
rect 1345 621 1411 655
rect 1345 587 1361 621
rect 1395 587 1411 621
rect 1345 553 1411 587
rect 1345 519 1361 553
rect 1395 519 1411 553
rect 1345 485 1411 519
rect 1033 441 1099 451
rect 1345 451 1361 485
rect 1395 451 1411 485
rect 1445 663 1623 695
rect 1445 629 1517 663
rect 1551 629 1623 663
rect 1445 595 1623 629
rect 1445 561 1517 595
rect 1551 561 1623 595
rect 1445 527 1623 561
rect 1445 493 1517 527
rect 1551 493 1623 527
rect 1445 477 1623 493
rect 1657 655 1673 689
rect 1707 655 1747 689
rect 1657 646 1747 655
rect 1827 663 1901 695
rect 1657 621 1793 646
rect 1657 587 1673 621
rect 1707 587 1793 621
rect 1657 553 1793 587
rect 1657 519 1673 553
rect 1707 519 1793 553
rect 1657 485 1793 519
rect 1345 441 1411 451
rect 1657 451 1673 485
rect 1707 451 1793 485
rect 1827 629 1829 663
rect 1863 629 1901 663
rect 1827 595 1901 629
rect 1827 561 1829 595
rect 1863 561 1901 595
rect 1827 527 1901 561
rect 1827 493 1829 527
rect 1863 493 1901 527
rect 1827 477 1901 493
rect 1657 441 1793 451
rect 721 424 1793 441
rect 721 391 1124 424
rect 485 375 676 391
rect 127 329 330 363
rect 364 329 449 363
rect 127 316 449 329
rect 485 341 642 375
rect 485 325 676 341
rect 733 390 1124 391
rect 1158 390 1196 424
rect 1230 390 1793 424
rect 733 325 1793 390
rect 49 279 91 295
rect 485 280 519 325
rect 49 245 57 279
rect 49 211 91 245
rect 49 177 57 211
rect 49 161 91 177
rect 135 273 385 277
rect 135 239 225 273
rect 259 239 385 273
rect 135 205 385 239
rect 135 171 225 205
rect 259 171 385 205
rect 135 110 385 171
rect 421 264 519 280
rect 421 230 425 264
rect 459 246 519 264
rect 553 273 699 289
rect 459 230 463 246
rect 421 196 463 230
rect 421 162 425 196
rect 459 162 463 196
rect 421 146 463 162
rect 553 239 581 273
rect 615 239 699 273
rect 553 205 699 239
rect 553 171 581 205
rect 615 171 699 205
rect 553 152 699 171
rect 733 279 775 325
rect 733 245 737 279
rect 771 245 775 279
rect 733 211 775 245
rect 733 177 737 211
rect 771 177 775 211
rect 733 161 775 177
rect 809 273 1011 289
rect 809 239 893 273
rect 927 239 1011 273
rect 809 205 1011 239
rect 809 171 893 205
rect 927 171 1011 205
rect 521 110 699 152
rect 809 110 1011 171
rect 1045 279 1087 325
rect 1045 245 1049 279
rect 1083 245 1087 279
rect 1045 211 1087 245
rect 1045 177 1049 211
rect 1083 177 1087 211
rect 1045 161 1087 177
rect 1121 273 1323 289
rect 1121 239 1205 273
rect 1239 239 1323 273
rect 1121 205 1323 239
rect 1121 171 1205 205
rect 1239 171 1323 205
rect 1121 110 1323 171
rect 1357 279 1399 325
rect 1357 245 1361 279
rect 1395 245 1399 279
rect 1357 211 1399 245
rect 1357 177 1361 211
rect 1395 177 1399 211
rect 1357 161 1399 177
rect 1433 273 1635 289
rect 1433 239 1517 273
rect 1551 239 1635 273
rect 1433 205 1635 239
rect 1433 171 1517 205
rect 1551 171 1635 205
rect 1433 110 1635 171
rect 1669 279 1793 325
rect 1669 245 1673 279
rect 1707 245 1793 279
rect 1669 211 1793 245
rect 1669 177 1673 211
rect 1707 177 1793 211
rect 1669 161 1793 177
rect 1827 273 1901 289
rect 1827 239 1833 273
rect 1867 239 1901 273
rect 1827 205 1901 239
rect 1827 171 1833 205
rect 1867 171 1901 205
rect 1827 120 1901 171
rect 1795 110 1901 120
rect 169 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1867 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 123 695 157 729
rect 195 697 213 729
rect 213 697 229 729
rect 195 695 229 697
rect 267 695 301 729
rect 339 695 373 729
rect 554 697 581 729
rect 581 697 588 729
rect 554 695 588 697
rect 626 695 660 729
rect 821 695 855 729
rect 893 697 927 729
rect 893 695 927 697
rect 965 695 999 729
rect 1133 695 1167 729
rect 1205 697 1239 729
rect 1205 695 1239 697
rect 1277 695 1311 729
rect 1446 695 1480 729
rect 1589 695 1623 729
rect 1781 695 1815 729
rect 1853 697 1863 729
rect 1863 697 1887 729
rect 1853 695 1887 697
rect 1124 390 1158 424
rect 1196 390 1230 424
rect 135 76 169 110
rect 207 76 241 110
rect 279 76 313 110
rect 351 76 385 110
rect 521 76 555 110
rect 593 76 627 110
rect 665 76 699 110
rect 814 76 848 110
rect 886 76 920 110
rect 958 76 992 110
rect 1134 76 1168 110
rect 1206 76 1240 110
rect 1278 76 1312 110
rect 1447 76 1481 110
rect 1519 76 1553 110
rect 1591 76 1625 110
rect 1795 76 1829 110
rect 1867 76 1901 110
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 831 1920 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 0 791 1920 797
rect 0 753 1920 763
rect 0 729 1862 753
rect 0 695 123 729
rect 157 695 195 729
rect 229 695 267 729
rect 301 695 339 729
rect 373 695 554 729
rect 588 695 626 729
rect 660 695 821 729
rect 855 695 893 729
rect 927 695 965 729
rect 999 695 1133 729
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 695 1446 729
rect 1480 695 1589 729
rect 1623 695 1781 729
rect 1815 695 1853 729
rect 1914 701 1926 753
rect 1978 701 1984 753
rect 1887 695 1920 701
rect 0 689 1920 695
rect 1112 381 1120 433
rect 1172 381 1184 433
rect 1236 381 1242 433
rect 0 113 1920 125
rect 0 110 1862 113
rect 0 76 135 110
rect 169 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1862 110
rect 0 61 1862 76
rect 1914 61 1926 113
rect 1978 61 1984 113
rect 0 51 1920 61
rect 0 17 1920 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -23 1920 -17
<< via1 >>
rect 1862 729 1914 753
rect 1862 701 1887 729
rect 1887 701 1914 729
rect 1926 701 1978 753
rect 1120 424 1172 433
rect 1120 390 1124 424
rect 1124 390 1158 424
rect 1158 390 1172 424
rect 1120 381 1172 390
rect 1184 424 1236 433
rect 1184 390 1196 424
rect 1196 390 1230 424
rect 1230 390 1236 424
rect 1184 381 1236 390
rect 1862 110 1914 113
rect 1862 76 1867 110
rect 1867 76 1901 110
rect 1901 76 1914 110
rect 1862 61 1914 76
rect 1926 61 1978 113
<< metal2 >>
rect 1843 701 1852 757
rect 1908 753 1932 757
rect 1914 701 1926 753
rect 1988 701 1997 757
rect 1088 379 1097 435
rect 1153 433 1177 435
rect 1233 433 1242 435
rect 1172 381 1177 433
rect 1236 381 1242 433
rect 1153 379 1177 381
rect 1233 379 1242 381
rect 1843 57 1852 113
rect 1914 61 1926 113
rect 1908 57 1932 61
rect 1988 57 1997 113
<< via2 >>
rect 1852 753 1908 757
rect 1932 753 1988 757
rect 1852 701 1862 753
rect 1862 701 1908 753
rect 1932 701 1978 753
rect 1978 701 1988 753
rect 1097 433 1153 435
rect 1177 433 1233 435
rect 1097 381 1120 433
rect 1120 381 1153 433
rect 1177 381 1184 433
rect 1184 381 1233 433
rect 1097 379 1153 381
rect 1177 379 1233 381
rect 1852 61 1862 113
rect 1862 61 1908 113
rect 1932 61 1978 113
rect 1978 61 1988 113
rect 1852 57 1908 61
rect 1932 57 1988 61
<< metal3 >>
rect 1842 761 1998 762
rect 1842 697 1848 761
rect 1912 697 1928 761
rect 1992 697 1998 761
rect 1842 696 1998 697
rect 1087 439 1243 440
rect 567 375 573 439
rect 637 375 653 439
rect 717 375 723 439
rect 1087 375 1093 439
rect 1157 375 1173 439
rect 1237 375 1243 439
rect 1087 374 1243 375
rect 1842 117 1998 118
rect 1842 53 1848 117
rect 1912 53 1928 117
rect 1992 53 1998 117
rect 1842 52 1998 53
<< via3 >>
rect 1848 757 1912 761
rect 1848 701 1852 757
rect 1852 701 1908 757
rect 1908 701 1912 757
rect 1848 697 1912 701
rect 1928 757 1992 761
rect 1928 701 1932 757
rect 1932 701 1988 757
rect 1988 701 1992 757
rect 1928 697 1992 701
rect 573 375 637 439
rect 653 375 717 439
rect 1093 435 1157 439
rect 1093 379 1097 435
rect 1097 379 1153 435
rect 1153 379 1157 435
rect 1093 375 1157 379
rect 1173 435 1237 439
rect 1173 379 1177 435
rect 1177 379 1233 435
rect 1233 379 1237 435
rect 1173 375 1237 379
rect 1848 113 1912 117
rect 1848 57 1852 113
rect 1852 57 1908 113
rect 1908 57 1912 113
rect 1848 53 1912 57
rect 1928 113 1992 117
rect 1928 57 1932 113
rect 1932 57 1988 113
rect 1988 57 1992 113
rect 1928 53 1992 57
<< via4 >>
rect 1802 761 2038 845
rect 1802 697 1848 761
rect 1848 697 1912 761
rect 1912 697 1928 761
rect 1928 697 1992 761
rect 1992 697 2038 761
rect 1802 609 2038 697
rect 482 439 718 525
rect 482 375 573 439
rect 573 375 637 439
rect 637 375 653 439
rect 653 375 717 439
rect 717 375 718 439
rect 482 289 718 375
rect 1002 439 1238 525
rect 1002 375 1093 439
rect 1093 375 1157 439
rect 1157 375 1173 439
rect 1173 375 1237 439
rect 1237 375 1238 439
rect 1002 289 1238 375
rect 1802 117 2038 205
rect 1802 53 1848 117
rect 1848 53 1912 117
rect 1912 53 1928 117
rect 1928 53 1992 117
rect 1992 53 2038 117
rect 1802 -31 2038 53
<< metal5 >>
rect 942 567 1262 887
rect 1582 845 2082 887
rect 1582 609 1802 845
rect 2038 609 2082 845
rect 1582 567 2082 609
rect 458 525 832 567
rect 458 289 482 525
rect 718 289 832 525
rect 458 247 832 289
rect 852 525 1262 567
rect 852 289 1002 525
rect 1238 289 1262 525
rect 852 247 1262 289
rect 942 -73 1262 247
rect 1582 205 2082 247
rect 1582 -31 1802 205
rect 2038 -31 2082 205
rect 1582 -73 2082 -31
<< rm5 >>
rect 832 247 852 567
<< labels >>
flabel metal3 s 584 375 648 439 0 FreeSans 600 0 0 0 X
port 6 nsew signal output
rlabel comment s 0 0 0 0 4 probec_p_8
flabel metal1 s 0 0 1920 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 1920 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 1920 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 960 802 960 802 0 FreeSans 340 0 0 0 VPB
flabel metal1 s 0 51 1920 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 960 11 960 11 0 FreeSans 340 0 0 0 VNB
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
rlabel metal1 s 1112 381 1242 433 1 X
port 6 nsew signal output
rlabel metal2 s 1088 379 1242 435 1 X
port 6 nsew signal output
rlabel metal3 s 567 375 723 439 1 X
port 6 nsew signal output
rlabel metal3 s 1087 374 1243 440 1 X
port 6 nsew signal output
rlabel metal4 s 482 289 718 525 1 X
port 6 nsew signal output
rlabel metal4 s 1002 289 1238 525 1 X
port 6 nsew signal output
rlabel metal5 s 942 567 1262 887 1 X
port 6 nsew signal output
rlabel metal5 s 942 -73 1262 247 1 X
port 6 nsew signal output
rlabel metal1 s 0 113 1920 125 1 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 61 1984 113 1 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 51 1920 61 1 VGND
port 2 nsew ground bidirectional
rlabel metal2 s 1843 57 1997 113 1 VGND
port 2 nsew ground bidirectional
rlabel metal3 s 1842 52 1998 118 1 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 1802 -31 2038 205 1 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1582 -73 2082 247 1 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 1920 23 1 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 1920 837 1 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 753 1920 763 1 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 0 701 1984 753 1 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 0 689 1920 701 1 VPWR
port 5 nsew power bidirectional
rlabel metal2 s 1843 701 1997 757 1 VPWR
port 5 nsew power bidirectional
rlabel metal3 s 1842 696 1998 762 1 VPWR
port 5 nsew power bidirectional
rlabel metal4 s 1802 609 2038 845 1 VPWR
port 5 nsew power bidirectional
rlabel metal5 s 1582 567 2082 887 1 VPWR
port 5 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 1920 814
string GDS_END 336350
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 313384
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string path 27.800 10.175 31.050 10.175 
<< end >>
