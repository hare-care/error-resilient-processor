magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2013 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 417
rect 271 333 340 417
rect 882 333 948 417
rect 1050 333 1116 417
rect 103 299 1116 333
rect 22 215 337 255
rect 371 181 407 299
rect 441 215 708 255
rect 754 215 1076 255
rect 1218 215 1452 255
rect 1658 215 2007 255
rect 103 131 676 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 18 451 408 493
rect 18 299 69 451
rect 203 367 237 451
rect 374 401 408 451
rect 442 435 508 527
rect 542 401 576 485
rect 610 435 676 527
rect 710 401 760 493
rect 374 367 760 401
rect 798 451 1536 493
rect 798 367 848 451
rect 982 367 1016 451
rect 1150 367 1184 451
rect 1218 333 1284 417
rect 1318 367 1352 451
rect 1386 333 1452 417
rect 1486 367 1536 451
rect 1574 367 1624 527
rect 1658 333 1724 493
rect 1758 367 1792 527
rect 1826 333 1892 493
rect 1218 299 1892 333
rect 1926 299 2007 527
rect 18 93 69 181
rect 710 147 2007 181
rect 710 93 760 147
rect 18 51 760 93
rect 794 17 828 109
rect 862 51 928 147
rect 962 17 1028 109
rect 1062 51 1196 147
rect 1234 17 1268 109
rect 1302 51 1368 147
rect 1402 17 1436 109
rect 1470 51 1608 147
rect 1674 17 1708 109
rect 1742 51 1808 147
rect 1842 17 1894 109
rect 1929 51 2007 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 1658 215 2007 255 6 A1
port 1 nsew signal input
rlabel locali s 1218 215 1452 255 6 A2
port 2 nsew signal input
rlabel locali s 754 215 1076 255 6 A3
port 3 nsew signal input
rlabel locali s 441 215 708 255 6 B1
port 4 nsew signal input
rlabel locali s 22 215 337 255 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 2013 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 131 676 181 6 Y
port 10 nsew signal output
rlabel locali s 371 181 407 299 6 Y
port 10 nsew signal output
rlabel locali s 103 299 1116 333 6 Y
port 10 nsew signal output
rlabel locali s 1050 333 1116 417 6 Y
port 10 nsew signal output
rlabel locali s 882 333 948 417 6 Y
port 10 nsew signal output
rlabel locali s 271 333 340 417 6 Y
port 10 nsew signal output
rlabel locali s 103 333 169 417 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1513622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1497644
<< end >>
