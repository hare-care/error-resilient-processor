magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 140 157 806 203
rect 35 21 806 157
rect 35 17 64 21
rect 30 -17 64 17
<< scnmos >>
rect 121 47 151 131
rect 269 47 299 177
rect 353 47 383 177
rect 449 47 479 177
rect 521 47 551 177
rect 607 47 637 177
rect 693 47 723 177
<< scpmoshvt >>
rect 80 378 110 462
rect 269 297 299 497
rect 353 297 383 497
rect 437 297 467 497
rect 521 297 551 497
rect 607 297 637 497
rect 693 297 723 497
<< ndiff >>
rect 166 161 269 177
rect 166 131 204 161
rect 61 106 121 131
rect 61 72 69 106
rect 103 72 121 106
rect 61 47 121 72
rect 151 127 204 131
rect 238 127 269 161
rect 151 93 269 127
rect 151 59 204 93
rect 238 59 269 93
rect 151 47 269 59
rect 299 169 353 177
rect 299 135 309 169
rect 343 135 353 169
rect 299 101 353 135
rect 299 67 309 101
rect 343 67 353 101
rect 299 47 353 67
rect 383 89 449 177
rect 383 55 404 89
rect 438 55 449 89
rect 383 47 449 55
rect 479 47 521 177
rect 551 157 607 177
rect 551 123 562 157
rect 596 123 607 157
rect 551 89 607 123
rect 551 55 562 89
rect 596 55 607 89
rect 551 47 607 55
rect 637 47 693 177
rect 723 157 780 177
rect 723 123 734 157
rect 768 123 780 157
rect 723 89 780 123
rect 723 55 734 89
rect 768 55 780 89
rect 723 47 780 55
<< pdiff >>
rect 217 477 269 497
rect 27 450 80 462
rect 27 416 35 450
rect 69 416 80 450
rect 27 378 80 416
rect 110 437 163 462
rect 110 403 121 437
rect 155 403 163 437
rect 110 378 163 403
rect 217 443 225 477
rect 259 443 269 477
rect 217 409 269 443
rect 217 375 225 409
rect 259 375 269 409
rect 217 297 269 375
rect 299 407 353 497
rect 299 373 309 407
rect 343 373 353 407
rect 299 339 353 373
rect 299 305 309 339
rect 343 305 353 339
rect 299 297 353 305
rect 383 489 437 497
rect 383 455 393 489
rect 427 455 437 489
rect 383 421 437 455
rect 383 387 393 421
rect 427 387 437 421
rect 383 297 437 387
rect 467 489 521 497
rect 467 455 477 489
rect 511 455 521 489
rect 467 297 521 455
rect 551 477 607 497
rect 551 443 562 477
rect 596 443 607 477
rect 551 405 607 443
rect 551 371 562 405
rect 596 371 607 405
rect 551 297 607 371
rect 637 489 693 497
rect 637 455 648 489
rect 682 455 693 489
rect 637 297 693 455
rect 723 477 780 497
rect 723 443 734 477
rect 768 443 780 477
rect 723 409 780 443
rect 723 375 734 409
rect 768 375 780 409
rect 723 297 780 375
<< ndiffc >>
rect 69 72 103 106
rect 204 127 238 161
rect 204 59 238 93
rect 309 135 343 169
rect 309 67 343 101
rect 404 55 438 89
rect 562 123 596 157
rect 562 55 596 89
rect 734 123 768 157
rect 734 55 768 89
<< pdiffc >>
rect 35 416 69 450
rect 121 403 155 437
rect 225 443 259 477
rect 225 375 259 409
rect 309 373 343 407
rect 309 305 343 339
rect 393 455 427 489
rect 393 387 427 421
rect 477 455 511 489
rect 562 443 596 477
rect 562 371 596 405
rect 648 455 682 489
rect 734 443 768 477
rect 734 375 768 409
<< poly >>
rect 269 497 299 523
rect 353 497 383 523
rect 437 497 467 523
rect 521 497 551 523
rect 607 497 637 523
rect 693 497 723 523
rect 80 462 110 488
rect 80 287 110 378
rect 35 271 110 287
rect 35 237 51 271
rect 85 237 110 271
rect 269 261 299 297
rect 353 261 383 297
rect 437 265 467 297
rect 521 265 551 297
rect 607 265 637 297
rect 35 203 110 237
rect 199 249 383 261
rect 199 215 215 249
rect 249 215 383 249
rect 199 203 383 215
rect 35 169 51 203
rect 85 176 110 203
rect 269 177 299 203
rect 353 177 383 203
rect 425 249 479 265
rect 425 215 435 249
rect 469 215 479 249
rect 425 199 479 215
rect 449 177 479 199
rect 521 249 643 265
rect 521 215 531 249
rect 565 215 599 249
rect 633 215 643 249
rect 521 199 643 215
rect 693 261 723 297
rect 693 249 759 261
rect 693 215 709 249
rect 743 215 759 249
rect 693 203 759 215
rect 521 177 551 199
rect 607 177 637 199
rect 693 177 723 203
rect 85 169 151 176
rect 35 146 151 169
rect 121 131 151 146
rect 121 21 151 47
rect 269 21 299 47
rect 353 21 383 47
rect 449 21 479 47
rect 521 21 551 47
rect 607 21 637 47
rect 693 21 723 47
<< polycont >>
rect 51 237 85 271
rect 215 215 249 249
rect 51 169 85 203
rect 435 215 469 249
rect 531 215 565 249
rect 599 215 633 249
rect 709 215 743 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 19 450 85 527
rect 209 489 443 493
rect 209 477 393 489
rect 19 416 35 450
rect 69 416 85 450
rect 119 437 171 453
rect 119 403 121 437
rect 155 403 171 437
rect 24 271 85 361
rect 24 237 51 271
rect 24 203 85 237
rect 24 169 51 203
rect 24 153 85 169
rect 119 257 171 403
rect 209 443 225 477
rect 259 457 393 477
rect 259 443 270 457
rect 209 409 270 443
rect 377 455 393 457
rect 427 455 443 489
rect 209 375 225 409
rect 259 375 270 409
rect 209 359 270 375
rect 304 407 343 423
rect 304 373 309 407
rect 304 339 343 373
rect 377 421 443 455
rect 477 489 511 527
rect 477 439 511 455
rect 562 477 596 493
rect 632 489 698 527
rect 632 455 648 489
rect 682 455 698 489
rect 732 477 784 493
rect 377 387 393 421
rect 427 405 443 421
rect 562 421 596 443
rect 732 443 734 477
rect 768 443 784 477
rect 732 421 784 443
rect 562 409 784 421
rect 562 405 734 409
rect 427 387 562 405
rect 377 371 562 387
rect 596 375 734 405
rect 768 375 784 409
rect 596 371 784 375
rect 304 305 309 339
rect 119 249 265 257
rect 119 215 215 249
rect 249 215 265 249
rect 119 214 265 215
rect 119 106 159 214
rect 53 72 69 106
rect 103 72 159 106
rect 197 161 245 177
rect 197 127 204 161
rect 238 127 245 161
rect 197 93 245 127
rect 197 59 204 93
rect 238 59 245 93
rect 197 17 245 59
rect 304 169 343 305
rect 420 299 735 335
rect 420 249 485 299
rect 419 215 435 249
rect 469 215 485 249
rect 521 249 643 265
rect 521 215 531 249
rect 565 215 599 249
rect 633 215 643 249
rect 521 199 643 215
rect 677 259 735 299
rect 677 249 759 259
rect 677 215 709 249
rect 743 215 759 249
rect 677 207 759 215
rect 304 135 309 169
rect 727 157 786 173
rect 343 135 562 157
rect 304 123 562 135
rect 596 123 612 157
rect 304 101 344 123
rect 304 67 309 101
rect 343 67 344 101
rect 546 89 612 123
rect 304 51 344 67
rect 388 55 404 89
rect 438 55 454 89
rect 388 17 454 55
rect 546 55 562 89
rect 596 55 612 89
rect 546 51 612 55
rect 727 123 734 157
rect 768 123 786 157
rect 727 89 786 123
rect 727 55 734 89
rect 768 55 786 89
rect 727 17 786 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 30 153 64 187 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 678 289 712 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 310 85 344 119 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
rlabel comment s 0 0 0 0 4 a21boi_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 4016510
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4009878
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 20.700 13.600 
<< end >>
