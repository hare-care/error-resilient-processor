magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 4002 897
rect 3185 343 3698 377
<< pwell >>
rect 1545 283 1967 290
rect 1041 217 1967 283
rect 2408 217 3435 283
rect 3666 217 3932 283
rect 86 43 3932 217
rect -26 -43 3962 43
<< locali >>
rect 113 350 179 444
rect 313 386 395 488
rect 485 350 551 549
rect 113 310 551 350
rect 833 235 935 430
rect 2137 379 2279 424
rect 3243 503 3309 691
rect 3191 405 3309 503
rect 3191 99 3257 405
rect 3844 99 3911 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3936 831
rect 126 735 244 741
rect 126 701 132 735
rect 166 701 204 735
rect 238 701 244 735
rect 22 511 88 603
rect 126 524 244 701
rect 280 619 314 751
rect 350 735 540 751
rect 350 701 356 735
rect 390 701 428 735
rect 462 701 500 735
rect 534 701 540 735
rect 350 667 540 701
rect 576 722 806 756
rect 576 655 642 722
rect 686 619 736 686
rect 280 585 736 619
rect 772 570 806 722
rect 842 727 1228 761
rect 842 606 908 727
rect 998 570 1048 686
rect 22 269 56 511
rect 772 536 1048 570
rect 702 466 1027 500
rect 613 269 666 369
rect 22 235 666 269
rect 108 99 174 235
rect 702 199 736 466
rect 210 113 400 199
rect 210 79 216 113
rect 250 79 288 113
rect 322 79 360 113
rect 394 79 400 113
rect 562 165 736 199
rect 562 99 628 165
rect 772 113 957 199
rect 210 73 400 79
rect 772 79 775 113
rect 809 79 847 113
rect 881 79 919 113
rect 953 79 957 113
rect 772 73 957 79
rect 993 87 1027 466
rect 1084 355 1158 691
rect 1194 657 1228 727
rect 1264 735 1442 751
rect 1298 701 1336 735
rect 1370 701 1408 735
rect 1264 693 1442 701
rect 2107 735 2225 741
rect 2107 701 2113 735
rect 2147 701 2185 735
rect 2219 701 2225 735
rect 1478 657 1887 691
rect 1194 623 1512 657
rect 1194 425 1228 623
rect 1548 571 1731 621
rect 1821 620 1887 657
rect 1548 511 1582 571
rect 1767 550 2071 584
rect 1767 535 1801 550
rect 1264 461 1582 511
rect 1618 497 1801 535
rect 1935 464 2001 514
rect 2037 494 2071 550
rect 2107 530 2225 701
rect 2357 727 2868 761
rect 2263 494 2313 622
rect 1548 427 1757 461
rect 1194 391 1494 425
rect 1063 321 1424 355
rect 1063 123 1129 321
rect 1460 285 1494 391
rect 1165 251 1633 285
rect 1165 87 1199 251
rect 993 53 1199 87
rect 1235 113 1413 215
rect 1449 152 1515 215
rect 1567 188 1633 251
rect 1723 272 1757 427
rect 1814 343 1880 443
rect 1935 343 1969 464
rect 2037 460 2313 494
rect 2037 428 2071 460
rect 2357 441 2423 727
rect 2462 657 2759 691
rect 2005 379 2071 428
rect 2360 343 2426 405
rect 1814 309 2426 343
rect 1723 188 1789 272
rect 1879 152 1945 272
rect 1449 118 1945 152
rect 1269 79 1307 113
rect 1341 79 1379 113
rect 1997 99 2063 309
rect 2360 289 2426 309
rect 2099 253 2165 273
rect 2099 219 2375 253
rect 2462 249 2496 657
rect 2532 441 2598 621
rect 2688 453 2759 657
rect 2802 539 2868 727
rect 2904 735 3085 747
rect 2904 701 2905 735
rect 2939 701 2977 735
rect 3011 701 3049 735
rect 3083 701 3085 735
rect 2904 539 3085 701
rect 3121 727 3379 761
rect 3121 539 3199 727
rect 3121 503 3155 539
rect 2893 453 3155 503
rect 2099 113 2289 183
rect 1235 73 1413 79
rect 2099 79 2105 113
rect 2139 79 2177 113
rect 2211 79 2249 113
rect 2283 79 2289 113
rect 2325 129 2375 219
rect 2430 165 2496 249
rect 2564 417 2598 441
rect 2564 383 3027 417
rect 2564 265 2598 383
rect 2656 301 2722 347
rect 2961 309 3027 383
rect 2564 165 2652 265
rect 2688 129 2722 301
rect 2325 95 2722 129
rect 2783 113 2973 265
rect 2099 73 2289 79
rect 2783 79 2789 113
rect 2823 79 2861 113
rect 2895 79 2933 113
rect 2967 79 2973 113
rect 3063 99 3155 453
rect 3345 367 3379 727
rect 3415 735 3533 741
rect 3415 701 3421 735
rect 3455 701 3493 735
rect 3527 701 3533 735
rect 3415 405 3533 701
rect 3676 735 3794 751
rect 3676 701 3682 735
rect 3716 701 3754 735
rect 3788 701 3794 735
rect 3574 405 3640 563
rect 3676 435 3794 701
rect 3606 367 3640 405
rect 3345 301 3411 367
rect 3606 335 3808 367
rect 3526 301 3808 335
rect 3293 113 3483 265
rect 2783 73 2973 79
rect 3293 79 3299 113
rect 3333 79 3371 113
rect 3405 79 3443 113
rect 3477 79 3483 113
rect 3526 99 3592 301
rect 3628 113 3808 265
rect 3293 73 3483 79
rect 3628 79 3629 113
rect 3663 79 3701 113
rect 3735 79 3773 113
rect 3807 79 3808 113
rect 3628 73 3808 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3936 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 132 701 166 735
rect 204 701 238 735
rect 356 701 390 735
rect 428 701 462 735
rect 500 701 534 735
rect 216 79 250 113
rect 288 79 322 113
rect 360 79 394 113
rect 775 79 809 113
rect 847 79 881 113
rect 919 79 953 113
rect 1264 701 1298 735
rect 1336 701 1370 735
rect 1408 701 1442 735
rect 2113 701 2147 735
rect 2185 701 2219 735
rect 1235 79 1269 113
rect 1307 79 1341 113
rect 1379 79 1413 113
rect 2905 701 2939 735
rect 2977 701 3011 735
rect 3049 701 3083 735
rect 2105 79 2139 113
rect 2177 79 2211 113
rect 2249 79 2283 113
rect 2789 79 2823 113
rect 2861 79 2895 113
rect 2933 79 2967 113
rect 3421 701 3455 735
rect 3493 701 3527 735
rect 3682 701 3716 735
rect 3754 701 3788 735
rect 3299 79 3333 113
rect 3371 79 3405 113
rect 3443 79 3477 113
rect 3629 79 3663 113
rect 3701 79 3735 113
rect 3773 79 3807 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
<< metal1 >>
rect 0 831 3936 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3936 831
rect 0 791 3936 797
rect 0 735 3936 763
rect 0 701 132 735
rect 166 701 204 735
rect 238 701 356 735
rect 390 701 428 735
rect 462 701 500 735
rect 534 701 1264 735
rect 1298 701 1336 735
rect 1370 701 1408 735
rect 1442 701 2113 735
rect 2147 701 2185 735
rect 2219 701 2905 735
rect 2939 701 2977 735
rect 3011 701 3049 735
rect 3083 701 3421 735
rect 3455 701 3493 735
rect 3527 701 3682 735
rect 3716 701 3754 735
rect 3788 701 3936 735
rect 0 689 3936 701
rect 0 113 3936 125
rect 0 79 216 113
rect 250 79 288 113
rect 322 79 360 113
rect 394 79 775 113
rect 809 79 847 113
rect 881 79 919 113
rect 953 79 1235 113
rect 1269 79 1307 113
rect 1341 79 1379 113
rect 1413 79 2105 113
rect 2139 79 2177 113
rect 2211 79 2249 113
rect 2283 79 2789 113
rect 2823 79 2861 113
rect 2895 79 2933 113
rect 2967 79 3299 113
rect 3333 79 3371 113
rect 3405 79 3443 113
rect 3477 79 3629 113
rect 3663 79 3701 113
rect 3735 79 3773 113
rect 3807 79 3936 113
rect 0 51 3936 79
rect 0 17 3936 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3936 17
rect 0 -23 3936 -17
<< obsm1 >>
rect 1075 643 1133 652
rect 2707 643 2765 652
rect 1075 615 2765 643
rect 1075 606 1133 615
rect 2707 606 2765 615
<< labels >>
rlabel locali s 2137 379 2279 424 6 CLK
port 1 nsew clock input
rlabel locali s 833 235 935 430 6 D
port 2 nsew signal input
rlabel locali s 313 386 395 488 6 SCD
port 3 nsew signal input
rlabel locali s 113 310 551 350 6 SCE
port 4 nsew signal input
rlabel locali s 485 350 551 549 6 SCE
port 4 nsew signal input
rlabel locali s 113 350 179 444 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 51 3936 125 6 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 3936 23 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s -26 -43 3962 43 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s 86 43 3932 217 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 3666 217 3932 283 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 2408 217 3435 283 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1041 217 1967 283 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1545 283 1967 290 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 791 3936 837 6 VPB
port 7 nsew power bidirectional
rlabel nwell s 3185 343 3698 377 6 VPB
port 7 nsew power bidirectional
rlabel nwell s -66 377 4002 897 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 689 3936 763 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 3191 99 3257 405 6 Q
port 9 nsew signal output
rlabel locali s 3191 405 3309 503 6 Q
port 9 nsew signal output
rlabel locali s 3243 503 3309 691 6 Q
port 9 nsew signal output
rlabel locali s 3844 99 3911 751 6 Q_N
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3936 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 643078
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 605408
<< end >>
