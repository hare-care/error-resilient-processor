magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 99 201 2483 203
rect 2 23 2483 201
rect 2 21 344 23
rect 614 21 1122 23
rect 2013 21 2483 23
rect 29 -17 63 21
<< locali >>
rect 190 215 268 255
rect 1342 335 1376 357
rect 1322 185 1376 335
rect 1322 151 1387 185
rect 1353 119 1387 151
rect 2402 357 2467 493
rect 2106 215 2195 255
rect 2427 165 2467 357
rect 2399 51 2467 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 402 86 493
rect 120 436 154 527
rect 475 477 708 493
rect 188 459 708 477
rect 745 459 1020 493
rect 188 443 509 459
rect 188 402 222 443
rect 17 368 222 402
rect 256 375 584 409
rect 17 300 88 368
rect 256 334 290 375
rect 122 300 290 334
rect 17 161 51 300
rect 122 265 156 300
rect 85 199 156 265
rect 122 181 156 199
rect 302 187 356 265
rect 17 147 86 161
rect 122 147 265 181
rect 20 51 86 147
rect 126 17 160 109
rect 199 93 265 147
rect 302 153 305 187
rect 339 153 356 187
rect 302 142 356 153
rect 393 127 494 341
rect 528 232 620 323
rect 528 215 595 232
rect 654 185 688 459
rect 745 264 779 459
rect 842 351 876 419
rect 975 413 1020 459
rect 1054 447 1120 527
rect 1167 459 1592 493
rect 1167 413 1201 459
rect 975 379 1201 413
rect 1242 391 1444 425
rect 1242 379 1308 391
rect 1242 345 1276 379
rect 940 277 1036 345
rect 1129 311 1276 345
rect 745 230 819 264
rect 611 181 750 185
rect 528 151 750 181
rect 528 147 632 151
rect 528 131 605 147
rect 648 93 682 117
rect 199 51 682 93
rect 716 85 750 151
rect 785 119 819 230
rect 853 187 903 265
rect 853 153 862 187
rect 896 153 903 187
rect 853 129 903 153
rect 968 199 1036 277
rect 968 102 1006 199
rect 1162 163 1196 311
rect 853 85 919 95
rect 716 51 919 85
rect 1040 17 1106 161
rect 1140 76 1196 163
rect 1230 148 1287 265
rect 1410 246 1444 391
rect 1478 306 1512 425
rect 1558 344 1592 459
rect 1646 459 1990 493
rect 1646 357 1680 459
rect 1924 443 1990 459
rect 2024 455 2091 527
rect 1558 310 1609 344
rect 1714 323 1780 425
rect 1478 272 1524 306
rect 1490 258 1524 272
rect 1410 212 1456 246
rect 1490 221 1540 258
rect 1422 185 1456 212
rect 1422 119 1472 185
rect 1253 85 1319 114
rect 1506 85 1540 221
rect 1575 199 1609 310
rect 1688 306 1780 323
rect 1814 409 1884 425
rect 1814 306 1890 409
rect 1688 289 1748 306
rect 1253 51 1540 85
rect 1587 85 1654 165
rect 1688 153 1722 289
rect 1756 199 1822 255
rect 1688 119 1780 153
rect 1856 85 1890 306
rect 1587 51 1890 85
rect 1930 307 1990 443
rect 2125 409 2167 493
rect 1930 165 1964 307
rect 2038 291 2167 409
rect 2217 291 2283 493
rect 2317 357 2368 527
rect 2038 265 2072 291
rect 1998 199 2072 265
rect 2038 181 2072 199
rect 1930 51 2004 165
rect 2038 147 2184 181
rect 2040 17 2074 113
rect 2108 57 2184 147
rect 2233 136 2283 291
rect 2331 199 2393 323
rect 2233 54 2267 136
rect 2307 17 2365 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 305 153 339 187
rect 862 153 896 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 293 187 351 193
rect 293 153 305 187
rect 339 184 351 187
rect 850 187 908 193
rect 850 184 862 187
rect 339 156 862 184
rect 339 153 351 156
rect 293 147 351 153
rect 850 153 862 156
rect 896 153 908 187
rect 850 147 908 153
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< obsm1 >>
rect 239 388 302 397
rect 830 388 888 397
rect 239 360 888 388
rect 239 351 302 360
rect 830 351 888 360
rect 1839 388 1902 397
rect 2026 388 2084 397
rect 1839 360 2084 388
rect 1839 351 1902 360
rect 2026 351 2084 360
rect 569 320 632 329
rect 942 320 1000 329
rect 569 292 1000 320
rect 569 283 632 292
rect 942 283 1000 292
rect 1678 320 1736 329
rect 2326 320 2384 329
rect 1678 292 2384 320
rect 1678 283 1736 292
rect 2326 283 2384 292
rect 385 252 443 261
rect 1218 252 1276 261
rect 1770 252 1828 261
rect 385 224 1828 252
rect 385 215 443 224
rect 1218 215 1276 224
rect 1770 215 1828 224
rect 1494 184 1552 193
rect 2234 184 2292 193
rect 1494 156 2292 184
rect 1494 147 1552 156
rect 2234 147 2292 156
<< labels >>
rlabel locali s 190 215 268 255 6 A
port 1 nsew signal input
rlabel metal1 s 850 147 908 156 6 B
port 2 nsew signal input
rlabel metal1 s 293 147 351 156 6 B
port 2 nsew signal input
rlabel metal1 s 293 156 908 184 6 B
port 2 nsew signal input
rlabel metal1 s 850 184 908 193 6 B
port 2 nsew signal input
rlabel metal1 s 293 184 351 193 6 B
port 2 nsew signal input
rlabel locali s 2106 215 2195 255 6 CI
port 3 nsew signal input
rlabel metal1 s 0 -48 2484 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2013 21 2483 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 614 21 1122 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2 21 344 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2 23 2483 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 99 201 2483 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2522 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1353 119 1387 151 6 COUT_N
port 8 nsew signal output
rlabel locali s 1322 151 1387 185 6 COUT_N
port 8 nsew signal output
rlabel locali s 1322 185 1376 335 6 COUT_N
port 8 nsew signal output
rlabel locali s 1342 335 1376 357 6 COUT_N
port 8 nsew signal output
rlabel locali s 2399 51 2467 165 6 SUM
port 9 nsew signal output
rlabel locali s 2427 165 2467 357 6 SUM
port 9 nsew signal output
rlabel locali s 2402 357 2467 493 6 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2484 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2151672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2132868
<< end >>
