magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 2082 897
<< pwell >>
rect 1736 281 1994 283
rect 1412 269 1994 281
rect 4 242 418 269
rect 848 242 1994 269
rect 4 43 1994 242
rect -26 -43 2042 43
<< mvnmos >>
rect 89 159 189 243
rect 239 159 339 243
rect 505 132 605 216
rect 661 132 761 216
rect 927 159 1027 243
rect 1069 159 1169 243
rect 1225 159 1325 243
rect 1491 171 1591 255
rect 1647 171 1747 255
rect 1815 107 1915 257
<< mvpmos >>
rect 89 445 189 595
rect 239 445 339 595
rect 505 457 605 607
rect 661 457 761 607
rect 927 457 1027 541
rect 1069 457 1169 541
rect 1225 457 1325 541
rect 1491 443 1591 593
rect 1647 443 1747 593
rect 1815 443 1915 743
<< mvndiff >>
rect 30 218 89 243
rect 30 184 44 218
rect 78 184 89 218
rect 30 159 89 184
rect 189 159 239 243
rect 339 218 392 243
rect 339 184 350 218
rect 384 184 392 218
rect 339 159 392 184
rect 1762 255 1815 257
rect 874 218 927 243
rect 452 191 505 216
rect 452 157 460 191
rect 494 157 505 191
rect 452 132 505 157
rect 605 191 661 216
rect 605 157 616 191
rect 650 157 661 191
rect 605 132 661 157
rect 761 191 814 216
rect 761 157 772 191
rect 806 157 814 191
rect 874 184 882 218
rect 916 184 927 218
rect 874 159 927 184
rect 1027 159 1069 243
rect 1169 205 1225 243
rect 1169 171 1180 205
rect 1214 171 1225 205
rect 1169 159 1225 171
rect 1325 218 1378 243
rect 1325 184 1336 218
rect 1370 184 1378 218
rect 1325 159 1378 184
rect 1438 227 1491 255
rect 1438 193 1446 227
rect 1480 193 1491 227
rect 1438 171 1491 193
rect 1591 171 1647 255
rect 1747 235 1815 255
rect 1747 201 1770 235
rect 1804 201 1815 235
rect 1747 171 1815 201
rect 761 132 814 157
rect 1762 153 1815 171
rect 1762 119 1770 153
rect 1804 119 1815 153
rect 1762 107 1815 119
rect 1915 227 1968 257
rect 1915 193 1926 227
rect 1960 193 1968 227
rect 1915 153 1968 193
rect 1915 119 1926 153
rect 1960 119 1968 153
rect 1915 107 1968 119
<< mvpdiff >>
rect 1762 731 1815 743
rect 452 595 505 607
rect 30 583 89 595
rect 30 549 44 583
rect 78 549 89 583
rect 30 491 89 549
rect 30 457 44 491
rect 78 457 89 491
rect 30 445 89 457
rect 189 445 239 595
rect 339 583 392 595
rect 339 549 350 583
rect 384 549 392 583
rect 339 491 392 549
rect 339 457 350 491
rect 384 457 392 491
rect 452 561 460 595
rect 494 561 505 595
rect 452 503 505 561
rect 452 469 460 503
rect 494 469 505 503
rect 452 457 505 469
rect 605 599 661 607
rect 605 565 616 599
rect 650 565 661 599
rect 605 531 661 565
rect 605 497 616 531
rect 650 497 661 531
rect 605 457 661 497
rect 761 595 814 607
rect 761 561 772 595
rect 806 561 814 595
rect 761 503 814 561
rect 761 469 772 503
rect 806 469 814 503
rect 761 457 814 469
rect 339 445 392 457
rect 1762 697 1770 731
rect 1804 697 1815 731
rect 1762 663 1815 697
rect 1762 629 1770 663
rect 1804 629 1815 663
rect 1762 593 1815 629
rect 1438 581 1491 593
rect 1438 547 1446 581
rect 1480 547 1491 581
rect 874 516 927 541
rect 874 482 882 516
rect 916 482 927 516
rect 874 457 927 482
rect 1027 457 1069 541
rect 1169 516 1225 541
rect 1169 482 1180 516
rect 1214 482 1225 516
rect 1169 457 1225 482
rect 1325 516 1378 541
rect 1325 482 1336 516
rect 1370 482 1378 516
rect 1325 457 1378 482
rect 1438 489 1491 547
rect 1438 455 1446 489
rect 1480 455 1491 489
rect 1438 443 1491 455
rect 1591 575 1647 593
rect 1591 541 1602 575
rect 1636 541 1647 575
rect 1591 489 1647 541
rect 1591 455 1602 489
rect 1636 455 1647 489
rect 1591 443 1647 455
rect 1747 557 1815 593
rect 1747 523 1770 557
rect 1804 523 1815 557
rect 1747 489 1815 523
rect 1747 455 1770 489
rect 1804 455 1815 489
rect 1747 443 1815 455
rect 1915 731 1968 743
rect 1915 697 1926 731
rect 1960 697 1968 731
rect 1915 663 1968 697
rect 1915 629 1926 663
rect 1960 629 1968 663
rect 1915 557 1968 629
rect 1915 523 1926 557
rect 1960 523 1968 557
rect 1915 489 1968 523
rect 1915 455 1926 489
rect 1960 455 1968 489
rect 1915 443 1968 455
<< mvndiffc >>
rect 44 184 78 218
rect 350 184 384 218
rect 460 157 494 191
rect 616 157 650 191
rect 772 157 806 191
rect 882 184 916 218
rect 1180 171 1214 205
rect 1336 184 1370 218
rect 1446 193 1480 227
rect 1770 201 1804 235
rect 1770 119 1804 153
rect 1926 193 1960 227
rect 1926 119 1960 153
<< mvpdiffc >>
rect 44 549 78 583
rect 44 457 78 491
rect 350 549 384 583
rect 350 457 384 491
rect 460 561 494 595
rect 460 469 494 503
rect 616 565 650 599
rect 616 497 650 531
rect 772 561 806 595
rect 772 469 806 503
rect 1770 697 1804 731
rect 1770 629 1804 663
rect 1446 547 1480 581
rect 882 482 916 516
rect 1180 482 1214 516
rect 1336 482 1370 516
rect 1446 455 1480 489
rect 1602 541 1636 575
rect 1602 455 1636 489
rect 1770 523 1804 557
rect 1770 455 1804 489
rect 1926 697 1960 731
rect 1926 629 1960 663
rect 1926 523 1960 557
rect 1926 455 1960 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2016 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
<< poly >>
rect 1815 743 1915 769
rect 829 701 1107 731
rect 239 677 373 693
rect 239 643 255 677
rect 289 643 323 677
rect 357 643 373 677
rect 239 627 373 643
rect 89 595 189 621
rect 239 595 339 627
rect 505 607 605 633
rect 661 607 761 633
rect 89 395 189 445
rect 239 419 339 445
rect 89 361 138 395
rect 172 361 189 395
rect 505 377 605 457
rect 89 327 189 361
rect 89 293 138 327
rect 172 293 189 327
rect 303 361 437 377
rect 303 327 319 361
rect 353 327 387 361
rect 421 327 437 361
rect 303 311 437 327
rect 89 243 189 293
rect 239 243 339 269
rect 89 133 189 159
rect 239 137 339 159
rect 231 121 365 137
rect 231 87 247 121
rect 281 87 315 121
rect 349 87 365 121
rect 231 71 365 87
rect 407 64 437 311
rect 505 343 544 377
rect 578 343 605 377
rect 505 309 605 343
rect 505 275 544 309
rect 578 275 605 309
rect 505 216 605 275
rect 661 442 761 457
rect 829 442 859 701
rect 1077 691 1107 701
rect 1077 675 1713 691
rect 1077 661 1663 675
rect 901 643 1035 659
rect 901 609 917 643
rect 951 609 985 643
rect 1019 609 1035 643
rect 1647 641 1663 661
rect 1697 641 1713 675
rect 1647 619 1713 641
rect 901 593 1035 609
rect 1491 593 1591 619
rect 1647 593 1747 619
rect 927 541 1027 593
rect 1069 541 1169 567
rect 1225 541 1325 567
rect 661 412 859 442
rect 927 431 1027 457
rect 1069 431 1169 457
rect 661 395 761 412
rect 661 361 688 395
rect 722 361 761 395
rect 1103 409 1169 431
rect 661 327 761 361
rect 661 293 688 327
rect 722 293 761 327
rect 661 216 761 293
rect 927 373 1061 389
rect 927 339 943 373
rect 977 339 1011 373
rect 1045 339 1061 373
rect 927 323 1061 339
rect 1103 375 1119 409
rect 1153 375 1169 409
rect 1103 341 1169 375
rect 927 243 1027 323
rect 1103 307 1119 341
rect 1153 307 1169 341
rect 1103 269 1169 307
rect 1069 243 1169 269
rect 1225 315 1325 457
rect 1225 281 1241 315
rect 1275 281 1325 315
rect 1225 243 1325 281
rect 1491 395 1591 443
rect 1491 361 1507 395
rect 1541 361 1591 395
rect 1491 327 1591 361
rect 1491 293 1507 327
rect 1541 293 1591 327
rect 1491 255 1591 293
rect 1647 395 1747 443
rect 1647 361 1686 395
rect 1720 361 1747 395
rect 1647 255 1747 361
rect 1815 345 1915 443
rect 1789 329 1923 345
rect 1789 295 1805 329
rect 1839 295 1873 329
rect 1907 295 1923 329
rect 1789 279 1923 295
rect 1815 257 1915 279
rect 927 133 1027 159
rect 1069 133 1169 159
rect 1225 137 1325 159
rect 1491 145 1591 171
rect 1647 145 1747 171
rect 505 106 605 132
rect 661 106 761 132
rect 1225 121 1382 137
rect 819 99 885 115
rect 819 65 835 99
rect 869 91 885 99
rect 1225 91 1264 121
rect 869 87 1264 91
rect 1298 87 1332 121
rect 1366 87 1382 121
rect 869 71 1382 87
rect 1815 81 1915 107
rect 869 65 1255 71
rect 819 64 1255 65
rect 407 61 1255 64
rect 407 49 885 61
rect 407 34 849 49
<< polycont >>
rect 255 643 289 677
rect 323 643 357 677
rect 138 361 172 395
rect 138 293 172 327
rect 319 327 353 361
rect 387 327 421 361
rect 247 87 281 121
rect 315 87 349 121
rect 544 343 578 377
rect 544 275 578 309
rect 917 609 951 643
rect 985 609 1019 643
rect 1663 641 1697 675
rect 688 361 722 395
rect 688 293 722 327
rect 943 339 977 373
rect 1011 339 1045 373
rect 1119 375 1153 409
rect 1119 307 1153 341
rect 1241 281 1275 315
rect 1507 361 1541 395
rect 1507 293 1541 327
rect 1686 361 1720 395
rect 1805 295 1839 329
rect 1873 295 1907 329
rect 835 65 869 99
rect 1264 87 1298 121
rect 1332 87 1366 121
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2016 831
rect 22 754 666 763
rect 22 729 172 754
rect 22 695 28 729
rect 62 695 100 729
rect 134 720 172 729
rect 206 720 244 754
rect 278 720 316 754
rect 350 720 399 754
rect 433 720 471 754
rect 505 729 666 754
rect 505 720 543 729
rect 134 711 543 720
rect 134 695 205 711
rect 22 689 205 695
rect 533 695 543 711
rect 577 695 615 729
rect 649 695 666 729
rect 1137 757 1892 763
rect 1137 743 1639 757
rect 1137 729 1287 743
rect 533 689 666 695
rect 22 583 88 689
rect 239 643 255 677
rect 289 643 323 677
rect 357 643 499 677
rect 239 633 499 643
rect 22 549 44 583
rect 78 549 88 583
rect 22 491 88 549
rect 22 457 44 491
rect 78 457 88 491
rect 22 440 88 457
rect 334 583 400 599
rect 334 549 350 583
rect 384 549 400 583
rect 334 491 400 549
rect 334 457 350 491
rect 384 457 400 491
rect 122 395 188 440
rect 122 361 138 395
rect 172 361 188 395
rect 334 377 400 457
rect 455 595 499 633
rect 455 561 460 595
rect 494 561 499 595
rect 455 503 499 561
rect 455 469 460 503
rect 494 469 499 503
rect 600 599 666 689
rect 600 565 616 599
rect 650 565 666 599
rect 600 531 666 565
rect 600 497 616 531
rect 650 497 666 531
rect 704 677 1103 711
rect 1137 695 1143 729
rect 1177 695 1215 729
rect 1249 709 1287 729
rect 1321 709 1359 743
rect 1393 729 1639 743
rect 1393 709 1431 729
rect 1249 695 1431 709
rect 1465 695 1503 729
rect 1537 723 1639 729
rect 1673 723 1711 757
rect 1745 731 1892 757
rect 1745 723 1770 731
rect 1804 729 1892 731
rect 1537 695 1613 723
rect 1137 689 1613 695
rect 1754 697 1770 723
rect 1754 695 1783 697
rect 1817 695 1855 729
rect 1889 695 1892 729
rect 1754 689 1892 695
rect 1926 731 1999 747
rect 1960 697 1999 731
rect 455 463 499 469
rect 704 463 738 677
rect 455 429 738 463
rect 772 609 917 643
rect 951 609 985 643
rect 1019 609 1035 643
rect 772 601 1035 609
rect 772 595 814 601
rect 806 561 814 595
rect 772 503 814 561
rect 806 469 814 503
rect 122 327 188 361
rect 122 293 138 327
rect 172 293 188 327
rect 319 361 421 377
rect 353 327 387 361
rect 319 311 421 327
rect 122 277 188 293
rect 28 218 94 234
rect 28 184 44 218
rect 78 184 94 218
rect 28 125 94 184
rect 334 218 400 311
rect 334 184 350 218
rect 384 184 400 218
rect 455 216 494 429
rect 334 168 400 184
rect 444 191 494 216
rect 444 157 460 191
rect 444 141 494 157
rect 528 377 594 393
rect 528 343 544 377
rect 578 343 594 377
rect 528 309 594 343
rect 528 275 544 309
rect 578 275 594 309
rect 672 361 688 395
rect 722 361 738 395
rect 672 327 738 361
rect 672 293 688 327
rect 722 293 738 327
rect 528 259 594 275
rect 772 259 814 469
rect 528 225 814 259
rect 28 119 153 125
rect 28 85 35 119
rect 69 85 107 119
rect 141 85 153 119
rect 28 73 153 85
rect 231 121 373 134
rect 231 87 247 121
rect 281 87 315 121
rect 349 107 373 121
rect 528 107 562 225
rect 764 191 814 225
rect 349 87 562 107
rect 231 73 562 87
rect 596 157 616 191
rect 650 157 666 191
rect 596 125 666 157
rect 764 157 772 191
rect 806 157 814 191
rect 764 141 814 157
rect 875 516 932 532
rect 1069 519 1103 677
rect 875 482 882 516
rect 916 482 932 516
rect 875 466 932 482
rect 1027 485 1103 519
rect 1164 516 1230 689
rect 1430 581 1496 689
rect 1647 675 1720 689
rect 1647 641 1663 675
rect 1697 641 1720 675
rect 1647 625 1720 641
rect 1430 547 1446 581
rect 1480 547 1496 581
rect 875 273 909 466
rect 1027 389 1061 485
rect 1164 482 1180 516
rect 1214 482 1230 516
rect 1164 466 1230 482
rect 1332 516 1386 532
rect 1332 482 1336 516
rect 1370 482 1386 516
rect 1332 417 1386 482
rect 1430 489 1496 547
rect 1430 455 1446 489
rect 1480 455 1496 489
rect 1430 445 1496 455
rect 1591 575 1636 591
rect 1591 541 1602 575
rect 1591 489 1636 541
rect 1591 455 1602 489
rect 943 373 1061 389
rect 977 339 1011 373
rect 1045 339 1061 373
rect 943 323 1061 339
rect 1103 409 1386 417
rect 1103 375 1119 409
rect 1153 375 1386 409
rect 1103 341 1169 375
rect 1103 307 1119 341
rect 1153 307 1169 341
rect 1332 365 1386 375
rect 1491 395 1557 411
rect 1491 365 1507 395
rect 1332 361 1507 365
rect 1541 361 1557 395
rect 1225 315 1298 331
rect 1225 281 1241 315
rect 1275 281 1298 315
rect 1225 273 1298 281
rect 875 239 1298 273
rect 875 218 932 239
rect 875 184 882 218
rect 916 184 932 218
rect 596 119 730 125
rect 596 85 599 119
rect 633 85 671 119
rect 705 107 730 119
rect 875 107 932 184
rect 1164 171 1180 205
rect 1214 171 1230 205
rect 1164 125 1230 171
rect 705 105 785 107
rect 705 85 743 105
rect 596 71 743 85
rect 777 71 785 105
rect 596 51 785 71
rect 819 99 932 107
rect 819 65 835 99
rect 869 65 932 99
rect 819 51 932 65
rect 966 119 1230 125
rect 966 105 1118 119
rect 966 71 974 105
rect 1008 71 1046 105
rect 1080 85 1118 105
rect 1152 85 1190 119
rect 1224 85 1230 119
rect 1080 71 1230 85
rect 1264 134 1298 239
rect 1332 327 1557 361
rect 1332 323 1507 327
rect 1332 218 1386 323
rect 1491 293 1507 323
rect 1541 293 1557 327
rect 1491 277 1557 293
rect 1591 311 1636 455
rect 1670 405 1720 625
rect 1754 663 1820 689
rect 1754 629 1770 663
rect 1804 629 1820 663
rect 1754 557 1820 629
rect 1754 523 1770 557
rect 1804 523 1820 557
rect 1754 489 1820 523
rect 1754 455 1770 489
rect 1804 455 1820 489
rect 1754 439 1820 455
rect 1926 663 1999 697
rect 1960 629 1999 663
rect 1926 557 1999 629
rect 1960 523 1999 557
rect 1926 489 1999 523
rect 1960 455 1999 489
rect 1670 395 1736 405
rect 1670 361 1686 395
rect 1720 361 1736 395
rect 1926 379 1999 455
rect 1670 345 1736 361
rect 1789 329 1911 345
rect 1789 311 1805 329
rect 1591 295 1805 311
rect 1839 295 1873 329
rect 1907 295 1911 329
rect 1591 277 1911 295
rect 1591 243 1636 277
rect 1945 243 1999 379
rect 1332 184 1336 218
rect 1370 184 1386 218
rect 1332 168 1386 184
rect 1430 227 1636 243
rect 1430 193 1446 227
rect 1480 193 1636 227
rect 1430 177 1636 193
rect 1754 235 1820 243
rect 1754 201 1770 235
rect 1804 201 1820 235
rect 1754 153 1820 201
rect 1264 121 1382 134
rect 1754 125 1770 153
rect 1298 87 1332 121
rect 1366 87 1382 121
rect 1264 71 1382 87
rect 1416 119 1770 125
rect 1804 125 1820 153
rect 1926 227 1999 243
rect 1960 193 1999 227
rect 1926 153 1999 193
rect 1804 119 1892 125
rect 1416 105 1708 119
rect 1416 71 1420 105
rect 1454 71 1492 105
rect 1526 71 1564 105
rect 1598 71 1636 105
rect 1670 85 1708 105
rect 1742 85 1780 119
rect 1814 85 1852 119
rect 1886 85 1892 119
rect 1960 119 1999 153
rect 1926 103 1999 119
rect 1670 71 1892 85
rect 966 51 1230 71
rect 1416 51 1892 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 28 695 62 729
rect 100 695 134 729
rect 172 720 206 754
rect 244 720 278 754
rect 316 720 350 754
rect 399 720 433 754
rect 471 720 505 754
rect 543 695 577 729
rect 615 695 649 729
rect 1143 695 1177 729
rect 1215 695 1249 729
rect 1287 709 1321 743
rect 1359 709 1393 743
rect 1431 695 1465 729
rect 1503 695 1537 729
rect 1639 723 1673 757
rect 1711 723 1745 757
rect 1783 697 1804 729
rect 1804 697 1817 729
rect 1783 695 1817 697
rect 1855 695 1889 729
rect 35 85 69 119
rect 107 85 141 119
rect 599 85 633 119
rect 671 85 705 119
rect 743 71 777 105
rect 974 71 1008 105
rect 1046 71 1080 105
rect 1118 85 1152 119
rect 1190 85 1224 119
rect 1420 71 1454 105
rect 1492 71 1526 105
rect 1564 71 1598 105
rect 1636 71 1670 105
rect 1708 85 1742 119
rect 1780 85 1814 119
rect 1852 85 1886 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 831 2016 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2016 831
rect 0 791 2016 797
rect 0 757 2016 763
rect 0 754 1639 757
rect 0 729 172 754
rect 0 695 28 729
rect 62 695 100 729
rect 134 720 172 729
rect 206 720 244 754
rect 278 720 316 754
rect 350 720 399 754
rect 433 720 471 754
rect 505 743 1639 754
rect 505 729 1287 743
rect 505 720 543 729
rect 134 695 543 720
rect 577 695 615 729
rect 649 695 1143 729
rect 1177 695 1215 729
rect 1249 709 1287 729
rect 1321 709 1359 743
rect 1393 729 1639 743
rect 1393 709 1431 729
rect 1249 695 1431 709
rect 1465 695 1503 729
rect 1537 723 1639 729
rect 1673 723 1711 757
rect 1745 729 2016 757
rect 1745 723 1783 729
rect 1537 695 1783 723
rect 1817 695 1855 729
rect 1889 695 2016 729
rect 0 689 2016 695
rect 0 119 2016 125
rect 0 85 35 119
rect 69 85 107 119
rect 141 85 599 119
rect 633 85 671 119
rect 705 105 1118 119
rect 705 85 743 105
rect 0 71 743 85
rect 777 71 974 105
rect 1008 71 1046 105
rect 1080 85 1118 105
rect 1152 85 1190 119
rect 1224 105 1708 119
rect 1224 85 1420 105
rect 1080 71 1420 85
rect 1454 71 1492 105
rect 1526 71 1564 105
rect 1598 71 1636 105
rect 1670 85 1708 105
rect 1742 85 1780 119
rect 1814 85 1852 119
rect 1886 85 2016 119
rect 1670 71 2016 85
rect 0 51 2016 71
rect 0 17 2016 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -23 2016 -17
<< labels >>
flabel comment s 978 303 978 303 0 FreeSans 200 0 0 0 clkneg
flabel comment s 556 234 556 234 0 FreeSans 200 0 0 0 clkpos
flabel comment s 978 446 978 446 0 FreeSans 200 0 0 0 clkpos
rlabel comment s 0 0 0 0 4 dlclkp_1
flabel comment s 474 352 474 352 0 FreeSans 200 90 0 0 clkneg
flabel comment s 290 259 290 259 0 FreeSans 200 0 0 0 clkpos
flabel comment s 786 352 786 352 0 FreeSans 200 90 0 0 clkpos
flabel comment s 290 434 290 434 0 FreeSans 200 0 0 0 clkneg
flabel comment s 629 53 629 53 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 51 2016 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 2016 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 2016 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 2016 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2016 814
string GDS_END 1183864
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1159928
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
