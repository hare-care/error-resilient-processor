magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< pwell >>
rect 10 10 290 392
<< nmoslvt >>
rect 92 36 122 366
rect 178 36 208 366
<< ndiff >>
rect 36 329 92 366
rect 36 295 47 329
rect 81 295 92 329
rect 36 257 92 295
rect 36 223 47 257
rect 81 223 92 257
rect 36 185 92 223
rect 36 151 47 185
rect 81 151 92 185
rect 36 113 92 151
rect 36 79 47 113
rect 81 79 92 113
rect 36 36 92 79
rect 122 329 178 366
rect 122 295 133 329
rect 167 295 178 329
rect 122 257 178 295
rect 122 223 133 257
rect 167 223 178 257
rect 122 185 178 223
rect 122 151 133 185
rect 167 151 178 185
rect 122 113 178 151
rect 122 79 133 113
rect 167 79 178 113
rect 122 36 178 79
rect 208 329 264 366
rect 208 295 219 329
rect 253 295 264 329
rect 208 257 264 295
rect 208 223 219 257
rect 253 223 264 257
rect 208 185 264 223
rect 208 151 219 185
rect 253 151 264 185
rect 208 113 264 151
rect 208 79 219 113
rect 253 79 264 113
rect 208 36 264 79
<< ndiffc >>
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
<< poly >>
rect 83 447 217 463
rect 83 413 99 447
rect 133 413 167 447
rect 201 413 217 447
rect 83 397 217 413
rect 92 392 208 397
rect 92 366 122 392
rect 178 366 208 392
rect 92 10 122 36
rect 178 10 208 36
<< polycont >>
rect 99 413 133 447
rect 167 413 201 447
<< locali >>
rect 83 447 217 463
rect 83 413 97 447
rect 133 413 167 447
rect 203 413 217 447
rect 83 397 217 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 329 167 357
rect 133 257 167 295
rect 133 185 167 223
rect 133 113 167 151
rect 133 51 167 79
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
<< viali >>
rect 97 413 99 447
rect 99 413 131 447
rect 169 413 201 447
rect 201 413 203 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
<< metal1 >>
rect 85 447 215 459
rect 85 413 97 447
rect 131 413 169 447
rect 203 413 215 447
rect 85 401 215 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 124 346 176 357
rect 124 282 176 294
rect 124 223 133 230
rect 167 223 176 230
rect 124 185 176 223
rect 124 151 133 185
rect 167 151 176 185
rect 124 113 176 151
rect 124 79 133 113
rect 167 79 176 113
rect 124 51 176 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 41 -89 259 -29
<< via1 >>
rect 124 329 176 346
rect 124 295 133 329
rect 133 295 167 329
rect 167 295 176 329
rect 124 294 176 295
rect 124 257 176 282
rect 124 230 133 257
rect 133 230 167 257
rect 167 230 176 257
<< metal2 >>
rect 124 346 176 352
rect 124 282 176 294
rect 124 224 176 230
<< labels >>
flabel metal2 s 124 224 176 352 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 41 -89 259 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 85 401 215 459 0 FreeSans 400 0 0 0 GATE
port 4 nsew
flabel pwell s 78 373 88 389 0 FreeSans 200 0 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 5769084
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5764462
string path 1.600 8.925 1.600 -2.225 
<< end >>
