magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1839 203
rect 30 -17 64 21
<< locali >>
rect 103 267 169 483
rect 271 313 337 483
rect 271 267 310 313
rect 103 213 310 267
rect 103 63 169 213
rect 271 165 310 213
rect 271 63 337 165
rect 842 301 1362 335
rect 842 249 876 301
rect 664 215 876 249
rect 910 233 944 265
rect 910 199 1091 233
rect 1125 199 1159 301
rect 1316 265 1362 301
rect 1057 175 1091 199
rect 1057 169 1099 175
rect 1057 165 1107 169
rect 1217 165 1263 265
rect 1316 199 1411 265
rect 1519 317 1553 483
rect 1681 317 1737 483
rect 1519 283 1737 317
rect 1057 146 1263 165
rect 1681 181 1737 283
rect 1059 144 1263 146
rect 1062 142 1263 144
rect 1064 139 1263 142
rect 1067 135 1263 139
rect 1069 131 1263 135
rect 1519 147 1737 181
rect 1519 63 1569 147
rect 1681 63 1737 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 27 299 69 527
rect 203 303 237 527
rect 371 299 473 527
rect 554 387 588 471
rect 638 421 672 527
rect 706 441 866 475
rect 1048 441 1114 527
rect 706 387 740 441
rect 1167 405 1201 471
rect 1235 441 1301 527
rect 1335 405 1369 471
rect 1411 441 1477 527
rect 516 353 740 387
rect 774 371 1479 405
rect 516 249 550 353
rect 774 319 808 371
rect 344 215 550 249
rect 27 17 69 177
rect 203 17 237 177
rect 371 17 419 177
rect 516 163 550 215
rect 584 285 808 319
rect 584 199 618 285
rect 1445 249 1479 371
rect 1587 351 1645 527
rect 1771 299 1813 527
rect 1445 215 1645 249
rect 516 129 609 163
rect 643 129 1023 163
rect 1445 163 1479 215
rect 643 95 677 129
rect 454 61 677 95
rect 711 17 782 93
rect 816 69 850 129
rect 984 117 1023 129
rect 1341 129 1479 163
rect 884 17 950 93
rect 984 51 1038 117
rect 1341 93 1375 129
rect 1077 17 1143 93
rect 1235 59 1375 93
rect 1411 17 1477 93
rect 1603 17 1645 113
rect 1771 17 1813 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
rlabel locali s 1316 199 1411 265 6 A
port 1 nsew signal input
rlabel locali s 1316 265 1362 301 6 A
port 1 nsew signal input
rlabel locali s 1125 199 1159 301 6 A
port 1 nsew signal input
rlabel locali s 664 215 876 249 6 A
port 1 nsew signal input
rlabel locali s 842 249 876 301 6 A
port 1 nsew signal input
rlabel locali s 842 301 1362 335 6 A
port 1 nsew signal input
rlabel locali s 1069 131 1263 135 6 B
port 2 nsew signal input
rlabel locali s 1067 135 1263 139 6 B
port 2 nsew signal input
rlabel locali s 1064 139 1263 142 6 B
port 2 nsew signal input
rlabel locali s 1062 142 1263 144 6 B
port 2 nsew signal input
rlabel locali s 1059 144 1263 146 6 B
port 2 nsew signal input
rlabel locali s 1057 146 1263 165 6 B
port 2 nsew signal input
rlabel locali s 1217 165 1263 265 6 B
port 2 nsew signal input
rlabel locali s 1057 165 1107 169 6 B
port 2 nsew signal input
rlabel locali s 1057 169 1099 175 6 B
port 2 nsew signal input
rlabel locali s 1057 175 1091 199 6 B
port 2 nsew signal input
rlabel locali s 910 199 1091 233 6 B
port 2 nsew signal input
rlabel locali s 910 233 944 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1840 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1839 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1878 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1681 63 1737 147 6 COUT
port 7 nsew signal output
rlabel locali s 1519 63 1569 147 6 COUT
port 7 nsew signal output
rlabel locali s 1519 147 1737 181 6 COUT
port 7 nsew signal output
rlabel locali s 1681 181 1737 283 6 COUT
port 7 nsew signal output
rlabel locali s 1519 283 1737 317 6 COUT
port 7 nsew signal output
rlabel locali s 1681 317 1737 483 6 COUT
port 7 nsew signal output
rlabel locali s 1519 317 1553 483 6 COUT
port 7 nsew signal output
rlabel locali s 271 63 337 165 6 SUM
port 8 nsew signal output
rlabel locali s 271 165 310 213 6 SUM
port 8 nsew signal output
rlabel locali s 103 63 169 213 6 SUM
port 8 nsew signal output
rlabel locali s 103 213 310 267 6 SUM
port 8 nsew signal output
rlabel locali s 271 267 310 313 6 SUM
port 8 nsew signal output
rlabel locali s 271 313 337 483 6 SUM
port 8 nsew signal output
rlabel locali s 103 267 169 483 6 SUM
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2190846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2176828
<< end >>
