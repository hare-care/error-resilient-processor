magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 975 203
rect 30 -17 64 21
<< locali >>
rect 459 349 493 425
rect 627 349 661 425
rect 459 289 661 349
rect 72 215 360 255
rect 459 181 525 289
rect 889 215 995 264
rect 107 145 677 181
rect 107 51 173 145
rect 275 51 341 145
rect 443 51 509 145
rect 611 51 677 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 333 73 493
rect 107 367 173 527
rect 207 333 241 493
rect 275 367 325 527
rect 359 459 771 493
rect 359 333 425 459
rect 17 291 425 333
rect 527 387 593 459
rect 695 315 771 459
rect 805 315 871 493
rect 805 255 855 315
rect 905 299 986 527
rect 559 215 855 255
rect 17 17 73 181
rect 207 17 241 111
rect 375 17 409 111
rect 543 17 577 111
rect 711 17 769 181
rect 805 163 855 215
rect 805 51 871 163
rect 905 17 963 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 72 215 360 255 6 A
port 1 nsew signal input
rlabel locali s 889 215 995 264 6 B_N
port 2 nsew signal input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 975 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 611 51 677 145 6 Y
port 7 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 7 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 7 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 7 nsew signal output
rlabel locali s 107 145 677 181 6 Y
port 7 nsew signal output
rlabel locali s 459 181 525 289 6 Y
port 7 nsew signal output
rlabel locali s 459 289 661 349 6 Y
port 7 nsew signal output
rlabel locali s 627 349 661 425 6 Y
port 7 nsew signal output
rlabel locali s 459 349 493 425 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1999856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1991350
<< end >>
