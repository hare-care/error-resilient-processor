magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -36 679 294 1471
<< poly >>
rect 114 721 144 1113
rect 48 705 144 721
rect 48 671 64 705
rect 98 671 144 705
rect 48 655 144 671
rect 114 225 144 655
<< polycont >>
rect 64 671 98 705
<< locali >>
rect 0 1397 258 1431
rect 62 1218 96 1397
rect 64 705 98 721
rect 64 655 98 671
rect 162 705 196 1284
rect 162 671 213 705
rect 162 92 196 671
rect 62 17 96 92
rect 0 -17 258 17
use contact_12  contact_12_0
timestamp 1694700623
transform 1 0 48 0 1 655
box 0 0 1 1
use nmos_m2_w0_740_sli_dli_da_p  nmos_m2_w0_740_sli_dli_da_p_0
timestamp 1694700623
transform 1 0 54 0 1 51
box -26 -26 176 174
use pmos_m2_w1_120_sli_dli_da_p  pmos_m2_w1_120_sli_dli_da_p_0
timestamp 1694700623
transform 1 0 54 0 1 1139
box -59 -54 209 278
<< labels >>
rlabel locali s 196 688 196 688 4 Z
port 2 nsew
rlabel locali s 81 688 81 688 4 A
port 1 nsew
rlabel locali s 129 1414 129 1414 4 vdd
port 3 nsew
rlabel locali s 129 0 129 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 258 1414
string GDS_END 4082448
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4081054
<< end >>
