magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 269 163 545 203
rect 4 27 545 163
rect 29 -17 63 27
rect 269 21 545 27
<< locali >>
rect 17 425 256 483
rect 121 265 166 323
rect 388 299 443 493
rect 17 199 87 265
rect 121 199 286 265
rect 409 152 443 299
rect 388 83 443 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 21 357 254 391
rect 290 367 346 527
rect 21 299 87 357
rect 220 333 254 357
rect 220 299 354 333
rect 320 265 354 299
rect 320 199 375 265
rect 320 165 354 199
rect 21 131 354 165
rect 477 286 535 527
rect 21 61 72 131
rect 106 17 172 97
rect 206 61 240 131
rect 274 17 350 97
rect 477 17 535 183
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 121 199 286 265 6 A
port 1 nsew signal input
rlabel locali s 121 265 166 323 6 A
port 1 nsew signal input
rlabel locali s 17 425 256 483 6 B
port 2 nsew signal input
rlabel locali s 17 199 87 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 269 21 545 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 -17 63 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 4 27 545 163 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 269 163 545 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 388 83 443 152 6 X
port 8 nsew signal output
rlabel locali s 409 152 443 299 6 X
port 8 nsew signal output
rlabel locali s 388 299 443 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1022512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1016898
<< end >>
