magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 4 43 668 299
rect -26 -43 698 43
<< locali >>
rect 489 391 562 508
rect 596 425 647 751
rect 103 301 261 350
rect 455 325 573 391
rect 489 232 562 325
rect 607 291 647 425
rect 596 115 647 291
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 166 735 560 751
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 35 420 130 601
rect 166 542 560 701
rect 166 456 455 542
rect 35 386 413 420
rect 35 267 69 386
rect 295 345 413 386
rect 35 181 76 267
rect 110 198 455 267
rect 110 147 560 198
rect 94 113 560 147
rect 128 79 166 113
rect 200 79 238 113
rect 272 79 310 113
rect 344 79 382 113
rect 416 79 454 113
rect 488 79 526 113
rect 94 73 560 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 166 701 200 735
rect 238 701 272 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 94 79 128 113
rect 166 79 200 113
rect 238 79 272 113
rect 310 79 344 113
rect 382 79 416 113
rect 454 79 488 113
rect 526 79 560 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 166 735
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 94 113
rect 128 79 166 113
rect 200 79 238 113
rect 272 79 310 113
rect 344 79 382 113
rect 416 79 454 113
rect 488 79 526 113
rect 560 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel locali s 489 232 562 325 6 A
port 1 nsew signal input
rlabel locali s 455 325 573 391 6 A
port 1 nsew signal input
rlabel locali s 489 391 562 508 6 A
port 1 nsew signal input
rlabel locali s 103 301 261 350 6 TE
port 2 nsew signal input
rlabel metal1 s 0 51 672 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 672 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 698 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 668 299 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 672 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 738 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 672 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 596 115 647 291 6 Z
port 7 nsew signal output
rlabel locali s 607 291 647 425 6 Z
port 7 nsew signal output
rlabel locali s 596 425 647 751 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1239596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1230040
<< end >>
