magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -36 538 512 1177
<< locali >>
rect 0 1103 476 1137
rect 64 501 98 567
rect 183 517 217 551
rect 0 -17 476 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_0
timestamp 1694700623
transform 1 0 0 0 1 0
box -36 -17 512 1177
<< labels >>
rlabel locali s 200 534 200 534 4 Z
rlabel locali s 81 534 81 534 4 A
rlabel locali s 238 0 238 0 4 gnd
rlabel locali s 238 1120 238 1120 4 vdd
<< properties >>
string FIXED_BBOX 0 0 476 1120
string GDS_END 64592
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 63764
<< end >>
