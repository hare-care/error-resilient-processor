magic
tech sky130B
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_0
timestamp 1694700623
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_1
timestamp 1694700623
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_2
timestamp 1694700623
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_1
timestamp 1694700623
transform 1 0 648 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 39943716
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39940852
<< end >>
