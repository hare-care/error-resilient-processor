magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1287 203
rect 29 -17 63 21
<< locali >>
rect 196 340 232 493
rect 368 340 406 493
rect 17 287 406 340
rect 17 161 73 287
rect 508 289 856 337
rect 508 199 566 289
rect 611 207 748 255
rect 790 207 856 289
rect 898 299 1258 337
rect 898 207 969 299
rect 1006 207 1141 265
rect 1178 207 1258 299
rect 17 127 321 161
rect 119 123 321 127
rect 119 51 153 123
rect 287 51 321 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 96 374 162 527
rect 268 374 334 527
rect 440 440 506 527
rect 540 405 612 493
rect 657 439 723 527
rect 757 405 824 493
rect 858 439 911 527
rect 1031 405 1097 493
rect 440 371 1097 405
rect 1203 383 1269 527
rect 440 253 474 371
rect 107 213 474 253
rect 440 163 474 213
rect 440 127 704 163
rect 834 139 1269 173
rect 19 17 85 93
rect 187 17 253 89
rect 834 93 900 139
rect 355 17 428 93
rect 466 51 900 93
rect 934 17 997 105
rect 1031 51 1097 139
rect 1131 17 1169 105
rect 1203 51 1269 139
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 1178 207 1258 299 6 A1
port 1 nsew signal input
rlabel locali s 898 207 969 299 6 A1
port 1 nsew signal input
rlabel locali s 898 299 1258 337 6 A1
port 1 nsew signal input
rlabel locali s 1006 207 1141 265 6 A2
port 2 nsew signal input
rlabel locali s 790 207 856 289 6 B1
port 3 nsew signal input
rlabel locali s 508 199 566 289 6 B1
port 3 nsew signal input
rlabel locali s 508 289 856 337 6 B1
port 3 nsew signal input
rlabel locali s 611 207 748 255 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1287 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 287 51 321 123 6 X
port 9 nsew signal output
rlabel locali s 119 51 153 123 6 X
port 9 nsew signal output
rlabel locali s 119 123 321 127 6 X
port 9 nsew signal output
rlabel locali s 17 127 321 161 6 X
port 9 nsew signal output
rlabel locali s 17 161 73 287 6 X
port 9 nsew signal output
rlabel locali s 17 287 406 340 6 X
port 9 nsew signal output
rlabel locali s 368 340 406 493 6 X
port 9 nsew signal output
rlabel locali s 196 340 232 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 770896
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 761900
<< end >>
