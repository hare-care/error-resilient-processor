magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< pwell >>
rect -1566 -5162 1566 5162
<< mvpsubdiff >>
rect -1540 5124 1540 5136
rect -1540 5090 -1351 5124
rect -1317 5090 -1283 5124
rect -1249 5090 -1215 5124
rect -1181 5090 -1147 5124
rect -1113 5090 -735 5124
rect -701 5090 -667 5124
rect -633 5090 -599 5124
rect -565 5090 -531 5124
rect -497 5090 -119 5124
rect -85 5090 -51 5124
rect -17 5090 17 5124
rect 51 5090 85 5124
rect 119 5090 497 5124
rect 531 5090 565 5124
rect 599 5090 633 5124
rect 667 5090 701 5124
rect 735 5090 1113 5124
rect 1147 5090 1181 5124
rect 1215 5090 1249 5124
rect 1283 5090 1317 5124
rect 1351 5090 1540 5124
rect -1540 5078 1540 5090
rect -1540 5015 -1410 5078
rect -1540 -5015 -1524 5015
rect -1422 -5015 -1410 5015
rect -1054 5015 -794 5078
rect -1054 4981 -1042 5015
rect -1008 4981 -946 5015
rect -912 4981 -840 5015
rect -806 4981 -794 5015
rect -438 5015 -178 5078
rect -1054 4947 -794 4981
rect -1054 4913 -1042 4947
rect -1008 4913 -946 4947
rect -912 4913 -840 4947
rect -806 4913 -794 4947
rect -1054 4879 -794 4913
rect -1054 4845 -1042 4879
rect -1008 4845 -946 4879
rect -912 4845 -840 4879
rect -806 4845 -794 4879
rect -1054 4811 -794 4845
rect -1054 4777 -1042 4811
rect -1008 4777 -946 4811
rect -912 4777 -840 4811
rect -806 4777 -794 4811
rect -1054 4743 -794 4777
rect -1054 4709 -1042 4743
rect -1008 4709 -946 4743
rect -912 4709 -840 4743
rect -806 4709 -794 4743
rect -1054 4675 -794 4709
rect -1054 4641 -1042 4675
rect -1008 4641 -946 4675
rect -912 4641 -840 4675
rect -806 4641 -794 4675
rect -1054 4607 -794 4641
rect -1054 4573 -1042 4607
rect -1008 4573 -946 4607
rect -912 4573 -840 4607
rect -806 4573 -794 4607
rect -1054 4539 -794 4573
rect -1054 4505 -1042 4539
rect -1008 4505 -946 4539
rect -912 4505 -840 4539
rect -806 4505 -794 4539
rect -1054 4471 -794 4505
rect -1054 4437 -1042 4471
rect -1008 4437 -946 4471
rect -912 4437 -840 4471
rect -806 4437 -794 4471
rect -1054 4403 -794 4437
rect -1054 4369 -1042 4403
rect -1008 4369 -946 4403
rect -912 4369 -840 4403
rect -806 4369 -794 4403
rect -1054 4335 -794 4369
rect -1054 4301 -1042 4335
rect -1008 4301 -946 4335
rect -912 4301 -840 4335
rect -806 4301 -794 4335
rect -1054 4267 -794 4301
rect -1054 4233 -1042 4267
rect -1008 4233 -946 4267
rect -912 4233 -840 4267
rect -806 4233 -794 4267
rect -1054 4199 -794 4233
rect -1054 4165 -1042 4199
rect -1008 4165 -946 4199
rect -912 4165 -840 4199
rect -806 4165 -794 4199
rect -1054 4131 -794 4165
rect -1054 4097 -1042 4131
rect -1008 4097 -946 4131
rect -912 4097 -840 4131
rect -806 4097 -794 4131
rect -1054 4063 -794 4097
rect -1054 4029 -1042 4063
rect -1008 4029 -946 4063
rect -912 4029 -840 4063
rect -806 4029 -794 4063
rect -1054 3995 -794 4029
rect -1054 3961 -1042 3995
rect -1008 3961 -946 3995
rect -912 3961 -840 3995
rect -806 3961 -794 3995
rect -1054 3927 -794 3961
rect -1054 3893 -1042 3927
rect -1008 3893 -946 3927
rect -912 3893 -840 3927
rect -806 3893 -794 3927
rect -1054 3859 -794 3893
rect -1054 3825 -1042 3859
rect -1008 3825 -946 3859
rect -912 3825 -840 3859
rect -806 3825 -794 3859
rect -1054 3791 -794 3825
rect -1054 3757 -1042 3791
rect -1008 3757 -946 3791
rect -912 3757 -840 3791
rect -806 3757 -794 3791
rect -1054 3723 -794 3757
rect -1054 3689 -1042 3723
rect -1008 3689 -946 3723
rect -912 3689 -840 3723
rect -806 3689 -794 3723
rect -1054 3655 -794 3689
rect -1054 3621 -1042 3655
rect -1008 3621 -946 3655
rect -912 3621 -840 3655
rect -806 3621 -794 3655
rect -1054 3587 -794 3621
rect -1054 3553 -1042 3587
rect -1008 3553 -946 3587
rect -912 3553 -840 3587
rect -806 3553 -794 3587
rect -1054 3519 -794 3553
rect -1054 3485 -1042 3519
rect -1008 3485 -946 3519
rect -912 3485 -840 3519
rect -806 3485 -794 3519
rect -1054 3451 -794 3485
rect -1054 3417 -1042 3451
rect -1008 3417 -946 3451
rect -912 3417 -840 3451
rect -806 3417 -794 3451
rect -1054 3383 -794 3417
rect -1054 3349 -1042 3383
rect -1008 3349 -946 3383
rect -912 3349 -840 3383
rect -806 3349 -794 3383
rect -1054 3315 -794 3349
rect -1054 3281 -1042 3315
rect -1008 3281 -946 3315
rect -912 3281 -840 3315
rect -806 3281 -794 3315
rect -1054 3247 -794 3281
rect -1054 3213 -1042 3247
rect -1008 3213 -946 3247
rect -912 3213 -840 3247
rect -806 3213 -794 3247
rect -1054 3179 -794 3213
rect -1054 3145 -1042 3179
rect -1008 3145 -946 3179
rect -912 3145 -840 3179
rect -806 3145 -794 3179
rect -1054 3111 -794 3145
rect -1054 3077 -1042 3111
rect -1008 3077 -946 3111
rect -912 3077 -840 3111
rect -806 3077 -794 3111
rect -1054 3043 -794 3077
rect -1054 3009 -1042 3043
rect -1008 3009 -946 3043
rect -912 3009 -840 3043
rect -806 3009 -794 3043
rect -1054 2975 -794 3009
rect -1054 2941 -1042 2975
rect -1008 2941 -946 2975
rect -912 2941 -840 2975
rect -806 2941 -794 2975
rect -1054 2907 -794 2941
rect -1054 2873 -1042 2907
rect -1008 2873 -946 2907
rect -912 2873 -840 2907
rect -806 2873 -794 2907
rect -1054 2839 -794 2873
rect -1054 2805 -1042 2839
rect -1008 2805 -946 2839
rect -912 2805 -840 2839
rect -806 2805 -794 2839
rect -1054 2771 -794 2805
rect -1054 2737 -1042 2771
rect -1008 2737 -946 2771
rect -912 2737 -840 2771
rect -806 2737 -794 2771
rect -1054 2703 -794 2737
rect -1054 2669 -1042 2703
rect -1008 2669 -946 2703
rect -912 2669 -840 2703
rect -806 2669 -794 2703
rect -1054 2635 -794 2669
rect -1054 2601 -1042 2635
rect -1008 2601 -946 2635
rect -912 2601 -840 2635
rect -806 2601 -794 2635
rect -1054 2567 -794 2601
rect -1054 2533 -1042 2567
rect -1008 2533 -946 2567
rect -912 2533 -840 2567
rect -806 2533 -794 2567
rect -1054 2499 -794 2533
rect -1054 2465 -1042 2499
rect -1008 2465 -946 2499
rect -912 2465 -840 2499
rect -806 2465 -794 2499
rect -1054 2431 -794 2465
rect -1054 2397 -1042 2431
rect -1008 2397 -946 2431
rect -912 2397 -840 2431
rect -806 2397 -794 2431
rect -1054 2363 -794 2397
rect -1054 2329 -1042 2363
rect -1008 2329 -946 2363
rect -912 2329 -840 2363
rect -806 2329 -794 2363
rect -1054 2295 -794 2329
rect -1054 2261 -1042 2295
rect -1008 2261 -946 2295
rect -912 2261 -840 2295
rect -806 2261 -794 2295
rect -1054 2227 -794 2261
rect -1054 2193 -1042 2227
rect -1008 2193 -946 2227
rect -912 2193 -840 2227
rect -806 2193 -794 2227
rect -1054 2159 -794 2193
rect -1054 2125 -1042 2159
rect -1008 2125 -946 2159
rect -912 2125 -840 2159
rect -806 2125 -794 2159
rect -1054 2091 -794 2125
rect -1054 2057 -1042 2091
rect -1008 2057 -946 2091
rect -912 2057 -840 2091
rect -806 2057 -794 2091
rect -1054 2023 -794 2057
rect -1054 1989 -1042 2023
rect -1008 1989 -946 2023
rect -912 1989 -840 2023
rect -806 1989 -794 2023
rect -1054 1955 -794 1989
rect -1054 1921 -1042 1955
rect -1008 1921 -946 1955
rect -912 1921 -840 1955
rect -806 1921 -794 1955
rect -1054 1887 -794 1921
rect -1054 1853 -1042 1887
rect -1008 1853 -946 1887
rect -912 1853 -840 1887
rect -806 1853 -794 1887
rect -1054 1819 -794 1853
rect -1054 1785 -1042 1819
rect -1008 1785 -946 1819
rect -912 1785 -840 1819
rect -806 1785 -794 1819
rect -1054 1751 -794 1785
rect -1054 1717 -1042 1751
rect -1008 1717 -946 1751
rect -912 1717 -840 1751
rect -806 1717 -794 1751
rect -1054 1683 -794 1717
rect -1054 1649 -1042 1683
rect -1008 1649 -946 1683
rect -912 1649 -840 1683
rect -806 1649 -794 1683
rect -1054 1615 -794 1649
rect -1054 1581 -1042 1615
rect -1008 1581 -946 1615
rect -912 1581 -840 1615
rect -806 1581 -794 1615
rect -1054 1547 -794 1581
rect -1054 1513 -1042 1547
rect -1008 1513 -946 1547
rect -912 1513 -840 1547
rect -806 1513 -794 1547
rect -1054 1479 -794 1513
rect -1054 1445 -1042 1479
rect -1008 1445 -946 1479
rect -912 1445 -840 1479
rect -806 1445 -794 1479
rect -1054 1411 -794 1445
rect -1054 1377 -1042 1411
rect -1008 1377 -946 1411
rect -912 1377 -840 1411
rect -806 1377 -794 1411
rect -1054 1343 -794 1377
rect -1054 1309 -1042 1343
rect -1008 1309 -946 1343
rect -912 1309 -840 1343
rect -806 1309 -794 1343
rect -1054 1275 -794 1309
rect -1054 1241 -1042 1275
rect -1008 1241 -946 1275
rect -912 1241 -840 1275
rect -806 1241 -794 1275
rect -1054 1207 -794 1241
rect -1054 1173 -1042 1207
rect -1008 1173 -946 1207
rect -912 1173 -840 1207
rect -806 1173 -794 1207
rect -1054 1139 -794 1173
rect -1054 1105 -1042 1139
rect -1008 1105 -946 1139
rect -912 1105 -840 1139
rect -806 1105 -794 1139
rect -1054 1071 -794 1105
rect -1054 1037 -1042 1071
rect -1008 1037 -946 1071
rect -912 1037 -840 1071
rect -806 1037 -794 1071
rect -1054 1003 -794 1037
rect -1054 969 -1042 1003
rect -1008 969 -946 1003
rect -912 969 -840 1003
rect -806 969 -794 1003
rect -1054 935 -794 969
rect -1054 901 -1042 935
rect -1008 901 -946 935
rect -912 901 -840 935
rect -806 901 -794 935
rect -1054 867 -794 901
rect -1054 833 -1042 867
rect -1008 833 -946 867
rect -912 833 -840 867
rect -806 833 -794 867
rect -1054 799 -794 833
rect -1054 765 -1042 799
rect -1008 765 -946 799
rect -912 765 -840 799
rect -806 765 -794 799
rect -1054 731 -794 765
rect -1054 697 -1042 731
rect -1008 697 -946 731
rect -912 697 -840 731
rect -806 697 -794 731
rect -1054 663 -794 697
rect -1054 629 -1042 663
rect -1008 629 -946 663
rect -912 629 -840 663
rect -806 629 -794 663
rect -1054 595 -794 629
rect -1054 561 -1042 595
rect -1008 561 -946 595
rect -912 561 -840 595
rect -806 561 -794 595
rect -1054 527 -794 561
rect -1054 493 -1042 527
rect -1008 493 -946 527
rect -912 493 -840 527
rect -806 493 -794 527
rect -1054 459 -794 493
rect -1054 425 -1042 459
rect -1008 425 -946 459
rect -912 425 -840 459
rect -806 425 -794 459
rect -1054 391 -794 425
rect -1054 357 -1042 391
rect -1008 357 -946 391
rect -912 357 -840 391
rect -806 357 -794 391
rect -1054 323 -794 357
rect -1054 289 -1042 323
rect -1008 289 -946 323
rect -912 289 -840 323
rect -806 289 -794 323
rect -1054 255 -794 289
rect -1054 221 -1042 255
rect -1008 221 -946 255
rect -912 221 -840 255
rect -806 221 -794 255
rect -1054 187 -794 221
rect -1054 153 -1042 187
rect -1008 153 -946 187
rect -912 153 -840 187
rect -806 153 -794 187
rect -1054 119 -794 153
rect -1054 85 -1042 119
rect -1008 85 -946 119
rect -912 85 -840 119
rect -806 85 -794 119
rect -1054 51 -794 85
rect -1054 17 -1042 51
rect -1008 17 -946 51
rect -912 17 -840 51
rect -806 17 -794 51
rect -1054 -17 -794 17
rect -1054 -51 -1042 -17
rect -1008 -51 -946 -17
rect -912 -51 -840 -17
rect -806 -51 -794 -17
rect -1054 -85 -794 -51
rect -1054 -119 -1042 -85
rect -1008 -119 -946 -85
rect -912 -119 -840 -85
rect -806 -119 -794 -85
rect -1054 -153 -794 -119
rect -1054 -187 -1042 -153
rect -1008 -187 -946 -153
rect -912 -187 -840 -153
rect -806 -187 -794 -153
rect -1054 -221 -794 -187
rect -1054 -255 -1042 -221
rect -1008 -255 -946 -221
rect -912 -255 -840 -221
rect -806 -255 -794 -221
rect -1054 -289 -794 -255
rect -1054 -323 -1042 -289
rect -1008 -323 -946 -289
rect -912 -323 -840 -289
rect -806 -323 -794 -289
rect -1054 -357 -794 -323
rect -1054 -391 -1042 -357
rect -1008 -391 -946 -357
rect -912 -391 -840 -357
rect -806 -391 -794 -357
rect -1054 -425 -794 -391
rect -1054 -459 -1042 -425
rect -1008 -459 -946 -425
rect -912 -459 -840 -425
rect -806 -459 -794 -425
rect -1054 -493 -794 -459
rect -1054 -527 -1042 -493
rect -1008 -527 -946 -493
rect -912 -527 -840 -493
rect -806 -527 -794 -493
rect -1054 -561 -794 -527
rect -1054 -595 -1042 -561
rect -1008 -595 -946 -561
rect -912 -595 -840 -561
rect -806 -595 -794 -561
rect -1054 -629 -794 -595
rect -1054 -663 -1042 -629
rect -1008 -663 -946 -629
rect -912 -663 -840 -629
rect -806 -663 -794 -629
rect -1054 -697 -794 -663
rect -1054 -731 -1042 -697
rect -1008 -731 -946 -697
rect -912 -731 -840 -697
rect -806 -731 -794 -697
rect -1054 -765 -794 -731
rect -1054 -799 -1042 -765
rect -1008 -799 -946 -765
rect -912 -799 -840 -765
rect -806 -799 -794 -765
rect -1054 -833 -794 -799
rect -1054 -867 -1042 -833
rect -1008 -867 -946 -833
rect -912 -867 -840 -833
rect -806 -867 -794 -833
rect -1054 -901 -794 -867
rect -1054 -935 -1042 -901
rect -1008 -935 -946 -901
rect -912 -935 -840 -901
rect -806 -935 -794 -901
rect -1054 -969 -794 -935
rect -1054 -1003 -1042 -969
rect -1008 -1003 -946 -969
rect -912 -1003 -840 -969
rect -806 -1003 -794 -969
rect -1054 -1037 -794 -1003
rect -1054 -1071 -1042 -1037
rect -1008 -1071 -946 -1037
rect -912 -1071 -840 -1037
rect -806 -1071 -794 -1037
rect -1054 -1105 -794 -1071
rect -1054 -1139 -1042 -1105
rect -1008 -1139 -946 -1105
rect -912 -1139 -840 -1105
rect -806 -1139 -794 -1105
rect -1054 -1173 -794 -1139
rect -1054 -1207 -1042 -1173
rect -1008 -1207 -946 -1173
rect -912 -1207 -840 -1173
rect -806 -1207 -794 -1173
rect -1054 -1241 -794 -1207
rect -1054 -1275 -1042 -1241
rect -1008 -1275 -946 -1241
rect -912 -1275 -840 -1241
rect -806 -1275 -794 -1241
rect -1054 -1309 -794 -1275
rect -1054 -1343 -1042 -1309
rect -1008 -1343 -946 -1309
rect -912 -1343 -840 -1309
rect -806 -1343 -794 -1309
rect -1054 -1377 -794 -1343
rect -1054 -1411 -1042 -1377
rect -1008 -1411 -946 -1377
rect -912 -1411 -840 -1377
rect -806 -1411 -794 -1377
rect -1054 -1445 -794 -1411
rect -1054 -1479 -1042 -1445
rect -1008 -1479 -946 -1445
rect -912 -1479 -840 -1445
rect -806 -1479 -794 -1445
rect -1054 -1513 -794 -1479
rect -1054 -1547 -1042 -1513
rect -1008 -1547 -946 -1513
rect -912 -1547 -840 -1513
rect -806 -1547 -794 -1513
rect -1054 -1581 -794 -1547
rect -1054 -1615 -1042 -1581
rect -1008 -1615 -946 -1581
rect -912 -1615 -840 -1581
rect -806 -1615 -794 -1581
rect -1054 -1649 -794 -1615
rect -1054 -1683 -1042 -1649
rect -1008 -1683 -946 -1649
rect -912 -1683 -840 -1649
rect -806 -1683 -794 -1649
rect -1054 -1717 -794 -1683
rect -1054 -1751 -1042 -1717
rect -1008 -1751 -946 -1717
rect -912 -1751 -840 -1717
rect -806 -1751 -794 -1717
rect -1054 -1785 -794 -1751
rect -1054 -1819 -1042 -1785
rect -1008 -1819 -946 -1785
rect -912 -1819 -840 -1785
rect -806 -1819 -794 -1785
rect -1054 -1853 -794 -1819
rect -1054 -1887 -1042 -1853
rect -1008 -1887 -946 -1853
rect -912 -1887 -840 -1853
rect -806 -1887 -794 -1853
rect -1054 -1921 -794 -1887
rect -1054 -1955 -1042 -1921
rect -1008 -1955 -946 -1921
rect -912 -1955 -840 -1921
rect -806 -1955 -794 -1921
rect -1054 -1989 -794 -1955
rect -1054 -2023 -1042 -1989
rect -1008 -2023 -946 -1989
rect -912 -2023 -840 -1989
rect -806 -2023 -794 -1989
rect -1054 -2057 -794 -2023
rect -1054 -2091 -1042 -2057
rect -1008 -2091 -946 -2057
rect -912 -2091 -840 -2057
rect -806 -2091 -794 -2057
rect -1054 -2125 -794 -2091
rect -1054 -2159 -1042 -2125
rect -1008 -2159 -946 -2125
rect -912 -2159 -840 -2125
rect -806 -2159 -794 -2125
rect -1054 -2193 -794 -2159
rect -1054 -2227 -1042 -2193
rect -1008 -2227 -946 -2193
rect -912 -2227 -840 -2193
rect -806 -2227 -794 -2193
rect -1054 -2261 -794 -2227
rect -1054 -2295 -1042 -2261
rect -1008 -2295 -946 -2261
rect -912 -2295 -840 -2261
rect -806 -2295 -794 -2261
rect -1054 -2329 -794 -2295
rect -1054 -2363 -1042 -2329
rect -1008 -2363 -946 -2329
rect -912 -2363 -840 -2329
rect -806 -2363 -794 -2329
rect -1054 -2397 -794 -2363
rect -1054 -2431 -1042 -2397
rect -1008 -2431 -946 -2397
rect -912 -2431 -840 -2397
rect -806 -2431 -794 -2397
rect -1054 -2465 -794 -2431
rect -1054 -2499 -1042 -2465
rect -1008 -2499 -946 -2465
rect -912 -2499 -840 -2465
rect -806 -2499 -794 -2465
rect -1054 -2533 -794 -2499
rect -1054 -2567 -1042 -2533
rect -1008 -2567 -946 -2533
rect -912 -2567 -840 -2533
rect -806 -2567 -794 -2533
rect -1054 -2601 -794 -2567
rect -1054 -2635 -1042 -2601
rect -1008 -2635 -946 -2601
rect -912 -2635 -840 -2601
rect -806 -2635 -794 -2601
rect -1054 -2669 -794 -2635
rect -1054 -2703 -1042 -2669
rect -1008 -2703 -946 -2669
rect -912 -2703 -840 -2669
rect -806 -2703 -794 -2669
rect -1054 -2737 -794 -2703
rect -1054 -2771 -1042 -2737
rect -1008 -2771 -946 -2737
rect -912 -2771 -840 -2737
rect -806 -2771 -794 -2737
rect -1054 -2805 -794 -2771
rect -1054 -2839 -1042 -2805
rect -1008 -2839 -946 -2805
rect -912 -2839 -840 -2805
rect -806 -2839 -794 -2805
rect -1054 -2873 -794 -2839
rect -1054 -2907 -1042 -2873
rect -1008 -2907 -946 -2873
rect -912 -2907 -840 -2873
rect -806 -2907 -794 -2873
rect -1054 -2941 -794 -2907
rect -1054 -2975 -1042 -2941
rect -1008 -2975 -946 -2941
rect -912 -2975 -840 -2941
rect -806 -2975 -794 -2941
rect -1054 -3009 -794 -2975
rect -1054 -3043 -1042 -3009
rect -1008 -3043 -946 -3009
rect -912 -3043 -840 -3009
rect -806 -3043 -794 -3009
rect -1054 -3077 -794 -3043
rect -1054 -3111 -1042 -3077
rect -1008 -3111 -946 -3077
rect -912 -3111 -840 -3077
rect -806 -3111 -794 -3077
rect -1054 -3145 -794 -3111
rect -1054 -3179 -1042 -3145
rect -1008 -3179 -946 -3145
rect -912 -3179 -840 -3145
rect -806 -3179 -794 -3145
rect -1054 -3213 -794 -3179
rect -1054 -3247 -1042 -3213
rect -1008 -3247 -946 -3213
rect -912 -3247 -840 -3213
rect -806 -3247 -794 -3213
rect -1054 -3281 -794 -3247
rect -1054 -3315 -1042 -3281
rect -1008 -3315 -946 -3281
rect -912 -3315 -840 -3281
rect -806 -3315 -794 -3281
rect -1054 -3349 -794 -3315
rect -1054 -3383 -1042 -3349
rect -1008 -3383 -946 -3349
rect -912 -3383 -840 -3349
rect -806 -3383 -794 -3349
rect -1054 -3417 -794 -3383
rect -1054 -3451 -1042 -3417
rect -1008 -3451 -946 -3417
rect -912 -3451 -840 -3417
rect -806 -3451 -794 -3417
rect -1054 -3485 -794 -3451
rect -1054 -3519 -1042 -3485
rect -1008 -3519 -946 -3485
rect -912 -3519 -840 -3485
rect -806 -3519 -794 -3485
rect -1054 -3553 -794 -3519
rect -1054 -3587 -1042 -3553
rect -1008 -3587 -946 -3553
rect -912 -3587 -840 -3553
rect -806 -3587 -794 -3553
rect -1054 -3621 -794 -3587
rect -1054 -3655 -1042 -3621
rect -1008 -3655 -946 -3621
rect -912 -3655 -840 -3621
rect -806 -3655 -794 -3621
rect -1054 -3689 -794 -3655
rect -1054 -3723 -1042 -3689
rect -1008 -3723 -946 -3689
rect -912 -3723 -840 -3689
rect -806 -3723 -794 -3689
rect -1054 -3757 -794 -3723
rect -1054 -3791 -1042 -3757
rect -1008 -3791 -946 -3757
rect -912 -3791 -840 -3757
rect -806 -3791 -794 -3757
rect -1054 -3825 -794 -3791
rect -1054 -3859 -1042 -3825
rect -1008 -3859 -946 -3825
rect -912 -3859 -840 -3825
rect -806 -3859 -794 -3825
rect -1054 -3893 -794 -3859
rect -1054 -3927 -1042 -3893
rect -1008 -3927 -946 -3893
rect -912 -3927 -840 -3893
rect -806 -3927 -794 -3893
rect -1054 -3961 -794 -3927
rect -1054 -3995 -1042 -3961
rect -1008 -3995 -946 -3961
rect -912 -3995 -840 -3961
rect -806 -3995 -794 -3961
rect -1054 -4029 -794 -3995
rect -1054 -4063 -1042 -4029
rect -1008 -4063 -946 -4029
rect -912 -4063 -840 -4029
rect -806 -4063 -794 -4029
rect -1054 -4097 -794 -4063
rect -1054 -4131 -1042 -4097
rect -1008 -4131 -946 -4097
rect -912 -4131 -840 -4097
rect -806 -4131 -794 -4097
rect -1054 -4165 -794 -4131
rect -1054 -4199 -1042 -4165
rect -1008 -4199 -946 -4165
rect -912 -4199 -840 -4165
rect -806 -4199 -794 -4165
rect -1054 -4233 -794 -4199
rect -1054 -4267 -1042 -4233
rect -1008 -4267 -946 -4233
rect -912 -4267 -840 -4233
rect -806 -4267 -794 -4233
rect -1054 -4301 -794 -4267
rect -1054 -4335 -1042 -4301
rect -1008 -4335 -946 -4301
rect -912 -4335 -840 -4301
rect -806 -4335 -794 -4301
rect -1054 -4369 -794 -4335
rect -1054 -4403 -1042 -4369
rect -1008 -4403 -946 -4369
rect -912 -4403 -840 -4369
rect -806 -4403 -794 -4369
rect -1054 -4437 -794 -4403
rect -1054 -4471 -1042 -4437
rect -1008 -4471 -946 -4437
rect -912 -4471 -840 -4437
rect -806 -4471 -794 -4437
rect -1054 -4505 -794 -4471
rect -1054 -4539 -1042 -4505
rect -1008 -4539 -946 -4505
rect -912 -4539 -840 -4505
rect -806 -4539 -794 -4505
rect -1054 -4573 -794 -4539
rect -1054 -4607 -1042 -4573
rect -1008 -4607 -946 -4573
rect -912 -4607 -840 -4573
rect -806 -4607 -794 -4573
rect -1054 -4641 -794 -4607
rect -1054 -4675 -1042 -4641
rect -1008 -4675 -946 -4641
rect -912 -4675 -840 -4641
rect -806 -4675 -794 -4641
rect -1054 -4709 -794 -4675
rect -1054 -4743 -1042 -4709
rect -1008 -4743 -946 -4709
rect -912 -4743 -840 -4709
rect -806 -4743 -794 -4709
rect -1054 -4777 -794 -4743
rect -1054 -4811 -1042 -4777
rect -1008 -4811 -946 -4777
rect -912 -4811 -840 -4777
rect -806 -4811 -794 -4777
rect -1054 -4845 -794 -4811
rect -1054 -4879 -1042 -4845
rect -1008 -4879 -946 -4845
rect -912 -4879 -840 -4845
rect -806 -4879 -794 -4845
rect -1054 -4913 -794 -4879
rect -1054 -4947 -1042 -4913
rect -1008 -4947 -946 -4913
rect -912 -4947 -840 -4913
rect -806 -4947 -794 -4913
rect -1054 -4981 -794 -4947
rect -1540 -5078 -1410 -5015
rect -1054 -5015 -1042 -4981
rect -1008 -5015 -946 -4981
rect -912 -5015 -840 -4981
rect -806 -5015 -794 -4981
rect -438 4981 -426 5015
rect -392 4981 -330 5015
rect -296 4981 -224 5015
rect -190 4981 -178 5015
rect 178 5015 438 5078
rect -438 4947 -178 4981
rect -438 4913 -426 4947
rect -392 4913 -330 4947
rect -296 4913 -224 4947
rect -190 4913 -178 4947
rect -438 4879 -178 4913
rect -438 4845 -426 4879
rect -392 4845 -330 4879
rect -296 4845 -224 4879
rect -190 4845 -178 4879
rect -438 4811 -178 4845
rect -438 4777 -426 4811
rect -392 4777 -330 4811
rect -296 4777 -224 4811
rect -190 4777 -178 4811
rect -438 4743 -178 4777
rect -438 4709 -426 4743
rect -392 4709 -330 4743
rect -296 4709 -224 4743
rect -190 4709 -178 4743
rect -438 4675 -178 4709
rect -438 4641 -426 4675
rect -392 4641 -330 4675
rect -296 4641 -224 4675
rect -190 4641 -178 4675
rect -438 4607 -178 4641
rect -438 4573 -426 4607
rect -392 4573 -330 4607
rect -296 4573 -224 4607
rect -190 4573 -178 4607
rect -438 4539 -178 4573
rect -438 4505 -426 4539
rect -392 4505 -330 4539
rect -296 4505 -224 4539
rect -190 4505 -178 4539
rect -438 4471 -178 4505
rect -438 4437 -426 4471
rect -392 4437 -330 4471
rect -296 4437 -224 4471
rect -190 4437 -178 4471
rect -438 4403 -178 4437
rect -438 4369 -426 4403
rect -392 4369 -330 4403
rect -296 4369 -224 4403
rect -190 4369 -178 4403
rect -438 4335 -178 4369
rect -438 4301 -426 4335
rect -392 4301 -330 4335
rect -296 4301 -224 4335
rect -190 4301 -178 4335
rect -438 4267 -178 4301
rect -438 4233 -426 4267
rect -392 4233 -330 4267
rect -296 4233 -224 4267
rect -190 4233 -178 4267
rect -438 4199 -178 4233
rect -438 4165 -426 4199
rect -392 4165 -330 4199
rect -296 4165 -224 4199
rect -190 4165 -178 4199
rect -438 4131 -178 4165
rect -438 4097 -426 4131
rect -392 4097 -330 4131
rect -296 4097 -224 4131
rect -190 4097 -178 4131
rect -438 4063 -178 4097
rect -438 4029 -426 4063
rect -392 4029 -330 4063
rect -296 4029 -224 4063
rect -190 4029 -178 4063
rect -438 3995 -178 4029
rect -438 3961 -426 3995
rect -392 3961 -330 3995
rect -296 3961 -224 3995
rect -190 3961 -178 3995
rect -438 3927 -178 3961
rect -438 3893 -426 3927
rect -392 3893 -330 3927
rect -296 3893 -224 3927
rect -190 3893 -178 3927
rect -438 3859 -178 3893
rect -438 3825 -426 3859
rect -392 3825 -330 3859
rect -296 3825 -224 3859
rect -190 3825 -178 3859
rect -438 3791 -178 3825
rect -438 3757 -426 3791
rect -392 3757 -330 3791
rect -296 3757 -224 3791
rect -190 3757 -178 3791
rect -438 3723 -178 3757
rect -438 3689 -426 3723
rect -392 3689 -330 3723
rect -296 3689 -224 3723
rect -190 3689 -178 3723
rect -438 3655 -178 3689
rect -438 3621 -426 3655
rect -392 3621 -330 3655
rect -296 3621 -224 3655
rect -190 3621 -178 3655
rect -438 3587 -178 3621
rect -438 3553 -426 3587
rect -392 3553 -330 3587
rect -296 3553 -224 3587
rect -190 3553 -178 3587
rect -438 3519 -178 3553
rect -438 3485 -426 3519
rect -392 3485 -330 3519
rect -296 3485 -224 3519
rect -190 3485 -178 3519
rect -438 3451 -178 3485
rect -438 3417 -426 3451
rect -392 3417 -330 3451
rect -296 3417 -224 3451
rect -190 3417 -178 3451
rect -438 3383 -178 3417
rect -438 3349 -426 3383
rect -392 3349 -330 3383
rect -296 3349 -224 3383
rect -190 3349 -178 3383
rect -438 3315 -178 3349
rect -438 3281 -426 3315
rect -392 3281 -330 3315
rect -296 3281 -224 3315
rect -190 3281 -178 3315
rect -438 3247 -178 3281
rect -438 3213 -426 3247
rect -392 3213 -330 3247
rect -296 3213 -224 3247
rect -190 3213 -178 3247
rect -438 3179 -178 3213
rect -438 3145 -426 3179
rect -392 3145 -330 3179
rect -296 3145 -224 3179
rect -190 3145 -178 3179
rect -438 3111 -178 3145
rect -438 3077 -426 3111
rect -392 3077 -330 3111
rect -296 3077 -224 3111
rect -190 3077 -178 3111
rect -438 3043 -178 3077
rect -438 3009 -426 3043
rect -392 3009 -330 3043
rect -296 3009 -224 3043
rect -190 3009 -178 3043
rect -438 2975 -178 3009
rect -438 2941 -426 2975
rect -392 2941 -330 2975
rect -296 2941 -224 2975
rect -190 2941 -178 2975
rect -438 2907 -178 2941
rect -438 2873 -426 2907
rect -392 2873 -330 2907
rect -296 2873 -224 2907
rect -190 2873 -178 2907
rect -438 2839 -178 2873
rect -438 2805 -426 2839
rect -392 2805 -330 2839
rect -296 2805 -224 2839
rect -190 2805 -178 2839
rect -438 2771 -178 2805
rect -438 2737 -426 2771
rect -392 2737 -330 2771
rect -296 2737 -224 2771
rect -190 2737 -178 2771
rect -438 2703 -178 2737
rect -438 2669 -426 2703
rect -392 2669 -330 2703
rect -296 2669 -224 2703
rect -190 2669 -178 2703
rect -438 2635 -178 2669
rect -438 2601 -426 2635
rect -392 2601 -330 2635
rect -296 2601 -224 2635
rect -190 2601 -178 2635
rect -438 2567 -178 2601
rect -438 2533 -426 2567
rect -392 2533 -330 2567
rect -296 2533 -224 2567
rect -190 2533 -178 2567
rect -438 2499 -178 2533
rect -438 2465 -426 2499
rect -392 2465 -330 2499
rect -296 2465 -224 2499
rect -190 2465 -178 2499
rect -438 2431 -178 2465
rect -438 2397 -426 2431
rect -392 2397 -330 2431
rect -296 2397 -224 2431
rect -190 2397 -178 2431
rect -438 2363 -178 2397
rect -438 2329 -426 2363
rect -392 2329 -330 2363
rect -296 2329 -224 2363
rect -190 2329 -178 2363
rect -438 2295 -178 2329
rect -438 2261 -426 2295
rect -392 2261 -330 2295
rect -296 2261 -224 2295
rect -190 2261 -178 2295
rect -438 2227 -178 2261
rect -438 2193 -426 2227
rect -392 2193 -330 2227
rect -296 2193 -224 2227
rect -190 2193 -178 2227
rect -438 2159 -178 2193
rect -438 2125 -426 2159
rect -392 2125 -330 2159
rect -296 2125 -224 2159
rect -190 2125 -178 2159
rect -438 2091 -178 2125
rect -438 2057 -426 2091
rect -392 2057 -330 2091
rect -296 2057 -224 2091
rect -190 2057 -178 2091
rect -438 2023 -178 2057
rect -438 1989 -426 2023
rect -392 1989 -330 2023
rect -296 1989 -224 2023
rect -190 1989 -178 2023
rect -438 1955 -178 1989
rect -438 1921 -426 1955
rect -392 1921 -330 1955
rect -296 1921 -224 1955
rect -190 1921 -178 1955
rect -438 1887 -178 1921
rect -438 1853 -426 1887
rect -392 1853 -330 1887
rect -296 1853 -224 1887
rect -190 1853 -178 1887
rect -438 1819 -178 1853
rect -438 1785 -426 1819
rect -392 1785 -330 1819
rect -296 1785 -224 1819
rect -190 1785 -178 1819
rect -438 1751 -178 1785
rect -438 1717 -426 1751
rect -392 1717 -330 1751
rect -296 1717 -224 1751
rect -190 1717 -178 1751
rect -438 1683 -178 1717
rect -438 1649 -426 1683
rect -392 1649 -330 1683
rect -296 1649 -224 1683
rect -190 1649 -178 1683
rect -438 1615 -178 1649
rect -438 1581 -426 1615
rect -392 1581 -330 1615
rect -296 1581 -224 1615
rect -190 1581 -178 1615
rect -438 1547 -178 1581
rect -438 1513 -426 1547
rect -392 1513 -330 1547
rect -296 1513 -224 1547
rect -190 1513 -178 1547
rect -438 1479 -178 1513
rect -438 1445 -426 1479
rect -392 1445 -330 1479
rect -296 1445 -224 1479
rect -190 1445 -178 1479
rect -438 1411 -178 1445
rect -438 1377 -426 1411
rect -392 1377 -330 1411
rect -296 1377 -224 1411
rect -190 1377 -178 1411
rect -438 1343 -178 1377
rect -438 1309 -426 1343
rect -392 1309 -330 1343
rect -296 1309 -224 1343
rect -190 1309 -178 1343
rect -438 1275 -178 1309
rect -438 1241 -426 1275
rect -392 1241 -330 1275
rect -296 1241 -224 1275
rect -190 1241 -178 1275
rect -438 1207 -178 1241
rect -438 1173 -426 1207
rect -392 1173 -330 1207
rect -296 1173 -224 1207
rect -190 1173 -178 1207
rect -438 1139 -178 1173
rect -438 1105 -426 1139
rect -392 1105 -330 1139
rect -296 1105 -224 1139
rect -190 1105 -178 1139
rect -438 1071 -178 1105
rect -438 1037 -426 1071
rect -392 1037 -330 1071
rect -296 1037 -224 1071
rect -190 1037 -178 1071
rect -438 1003 -178 1037
rect -438 969 -426 1003
rect -392 969 -330 1003
rect -296 969 -224 1003
rect -190 969 -178 1003
rect -438 935 -178 969
rect -438 901 -426 935
rect -392 901 -330 935
rect -296 901 -224 935
rect -190 901 -178 935
rect -438 867 -178 901
rect -438 833 -426 867
rect -392 833 -330 867
rect -296 833 -224 867
rect -190 833 -178 867
rect -438 799 -178 833
rect -438 765 -426 799
rect -392 765 -330 799
rect -296 765 -224 799
rect -190 765 -178 799
rect -438 731 -178 765
rect -438 697 -426 731
rect -392 697 -330 731
rect -296 697 -224 731
rect -190 697 -178 731
rect -438 663 -178 697
rect -438 629 -426 663
rect -392 629 -330 663
rect -296 629 -224 663
rect -190 629 -178 663
rect -438 595 -178 629
rect -438 561 -426 595
rect -392 561 -330 595
rect -296 561 -224 595
rect -190 561 -178 595
rect -438 527 -178 561
rect -438 493 -426 527
rect -392 493 -330 527
rect -296 493 -224 527
rect -190 493 -178 527
rect -438 459 -178 493
rect -438 425 -426 459
rect -392 425 -330 459
rect -296 425 -224 459
rect -190 425 -178 459
rect -438 391 -178 425
rect -438 357 -426 391
rect -392 357 -330 391
rect -296 357 -224 391
rect -190 357 -178 391
rect -438 323 -178 357
rect -438 289 -426 323
rect -392 289 -330 323
rect -296 289 -224 323
rect -190 289 -178 323
rect -438 255 -178 289
rect -438 221 -426 255
rect -392 221 -330 255
rect -296 221 -224 255
rect -190 221 -178 255
rect -438 187 -178 221
rect -438 153 -426 187
rect -392 153 -330 187
rect -296 153 -224 187
rect -190 153 -178 187
rect -438 119 -178 153
rect -438 85 -426 119
rect -392 85 -330 119
rect -296 85 -224 119
rect -190 85 -178 119
rect -438 51 -178 85
rect -438 17 -426 51
rect -392 17 -330 51
rect -296 17 -224 51
rect -190 17 -178 51
rect -438 -17 -178 17
rect -438 -51 -426 -17
rect -392 -51 -330 -17
rect -296 -51 -224 -17
rect -190 -51 -178 -17
rect -438 -85 -178 -51
rect -438 -119 -426 -85
rect -392 -119 -330 -85
rect -296 -119 -224 -85
rect -190 -119 -178 -85
rect -438 -153 -178 -119
rect -438 -187 -426 -153
rect -392 -187 -330 -153
rect -296 -187 -224 -153
rect -190 -187 -178 -153
rect -438 -221 -178 -187
rect -438 -255 -426 -221
rect -392 -255 -330 -221
rect -296 -255 -224 -221
rect -190 -255 -178 -221
rect -438 -289 -178 -255
rect -438 -323 -426 -289
rect -392 -323 -330 -289
rect -296 -323 -224 -289
rect -190 -323 -178 -289
rect -438 -357 -178 -323
rect -438 -391 -426 -357
rect -392 -391 -330 -357
rect -296 -391 -224 -357
rect -190 -391 -178 -357
rect -438 -425 -178 -391
rect -438 -459 -426 -425
rect -392 -459 -330 -425
rect -296 -459 -224 -425
rect -190 -459 -178 -425
rect -438 -493 -178 -459
rect -438 -527 -426 -493
rect -392 -527 -330 -493
rect -296 -527 -224 -493
rect -190 -527 -178 -493
rect -438 -561 -178 -527
rect -438 -595 -426 -561
rect -392 -595 -330 -561
rect -296 -595 -224 -561
rect -190 -595 -178 -561
rect -438 -629 -178 -595
rect -438 -663 -426 -629
rect -392 -663 -330 -629
rect -296 -663 -224 -629
rect -190 -663 -178 -629
rect -438 -697 -178 -663
rect -438 -731 -426 -697
rect -392 -731 -330 -697
rect -296 -731 -224 -697
rect -190 -731 -178 -697
rect -438 -765 -178 -731
rect -438 -799 -426 -765
rect -392 -799 -330 -765
rect -296 -799 -224 -765
rect -190 -799 -178 -765
rect -438 -833 -178 -799
rect -438 -867 -426 -833
rect -392 -867 -330 -833
rect -296 -867 -224 -833
rect -190 -867 -178 -833
rect -438 -901 -178 -867
rect -438 -935 -426 -901
rect -392 -935 -330 -901
rect -296 -935 -224 -901
rect -190 -935 -178 -901
rect -438 -969 -178 -935
rect -438 -1003 -426 -969
rect -392 -1003 -330 -969
rect -296 -1003 -224 -969
rect -190 -1003 -178 -969
rect -438 -1037 -178 -1003
rect -438 -1071 -426 -1037
rect -392 -1071 -330 -1037
rect -296 -1071 -224 -1037
rect -190 -1071 -178 -1037
rect -438 -1105 -178 -1071
rect -438 -1139 -426 -1105
rect -392 -1139 -330 -1105
rect -296 -1139 -224 -1105
rect -190 -1139 -178 -1105
rect -438 -1173 -178 -1139
rect -438 -1207 -426 -1173
rect -392 -1207 -330 -1173
rect -296 -1207 -224 -1173
rect -190 -1207 -178 -1173
rect -438 -1241 -178 -1207
rect -438 -1275 -426 -1241
rect -392 -1275 -330 -1241
rect -296 -1275 -224 -1241
rect -190 -1275 -178 -1241
rect -438 -1309 -178 -1275
rect -438 -1343 -426 -1309
rect -392 -1343 -330 -1309
rect -296 -1343 -224 -1309
rect -190 -1343 -178 -1309
rect -438 -1377 -178 -1343
rect -438 -1411 -426 -1377
rect -392 -1411 -330 -1377
rect -296 -1411 -224 -1377
rect -190 -1411 -178 -1377
rect -438 -1445 -178 -1411
rect -438 -1479 -426 -1445
rect -392 -1479 -330 -1445
rect -296 -1479 -224 -1445
rect -190 -1479 -178 -1445
rect -438 -1513 -178 -1479
rect -438 -1547 -426 -1513
rect -392 -1547 -330 -1513
rect -296 -1547 -224 -1513
rect -190 -1547 -178 -1513
rect -438 -1581 -178 -1547
rect -438 -1615 -426 -1581
rect -392 -1615 -330 -1581
rect -296 -1615 -224 -1581
rect -190 -1615 -178 -1581
rect -438 -1649 -178 -1615
rect -438 -1683 -426 -1649
rect -392 -1683 -330 -1649
rect -296 -1683 -224 -1649
rect -190 -1683 -178 -1649
rect -438 -1717 -178 -1683
rect -438 -1751 -426 -1717
rect -392 -1751 -330 -1717
rect -296 -1751 -224 -1717
rect -190 -1751 -178 -1717
rect -438 -1785 -178 -1751
rect -438 -1819 -426 -1785
rect -392 -1819 -330 -1785
rect -296 -1819 -224 -1785
rect -190 -1819 -178 -1785
rect -438 -1853 -178 -1819
rect -438 -1887 -426 -1853
rect -392 -1887 -330 -1853
rect -296 -1887 -224 -1853
rect -190 -1887 -178 -1853
rect -438 -1921 -178 -1887
rect -438 -1955 -426 -1921
rect -392 -1955 -330 -1921
rect -296 -1955 -224 -1921
rect -190 -1955 -178 -1921
rect -438 -1989 -178 -1955
rect -438 -2023 -426 -1989
rect -392 -2023 -330 -1989
rect -296 -2023 -224 -1989
rect -190 -2023 -178 -1989
rect -438 -2057 -178 -2023
rect -438 -2091 -426 -2057
rect -392 -2091 -330 -2057
rect -296 -2091 -224 -2057
rect -190 -2091 -178 -2057
rect -438 -2125 -178 -2091
rect -438 -2159 -426 -2125
rect -392 -2159 -330 -2125
rect -296 -2159 -224 -2125
rect -190 -2159 -178 -2125
rect -438 -2193 -178 -2159
rect -438 -2227 -426 -2193
rect -392 -2227 -330 -2193
rect -296 -2227 -224 -2193
rect -190 -2227 -178 -2193
rect -438 -2261 -178 -2227
rect -438 -2295 -426 -2261
rect -392 -2295 -330 -2261
rect -296 -2295 -224 -2261
rect -190 -2295 -178 -2261
rect -438 -2329 -178 -2295
rect -438 -2363 -426 -2329
rect -392 -2363 -330 -2329
rect -296 -2363 -224 -2329
rect -190 -2363 -178 -2329
rect -438 -2397 -178 -2363
rect -438 -2431 -426 -2397
rect -392 -2431 -330 -2397
rect -296 -2431 -224 -2397
rect -190 -2431 -178 -2397
rect -438 -2465 -178 -2431
rect -438 -2499 -426 -2465
rect -392 -2499 -330 -2465
rect -296 -2499 -224 -2465
rect -190 -2499 -178 -2465
rect -438 -2533 -178 -2499
rect -438 -2567 -426 -2533
rect -392 -2567 -330 -2533
rect -296 -2567 -224 -2533
rect -190 -2567 -178 -2533
rect -438 -2601 -178 -2567
rect -438 -2635 -426 -2601
rect -392 -2635 -330 -2601
rect -296 -2635 -224 -2601
rect -190 -2635 -178 -2601
rect -438 -2669 -178 -2635
rect -438 -2703 -426 -2669
rect -392 -2703 -330 -2669
rect -296 -2703 -224 -2669
rect -190 -2703 -178 -2669
rect -438 -2737 -178 -2703
rect -438 -2771 -426 -2737
rect -392 -2771 -330 -2737
rect -296 -2771 -224 -2737
rect -190 -2771 -178 -2737
rect -438 -2805 -178 -2771
rect -438 -2839 -426 -2805
rect -392 -2839 -330 -2805
rect -296 -2839 -224 -2805
rect -190 -2839 -178 -2805
rect -438 -2873 -178 -2839
rect -438 -2907 -426 -2873
rect -392 -2907 -330 -2873
rect -296 -2907 -224 -2873
rect -190 -2907 -178 -2873
rect -438 -2941 -178 -2907
rect -438 -2975 -426 -2941
rect -392 -2975 -330 -2941
rect -296 -2975 -224 -2941
rect -190 -2975 -178 -2941
rect -438 -3009 -178 -2975
rect -438 -3043 -426 -3009
rect -392 -3043 -330 -3009
rect -296 -3043 -224 -3009
rect -190 -3043 -178 -3009
rect -438 -3077 -178 -3043
rect -438 -3111 -426 -3077
rect -392 -3111 -330 -3077
rect -296 -3111 -224 -3077
rect -190 -3111 -178 -3077
rect -438 -3145 -178 -3111
rect -438 -3179 -426 -3145
rect -392 -3179 -330 -3145
rect -296 -3179 -224 -3145
rect -190 -3179 -178 -3145
rect -438 -3213 -178 -3179
rect -438 -3247 -426 -3213
rect -392 -3247 -330 -3213
rect -296 -3247 -224 -3213
rect -190 -3247 -178 -3213
rect -438 -3281 -178 -3247
rect -438 -3315 -426 -3281
rect -392 -3315 -330 -3281
rect -296 -3315 -224 -3281
rect -190 -3315 -178 -3281
rect -438 -3349 -178 -3315
rect -438 -3383 -426 -3349
rect -392 -3383 -330 -3349
rect -296 -3383 -224 -3349
rect -190 -3383 -178 -3349
rect -438 -3417 -178 -3383
rect -438 -3451 -426 -3417
rect -392 -3451 -330 -3417
rect -296 -3451 -224 -3417
rect -190 -3451 -178 -3417
rect -438 -3485 -178 -3451
rect -438 -3519 -426 -3485
rect -392 -3519 -330 -3485
rect -296 -3519 -224 -3485
rect -190 -3519 -178 -3485
rect -438 -3553 -178 -3519
rect -438 -3587 -426 -3553
rect -392 -3587 -330 -3553
rect -296 -3587 -224 -3553
rect -190 -3587 -178 -3553
rect -438 -3621 -178 -3587
rect -438 -3655 -426 -3621
rect -392 -3655 -330 -3621
rect -296 -3655 -224 -3621
rect -190 -3655 -178 -3621
rect -438 -3689 -178 -3655
rect -438 -3723 -426 -3689
rect -392 -3723 -330 -3689
rect -296 -3723 -224 -3689
rect -190 -3723 -178 -3689
rect -438 -3757 -178 -3723
rect -438 -3791 -426 -3757
rect -392 -3791 -330 -3757
rect -296 -3791 -224 -3757
rect -190 -3791 -178 -3757
rect -438 -3825 -178 -3791
rect -438 -3859 -426 -3825
rect -392 -3859 -330 -3825
rect -296 -3859 -224 -3825
rect -190 -3859 -178 -3825
rect -438 -3893 -178 -3859
rect -438 -3927 -426 -3893
rect -392 -3927 -330 -3893
rect -296 -3927 -224 -3893
rect -190 -3927 -178 -3893
rect -438 -3961 -178 -3927
rect -438 -3995 -426 -3961
rect -392 -3995 -330 -3961
rect -296 -3995 -224 -3961
rect -190 -3995 -178 -3961
rect -438 -4029 -178 -3995
rect -438 -4063 -426 -4029
rect -392 -4063 -330 -4029
rect -296 -4063 -224 -4029
rect -190 -4063 -178 -4029
rect -438 -4097 -178 -4063
rect -438 -4131 -426 -4097
rect -392 -4131 -330 -4097
rect -296 -4131 -224 -4097
rect -190 -4131 -178 -4097
rect -438 -4165 -178 -4131
rect -438 -4199 -426 -4165
rect -392 -4199 -330 -4165
rect -296 -4199 -224 -4165
rect -190 -4199 -178 -4165
rect -438 -4233 -178 -4199
rect -438 -4267 -426 -4233
rect -392 -4267 -330 -4233
rect -296 -4267 -224 -4233
rect -190 -4267 -178 -4233
rect -438 -4301 -178 -4267
rect -438 -4335 -426 -4301
rect -392 -4335 -330 -4301
rect -296 -4335 -224 -4301
rect -190 -4335 -178 -4301
rect -438 -4369 -178 -4335
rect -438 -4403 -426 -4369
rect -392 -4403 -330 -4369
rect -296 -4403 -224 -4369
rect -190 -4403 -178 -4369
rect -438 -4437 -178 -4403
rect -438 -4471 -426 -4437
rect -392 -4471 -330 -4437
rect -296 -4471 -224 -4437
rect -190 -4471 -178 -4437
rect -438 -4505 -178 -4471
rect -438 -4539 -426 -4505
rect -392 -4539 -330 -4505
rect -296 -4539 -224 -4505
rect -190 -4539 -178 -4505
rect -438 -4573 -178 -4539
rect -438 -4607 -426 -4573
rect -392 -4607 -330 -4573
rect -296 -4607 -224 -4573
rect -190 -4607 -178 -4573
rect -438 -4641 -178 -4607
rect -438 -4675 -426 -4641
rect -392 -4675 -330 -4641
rect -296 -4675 -224 -4641
rect -190 -4675 -178 -4641
rect -438 -4709 -178 -4675
rect -438 -4743 -426 -4709
rect -392 -4743 -330 -4709
rect -296 -4743 -224 -4709
rect -190 -4743 -178 -4709
rect -438 -4777 -178 -4743
rect -438 -4811 -426 -4777
rect -392 -4811 -330 -4777
rect -296 -4811 -224 -4777
rect -190 -4811 -178 -4777
rect -438 -4845 -178 -4811
rect -438 -4879 -426 -4845
rect -392 -4879 -330 -4845
rect -296 -4879 -224 -4845
rect -190 -4879 -178 -4845
rect -438 -4913 -178 -4879
rect -438 -4947 -426 -4913
rect -392 -4947 -330 -4913
rect -296 -4947 -224 -4913
rect -190 -4947 -178 -4913
rect -438 -4981 -178 -4947
rect -1054 -5078 -794 -5015
rect -438 -5015 -426 -4981
rect -392 -5015 -330 -4981
rect -296 -5015 -224 -4981
rect -190 -5015 -178 -4981
rect 178 4981 190 5015
rect 224 4981 286 5015
rect 320 4981 392 5015
rect 426 4981 438 5015
rect 794 5015 1054 5078
rect 178 4947 438 4981
rect 178 4913 190 4947
rect 224 4913 286 4947
rect 320 4913 392 4947
rect 426 4913 438 4947
rect 178 4879 438 4913
rect 178 4845 190 4879
rect 224 4845 286 4879
rect 320 4845 392 4879
rect 426 4845 438 4879
rect 178 4811 438 4845
rect 178 4777 190 4811
rect 224 4777 286 4811
rect 320 4777 392 4811
rect 426 4777 438 4811
rect 178 4743 438 4777
rect 178 4709 190 4743
rect 224 4709 286 4743
rect 320 4709 392 4743
rect 426 4709 438 4743
rect 178 4675 438 4709
rect 178 4641 190 4675
rect 224 4641 286 4675
rect 320 4641 392 4675
rect 426 4641 438 4675
rect 178 4607 438 4641
rect 178 4573 190 4607
rect 224 4573 286 4607
rect 320 4573 392 4607
rect 426 4573 438 4607
rect 178 4539 438 4573
rect 178 4505 190 4539
rect 224 4505 286 4539
rect 320 4505 392 4539
rect 426 4505 438 4539
rect 178 4471 438 4505
rect 178 4437 190 4471
rect 224 4437 286 4471
rect 320 4437 392 4471
rect 426 4437 438 4471
rect 178 4403 438 4437
rect 178 4369 190 4403
rect 224 4369 286 4403
rect 320 4369 392 4403
rect 426 4369 438 4403
rect 178 4335 438 4369
rect 178 4301 190 4335
rect 224 4301 286 4335
rect 320 4301 392 4335
rect 426 4301 438 4335
rect 178 4267 438 4301
rect 178 4233 190 4267
rect 224 4233 286 4267
rect 320 4233 392 4267
rect 426 4233 438 4267
rect 178 4199 438 4233
rect 178 4165 190 4199
rect 224 4165 286 4199
rect 320 4165 392 4199
rect 426 4165 438 4199
rect 178 4131 438 4165
rect 178 4097 190 4131
rect 224 4097 286 4131
rect 320 4097 392 4131
rect 426 4097 438 4131
rect 178 4063 438 4097
rect 178 4029 190 4063
rect 224 4029 286 4063
rect 320 4029 392 4063
rect 426 4029 438 4063
rect 178 3995 438 4029
rect 178 3961 190 3995
rect 224 3961 286 3995
rect 320 3961 392 3995
rect 426 3961 438 3995
rect 178 3927 438 3961
rect 178 3893 190 3927
rect 224 3893 286 3927
rect 320 3893 392 3927
rect 426 3893 438 3927
rect 178 3859 438 3893
rect 178 3825 190 3859
rect 224 3825 286 3859
rect 320 3825 392 3859
rect 426 3825 438 3859
rect 178 3791 438 3825
rect 178 3757 190 3791
rect 224 3757 286 3791
rect 320 3757 392 3791
rect 426 3757 438 3791
rect 178 3723 438 3757
rect 178 3689 190 3723
rect 224 3689 286 3723
rect 320 3689 392 3723
rect 426 3689 438 3723
rect 178 3655 438 3689
rect 178 3621 190 3655
rect 224 3621 286 3655
rect 320 3621 392 3655
rect 426 3621 438 3655
rect 178 3587 438 3621
rect 178 3553 190 3587
rect 224 3553 286 3587
rect 320 3553 392 3587
rect 426 3553 438 3587
rect 178 3519 438 3553
rect 178 3485 190 3519
rect 224 3485 286 3519
rect 320 3485 392 3519
rect 426 3485 438 3519
rect 178 3451 438 3485
rect 178 3417 190 3451
rect 224 3417 286 3451
rect 320 3417 392 3451
rect 426 3417 438 3451
rect 178 3383 438 3417
rect 178 3349 190 3383
rect 224 3349 286 3383
rect 320 3349 392 3383
rect 426 3349 438 3383
rect 178 3315 438 3349
rect 178 3281 190 3315
rect 224 3281 286 3315
rect 320 3281 392 3315
rect 426 3281 438 3315
rect 178 3247 438 3281
rect 178 3213 190 3247
rect 224 3213 286 3247
rect 320 3213 392 3247
rect 426 3213 438 3247
rect 178 3179 438 3213
rect 178 3145 190 3179
rect 224 3145 286 3179
rect 320 3145 392 3179
rect 426 3145 438 3179
rect 178 3111 438 3145
rect 178 3077 190 3111
rect 224 3077 286 3111
rect 320 3077 392 3111
rect 426 3077 438 3111
rect 178 3043 438 3077
rect 178 3009 190 3043
rect 224 3009 286 3043
rect 320 3009 392 3043
rect 426 3009 438 3043
rect 178 2975 438 3009
rect 178 2941 190 2975
rect 224 2941 286 2975
rect 320 2941 392 2975
rect 426 2941 438 2975
rect 178 2907 438 2941
rect 178 2873 190 2907
rect 224 2873 286 2907
rect 320 2873 392 2907
rect 426 2873 438 2907
rect 178 2839 438 2873
rect 178 2805 190 2839
rect 224 2805 286 2839
rect 320 2805 392 2839
rect 426 2805 438 2839
rect 178 2771 438 2805
rect 178 2737 190 2771
rect 224 2737 286 2771
rect 320 2737 392 2771
rect 426 2737 438 2771
rect 178 2703 438 2737
rect 178 2669 190 2703
rect 224 2669 286 2703
rect 320 2669 392 2703
rect 426 2669 438 2703
rect 178 2635 438 2669
rect 178 2601 190 2635
rect 224 2601 286 2635
rect 320 2601 392 2635
rect 426 2601 438 2635
rect 178 2567 438 2601
rect 178 2533 190 2567
rect 224 2533 286 2567
rect 320 2533 392 2567
rect 426 2533 438 2567
rect 178 2499 438 2533
rect 178 2465 190 2499
rect 224 2465 286 2499
rect 320 2465 392 2499
rect 426 2465 438 2499
rect 178 2431 438 2465
rect 178 2397 190 2431
rect 224 2397 286 2431
rect 320 2397 392 2431
rect 426 2397 438 2431
rect 178 2363 438 2397
rect 178 2329 190 2363
rect 224 2329 286 2363
rect 320 2329 392 2363
rect 426 2329 438 2363
rect 178 2295 438 2329
rect 178 2261 190 2295
rect 224 2261 286 2295
rect 320 2261 392 2295
rect 426 2261 438 2295
rect 178 2227 438 2261
rect 178 2193 190 2227
rect 224 2193 286 2227
rect 320 2193 392 2227
rect 426 2193 438 2227
rect 178 2159 438 2193
rect 178 2125 190 2159
rect 224 2125 286 2159
rect 320 2125 392 2159
rect 426 2125 438 2159
rect 178 2091 438 2125
rect 178 2057 190 2091
rect 224 2057 286 2091
rect 320 2057 392 2091
rect 426 2057 438 2091
rect 178 2023 438 2057
rect 178 1989 190 2023
rect 224 1989 286 2023
rect 320 1989 392 2023
rect 426 1989 438 2023
rect 178 1955 438 1989
rect 178 1921 190 1955
rect 224 1921 286 1955
rect 320 1921 392 1955
rect 426 1921 438 1955
rect 178 1887 438 1921
rect 178 1853 190 1887
rect 224 1853 286 1887
rect 320 1853 392 1887
rect 426 1853 438 1887
rect 178 1819 438 1853
rect 178 1785 190 1819
rect 224 1785 286 1819
rect 320 1785 392 1819
rect 426 1785 438 1819
rect 178 1751 438 1785
rect 178 1717 190 1751
rect 224 1717 286 1751
rect 320 1717 392 1751
rect 426 1717 438 1751
rect 178 1683 438 1717
rect 178 1649 190 1683
rect 224 1649 286 1683
rect 320 1649 392 1683
rect 426 1649 438 1683
rect 178 1615 438 1649
rect 178 1581 190 1615
rect 224 1581 286 1615
rect 320 1581 392 1615
rect 426 1581 438 1615
rect 178 1547 438 1581
rect 178 1513 190 1547
rect 224 1513 286 1547
rect 320 1513 392 1547
rect 426 1513 438 1547
rect 178 1479 438 1513
rect 178 1445 190 1479
rect 224 1445 286 1479
rect 320 1445 392 1479
rect 426 1445 438 1479
rect 178 1411 438 1445
rect 178 1377 190 1411
rect 224 1377 286 1411
rect 320 1377 392 1411
rect 426 1377 438 1411
rect 178 1343 438 1377
rect 178 1309 190 1343
rect 224 1309 286 1343
rect 320 1309 392 1343
rect 426 1309 438 1343
rect 178 1275 438 1309
rect 178 1241 190 1275
rect 224 1241 286 1275
rect 320 1241 392 1275
rect 426 1241 438 1275
rect 178 1207 438 1241
rect 178 1173 190 1207
rect 224 1173 286 1207
rect 320 1173 392 1207
rect 426 1173 438 1207
rect 178 1139 438 1173
rect 178 1105 190 1139
rect 224 1105 286 1139
rect 320 1105 392 1139
rect 426 1105 438 1139
rect 178 1071 438 1105
rect 178 1037 190 1071
rect 224 1037 286 1071
rect 320 1037 392 1071
rect 426 1037 438 1071
rect 178 1003 438 1037
rect 178 969 190 1003
rect 224 969 286 1003
rect 320 969 392 1003
rect 426 969 438 1003
rect 178 935 438 969
rect 178 901 190 935
rect 224 901 286 935
rect 320 901 392 935
rect 426 901 438 935
rect 178 867 438 901
rect 178 833 190 867
rect 224 833 286 867
rect 320 833 392 867
rect 426 833 438 867
rect 178 799 438 833
rect 178 765 190 799
rect 224 765 286 799
rect 320 765 392 799
rect 426 765 438 799
rect 178 731 438 765
rect 178 697 190 731
rect 224 697 286 731
rect 320 697 392 731
rect 426 697 438 731
rect 178 663 438 697
rect 178 629 190 663
rect 224 629 286 663
rect 320 629 392 663
rect 426 629 438 663
rect 178 595 438 629
rect 178 561 190 595
rect 224 561 286 595
rect 320 561 392 595
rect 426 561 438 595
rect 178 527 438 561
rect 178 493 190 527
rect 224 493 286 527
rect 320 493 392 527
rect 426 493 438 527
rect 178 459 438 493
rect 178 425 190 459
rect 224 425 286 459
rect 320 425 392 459
rect 426 425 438 459
rect 178 391 438 425
rect 178 357 190 391
rect 224 357 286 391
rect 320 357 392 391
rect 426 357 438 391
rect 178 323 438 357
rect 178 289 190 323
rect 224 289 286 323
rect 320 289 392 323
rect 426 289 438 323
rect 178 255 438 289
rect 178 221 190 255
rect 224 221 286 255
rect 320 221 392 255
rect 426 221 438 255
rect 178 187 438 221
rect 178 153 190 187
rect 224 153 286 187
rect 320 153 392 187
rect 426 153 438 187
rect 178 119 438 153
rect 178 85 190 119
rect 224 85 286 119
rect 320 85 392 119
rect 426 85 438 119
rect 178 51 438 85
rect 178 17 190 51
rect 224 17 286 51
rect 320 17 392 51
rect 426 17 438 51
rect 178 -17 438 17
rect 178 -51 190 -17
rect 224 -51 286 -17
rect 320 -51 392 -17
rect 426 -51 438 -17
rect 178 -85 438 -51
rect 178 -119 190 -85
rect 224 -119 286 -85
rect 320 -119 392 -85
rect 426 -119 438 -85
rect 178 -153 438 -119
rect 178 -187 190 -153
rect 224 -187 286 -153
rect 320 -187 392 -153
rect 426 -187 438 -153
rect 178 -221 438 -187
rect 178 -255 190 -221
rect 224 -255 286 -221
rect 320 -255 392 -221
rect 426 -255 438 -221
rect 178 -289 438 -255
rect 178 -323 190 -289
rect 224 -323 286 -289
rect 320 -323 392 -289
rect 426 -323 438 -289
rect 178 -357 438 -323
rect 178 -391 190 -357
rect 224 -391 286 -357
rect 320 -391 392 -357
rect 426 -391 438 -357
rect 178 -425 438 -391
rect 178 -459 190 -425
rect 224 -459 286 -425
rect 320 -459 392 -425
rect 426 -459 438 -425
rect 178 -493 438 -459
rect 178 -527 190 -493
rect 224 -527 286 -493
rect 320 -527 392 -493
rect 426 -527 438 -493
rect 178 -561 438 -527
rect 178 -595 190 -561
rect 224 -595 286 -561
rect 320 -595 392 -561
rect 426 -595 438 -561
rect 178 -629 438 -595
rect 178 -663 190 -629
rect 224 -663 286 -629
rect 320 -663 392 -629
rect 426 -663 438 -629
rect 178 -697 438 -663
rect 178 -731 190 -697
rect 224 -731 286 -697
rect 320 -731 392 -697
rect 426 -731 438 -697
rect 178 -765 438 -731
rect 178 -799 190 -765
rect 224 -799 286 -765
rect 320 -799 392 -765
rect 426 -799 438 -765
rect 178 -833 438 -799
rect 178 -867 190 -833
rect 224 -867 286 -833
rect 320 -867 392 -833
rect 426 -867 438 -833
rect 178 -901 438 -867
rect 178 -935 190 -901
rect 224 -935 286 -901
rect 320 -935 392 -901
rect 426 -935 438 -901
rect 178 -969 438 -935
rect 178 -1003 190 -969
rect 224 -1003 286 -969
rect 320 -1003 392 -969
rect 426 -1003 438 -969
rect 178 -1037 438 -1003
rect 178 -1071 190 -1037
rect 224 -1071 286 -1037
rect 320 -1071 392 -1037
rect 426 -1071 438 -1037
rect 178 -1105 438 -1071
rect 178 -1139 190 -1105
rect 224 -1139 286 -1105
rect 320 -1139 392 -1105
rect 426 -1139 438 -1105
rect 178 -1173 438 -1139
rect 178 -1207 190 -1173
rect 224 -1207 286 -1173
rect 320 -1207 392 -1173
rect 426 -1207 438 -1173
rect 178 -1241 438 -1207
rect 178 -1275 190 -1241
rect 224 -1275 286 -1241
rect 320 -1275 392 -1241
rect 426 -1275 438 -1241
rect 178 -1309 438 -1275
rect 178 -1343 190 -1309
rect 224 -1343 286 -1309
rect 320 -1343 392 -1309
rect 426 -1343 438 -1309
rect 178 -1377 438 -1343
rect 178 -1411 190 -1377
rect 224 -1411 286 -1377
rect 320 -1411 392 -1377
rect 426 -1411 438 -1377
rect 178 -1445 438 -1411
rect 178 -1479 190 -1445
rect 224 -1479 286 -1445
rect 320 -1479 392 -1445
rect 426 -1479 438 -1445
rect 178 -1513 438 -1479
rect 178 -1547 190 -1513
rect 224 -1547 286 -1513
rect 320 -1547 392 -1513
rect 426 -1547 438 -1513
rect 178 -1581 438 -1547
rect 178 -1615 190 -1581
rect 224 -1615 286 -1581
rect 320 -1615 392 -1581
rect 426 -1615 438 -1581
rect 178 -1649 438 -1615
rect 178 -1683 190 -1649
rect 224 -1683 286 -1649
rect 320 -1683 392 -1649
rect 426 -1683 438 -1649
rect 178 -1717 438 -1683
rect 178 -1751 190 -1717
rect 224 -1751 286 -1717
rect 320 -1751 392 -1717
rect 426 -1751 438 -1717
rect 178 -1785 438 -1751
rect 178 -1819 190 -1785
rect 224 -1819 286 -1785
rect 320 -1819 392 -1785
rect 426 -1819 438 -1785
rect 178 -1853 438 -1819
rect 178 -1887 190 -1853
rect 224 -1887 286 -1853
rect 320 -1887 392 -1853
rect 426 -1887 438 -1853
rect 178 -1921 438 -1887
rect 178 -1955 190 -1921
rect 224 -1955 286 -1921
rect 320 -1955 392 -1921
rect 426 -1955 438 -1921
rect 178 -1989 438 -1955
rect 178 -2023 190 -1989
rect 224 -2023 286 -1989
rect 320 -2023 392 -1989
rect 426 -2023 438 -1989
rect 178 -2057 438 -2023
rect 178 -2091 190 -2057
rect 224 -2091 286 -2057
rect 320 -2091 392 -2057
rect 426 -2091 438 -2057
rect 178 -2125 438 -2091
rect 178 -2159 190 -2125
rect 224 -2159 286 -2125
rect 320 -2159 392 -2125
rect 426 -2159 438 -2125
rect 178 -2193 438 -2159
rect 178 -2227 190 -2193
rect 224 -2227 286 -2193
rect 320 -2227 392 -2193
rect 426 -2227 438 -2193
rect 178 -2261 438 -2227
rect 178 -2295 190 -2261
rect 224 -2295 286 -2261
rect 320 -2295 392 -2261
rect 426 -2295 438 -2261
rect 178 -2329 438 -2295
rect 178 -2363 190 -2329
rect 224 -2363 286 -2329
rect 320 -2363 392 -2329
rect 426 -2363 438 -2329
rect 178 -2397 438 -2363
rect 178 -2431 190 -2397
rect 224 -2431 286 -2397
rect 320 -2431 392 -2397
rect 426 -2431 438 -2397
rect 178 -2465 438 -2431
rect 178 -2499 190 -2465
rect 224 -2499 286 -2465
rect 320 -2499 392 -2465
rect 426 -2499 438 -2465
rect 178 -2533 438 -2499
rect 178 -2567 190 -2533
rect 224 -2567 286 -2533
rect 320 -2567 392 -2533
rect 426 -2567 438 -2533
rect 178 -2601 438 -2567
rect 178 -2635 190 -2601
rect 224 -2635 286 -2601
rect 320 -2635 392 -2601
rect 426 -2635 438 -2601
rect 178 -2669 438 -2635
rect 178 -2703 190 -2669
rect 224 -2703 286 -2669
rect 320 -2703 392 -2669
rect 426 -2703 438 -2669
rect 178 -2737 438 -2703
rect 178 -2771 190 -2737
rect 224 -2771 286 -2737
rect 320 -2771 392 -2737
rect 426 -2771 438 -2737
rect 178 -2805 438 -2771
rect 178 -2839 190 -2805
rect 224 -2839 286 -2805
rect 320 -2839 392 -2805
rect 426 -2839 438 -2805
rect 178 -2873 438 -2839
rect 178 -2907 190 -2873
rect 224 -2907 286 -2873
rect 320 -2907 392 -2873
rect 426 -2907 438 -2873
rect 178 -2941 438 -2907
rect 178 -2975 190 -2941
rect 224 -2975 286 -2941
rect 320 -2975 392 -2941
rect 426 -2975 438 -2941
rect 178 -3009 438 -2975
rect 178 -3043 190 -3009
rect 224 -3043 286 -3009
rect 320 -3043 392 -3009
rect 426 -3043 438 -3009
rect 178 -3077 438 -3043
rect 178 -3111 190 -3077
rect 224 -3111 286 -3077
rect 320 -3111 392 -3077
rect 426 -3111 438 -3077
rect 178 -3145 438 -3111
rect 178 -3179 190 -3145
rect 224 -3179 286 -3145
rect 320 -3179 392 -3145
rect 426 -3179 438 -3145
rect 178 -3213 438 -3179
rect 178 -3247 190 -3213
rect 224 -3247 286 -3213
rect 320 -3247 392 -3213
rect 426 -3247 438 -3213
rect 178 -3281 438 -3247
rect 178 -3315 190 -3281
rect 224 -3315 286 -3281
rect 320 -3315 392 -3281
rect 426 -3315 438 -3281
rect 178 -3349 438 -3315
rect 178 -3383 190 -3349
rect 224 -3383 286 -3349
rect 320 -3383 392 -3349
rect 426 -3383 438 -3349
rect 178 -3417 438 -3383
rect 178 -3451 190 -3417
rect 224 -3451 286 -3417
rect 320 -3451 392 -3417
rect 426 -3451 438 -3417
rect 178 -3485 438 -3451
rect 178 -3519 190 -3485
rect 224 -3519 286 -3485
rect 320 -3519 392 -3485
rect 426 -3519 438 -3485
rect 178 -3553 438 -3519
rect 178 -3587 190 -3553
rect 224 -3587 286 -3553
rect 320 -3587 392 -3553
rect 426 -3587 438 -3553
rect 178 -3621 438 -3587
rect 178 -3655 190 -3621
rect 224 -3655 286 -3621
rect 320 -3655 392 -3621
rect 426 -3655 438 -3621
rect 178 -3689 438 -3655
rect 178 -3723 190 -3689
rect 224 -3723 286 -3689
rect 320 -3723 392 -3689
rect 426 -3723 438 -3689
rect 178 -3757 438 -3723
rect 178 -3791 190 -3757
rect 224 -3791 286 -3757
rect 320 -3791 392 -3757
rect 426 -3791 438 -3757
rect 178 -3825 438 -3791
rect 178 -3859 190 -3825
rect 224 -3859 286 -3825
rect 320 -3859 392 -3825
rect 426 -3859 438 -3825
rect 178 -3893 438 -3859
rect 178 -3927 190 -3893
rect 224 -3927 286 -3893
rect 320 -3927 392 -3893
rect 426 -3927 438 -3893
rect 178 -3961 438 -3927
rect 178 -3995 190 -3961
rect 224 -3995 286 -3961
rect 320 -3995 392 -3961
rect 426 -3995 438 -3961
rect 178 -4029 438 -3995
rect 178 -4063 190 -4029
rect 224 -4063 286 -4029
rect 320 -4063 392 -4029
rect 426 -4063 438 -4029
rect 178 -4097 438 -4063
rect 178 -4131 190 -4097
rect 224 -4131 286 -4097
rect 320 -4131 392 -4097
rect 426 -4131 438 -4097
rect 178 -4165 438 -4131
rect 178 -4199 190 -4165
rect 224 -4199 286 -4165
rect 320 -4199 392 -4165
rect 426 -4199 438 -4165
rect 178 -4233 438 -4199
rect 178 -4267 190 -4233
rect 224 -4267 286 -4233
rect 320 -4267 392 -4233
rect 426 -4267 438 -4233
rect 178 -4301 438 -4267
rect 178 -4335 190 -4301
rect 224 -4335 286 -4301
rect 320 -4335 392 -4301
rect 426 -4335 438 -4301
rect 178 -4369 438 -4335
rect 178 -4403 190 -4369
rect 224 -4403 286 -4369
rect 320 -4403 392 -4369
rect 426 -4403 438 -4369
rect 178 -4437 438 -4403
rect 178 -4471 190 -4437
rect 224 -4471 286 -4437
rect 320 -4471 392 -4437
rect 426 -4471 438 -4437
rect 178 -4505 438 -4471
rect 178 -4539 190 -4505
rect 224 -4539 286 -4505
rect 320 -4539 392 -4505
rect 426 -4539 438 -4505
rect 178 -4573 438 -4539
rect 178 -4607 190 -4573
rect 224 -4607 286 -4573
rect 320 -4607 392 -4573
rect 426 -4607 438 -4573
rect 178 -4641 438 -4607
rect 178 -4675 190 -4641
rect 224 -4675 286 -4641
rect 320 -4675 392 -4641
rect 426 -4675 438 -4641
rect 178 -4709 438 -4675
rect 178 -4743 190 -4709
rect 224 -4743 286 -4709
rect 320 -4743 392 -4709
rect 426 -4743 438 -4709
rect 178 -4777 438 -4743
rect 178 -4811 190 -4777
rect 224 -4811 286 -4777
rect 320 -4811 392 -4777
rect 426 -4811 438 -4777
rect 178 -4845 438 -4811
rect 178 -4879 190 -4845
rect 224 -4879 286 -4845
rect 320 -4879 392 -4845
rect 426 -4879 438 -4845
rect 178 -4913 438 -4879
rect 178 -4947 190 -4913
rect 224 -4947 286 -4913
rect 320 -4947 392 -4913
rect 426 -4947 438 -4913
rect 178 -4981 438 -4947
rect -438 -5078 -178 -5015
rect 178 -5015 190 -4981
rect 224 -5015 286 -4981
rect 320 -5015 392 -4981
rect 426 -5015 438 -4981
rect 794 4981 806 5015
rect 840 4981 902 5015
rect 936 4981 1008 5015
rect 1042 4981 1054 5015
rect 1410 5015 1540 5078
rect 794 4947 1054 4981
rect 794 4913 806 4947
rect 840 4913 902 4947
rect 936 4913 1008 4947
rect 1042 4913 1054 4947
rect 794 4879 1054 4913
rect 794 4845 806 4879
rect 840 4845 902 4879
rect 936 4845 1008 4879
rect 1042 4845 1054 4879
rect 794 4811 1054 4845
rect 794 4777 806 4811
rect 840 4777 902 4811
rect 936 4777 1008 4811
rect 1042 4777 1054 4811
rect 794 4743 1054 4777
rect 794 4709 806 4743
rect 840 4709 902 4743
rect 936 4709 1008 4743
rect 1042 4709 1054 4743
rect 794 4675 1054 4709
rect 794 4641 806 4675
rect 840 4641 902 4675
rect 936 4641 1008 4675
rect 1042 4641 1054 4675
rect 794 4607 1054 4641
rect 794 4573 806 4607
rect 840 4573 902 4607
rect 936 4573 1008 4607
rect 1042 4573 1054 4607
rect 794 4539 1054 4573
rect 794 4505 806 4539
rect 840 4505 902 4539
rect 936 4505 1008 4539
rect 1042 4505 1054 4539
rect 794 4471 1054 4505
rect 794 4437 806 4471
rect 840 4437 902 4471
rect 936 4437 1008 4471
rect 1042 4437 1054 4471
rect 794 4403 1054 4437
rect 794 4369 806 4403
rect 840 4369 902 4403
rect 936 4369 1008 4403
rect 1042 4369 1054 4403
rect 794 4335 1054 4369
rect 794 4301 806 4335
rect 840 4301 902 4335
rect 936 4301 1008 4335
rect 1042 4301 1054 4335
rect 794 4267 1054 4301
rect 794 4233 806 4267
rect 840 4233 902 4267
rect 936 4233 1008 4267
rect 1042 4233 1054 4267
rect 794 4199 1054 4233
rect 794 4165 806 4199
rect 840 4165 902 4199
rect 936 4165 1008 4199
rect 1042 4165 1054 4199
rect 794 4131 1054 4165
rect 794 4097 806 4131
rect 840 4097 902 4131
rect 936 4097 1008 4131
rect 1042 4097 1054 4131
rect 794 4063 1054 4097
rect 794 4029 806 4063
rect 840 4029 902 4063
rect 936 4029 1008 4063
rect 1042 4029 1054 4063
rect 794 3995 1054 4029
rect 794 3961 806 3995
rect 840 3961 902 3995
rect 936 3961 1008 3995
rect 1042 3961 1054 3995
rect 794 3927 1054 3961
rect 794 3893 806 3927
rect 840 3893 902 3927
rect 936 3893 1008 3927
rect 1042 3893 1054 3927
rect 794 3859 1054 3893
rect 794 3825 806 3859
rect 840 3825 902 3859
rect 936 3825 1008 3859
rect 1042 3825 1054 3859
rect 794 3791 1054 3825
rect 794 3757 806 3791
rect 840 3757 902 3791
rect 936 3757 1008 3791
rect 1042 3757 1054 3791
rect 794 3723 1054 3757
rect 794 3689 806 3723
rect 840 3689 902 3723
rect 936 3689 1008 3723
rect 1042 3689 1054 3723
rect 794 3655 1054 3689
rect 794 3621 806 3655
rect 840 3621 902 3655
rect 936 3621 1008 3655
rect 1042 3621 1054 3655
rect 794 3587 1054 3621
rect 794 3553 806 3587
rect 840 3553 902 3587
rect 936 3553 1008 3587
rect 1042 3553 1054 3587
rect 794 3519 1054 3553
rect 794 3485 806 3519
rect 840 3485 902 3519
rect 936 3485 1008 3519
rect 1042 3485 1054 3519
rect 794 3451 1054 3485
rect 794 3417 806 3451
rect 840 3417 902 3451
rect 936 3417 1008 3451
rect 1042 3417 1054 3451
rect 794 3383 1054 3417
rect 794 3349 806 3383
rect 840 3349 902 3383
rect 936 3349 1008 3383
rect 1042 3349 1054 3383
rect 794 3315 1054 3349
rect 794 3281 806 3315
rect 840 3281 902 3315
rect 936 3281 1008 3315
rect 1042 3281 1054 3315
rect 794 3247 1054 3281
rect 794 3213 806 3247
rect 840 3213 902 3247
rect 936 3213 1008 3247
rect 1042 3213 1054 3247
rect 794 3179 1054 3213
rect 794 3145 806 3179
rect 840 3145 902 3179
rect 936 3145 1008 3179
rect 1042 3145 1054 3179
rect 794 3111 1054 3145
rect 794 3077 806 3111
rect 840 3077 902 3111
rect 936 3077 1008 3111
rect 1042 3077 1054 3111
rect 794 3043 1054 3077
rect 794 3009 806 3043
rect 840 3009 902 3043
rect 936 3009 1008 3043
rect 1042 3009 1054 3043
rect 794 2975 1054 3009
rect 794 2941 806 2975
rect 840 2941 902 2975
rect 936 2941 1008 2975
rect 1042 2941 1054 2975
rect 794 2907 1054 2941
rect 794 2873 806 2907
rect 840 2873 902 2907
rect 936 2873 1008 2907
rect 1042 2873 1054 2907
rect 794 2839 1054 2873
rect 794 2805 806 2839
rect 840 2805 902 2839
rect 936 2805 1008 2839
rect 1042 2805 1054 2839
rect 794 2771 1054 2805
rect 794 2737 806 2771
rect 840 2737 902 2771
rect 936 2737 1008 2771
rect 1042 2737 1054 2771
rect 794 2703 1054 2737
rect 794 2669 806 2703
rect 840 2669 902 2703
rect 936 2669 1008 2703
rect 1042 2669 1054 2703
rect 794 2635 1054 2669
rect 794 2601 806 2635
rect 840 2601 902 2635
rect 936 2601 1008 2635
rect 1042 2601 1054 2635
rect 794 2567 1054 2601
rect 794 2533 806 2567
rect 840 2533 902 2567
rect 936 2533 1008 2567
rect 1042 2533 1054 2567
rect 794 2499 1054 2533
rect 794 2465 806 2499
rect 840 2465 902 2499
rect 936 2465 1008 2499
rect 1042 2465 1054 2499
rect 794 2431 1054 2465
rect 794 2397 806 2431
rect 840 2397 902 2431
rect 936 2397 1008 2431
rect 1042 2397 1054 2431
rect 794 2363 1054 2397
rect 794 2329 806 2363
rect 840 2329 902 2363
rect 936 2329 1008 2363
rect 1042 2329 1054 2363
rect 794 2295 1054 2329
rect 794 2261 806 2295
rect 840 2261 902 2295
rect 936 2261 1008 2295
rect 1042 2261 1054 2295
rect 794 2227 1054 2261
rect 794 2193 806 2227
rect 840 2193 902 2227
rect 936 2193 1008 2227
rect 1042 2193 1054 2227
rect 794 2159 1054 2193
rect 794 2125 806 2159
rect 840 2125 902 2159
rect 936 2125 1008 2159
rect 1042 2125 1054 2159
rect 794 2091 1054 2125
rect 794 2057 806 2091
rect 840 2057 902 2091
rect 936 2057 1008 2091
rect 1042 2057 1054 2091
rect 794 2023 1054 2057
rect 794 1989 806 2023
rect 840 1989 902 2023
rect 936 1989 1008 2023
rect 1042 1989 1054 2023
rect 794 1955 1054 1989
rect 794 1921 806 1955
rect 840 1921 902 1955
rect 936 1921 1008 1955
rect 1042 1921 1054 1955
rect 794 1887 1054 1921
rect 794 1853 806 1887
rect 840 1853 902 1887
rect 936 1853 1008 1887
rect 1042 1853 1054 1887
rect 794 1819 1054 1853
rect 794 1785 806 1819
rect 840 1785 902 1819
rect 936 1785 1008 1819
rect 1042 1785 1054 1819
rect 794 1751 1054 1785
rect 794 1717 806 1751
rect 840 1717 902 1751
rect 936 1717 1008 1751
rect 1042 1717 1054 1751
rect 794 1683 1054 1717
rect 794 1649 806 1683
rect 840 1649 902 1683
rect 936 1649 1008 1683
rect 1042 1649 1054 1683
rect 794 1615 1054 1649
rect 794 1581 806 1615
rect 840 1581 902 1615
rect 936 1581 1008 1615
rect 1042 1581 1054 1615
rect 794 1547 1054 1581
rect 794 1513 806 1547
rect 840 1513 902 1547
rect 936 1513 1008 1547
rect 1042 1513 1054 1547
rect 794 1479 1054 1513
rect 794 1445 806 1479
rect 840 1445 902 1479
rect 936 1445 1008 1479
rect 1042 1445 1054 1479
rect 794 1411 1054 1445
rect 794 1377 806 1411
rect 840 1377 902 1411
rect 936 1377 1008 1411
rect 1042 1377 1054 1411
rect 794 1343 1054 1377
rect 794 1309 806 1343
rect 840 1309 902 1343
rect 936 1309 1008 1343
rect 1042 1309 1054 1343
rect 794 1275 1054 1309
rect 794 1241 806 1275
rect 840 1241 902 1275
rect 936 1241 1008 1275
rect 1042 1241 1054 1275
rect 794 1207 1054 1241
rect 794 1173 806 1207
rect 840 1173 902 1207
rect 936 1173 1008 1207
rect 1042 1173 1054 1207
rect 794 1139 1054 1173
rect 794 1105 806 1139
rect 840 1105 902 1139
rect 936 1105 1008 1139
rect 1042 1105 1054 1139
rect 794 1071 1054 1105
rect 794 1037 806 1071
rect 840 1037 902 1071
rect 936 1037 1008 1071
rect 1042 1037 1054 1071
rect 794 1003 1054 1037
rect 794 969 806 1003
rect 840 969 902 1003
rect 936 969 1008 1003
rect 1042 969 1054 1003
rect 794 935 1054 969
rect 794 901 806 935
rect 840 901 902 935
rect 936 901 1008 935
rect 1042 901 1054 935
rect 794 867 1054 901
rect 794 833 806 867
rect 840 833 902 867
rect 936 833 1008 867
rect 1042 833 1054 867
rect 794 799 1054 833
rect 794 765 806 799
rect 840 765 902 799
rect 936 765 1008 799
rect 1042 765 1054 799
rect 794 731 1054 765
rect 794 697 806 731
rect 840 697 902 731
rect 936 697 1008 731
rect 1042 697 1054 731
rect 794 663 1054 697
rect 794 629 806 663
rect 840 629 902 663
rect 936 629 1008 663
rect 1042 629 1054 663
rect 794 595 1054 629
rect 794 561 806 595
rect 840 561 902 595
rect 936 561 1008 595
rect 1042 561 1054 595
rect 794 527 1054 561
rect 794 493 806 527
rect 840 493 902 527
rect 936 493 1008 527
rect 1042 493 1054 527
rect 794 459 1054 493
rect 794 425 806 459
rect 840 425 902 459
rect 936 425 1008 459
rect 1042 425 1054 459
rect 794 391 1054 425
rect 794 357 806 391
rect 840 357 902 391
rect 936 357 1008 391
rect 1042 357 1054 391
rect 794 323 1054 357
rect 794 289 806 323
rect 840 289 902 323
rect 936 289 1008 323
rect 1042 289 1054 323
rect 794 255 1054 289
rect 794 221 806 255
rect 840 221 902 255
rect 936 221 1008 255
rect 1042 221 1054 255
rect 794 187 1054 221
rect 794 153 806 187
rect 840 153 902 187
rect 936 153 1008 187
rect 1042 153 1054 187
rect 794 119 1054 153
rect 794 85 806 119
rect 840 85 902 119
rect 936 85 1008 119
rect 1042 85 1054 119
rect 794 51 1054 85
rect 794 17 806 51
rect 840 17 902 51
rect 936 17 1008 51
rect 1042 17 1054 51
rect 794 -17 1054 17
rect 794 -51 806 -17
rect 840 -51 902 -17
rect 936 -51 1008 -17
rect 1042 -51 1054 -17
rect 794 -85 1054 -51
rect 794 -119 806 -85
rect 840 -119 902 -85
rect 936 -119 1008 -85
rect 1042 -119 1054 -85
rect 794 -153 1054 -119
rect 794 -187 806 -153
rect 840 -187 902 -153
rect 936 -187 1008 -153
rect 1042 -187 1054 -153
rect 794 -221 1054 -187
rect 794 -255 806 -221
rect 840 -255 902 -221
rect 936 -255 1008 -221
rect 1042 -255 1054 -221
rect 794 -289 1054 -255
rect 794 -323 806 -289
rect 840 -323 902 -289
rect 936 -323 1008 -289
rect 1042 -323 1054 -289
rect 794 -357 1054 -323
rect 794 -391 806 -357
rect 840 -391 902 -357
rect 936 -391 1008 -357
rect 1042 -391 1054 -357
rect 794 -425 1054 -391
rect 794 -459 806 -425
rect 840 -459 902 -425
rect 936 -459 1008 -425
rect 1042 -459 1054 -425
rect 794 -493 1054 -459
rect 794 -527 806 -493
rect 840 -527 902 -493
rect 936 -527 1008 -493
rect 1042 -527 1054 -493
rect 794 -561 1054 -527
rect 794 -595 806 -561
rect 840 -595 902 -561
rect 936 -595 1008 -561
rect 1042 -595 1054 -561
rect 794 -629 1054 -595
rect 794 -663 806 -629
rect 840 -663 902 -629
rect 936 -663 1008 -629
rect 1042 -663 1054 -629
rect 794 -697 1054 -663
rect 794 -731 806 -697
rect 840 -731 902 -697
rect 936 -731 1008 -697
rect 1042 -731 1054 -697
rect 794 -765 1054 -731
rect 794 -799 806 -765
rect 840 -799 902 -765
rect 936 -799 1008 -765
rect 1042 -799 1054 -765
rect 794 -833 1054 -799
rect 794 -867 806 -833
rect 840 -867 902 -833
rect 936 -867 1008 -833
rect 1042 -867 1054 -833
rect 794 -901 1054 -867
rect 794 -935 806 -901
rect 840 -935 902 -901
rect 936 -935 1008 -901
rect 1042 -935 1054 -901
rect 794 -969 1054 -935
rect 794 -1003 806 -969
rect 840 -1003 902 -969
rect 936 -1003 1008 -969
rect 1042 -1003 1054 -969
rect 794 -1037 1054 -1003
rect 794 -1071 806 -1037
rect 840 -1071 902 -1037
rect 936 -1071 1008 -1037
rect 1042 -1071 1054 -1037
rect 794 -1105 1054 -1071
rect 794 -1139 806 -1105
rect 840 -1139 902 -1105
rect 936 -1139 1008 -1105
rect 1042 -1139 1054 -1105
rect 794 -1173 1054 -1139
rect 794 -1207 806 -1173
rect 840 -1207 902 -1173
rect 936 -1207 1008 -1173
rect 1042 -1207 1054 -1173
rect 794 -1241 1054 -1207
rect 794 -1275 806 -1241
rect 840 -1275 902 -1241
rect 936 -1275 1008 -1241
rect 1042 -1275 1054 -1241
rect 794 -1309 1054 -1275
rect 794 -1343 806 -1309
rect 840 -1343 902 -1309
rect 936 -1343 1008 -1309
rect 1042 -1343 1054 -1309
rect 794 -1377 1054 -1343
rect 794 -1411 806 -1377
rect 840 -1411 902 -1377
rect 936 -1411 1008 -1377
rect 1042 -1411 1054 -1377
rect 794 -1445 1054 -1411
rect 794 -1479 806 -1445
rect 840 -1479 902 -1445
rect 936 -1479 1008 -1445
rect 1042 -1479 1054 -1445
rect 794 -1513 1054 -1479
rect 794 -1547 806 -1513
rect 840 -1547 902 -1513
rect 936 -1547 1008 -1513
rect 1042 -1547 1054 -1513
rect 794 -1581 1054 -1547
rect 794 -1615 806 -1581
rect 840 -1615 902 -1581
rect 936 -1615 1008 -1581
rect 1042 -1615 1054 -1581
rect 794 -1649 1054 -1615
rect 794 -1683 806 -1649
rect 840 -1683 902 -1649
rect 936 -1683 1008 -1649
rect 1042 -1683 1054 -1649
rect 794 -1717 1054 -1683
rect 794 -1751 806 -1717
rect 840 -1751 902 -1717
rect 936 -1751 1008 -1717
rect 1042 -1751 1054 -1717
rect 794 -1785 1054 -1751
rect 794 -1819 806 -1785
rect 840 -1819 902 -1785
rect 936 -1819 1008 -1785
rect 1042 -1819 1054 -1785
rect 794 -1853 1054 -1819
rect 794 -1887 806 -1853
rect 840 -1887 902 -1853
rect 936 -1887 1008 -1853
rect 1042 -1887 1054 -1853
rect 794 -1921 1054 -1887
rect 794 -1955 806 -1921
rect 840 -1955 902 -1921
rect 936 -1955 1008 -1921
rect 1042 -1955 1054 -1921
rect 794 -1989 1054 -1955
rect 794 -2023 806 -1989
rect 840 -2023 902 -1989
rect 936 -2023 1008 -1989
rect 1042 -2023 1054 -1989
rect 794 -2057 1054 -2023
rect 794 -2091 806 -2057
rect 840 -2091 902 -2057
rect 936 -2091 1008 -2057
rect 1042 -2091 1054 -2057
rect 794 -2125 1054 -2091
rect 794 -2159 806 -2125
rect 840 -2159 902 -2125
rect 936 -2159 1008 -2125
rect 1042 -2159 1054 -2125
rect 794 -2193 1054 -2159
rect 794 -2227 806 -2193
rect 840 -2227 902 -2193
rect 936 -2227 1008 -2193
rect 1042 -2227 1054 -2193
rect 794 -2261 1054 -2227
rect 794 -2295 806 -2261
rect 840 -2295 902 -2261
rect 936 -2295 1008 -2261
rect 1042 -2295 1054 -2261
rect 794 -2329 1054 -2295
rect 794 -2363 806 -2329
rect 840 -2363 902 -2329
rect 936 -2363 1008 -2329
rect 1042 -2363 1054 -2329
rect 794 -2397 1054 -2363
rect 794 -2431 806 -2397
rect 840 -2431 902 -2397
rect 936 -2431 1008 -2397
rect 1042 -2431 1054 -2397
rect 794 -2465 1054 -2431
rect 794 -2499 806 -2465
rect 840 -2499 902 -2465
rect 936 -2499 1008 -2465
rect 1042 -2499 1054 -2465
rect 794 -2533 1054 -2499
rect 794 -2567 806 -2533
rect 840 -2567 902 -2533
rect 936 -2567 1008 -2533
rect 1042 -2567 1054 -2533
rect 794 -2601 1054 -2567
rect 794 -2635 806 -2601
rect 840 -2635 902 -2601
rect 936 -2635 1008 -2601
rect 1042 -2635 1054 -2601
rect 794 -2669 1054 -2635
rect 794 -2703 806 -2669
rect 840 -2703 902 -2669
rect 936 -2703 1008 -2669
rect 1042 -2703 1054 -2669
rect 794 -2737 1054 -2703
rect 794 -2771 806 -2737
rect 840 -2771 902 -2737
rect 936 -2771 1008 -2737
rect 1042 -2771 1054 -2737
rect 794 -2805 1054 -2771
rect 794 -2839 806 -2805
rect 840 -2839 902 -2805
rect 936 -2839 1008 -2805
rect 1042 -2839 1054 -2805
rect 794 -2873 1054 -2839
rect 794 -2907 806 -2873
rect 840 -2907 902 -2873
rect 936 -2907 1008 -2873
rect 1042 -2907 1054 -2873
rect 794 -2941 1054 -2907
rect 794 -2975 806 -2941
rect 840 -2975 902 -2941
rect 936 -2975 1008 -2941
rect 1042 -2975 1054 -2941
rect 794 -3009 1054 -2975
rect 794 -3043 806 -3009
rect 840 -3043 902 -3009
rect 936 -3043 1008 -3009
rect 1042 -3043 1054 -3009
rect 794 -3077 1054 -3043
rect 794 -3111 806 -3077
rect 840 -3111 902 -3077
rect 936 -3111 1008 -3077
rect 1042 -3111 1054 -3077
rect 794 -3145 1054 -3111
rect 794 -3179 806 -3145
rect 840 -3179 902 -3145
rect 936 -3179 1008 -3145
rect 1042 -3179 1054 -3145
rect 794 -3213 1054 -3179
rect 794 -3247 806 -3213
rect 840 -3247 902 -3213
rect 936 -3247 1008 -3213
rect 1042 -3247 1054 -3213
rect 794 -3281 1054 -3247
rect 794 -3315 806 -3281
rect 840 -3315 902 -3281
rect 936 -3315 1008 -3281
rect 1042 -3315 1054 -3281
rect 794 -3349 1054 -3315
rect 794 -3383 806 -3349
rect 840 -3383 902 -3349
rect 936 -3383 1008 -3349
rect 1042 -3383 1054 -3349
rect 794 -3417 1054 -3383
rect 794 -3451 806 -3417
rect 840 -3451 902 -3417
rect 936 -3451 1008 -3417
rect 1042 -3451 1054 -3417
rect 794 -3485 1054 -3451
rect 794 -3519 806 -3485
rect 840 -3519 902 -3485
rect 936 -3519 1008 -3485
rect 1042 -3519 1054 -3485
rect 794 -3553 1054 -3519
rect 794 -3587 806 -3553
rect 840 -3587 902 -3553
rect 936 -3587 1008 -3553
rect 1042 -3587 1054 -3553
rect 794 -3621 1054 -3587
rect 794 -3655 806 -3621
rect 840 -3655 902 -3621
rect 936 -3655 1008 -3621
rect 1042 -3655 1054 -3621
rect 794 -3689 1054 -3655
rect 794 -3723 806 -3689
rect 840 -3723 902 -3689
rect 936 -3723 1008 -3689
rect 1042 -3723 1054 -3689
rect 794 -3757 1054 -3723
rect 794 -3791 806 -3757
rect 840 -3791 902 -3757
rect 936 -3791 1008 -3757
rect 1042 -3791 1054 -3757
rect 794 -3825 1054 -3791
rect 794 -3859 806 -3825
rect 840 -3859 902 -3825
rect 936 -3859 1008 -3825
rect 1042 -3859 1054 -3825
rect 794 -3893 1054 -3859
rect 794 -3927 806 -3893
rect 840 -3927 902 -3893
rect 936 -3927 1008 -3893
rect 1042 -3927 1054 -3893
rect 794 -3961 1054 -3927
rect 794 -3995 806 -3961
rect 840 -3995 902 -3961
rect 936 -3995 1008 -3961
rect 1042 -3995 1054 -3961
rect 794 -4029 1054 -3995
rect 794 -4063 806 -4029
rect 840 -4063 902 -4029
rect 936 -4063 1008 -4029
rect 1042 -4063 1054 -4029
rect 794 -4097 1054 -4063
rect 794 -4131 806 -4097
rect 840 -4131 902 -4097
rect 936 -4131 1008 -4097
rect 1042 -4131 1054 -4097
rect 794 -4165 1054 -4131
rect 794 -4199 806 -4165
rect 840 -4199 902 -4165
rect 936 -4199 1008 -4165
rect 1042 -4199 1054 -4165
rect 794 -4233 1054 -4199
rect 794 -4267 806 -4233
rect 840 -4267 902 -4233
rect 936 -4267 1008 -4233
rect 1042 -4267 1054 -4233
rect 794 -4301 1054 -4267
rect 794 -4335 806 -4301
rect 840 -4335 902 -4301
rect 936 -4335 1008 -4301
rect 1042 -4335 1054 -4301
rect 794 -4369 1054 -4335
rect 794 -4403 806 -4369
rect 840 -4403 902 -4369
rect 936 -4403 1008 -4369
rect 1042 -4403 1054 -4369
rect 794 -4437 1054 -4403
rect 794 -4471 806 -4437
rect 840 -4471 902 -4437
rect 936 -4471 1008 -4437
rect 1042 -4471 1054 -4437
rect 794 -4505 1054 -4471
rect 794 -4539 806 -4505
rect 840 -4539 902 -4505
rect 936 -4539 1008 -4505
rect 1042 -4539 1054 -4505
rect 794 -4573 1054 -4539
rect 794 -4607 806 -4573
rect 840 -4607 902 -4573
rect 936 -4607 1008 -4573
rect 1042 -4607 1054 -4573
rect 794 -4641 1054 -4607
rect 794 -4675 806 -4641
rect 840 -4675 902 -4641
rect 936 -4675 1008 -4641
rect 1042 -4675 1054 -4641
rect 794 -4709 1054 -4675
rect 794 -4743 806 -4709
rect 840 -4743 902 -4709
rect 936 -4743 1008 -4709
rect 1042 -4743 1054 -4709
rect 794 -4777 1054 -4743
rect 794 -4811 806 -4777
rect 840 -4811 902 -4777
rect 936 -4811 1008 -4777
rect 1042 -4811 1054 -4777
rect 794 -4845 1054 -4811
rect 794 -4879 806 -4845
rect 840 -4879 902 -4845
rect 936 -4879 1008 -4845
rect 1042 -4879 1054 -4845
rect 794 -4913 1054 -4879
rect 794 -4947 806 -4913
rect 840 -4947 902 -4913
rect 936 -4947 1008 -4913
rect 1042 -4947 1054 -4913
rect 794 -4981 1054 -4947
rect 178 -5078 438 -5015
rect 794 -5015 806 -4981
rect 840 -5015 902 -4981
rect 936 -5015 1008 -4981
rect 1042 -5015 1054 -4981
rect 794 -5078 1054 -5015
rect 1410 -5015 1422 5015
rect 1524 -5015 1540 5015
rect 1410 -5078 1540 -5015
rect -1540 -5090 1540 -5078
rect -1540 -5124 -1351 -5090
rect -1317 -5124 -1283 -5090
rect -1249 -5124 -1215 -5090
rect -1181 -5124 -1147 -5090
rect -1113 -5124 -735 -5090
rect -701 -5124 -667 -5090
rect -633 -5124 -599 -5090
rect -565 -5124 -531 -5090
rect -497 -5124 -119 -5090
rect -85 -5124 -51 -5090
rect -17 -5124 17 -5090
rect 51 -5124 85 -5090
rect 119 -5124 497 -5090
rect 531 -5124 565 -5090
rect 599 -5124 633 -5090
rect 667 -5124 701 -5090
rect 735 -5124 1113 -5090
rect 1147 -5124 1181 -5090
rect 1215 -5124 1249 -5090
rect 1283 -5124 1317 -5090
rect 1351 -5124 1540 -5090
rect -1540 -5136 1540 -5124
<< mvpsubdiffcont >>
rect -1351 5090 -1317 5124
rect -1283 5090 -1249 5124
rect -1215 5090 -1181 5124
rect -1147 5090 -1113 5124
rect -735 5090 -701 5124
rect -667 5090 -633 5124
rect -599 5090 -565 5124
rect -531 5090 -497 5124
rect -119 5090 -85 5124
rect -51 5090 -17 5124
rect 17 5090 51 5124
rect 85 5090 119 5124
rect 497 5090 531 5124
rect 565 5090 599 5124
rect 633 5090 667 5124
rect 701 5090 735 5124
rect 1113 5090 1147 5124
rect 1181 5090 1215 5124
rect 1249 5090 1283 5124
rect 1317 5090 1351 5124
rect -1524 -5015 -1422 5015
rect -1042 4981 -1008 5015
rect -946 4981 -912 5015
rect -840 4981 -806 5015
rect -1042 4913 -1008 4947
rect -946 4913 -912 4947
rect -840 4913 -806 4947
rect -1042 4845 -1008 4879
rect -946 4845 -912 4879
rect -840 4845 -806 4879
rect -1042 4777 -1008 4811
rect -946 4777 -912 4811
rect -840 4777 -806 4811
rect -1042 4709 -1008 4743
rect -946 4709 -912 4743
rect -840 4709 -806 4743
rect -1042 4641 -1008 4675
rect -946 4641 -912 4675
rect -840 4641 -806 4675
rect -1042 4573 -1008 4607
rect -946 4573 -912 4607
rect -840 4573 -806 4607
rect -1042 4505 -1008 4539
rect -946 4505 -912 4539
rect -840 4505 -806 4539
rect -1042 4437 -1008 4471
rect -946 4437 -912 4471
rect -840 4437 -806 4471
rect -1042 4369 -1008 4403
rect -946 4369 -912 4403
rect -840 4369 -806 4403
rect -1042 4301 -1008 4335
rect -946 4301 -912 4335
rect -840 4301 -806 4335
rect -1042 4233 -1008 4267
rect -946 4233 -912 4267
rect -840 4233 -806 4267
rect -1042 4165 -1008 4199
rect -946 4165 -912 4199
rect -840 4165 -806 4199
rect -1042 4097 -1008 4131
rect -946 4097 -912 4131
rect -840 4097 -806 4131
rect -1042 4029 -1008 4063
rect -946 4029 -912 4063
rect -840 4029 -806 4063
rect -1042 3961 -1008 3995
rect -946 3961 -912 3995
rect -840 3961 -806 3995
rect -1042 3893 -1008 3927
rect -946 3893 -912 3927
rect -840 3893 -806 3927
rect -1042 3825 -1008 3859
rect -946 3825 -912 3859
rect -840 3825 -806 3859
rect -1042 3757 -1008 3791
rect -946 3757 -912 3791
rect -840 3757 -806 3791
rect -1042 3689 -1008 3723
rect -946 3689 -912 3723
rect -840 3689 -806 3723
rect -1042 3621 -1008 3655
rect -946 3621 -912 3655
rect -840 3621 -806 3655
rect -1042 3553 -1008 3587
rect -946 3553 -912 3587
rect -840 3553 -806 3587
rect -1042 3485 -1008 3519
rect -946 3485 -912 3519
rect -840 3485 -806 3519
rect -1042 3417 -1008 3451
rect -946 3417 -912 3451
rect -840 3417 -806 3451
rect -1042 3349 -1008 3383
rect -946 3349 -912 3383
rect -840 3349 -806 3383
rect -1042 3281 -1008 3315
rect -946 3281 -912 3315
rect -840 3281 -806 3315
rect -1042 3213 -1008 3247
rect -946 3213 -912 3247
rect -840 3213 -806 3247
rect -1042 3145 -1008 3179
rect -946 3145 -912 3179
rect -840 3145 -806 3179
rect -1042 3077 -1008 3111
rect -946 3077 -912 3111
rect -840 3077 -806 3111
rect -1042 3009 -1008 3043
rect -946 3009 -912 3043
rect -840 3009 -806 3043
rect -1042 2941 -1008 2975
rect -946 2941 -912 2975
rect -840 2941 -806 2975
rect -1042 2873 -1008 2907
rect -946 2873 -912 2907
rect -840 2873 -806 2907
rect -1042 2805 -1008 2839
rect -946 2805 -912 2839
rect -840 2805 -806 2839
rect -1042 2737 -1008 2771
rect -946 2737 -912 2771
rect -840 2737 -806 2771
rect -1042 2669 -1008 2703
rect -946 2669 -912 2703
rect -840 2669 -806 2703
rect -1042 2601 -1008 2635
rect -946 2601 -912 2635
rect -840 2601 -806 2635
rect -1042 2533 -1008 2567
rect -946 2533 -912 2567
rect -840 2533 -806 2567
rect -1042 2465 -1008 2499
rect -946 2465 -912 2499
rect -840 2465 -806 2499
rect -1042 2397 -1008 2431
rect -946 2397 -912 2431
rect -840 2397 -806 2431
rect -1042 2329 -1008 2363
rect -946 2329 -912 2363
rect -840 2329 -806 2363
rect -1042 2261 -1008 2295
rect -946 2261 -912 2295
rect -840 2261 -806 2295
rect -1042 2193 -1008 2227
rect -946 2193 -912 2227
rect -840 2193 -806 2227
rect -1042 2125 -1008 2159
rect -946 2125 -912 2159
rect -840 2125 -806 2159
rect -1042 2057 -1008 2091
rect -946 2057 -912 2091
rect -840 2057 -806 2091
rect -1042 1989 -1008 2023
rect -946 1989 -912 2023
rect -840 1989 -806 2023
rect -1042 1921 -1008 1955
rect -946 1921 -912 1955
rect -840 1921 -806 1955
rect -1042 1853 -1008 1887
rect -946 1853 -912 1887
rect -840 1853 -806 1887
rect -1042 1785 -1008 1819
rect -946 1785 -912 1819
rect -840 1785 -806 1819
rect -1042 1717 -1008 1751
rect -946 1717 -912 1751
rect -840 1717 -806 1751
rect -1042 1649 -1008 1683
rect -946 1649 -912 1683
rect -840 1649 -806 1683
rect -1042 1581 -1008 1615
rect -946 1581 -912 1615
rect -840 1581 -806 1615
rect -1042 1513 -1008 1547
rect -946 1513 -912 1547
rect -840 1513 -806 1547
rect -1042 1445 -1008 1479
rect -946 1445 -912 1479
rect -840 1445 -806 1479
rect -1042 1377 -1008 1411
rect -946 1377 -912 1411
rect -840 1377 -806 1411
rect -1042 1309 -1008 1343
rect -946 1309 -912 1343
rect -840 1309 -806 1343
rect -1042 1241 -1008 1275
rect -946 1241 -912 1275
rect -840 1241 -806 1275
rect -1042 1173 -1008 1207
rect -946 1173 -912 1207
rect -840 1173 -806 1207
rect -1042 1105 -1008 1139
rect -946 1105 -912 1139
rect -840 1105 -806 1139
rect -1042 1037 -1008 1071
rect -946 1037 -912 1071
rect -840 1037 -806 1071
rect -1042 969 -1008 1003
rect -946 969 -912 1003
rect -840 969 -806 1003
rect -1042 901 -1008 935
rect -946 901 -912 935
rect -840 901 -806 935
rect -1042 833 -1008 867
rect -946 833 -912 867
rect -840 833 -806 867
rect -1042 765 -1008 799
rect -946 765 -912 799
rect -840 765 -806 799
rect -1042 697 -1008 731
rect -946 697 -912 731
rect -840 697 -806 731
rect -1042 629 -1008 663
rect -946 629 -912 663
rect -840 629 -806 663
rect -1042 561 -1008 595
rect -946 561 -912 595
rect -840 561 -806 595
rect -1042 493 -1008 527
rect -946 493 -912 527
rect -840 493 -806 527
rect -1042 425 -1008 459
rect -946 425 -912 459
rect -840 425 -806 459
rect -1042 357 -1008 391
rect -946 357 -912 391
rect -840 357 -806 391
rect -1042 289 -1008 323
rect -946 289 -912 323
rect -840 289 -806 323
rect -1042 221 -1008 255
rect -946 221 -912 255
rect -840 221 -806 255
rect -1042 153 -1008 187
rect -946 153 -912 187
rect -840 153 -806 187
rect -1042 85 -1008 119
rect -946 85 -912 119
rect -840 85 -806 119
rect -1042 17 -1008 51
rect -946 17 -912 51
rect -840 17 -806 51
rect -1042 -51 -1008 -17
rect -946 -51 -912 -17
rect -840 -51 -806 -17
rect -1042 -119 -1008 -85
rect -946 -119 -912 -85
rect -840 -119 -806 -85
rect -1042 -187 -1008 -153
rect -946 -187 -912 -153
rect -840 -187 -806 -153
rect -1042 -255 -1008 -221
rect -946 -255 -912 -221
rect -840 -255 -806 -221
rect -1042 -323 -1008 -289
rect -946 -323 -912 -289
rect -840 -323 -806 -289
rect -1042 -391 -1008 -357
rect -946 -391 -912 -357
rect -840 -391 -806 -357
rect -1042 -459 -1008 -425
rect -946 -459 -912 -425
rect -840 -459 -806 -425
rect -1042 -527 -1008 -493
rect -946 -527 -912 -493
rect -840 -527 -806 -493
rect -1042 -595 -1008 -561
rect -946 -595 -912 -561
rect -840 -595 -806 -561
rect -1042 -663 -1008 -629
rect -946 -663 -912 -629
rect -840 -663 -806 -629
rect -1042 -731 -1008 -697
rect -946 -731 -912 -697
rect -840 -731 -806 -697
rect -1042 -799 -1008 -765
rect -946 -799 -912 -765
rect -840 -799 -806 -765
rect -1042 -867 -1008 -833
rect -946 -867 -912 -833
rect -840 -867 -806 -833
rect -1042 -935 -1008 -901
rect -946 -935 -912 -901
rect -840 -935 -806 -901
rect -1042 -1003 -1008 -969
rect -946 -1003 -912 -969
rect -840 -1003 -806 -969
rect -1042 -1071 -1008 -1037
rect -946 -1071 -912 -1037
rect -840 -1071 -806 -1037
rect -1042 -1139 -1008 -1105
rect -946 -1139 -912 -1105
rect -840 -1139 -806 -1105
rect -1042 -1207 -1008 -1173
rect -946 -1207 -912 -1173
rect -840 -1207 -806 -1173
rect -1042 -1275 -1008 -1241
rect -946 -1275 -912 -1241
rect -840 -1275 -806 -1241
rect -1042 -1343 -1008 -1309
rect -946 -1343 -912 -1309
rect -840 -1343 -806 -1309
rect -1042 -1411 -1008 -1377
rect -946 -1411 -912 -1377
rect -840 -1411 -806 -1377
rect -1042 -1479 -1008 -1445
rect -946 -1479 -912 -1445
rect -840 -1479 -806 -1445
rect -1042 -1547 -1008 -1513
rect -946 -1547 -912 -1513
rect -840 -1547 -806 -1513
rect -1042 -1615 -1008 -1581
rect -946 -1615 -912 -1581
rect -840 -1615 -806 -1581
rect -1042 -1683 -1008 -1649
rect -946 -1683 -912 -1649
rect -840 -1683 -806 -1649
rect -1042 -1751 -1008 -1717
rect -946 -1751 -912 -1717
rect -840 -1751 -806 -1717
rect -1042 -1819 -1008 -1785
rect -946 -1819 -912 -1785
rect -840 -1819 -806 -1785
rect -1042 -1887 -1008 -1853
rect -946 -1887 -912 -1853
rect -840 -1887 -806 -1853
rect -1042 -1955 -1008 -1921
rect -946 -1955 -912 -1921
rect -840 -1955 -806 -1921
rect -1042 -2023 -1008 -1989
rect -946 -2023 -912 -1989
rect -840 -2023 -806 -1989
rect -1042 -2091 -1008 -2057
rect -946 -2091 -912 -2057
rect -840 -2091 -806 -2057
rect -1042 -2159 -1008 -2125
rect -946 -2159 -912 -2125
rect -840 -2159 -806 -2125
rect -1042 -2227 -1008 -2193
rect -946 -2227 -912 -2193
rect -840 -2227 -806 -2193
rect -1042 -2295 -1008 -2261
rect -946 -2295 -912 -2261
rect -840 -2295 -806 -2261
rect -1042 -2363 -1008 -2329
rect -946 -2363 -912 -2329
rect -840 -2363 -806 -2329
rect -1042 -2431 -1008 -2397
rect -946 -2431 -912 -2397
rect -840 -2431 -806 -2397
rect -1042 -2499 -1008 -2465
rect -946 -2499 -912 -2465
rect -840 -2499 -806 -2465
rect -1042 -2567 -1008 -2533
rect -946 -2567 -912 -2533
rect -840 -2567 -806 -2533
rect -1042 -2635 -1008 -2601
rect -946 -2635 -912 -2601
rect -840 -2635 -806 -2601
rect -1042 -2703 -1008 -2669
rect -946 -2703 -912 -2669
rect -840 -2703 -806 -2669
rect -1042 -2771 -1008 -2737
rect -946 -2771 -912 -2737
rect -840 -2771 -806 -2737
rect -1042 -2839 -1008 -2805
rect -946 -2839 -912 -2805
rect -840 -2839 -806 -2805
rect -1042 -2907 -1008 -2873
rect -946 -2907 -912 -2873
rect -840 -2907 -806 -2873
rect -1042 -2975 -1008 -2941
rect -946 -2975 -912 -2941
rect -840 -2975 -806 -2941
rect -1042 -3043 -1008 -3009
rect -946 -3043 -912 -3009
rect -840 -3043 -806 -3009
rect -1042 -3111 -1008 -3077
rect -946 -3111 -912 -3077
rect -840 -3111 -806 -3077
rect -1042 -3179 -1008 -3145
rect -946 -3179 -912 -3145
rect -840 -3179 -806 -3145
rect -1042 -3247 -1008 -3213
rect -946 -3247 -912 -3213
rect -840 -3247 -806 -3213
rect -1042 -3315 -1008 -3281
rect -946 -3315 -912 -3281
rect -840 -3315 -806 -3281
rect -1042 -3383 -1008 -3349
rect -946 -3383 -912 -3349
rect -840 -3383 -806 -3349
rect -1042 -3451 -1008 -3417
rect -946 -3451 -912 -3417
rect -840 -3451 -806 -3417
rect -1042 -3519 -1008 -3485
rect -946 -3519 -912 -3485
rect -840 -3519 -806 -3485
rect -1042 -3587 -1008 -3553
rect -946 -3587 -912 -3553
rect -840 -3587 -806 -3553
rect -1042 -3655 -1008 -3621
rect -946 -3655 -912 -3621
rect -840 -3655 -806 -3621
rect -1042 -3723 -1008 -3689
rect -946 -3723 -912 -3689
rect -840 -3723 -806 -3689
rect -1042 -3791 -1008 -3757
rect -946 -3791 -912 -3757
rect -840 -3791 -806 -3757
rect -1042 -3859 -1008 -3825
rect -946 -3859 -912 -3825
rect -840 -3859 -806 -3825
rect -1042 -3927 -1008 -3893
rect -946 -3927 -912 -3893
rect -840 -3927 -806 -3893
rect -1042 -3995 -1008 -3961
rect -946 -3995 -912 -3961
rect -840 -3995 -806 -3961
rect -1042 -4063 -1008 -4029
rect -946 -4063 -912 -4029
rect -840 -4063 -806 -4029
rect -1042 -4131 -1008 -4097
rect -946 -4131 -912 -4097
rect -840 -4131 -806 -4097
rect -1042 -4199 -1008 -4165
rect -946 -4199 -912 -4165
rect -840 -4199 -806 -4165
rect -1042 -4267 -1008 -4233
rect -946 -4267 -912 -4233
rect -840 -4267 -806 -4233
rect -1042 -4335 -1008 -4301
rect -946 -4335 -912 -4301
rect -840 -4335 -806 -4301
rect -1042 -4403 -1008 -4369
rect -946 -4403 -912 -4369
rect -840 -4403 -806 -4369
rect -1042 -4471 -1008 -4437
rect -946 -4471 -912 -4437
rect -840 -4471 -806 -4437
rect -1042 -4539 -1008 -4505
rect -946 -4539 -912 -4505
rect -840 -4539 -806 -4505
rect -1042 -4607 -1008 -4573
rect -946 -4607 -912 -4573
rect -840 -4607 -806 -4573
rect -1042 -4675 -1008 -4641
rect -946 -4675 -912 -4641
rect -840 -4675 -806 -4641
rect -1042 -4743 -1008 -4709
rect -946 -4743 -912 -4709
rect -840 -4743 -806 -4709
rect -1042 -4811 -1008 -4777
rect -946 -4811 -912 -4777
rect -840 -4811 -806 -4777
rect -1042 -4879 -1008 -4845
rect -946 -4879 -912 -4845
rect -840 -4879 -806 -4845
rect -1042 -4947 -1008 -4913
rect -946 -4947 -912 -4913
rect -840 -4947 -806 -4913
rect -1042 -5015 -1008 -4981
rect -946 -5015 -912 -4981
rect -840 -5015 -806 -4981
rect -426 4981 -392 5015
rect -330 4981 -296 5015
rect -224 4981 -190 5015
rect -426 4913 -392 4947
rect -330 4913 -296 4947
rect -224 4913 -190 4947
rect -426 4845 -392 4879
rect -330 4845 -296 4879
rect -224 4845 -190 4879
rect -426 4777 -392 4811
rect -330 4777 -296 4811
rect -224 4777 -190 4811
rect -426 4709 -392 4743
rect -330 4709 -296 4743
rect -224 4709 -190 4743
rect -426 4641 -392 4675
rect -330 4641 -296 4675
rect -224 4641 -190 4675
rect -426 4573 -392 4607
rect -330 4573 -296 4607
rect -224 4573 -190 4607
rect -426 4505 -392 4539
rect -330 4505 -296 4539
rect -224 4505 -190 4539
rect -426 4437 -392 4471
rect -330 4437 -296 4471
rect -224 4437 -190 4471
rect -426 4369 -392 4403
rect -330 4369 -296 4403
rect -224 4369 -190 4403
rect -426 4301 -392 4335
rect -330 4301 -296 4335
rect -224 4301 -190 4335
rect -426 4233 -392 4267
rect -330 4233 -296 4267
rect -224 4233 -190 4267
rect -426 4165 -392 4199
rect -330 4165 -296 4199
rect -224 4165 -190 4199
rect -426 4097 -392 4131
rect -330 4097 -296 4131
rect -224 4097 -190 4131
rect -426 4029 -392 4063
rect -330 4029 -296 4063
rect -224 4029 -190 4063
rect -426 3961 -392 3995
rect -330 3961 -296 3995
rect -224 3961 -190 3995
rect -426 3893 -392 3927
rect -330 3893 -296 3927
rect -224 3893 -190 3927
rect -426 3825 -392 3859
rect -330 3825 -296 3859
rect -224 3825 -190 3859
rect -426 3757 -392 3791
rect -330 3757 -296 3791
rect -224 3757 -190 3791
rect -426 3689 -392 3723
rect -330 3689 -296 3723
rect -224 3689 -190 3723
rect -426 3621 -392 3655
rect -330 3621 -296 3655
rect -224 3621 -190 3655
rect -426 3553 -392 3587
rect -330 3553 -296 3587
rect -224 3553 -190 3587
rect -426 3485 -392 3519
rect -330 3485 -296 3519
rect -224 3485 -190 3519
rect -426 3417 -392 3451
rect -330 3417 -296 3451
rect -224 3417 -190 3451
rect -426 3349 -392 3383
rect -330 3349 -296 3383
rect -224 3349 -190 3383
rect -426 3281 -392 3315
rect -330 3281 -296 3315
rect -224 3281 -190 3315
rect -426 3213 -392 3247
rect -330 3213 -296 3247
rect -224 3213 -190 3247
rect -426 3145 -392 3179
rect -330 3145 -296 3179
rect -224 3145 -190 3179
rect -426 3077 -392 3111
rect -330 3077 -296 3111
rect -224 3077 -190 3111
rect -426 3009 -392 3043
rect -330 3009 -296 3043
rect -224 3009 -190 3043
rect -426 2941 -392 2975
rect -330 2941 -296 2975
rect -224 2941 -190 2975
rect -426 2873 -392 2907
rect -330 2873 -296 2907
rect -224 2873 -190 2907
rect -426 2805 -392 2839
rect -330 2805 -296 2839
rect -224 2805 -190 2839
rect -426 2737 -392 2771
rect -330 2737 -296 2771
rect -224 2737 -190 2771
rect -426 2669 -392 2703
rect -330 2669 -296 2703
rect -224 2669 -190 2703
rect -426 2601 -392 2635
rect -330 2601 -296 2635
rect -224 2601 -190 2635
rect -426 2533 -392 2567
rect -330 2533 -296 2567
rect -224 2533 -190 2567
rect -426 2465 -392 2499
rect -330 2465 -296 2499
rect -224 2465 -190 2499
rect -426 2397 -392 2431
rect -330 2397 -296 2431
rect -224 2397 -190 2431
rect -426 2329 -392 2363
rect -330 2329 -296 2363
rect -224 2329 -190 2363
rect -426 2261 -392 2295
rect -330 2261 -296 2295
rect -224 2261 -190 2295
rect -426 2193 -392 2227
rect -330 2193 -296 2227
rect -224 2193 -190 2227
rect -426 2125 -392 2159
rect -330 2125 -296 2159
rect -224 2125 -190 2159
rect -426 2057 -392 2091
rect -330 2057 -296 2091
rect -224 2057 -190 2091
rect -426 1989 -392 2023
rect -330 1989 -296 2023
rect -224 1989 -190 2023
rect -426 1921 -392 1955
rect -330 1921 -296 1955
rect -224 1921 -190 1955
rect -426 1853 -392 1887
rect -330 1853 -296 1887
rect -224 1853 -190 1887
rect -426 1785 -392 1819
rect -330 1785 -296 1819
rect -224 1785 -190 1819
rect -426 1717 -392 1751
rect -330 1717 -296 1751
rect -224 1717 -190 1751
rect -426 1649 -392 1683
rect -330 1649 -296 1683
rect -224 1649 -190 1683
rect -426 1581 -392 1615
rect -330 1581 -296 1615
rect -224 1581 -190 1615
rect -426 1513 -392 1547
rect -330 1513 -296 1547
rect -224 1513 -190 1547
rect -426 1445 -392 1479
rect -330 1445 -296 1479
rect -224 1445 -190 1479
rect -426 1377 -392 1411
rect -330 1377 -296 1411
rect -224 1377 -190 1411
rect -426 1309 -392 1343
rect -330 1309 -296 1343
rect -224 1309 -190 1343
rect -426 1241 -392 1275
rect -330 1241 -296 1275
rect -224 1241 -190 1275
rect -426 1173 -392 1207
rect -330 1173 -296 1207
rect -224 1173 -190 1207
rect -426 1105 -392 1139
rect -330 1105 -296 1139
rect -224 1105 -190 1139
rect -426 1037 -392 1071
rect -330 1037 -296 1071
rect -224 1037 -190 1071
rect -426 969 -392 1003
rect -330 969 -296 1003
rect -224 969 -190 1003
rect -426 901 -392 935
rect -330 901 -296 935
rect -224 901 -190 935
rect -426 833 -392 867
rect -330 833 -296 867
rect -224 833 -190 867
rect -426 765 -392 799
rect -330 765 -296 799
rect -224 765 -190 799
rect -426 697 -392 731
rect -330 697 -296 731
rect -224 697 -190 731
rect -426 629 -392 663
rect -330 629 -296 663
rect -224 629 -190 663
rect -426 561 -392 595
rect -330 561 -296 595
rect -224 561 -190 595
rect -426 493 -392 527
rect -330 493 -296 527
rect -224 493 -190 527
rect -426 425 -392 459
rect -330 425 -296 459
rect -224 425 -190 459
rect -426 357 -392 391
rect -330 357 -296 391
rect -224 357 -190 391
rect -426 289 -392 323
rect -330 289 -296 323
rect -224 289 -190 323
rect -426 221 -392 255
rect -330 221 -296 255
rect -224 221 -190 255
rect -426 153 -392 187
rect -330 153 -296 187
rect -224 153 -190 187
rect -426 85 -392 119
rect -330 85 -296 119
rect -224 85 -190 119
rect -426 17 -392 51
rect -330 17 -296 51
rect -224 17 -190 51
rect -426 -51 -392 -17
rect -330 -51 -296 -17
rect -224 -51 -190 -17
rect -426 -119 -392 -85
rect -330 -119 -296 -85
rect -224 -119 -190 -85
rect -426 -187 -392 -153
rect -330 -187 -296 -153
rect -224 -187 -190 -153
rect -426 -255 -392 -221
rect -330 -255 -296 -221
rect -224 -255 -190 -221
rect -426 -323 -392 -289
rect -330 -323 -296 -289
rect -224 -323 -190 -289
rect -426 -391 -392 -357
rect -330 -391 -296 -357
rect -224 -391 -190 -357
rect -426 -459 -392 -425
rect -330 -459 -296 -425
rect -224 -459 -190 -425
rect -426 -527 -392 -493
rect -330 -527 -296 -493
rect -224 -527 -190 -493
rect -426 -595 -392 -561
rect -330 -595 -296 -561
rect -224 -595 -190 -561
rect -426 -663 -392 -629
rect -330 -663 -296 -629
rect -224 -663 -190 -629
rect -426 -731 -392 -697
rect -330 -731 -296 -697
rect -224 -731 -190 -697
rect -426 -799 -392 -765
rect -330 -799 -296 -765
rect -224 -799 -190 -765
rect -426 -867 -392 -833
rect -330 -867 -296 -833
rect -224 -867 -190 -833
rect -426 -935 -392 -901
rect -330 -935 -296 -901
rect -224 -935 -190 -901
rect -426 -1003 -392 -969
rect -330 -1003 -296 -969
rect -224 -1003 -190 -969
rect -426 -1071 -392 -1037
rect -330 -1071 -296 -1037
rect -224 -1071 -190 -1037
rect -426 -1139 -392 -1105
rect -330 -1139 -296 -1105
rect -224 -1139 -190 -1105
rect -426 -1207 -392 -1173
rect -330 -1207 -296 -1173
rect -224 -1207 -190 -1173
rect -426 -1275 -392 -1241
rect -330 -1275 -296 -1241
rect -224 -1275 -190 -1241
rect -426 -1343 -392 -1309
rect -330 -1343 -296 -1309
rect -224 -1343 -190 -1309
rect -426 -1411 -392 -1377
rect -330 -1411 -296 -1377
rect -224 -1411 -190 -1377
rect -426 -1479 -392 -1445
rect -330 -1479 -296 -1445
rect -224 -1479 -190 -1445
rect -426 -1547 -392 -1513
rect -330 -1547 -296 -1513
rect -224 -1547 -190 -1513
rect -426 -1615 -392 -1581
rect -330 -1615 -296 -1581
rect -224 -1615 -190 -1581
rect -426 -1683 -392 -1649
rect -330 -1683 -296 -1649
rect -224 -1683 -190 -1649
rect -426 -1751 -392 -1717
rect -330 -1751 -296 -1717
rect -224 -1751 -190 -1717
rect -426 -1819 -392 -1785
rect -330 -1819 -296 -1785
rect -224 -1819 -190 -1785
rect -426 -1887 -392 -1853
rect -330 -1887 -296 -1853
rect -224 -1887 -190 -1853
rect -426 -1955 -392 -1921
rect -330 -1955 -296 -1921
rect -224 -1955 -190 -1921
rect -426 -2023 -392 -1989
rect -330 -2023 -296 -1989
rect -224 -2023 -190 -1989
rect -426 -2091 -392 -2057
rect -330 -2091 -296 -2057
rect -224 -2091 -190 -2057
rect -426 -2159 -392 -2125
rect -330 -2159 -296 -2125
rect -224 -2159 -190 -2125
rect -426 -2227 -392 -2193
rect -330 -2227 -296 -2193
rect -224 -2227 -190 -2193
rect -426 -2295 -392 -2261
rect -330 -2295 -296 -2261
rect -224 -2295 -190 -2261
rect -426 -2363 -392 -2329
rect -330 -2363 -296 -2329
rect -224 -2363 -190 -2329
rect -426 -2431 -392 -2397
rect -330 -2431 -296 -2397
rect -224 -2431 -190 -2397
rect -426 -2499 -392 -2465
rect -330 -2499 -296 -2465
rect -224 -2499 -190 -2465
rect -426 -2567 -392 -2533
rect -330 -2567 -296 -2533
rect -224 -2567 -190 -2533
rect -426 -2635 -392 -2601
rect -330 -2635 -296 -2601
rect -224 -2635 -190 -2601
rect -426 -2703 -392 -2669
rect -330 -2703 -296 -2669
rect -224 -2703 -190 -2669
rect -426 -2771 -392 -2737
rect -330 -2771 -296 -2737
rect -224 -2771 -190 -2737
rect -426 -2839 -392 -2805
rect -330 -2839 -296 -2805
rect -224 -2839 -190 -2805
rect -426 -2907 -392 -2873
rect -330 -2907 -296 -2873
rect -224 -2907 -190 -2873
rect -426 -2975 -392 -2941
rect -330 -2975 -296 -2941
rect -224 -2975 -190 -2941
rect -426 -3043 -392 -3009
rect -330 -3043 -296 -3009
rect -224 -3043 -190 -3009
rect -426 -3111 -392 -3077
rect -330 -3111 -296 -3077
rect -224 -3111 -190 -3077
rect -426 -3179 -392 -3145
rect -330 -3179 -296 -3145
rect -224 -3179 -190 -3145
rect -426 -3247 -392 -3213
rect -330 -3247 -296 -3213
rect -224 -3247 -190 -3213
rect -426 -3315 -392 -3281
rect -330 -3315 -296 -3281
rect -224 -3315 -190 -3281
rect -426 -3383 -392 -3349
rect -330 -3383 -296 -3349
rect -224 -3383 -190 -3349
rect -426 -3451 -392 -3417
rect -330 -3451 -296 -3417
rect -224 -3451 -190 -3417
rect -426 -3519 -392 -3485
rect -330 -3519 -296 -3485
rect -224 -3519 -190 -3485
rect -426 -3587 -392 -3553
rect -330 -3587 -296 -3553
rect -224 -3587 -190 -3553
rect -426 -3655 -392 -3621
rect -330 -3655 -296 -3621
rect -224 -3655 -190 -3621
rect -426 -3723 -392 -3689
rect -330 -3723 -296 -3689
rect -224 -3723 -190 -3689
rect -426 -3791 -392 -3757
rect -330 -3791 -296 -3757
rect -224 -3791 -190 -3757
rect -426 -3859 -392 -3825
rect -330 -3859 -296 -3825
rect -224 -3859 -190 -3825
rect -426 -3927 -392 -3893
rect -330 -3927 -296 -3893
rect -224 -3927 -190 -3893
rect -426 -3995 -392 -3961
rect -330 -3995 -296 -3961
rect -224 -3995 -190 -3961
rect -426 -4063 -392 -4029
rect -330 -4063 -296 -4029
rect -224 -4063 -190 -4029
rect -426 -4131 -392 -4097
rect -330 -4131 -296 -4097
rect -224 -4131 -190 -4097
rect -426 -4199 -392 -4165
rect -330 -4199 -296 -4165
rect -224 -4199 -190 -4165
rect -426 -4267 -392 -4233
rect -330 -4267 -296 -4233
rect -224 -4267 -190 -4233
rect -426 -4335 -392 -4301
rect -330 -4335 -296 -4301
rect -224 -4335 -190 -4301
rect -426 -4403 -392 -4369
rect -330 -4403 -296 -4369
rect -224 -4403 -190 -4369
rect -426 -4471 -392 -4437
rect -330 -4471 -296 -4437
rect -224 -4471 -190 -4437
rect -426 -4539 -392 -4505
rect -330 -4539 -296 -4505
rect -224 -4539 -190 -4505
rect -426 -4607 -392 -4573
rect -330 -4607 -296 -4573
rect -224 -4607 -190 -4573
rect -426 -4675 -392 -4641
rect -330 -4675 -296 -4641
rect -224 -4675 -190 -4641
rect -426 -4743 -392 -4709
rect -330 -4743 -296 -4709
rect -224 -4743 -190 -4709
rect -426 -4811 -392 -4777
rect -330 -4811 -296 -4777
rect -224 -4811 -190 -4777
rect -426 -4879 -392 -4845
rect -330 -4879 -296 -4845
rect -224 -4879 -190 -4845
rect -426 -4947 -392 -4913
rect -330 -4947 -296 -4913
rect -224 -4947 -190 -4913
rect -426 -5015 -392 -4981
rect -330 -5015 -296 -4981
rect -224 -5015 -190 -4981
rect 190 4981 224 5015
rect 286 4981 320 5015
rect 392 4981 426 5015
rect 190 4913 224 4947
rect 286 4913 320 4947
rect 392 4913 426 4947
rect 190 4845 224 4879
rect 286 4845 320 4879
rect 392 4845 426 4879
rect 190 4777 224 4811
rect 286 4777 320 4811
rect 392 4777 426 4811
rect 190 4709 224 4743
rect 286 4709 320 4743
rect 392 4709 426 4743
rect 190 4641 224 4675
rect 286 4641 320 4675
rect 392 4641 426 4675
rect 190 4573 224 4607
rect 286 4573 320 4607
rect 392 4573 426 4607
rect 190 4505 224 4539
rect 286 4505 320 4539
rect 392 4505 426 4539
rect 190 4437 224 4471
rect 286 4437 320 4471
rect 392 4437 426 4471
rect 190 4369 224 4403
rect 286 4369 320 4403
rect 392 4369 426 4403
rect 190 4301 224 4335
rect 286 4301 320 4335
rect 392 4301 426 4335
rect 190 4233 224 4267
rect 286 4233 320 4267
rect 392 4233 426 4267
rect 190 4165 224 4199
rect 286 4165 320 4199
rect 392 4165 426 4199
rect 190 4097 224 4131
rect 286 4097 320 4131
rect 392 4097 426 4131
rect 190 4029 224 4063
rect 286 4029 320 4063
rect 392 4029 426 4063
rect 190 3961 224 3995
rect 286 3961 320 3995
rect 392 3961 426 3995
rect 190 3893 224 3927
rect 286 3893 320 3927
rect 392 3893 426 3927
rect 190 3825 224 3859
rect 286 3825 320 3859
rect 392 3825 426 3859
rect 190 3757 224 3791
rect 286 3757 320 3791
rect 392 3757 426 3791
rect 190 3689 224 3723
rect 286 3689 320 3723
rect 392 3689 426 3723
rect 190 3621 224 3655
rect 286 3621 320 3655
rect 392 3621 426 3655
rect 190 3553 224 3587
rect 286 3553 320 3587
rect 392 3553 426 3587
rect 190 3485 224 3519
rect 286 3485 320 3519
rect 392 3485 426 3519
rect 190 3417 224 3451
rect 286 3417 320 3451
rect 392 3417 426 3451
rect 190 3349 224 3383
rect 286 3349 320 3383
rect 392 3349 426 3383
rect 190 3281 224 3315
rect 286 3281 320 3315
rect 392 3281 426 3315
rect 190 3213 224 3247
rect 286 3213 320 3247
rect 392 3213 426 3247
rect 190 3145 224 3179
rect 286 3145 320 3179
rect 392 3145 426 3179
rect 190 3077 224 3111
rect 286 3077 320 3111
rect 392 3077 426 3111
rect 190 3009 224 3043
rect 286 3009 320 3043
rect 392 3009 426 3043
rect 190 2941 224 2975
rect 286 2941 320 2975
rect 392 2941 426 2975
rect 190 2873 224 2907
rect 286 2873 320 2907
rect 392 2873 426 2907
rect 190 2805 224 2839
rect 286 2805 320 2839
rect 392 2805 426 2839
rect 190 2737 224 2771
rect 286 2737 320 2771
rect 392 2737 426 2771
rect 190 2669 224 2703
rect 286 2669 320 2703
rect 392 2669 426 2703
rect 190 2601 224 2635
rect 286 2601 320 2635
rect 392 2601 426 2635
rect 190 2533 224 2567
rect 286 2533 320 2567
rect 392 2533 426 2567
rect 190 2465 224 2499
rect 286 2465 320 2499
rect 392 2465 426 2499
rect 190 2397 224 2431
rect 286 2397 320 2431
rect 392 2397 426 2431
rect 190 2329 224 2363
rect 286 2329 320 2363
rect 392 2329 426 2363
rect 190 2261 224 2295
rect 286 2261 320 2295
rect 392 2261 426 2295
rect 190 2193 224 2227
rect 286 2193 320 2227
rect 392 2193 426 2227
rect 190 2125 224 2159
rect 286 2125 320 2159
rect 392 2125 426 2159
rect 190 2057 224 2091
rect 286 2057 320 2091
rect 392 2057 426 2091
rect 190 1989 224 2023
rect 286 1989 320 2023
rect 392 1989 426 2023
rect 190 1921 224 1955
rect 286 1921 320 1955
rect 392 1921 426 1955
rect 190 1853 224 1887
rect 286 1853 320 1887
rect 392 1853 426 1887
rect 190 1785 224 1819
rect 286 1785 320 1819
rect 392 1785 426 1819
rect 190 1717 224 1751
rect 286 1717 320 1751
rect 392 1717 426 1751
rect 190 1649 224 1683
rect 286 1649 320 1683
rect 392 1649 426 1683
rect 190 1581 224 1615
rect 286 1581 320 1615
rect 392 1581 426 1615
rect 190 1513 224 1547
rect 286 1513 320 1547
rect 392 1513 426 1547
rect 190 1445 224 1479
rect 286 1445 320 1479
rect 392 1445 426 1479
rect 190 1377 224 1411
rect 286 1377 320 1411
rect 392 1377 426 1411
rect 190 1309 224 1343
rect 286 1309 320 1343
rect 392 1309 426 1343
rect 190 1241 224 1275
rect 286 1241 320 1275
rect 392 1241 426 1275
rect 190 1173 224 1207
rect 286 1173 320 1207
rect 392 1173 426 1207
rect 190 1105 224 1139
rect 286 1105 320 1139
rect 392 1105 426 1139
rect 190 1037 224 1071
rect 286 1037 320 1071
rect 392 1037 426 1071
rect 190 969 224 1003
rect 286 969 320 1003
rect 392 969 426 1003
rect 190 901 224 935
rect 286 901 320 935
rect 392 901 426 935
rect 190 833 224 867
rect 286 833 320 867
rect 392 833 426 867
rect 190 765 224 799
rect 286 765 320 799
rect 392 765 426 799
rect 190 697 224 731
rect 286 697 320 731
rect 392 697 426 731
rect 190 629 224 663
rect 286 629 320 663
rect 392 629 426 663
rect 190 561 224 595
rect 286 561 320 595
rect 392 561 426 595
rect 190 493 224 527
rect 286 493 320 527
rect 392 493 426 527
rect 190 425 224 459
rect 286 425 320 459
rect 392 425 426 459
rect 190 357 224 391
rect 286 357 320 391
rect 392 357 426 391
rect 190 289 224 323
rect 286 289 320 323
rect 392 289 426 323
rect 190 221 224 255
rect 286 221 320 255
rect 392 221 426 255
rect 190 153 224 187
rect 286 153 320 187
rect 392 153 426 187
rect 190 85 224 119
rect 286 85 320 119
rect 392 85 426 119
rect 190 17 224 51
rect 286 17 320 51
rect 392 17 426 51
rect 190 -51 224 -17
rect 286 -51 320 -17
rect 392 -51 426 -17
rect 190 -119 224 -85
rect 286 -119 320 -85
rect 392 -119 426 -85
rect 190 -187 224 -153
rect 286 -187 320 -153
rect 392 -187 426 -153
rect 190 -255 224 -221
rect 286 -255 320 -221
rect 392 -255 426 -221
rect 190 -323 224 -289
rect 286 -323 320 -289
rect 392 -323 426 -289
rect 190 -391 224 -357
rect 286 -391 320 -357
rect 392 -391 426 -357
rect 190 -459 224 -425
rect 286 -459 320 -425
rect 392 -459 426 -425
rect 190 -527 224 -493
rect 286 -527 320 -493
rect 392 -527 426 -493
rect 190 -595 224 -561
rect 286 -595 320 -561
rect 392 -595 426 -561
rect 190 -663 224 -629
rect 286 -663 320 -629
rect 392 -663 426 -629
rect 190 -731 224 -697
rect 286 -731 320 -697
rect 392 -731 426 -697
rect 190 -799 224 -765
rect 286 -799 320 -765
rect 392 -799 426 -765
rect 190 -867 224 -833
rect 286 -867 320 -833
rect 392 -867 426 -833
rect 190 -935 224 -901
rect 286 -935 320 -901
rect 392 -935 426 -901
rect 190 -1003 224 -969
rect 286 -1003 320 -969
rect 392 -1003 426 -969
rect 190 -1071 224 -1037
rect 286 -1071 320 -1037
rect 392 -1071 426 -1037
rect 190 -1139 224 -1105
rect 286 -1139 320 -1105
rect 392 -1139 426 -1105
rect 190 -1207 224 -1173
rect 286 -1207 320 -1173
rect 392 -1207 426 -1173
rect 190 -1275 224 -1241
rect 286 -1275 320 -1241
rect 392 -1275 426 -1241
rect 190 -1343 224 -1309
rect 286 -1343 320 -1309
rect 392 -1343 426 -1309
rect 190 -1411 224 -1377
rect 286 -1411 320 -1377
rect 392 -1411 426 -1377
rect 190 -1479 224 -1445
rect 286 -1479 320 -1445
rect 392 -1479 426 -1445
rect 190 -1547 224 -1513
rect 286 -1547 320 -1513
rect 392 -1547 426 -1513
rect 190 -1615 224 -1581
rect 286 -1615 320 -1581
rect 392 -1615 426 -1581
rect 190 -1683 224 -1649
rect 286 -1683 320 -1649
rect 392 -1683 426 -1649
rect 190 -1751 224 -1717
rect 286 -1751 320 -1717
rect 392 -1751 426 -1717
rect 190 -1819 224 -1785
rect 286 -1819 320 -1785
rect 392 -1819 426 -1785
rect 190 -1887 224 -1853
rect 286 -1887 320 -1853
rect 392 -1887 426 -1853
rect 190 -1955 224 -1921
rect 286 -1955 320 -1921
rect 392 -1955 426 -1921
rect 190 -2023 224 -1989
rect 286 -2023 320 -1989
rect 392 -2023 426 -1989
rect 190 -2091 224 -2057
rect 286 -2091 320 -2057
rect 392 -2091 426 -2057
rect 190 -2159 224 -2125
rect 286 -2159 320 -2125
rect 392 -2159 426 -2125
rect 190 -2227 224 -2193
rect 286 -2227 320 -2193
rect 392 -2227 426 -2193
rect 190 -2295 224 -2261
rect 286 -2295 320 -2261
rect 392 -2295 426 -2261
rect 190 -2363 224 -2329
rect 286 -2363 320 -2329
rect 392 -2363 426 -2329
rect 190 -2431 224 -2397
rect 286 -2431 320 -2397
rect 392 -2431 426 -2397
rect 190 -2499 224 -2465
rect 286 -2499 320 -2465
rect 392 -2499 426 -2465
rect 190 -2567 224 -2533
rect 286 -2567 320 -2533
rect 392 -2567 426 -2533
rect 190 -2635 224 -2601
rect 286 -2635 320 -2601
rect 392 -2635 426 -2601
rect 190 -2703 224 -2669
rect 286 -2703 320 -2669
rect 392 -2703 426 -2669
rect 190 -2771 224 -2737
rect 286 -2771 320 -2737
rect 392 -2771 426 -2737
rect 190 -2839 224 -2805
rect 286 -2839 320 -2805
rect 392 -2839 426 -2805
rect 190 -2907 224 -2873
rect 286 -2907 320 -2873
rect 392 -2907 426 -2873
rect 190 -2975 224 -2941
rect 286 -2975 320 -2941
rect 392 -2975 426 -2941
rect 190 -3043 224 -3009
rect 286 -3043 320 -3009
rect 392 -3043 426 -3009
rect 190 -3111 224 -3077
rect 286 -3111 320 -3077
rect 392 -3111 426 -3077
rect 190 -3179 224 -3145
rect 286 -3179 320 -3145
rect 392 -3179 426 -3145
rect 190 -3247 224 -3213
rect 286 -3247 320 -3213
rect 392 -3247 426 -3213
rect 190 -3315 224 -3281
rect 286 -3315 320 -3281
rect 392 -3315 426 -3281
rect 190 -3383 224 -3349
rect 286 -3383 320 -3349
rect 392 -3383 426 -3349
rect 190 -3451 224 -3417
rect 286 -3451 320 -3417
rect 392 -3451 426 -3417
rect 190 -3519 224 -3485
rect 286 -3519 320 -3485
rect 392 -3519 426 -3485
rect 190 -3587 224 -3553
rect 286 -3587 320 -3553
rect 392 -3587 426 -3553
rect 190 -3655 224 -3621
rect 286 -3655 320 -3621
rect 392 -3655 426 -3621
rect 190 -3723 224 -3689
rect 286 -3723 320 -3689
rect 392 -3723 426 -3689
rect 190 -3791 224 -3757
rect 286 -3791 320 -3757
rect 392 -3791 426 -3757
rect 190 -3859 224 -3825
rect 286 -3859 320 -3825
rect 392 -3859 426 -3825
rect 190 -3927 224 -3893
rect 286 -3927 320 -3893
rect 392 -3927 426 -3893
rect 190 -3995 224 -3961
rect 286 -3995 320 -3961
rect 392 -3995 426 -3961
rect 190 -4063 224 -4029
rect 286 -4063 320 -4029
rect 392 -4063 426 -4029
rect 190 -4131 224 -4097
rect 286 -4131 320 -4097
rect 392 -4131 426 -4097
rect 190 -4199 224 -4165
rect 286 -4199 320 -4165
rect 392 -4199 426 -4165
rect 190 -4267 224 -4233
rect 286 -4267 320 -4233
rect 392 -4267 426 -4233
rect 190 -4335 224 -4301
rect 286 -4335 320 -4301
rect 392 -4335 426 -4301
rect 190 -4403 224 -4369
rect 286 -4403 320 -4369
rect 392 -4403 426 -4369
rect 190 -4471 224 -4437
rect 286 -4471 320 -4437
rect 392 -4471 426 -4437
rect 190 -4539 224 -4505
rect 286 -4539 320 -4505
rect 392 -4539 426 -4505
rect 190 -4607 224 -4573
rect 286 -4607 320 -4573
rect 392 -4607 426 -4573
rect 190 -4675 224 -4641
rect 286 -4675 320 -4641
rect 392 -4675 426 -4641
rect 190 -4743 224 -4709
rect 286 -4743 320 -4709
rect 392 -4743 426 -4709
rect 190 -4811 224 -4777
rect 286 -4811 320 -4777
rect 392 -4811 426 -4777
rect 190 -4879 224 -4845
rect 286 -4879 320 -4845
rect 392 -4879 426 -4845
rect 190 -4947 224 -4913
rect 286 -4947 320 -4913
rect 392 -4947 426 -4913
rect 190 -5015 224 -4981
rect 286 -5015 320 -4981
rect 392 -5015 426 -4981
rect 806 4981 840 5015
rect 902 4981 936 5015
rect 1008 4981 1042 5015
rect 806 4913 840 4947
rect 902 4913 936 4947
rect 1008 4913 1042 4947
rect 806 4845 840 4879
rect 902 4845 936 4879
rect 1008 4845 1042 4879
rect 806 4777 840 4811
rect 902 4777 936 4811
rect 1008 4777 1042 4811
rect 806 4709 840 4743
rect 902 4709 936 4743
rect 1008 4709 1042 4743
rect 806 4641 840 4675
rect 902 4641 936 4675
rect 1008 4641 1042 4675
rect 806 4573 840 4607
rect 902 4573 936 4607
rect 1008 4573 1042 4607
rect 806 4505 840 4539
rect 902 4505 936 4539
rect 1008 4505 1042 4539
rect 806 4437 840 4471
rect 902 4437 936 4471
rect 1008 4437 1042 4471
rect 806 4369 840 4403
rect 902 4369 936 4403
rect 1008 4369 1042 4403
rect 806 4301 840 4335
rect 902 4301 936 4335
rect 1008 4301 1042 4335
rect 806 4233 840 4267
rect 902 4233 936 4267
rect 1008 4233 1042 4267
rect 806 4165 840 4199
rect 902 4165 936 4199
rect 1008 4165 1042 4199
rect 806 4097 840 4131
rect 902 4097 936 4131
rect 1008 4097 1042 4131
rect 806 4029 840 4063
rect 902 4029 936 4063
rect 1008 4029 1042 4063
rect 806 3961 840 3995
rect 902 3961 936 3995
rect 1008 3961 1042 3995
rect 806 3893 840 3927
rect 902 3893 936 3927
rect 1008 3893 1042 3927
rect 806 3825 840 3859
rect 902 3825 936 3859
rect 1008 3825 1042 3859
rect 806 3757 840 3791
rect 902 3757 936 3791
rect 1008 3757 1042 3791
rect 806 3689 840 3723
rect 902 3689 936 3723
rect 1008 3689 1042 3723
rect 806 3621 840 3655
rect 902 3621 936 3655
rect 1008 3621 1042 3655
rect 806 3553 840 3587
rect 902 3553 936 3587
rect 1008 3553 1042 3587
rect 806 3485 840 3519
rect 902 3485 936 3519
rect 1008 3485 1042 3519
rect 806 3417 840 3451
rect 902 3417 936 3451
rect 1008 3417 1042 3451
rect 806 3349 840 3383
rect 902 3349 936 3383
rect 1008 3349 1042 3383
rect 806 3281 840 3315
rect 902 3281 936 3315
rect 1008 3281 1042 3315
rect 806 3213 840 3247
rect 902 3213 936 3247
rect 1008 3213 1042 3247
rect 806 3145 840 3179
rect 902 3145 936 3179
rect 1008 3145 1042 3179
rect 806 3077 840 3111
rect 902 3077 936 3111
rect 1008 3077 1042 3111
rect 806 3009 840 3043
rect 902 3009 936 3043
rect 1008 3009 1042 3043
rect 806 2941 840 2975
rect 902 2941 936 2975
rect 1008 2941 1042 2975
rect 806 2873 840 2907
rect 902 2873 936 2907
rect 1008 2873 1042 2907
rect 806 2805 840 2839
rect 902 2805 936 2839
rect 1008 2805 1042 2839
rect 806 2737 840 2771
rect 902 2737 936 2771
rect 1008 2737 1042 2771
rect 806 2669 840 2703
rect 902 2669 936 2703
rect 1008 2669 1042 2703
rect 806 2601 840 2635
rect 902 2601 936 2635
rect 1008 2601 1042 2635
rect 806 2533 840 2567
rect 902 2533 936 2567
rect 1008 2533 1042 2567
rect 806 2465 840 2499
rect 902 2465 936 2499
rect 1008 2465 1042 2499
rect 806 2397 840 2431
rect 902 2397 936 2431
rect 1008 2397 1042 2431
rect 806 2329 840 2363
rect 902 2329 936 2363
rect 1008 2329 1042 2363
rect 806 2261 840 2295
rect 902 2261 936 2295
rect 1008 2261 1042 2295
rect 806 2193 840 2227
rect 902 2193 936 2227
rect 1008 2193 1042 2227
rect 806 2125 840 2159
rect 902 2125 936 2159
rect 1008 2125 1042 2159
rect 806 2057 840 2091
rect 902 2057 936 2091
rect 1008 2057 1042 2091
rect 806 1989 840 2023
rect 902 1989 936 2023
rect 1008 1989 1042 2023
rect 806 1921 840 1955
rect 902 1921 936 1955
rect 1008 1921 1042 1955
rect 806 1853 840 1887
rect 902 1853 936 1887
rect 1008 1853 1042 1887
rect 806 1785 840 1819
rect 902 1785 936 1819
rect 1008 1785 1042 1819
rect 806 1717 840 1751
rect 902 1717 936 1751
rect 1008 1717 1042 1751
rect 806 1649 840 1683
rect 902 1649 936 1683
rect 1008 1649 1042 1683
rect 806 1581 840 1615
rect 902 1581 936 1615
rect 1008 1581 1042 1615
rect 806 1513 840 1547
rect 902 1513 936 1547
rect 1008 1513 1042 1547
rect 806 1445 840 1479
rect 902 1445 936 1479
rect 1008 1445 1042 1479
rect 806 1377 840 1411
rect 902 1377 936 1411
rect 1008 1377 1042 1411
rect 806 1309 840 1343
rect 902 1309 936 1343
rect 1008 1309 1042 1343
rect 806 1241 840 1275
rect 902 1241 936 1275
rect 1008 1241 1042 1275
rect 806 1173 840 1207
rect 902 1173 936 1207
rect 1008 1173 1042 1207
rect 806 1105 840 1139
rect 902 1105 936 1139
rect 1008 1105 1042 1139
rect 806 1037 840 1071
rect 902 1037 936 1071
rect 1008 1037 1042 1071
rect 806 969 840 1003
rect 902 969 936 1003
rect 1008 969 1042 1003
rect 806 901 840 935
rect 902 901 936 935
rect 1008 901 1042 935
rect 806 833 840 867
rect 902 833 936 867
rect 1008 833 1042 867
rect 806 765 840 799
rect 902 765 936 799
rect 1008 765 1042 799
rect 806 697 840 731
rect 902 697 936 731
rect 1008 697 1042 731
rect 806 629 840 663
rect 902 629 936 663
rect 1008 629 1042 663
rect 806 561 840 595
rect 902 561 936 595
rect 1008 561 1042 595
rect 806 493 840 527
rect 902 493 936 527
rect 1008 493 1042 527
rect 806 425 840 459
rect 902 425 936 459
rect 1008 425 1042 459
rect 806 357 840 391
rect 902 357 936 391
rect 1008 357 1042 391
rect 806 289 840 323
rect 902 289 936 323
rect 1008 289 1042 323
rect 806 221 840 255
rect 902 221 936 255
rect 1008 221 1042 255
rect 806 153 840 187
rect 902 153 936 187
rect 1008 153 1042 187
rect 806 85 840 119
rect 902 85 936 119
rect 1008 85 1042 119
rect 806 17 840 51
rect 902 17 936 51
rect 1008 17 1042 51
rect 806 -51 840 -17
rect 902 -51 936 -17
rect 1008 -51 1042 -17
rect 806 -119 840 -85
rect 902 -119 936 -85
rect 1008 -119 1042 -85
rect 806 -187 840 -153
rect 902 -187 936 -153
rect 1008 -187 1042 -153
rect 806 -255 840 -221
rect 902 -255 936 -221
rect 1008 -255 1042 -221
rect 806 -323 840 -289
rect 902 -323 936 -289
rect 1008 -323 1042 -289
rect 806 -391 840 -357
rect 902 -391 936 -357
rect 1008 -391 1042 -357
rect 806 -459 840 -425
rect 902 -459 936 -425
rect 1008 -459 1042 -425
rect 806 -527 840 -493
rect 902 -527 936 -493
rect 1008 -527 1042 -493
rect 806 -595 840 -561
rect 902 -595 936 -561
rect 1008 -595 1042 -561
rect 806 -663 840 -629
rect 902 -663 936 -629
rect 1008 -663 1042 -629
rect 806 -731 840 -697
rect 902 -731 936 -697
rect 1008 -731 1042 -697
rect 806 -799 840 -765
rect 902 -799 936 -765
rect 1008 -799 1042 -765
rect 806 -867 840 -833
rect 902 -867 936 -833
rect 1008 -867 1042 -833
rect 806 -935 840 -901
rect 902 -935 936 -901
rect 1008 -935 1042 -901
rect 806 -1003 840 -969
rect 902 -1003 936 -969
rect 1008 -1003 1042 -969
rect 806 -1071 840 -1037
rect 902 -1071 936 -1037
rect 1008 -1071 1042 -1037
rect 806 -1139 840 -1105
rect 902 -1139 936 -1105
rect 1008 -1139 1042 -1105
rect 806 -1207 840 -1173
rect 902 -1207 936 -1173
rect 1008 -1207 1042 -1173
rect 806 -1275 840 -1241
rect 902 -1275 936 -1241
rect 1008 -1275 1042 -1241
rect 806 -1343 840 -1309
rect 902 -1343 936 -1309
rect 1008 -1343 1042 -1309
rect 806 -1411 840 -1377
rect 902 -1411 936 -1377
rect 1008 -1411 1042 -1377
rect 806 -1479 840 -1445
rect 902 -1479 936 -1445
rect 1008 -1479 1042 -1445
rect 806 -1547 840 -1513
rect 902 -1547 936 -1513
rect 1008 -1547 1042 -1513
rect 806 -1615 840 -1581
rect 902 -1615 936 -1581
rect 1008 -1615 1042 -1581
rect 806 -1683 840 -1649
rect 902 -1683 936 -1649
rect 1008 -1683 1042 -1649
rect 806 -1751 840 -1717
rect 902 -1751 936 -1717
rect 1008 -1751 1042 -1717
rect 806 -1819 840 -1785
rect 902 -1819 936 -1785
rect 1008 -1819 1042 -1785
rect 806 -1887 840 -1853
rect 902 -1887 936 -1853
rect 1008 -1887 1042 -1853
rect 806 -1955 840 -1921
rect 902 -1955 936 -1921
rect 1008 -1955 1042 -1921
rect 806 -2023 840 -1989
rect 902 -2023 936 -1989
rect 1008 -2023 1042 -1989
rect 806 -2091 840 -2057
rect 902 -2091 936 -2057
rect 1008 -2091 1042 -2057
rect 806 -2159 840 -2125
rect 902 -2159 936 -2125
rect 1008 -2159 1042 -2125
rect 806 -2227 840 -2193
rect 902 -2227 936 -2193
rect 1008 -2227 1042 -2193
rect 806 -2295 840 -2261
rect 902 -2295 936 -2261
rect 1008 -2295 1042 -2261
rect 806 -2363 840 -2329
rect 902 -2363 936 -2329
rect 1008 -2363 1042 -2329
rect 806 -2431 840 -2397
rect 902 -2431 936 -2397
rect 1008 -2431 1042 -2397
rect 806 -2499 840 -2465
rect 902 -2499 936 -2465
rect 1008 -2499 1042 -2465
rect 806 -2567 840 -2533
rect 902 -2567 936 -2533
rect 1008 -2567 1042 -2533
rect 806 -2635 840 -2601
rect 902 -2635 936 -2601
rect 1008 -2635 1042 -2601
rect 806 -2703 840 -2669
rect 902 -2703 936 -2669
rect 1008 -2703 1042 -2669
rect 806 -2771 840 -2737
rect 902 -2771 936 -2737
rect 1008 -2771 1042 -2737
rect 806 -2839 840 -2805
rect 902 -2839 936 -2805
rect 1008 -2839 1042 -2805
rect 806 -2907 840 -2873
rect 902 -2907 936 -2873
rect 1008 -2907 1042 -2873
rect 806 -2975 840 -2941
rect 902 -2975 936 -2941
rect 1008 -2975 1042 -2941
rect 806 -3043 840 -3009
rect 902 -3043 936 -3009
rect 1008 -3043 1042 -3009
rect 806 -3111 840 -3077
rect 902 -3111 936 -3077
rect 1008 -3111 1042 -3077
rect 806 -3179 840 -3145
rect 902 -3179 936 -3145
rect 1008 -3179 1042 -3145
rect 806 -3247 840 -3213
rect 902 -3247 936 -3213
rect 1008 -3247 1042 -3213
rect 806 -3315 840 -3281
rect 902 -3315 936 -3281
rect 1008 -3315 1042 -3281
rect 806 -3383 840 -3349
rect 902 -3383 936 -3349
rect 1008 -3383 1042 -3349
rect 806 -3451 840 -3417
rect 902 -3451 936 -3417
rect 1008 -3451 1042 -3417
rect 806 -3519 840 -3485
rect 902 -3519 936 -3485
rect 1008 -3519 1042 -3485
rect 806 -3587 840 -3553
rect 902 -3587 936 -3553
rect 1008 -3587 1042 -3553
rect 806 -3655 840 -3621
rect 902 -3655 936 -3621
rect 1008 -3655 1042 -3621
rect 806 -3723 840 -3689
rect 902 -3723 936 -3689
rect 1008 -3723 1042 -3689
rect 806 -3791 840 -3757
rect 902 -3791 936 -3757
rect 1008 -3791 1042 -3757
rect 806 -3859 840 -3825
rect 902 -3859 936 -3825
rect 1008 -3859 1042 -3825
rect 806 -3927 840 -3893
rect 902 -3927 936 -3893
rect 1008 -3927 1042 -3893
rect 806 -3995 840 -3961
rect 902 -3995 936 -3961
rect 1008 -3995 1042 -3961
rect 806 -4063 840 -4029
rect 902 -4063 936 -4029
rect 1008 -4063 1042 -4029
rect 806 -4131 840 -4097
rect 902 -4131 936 -4097
rect 1008 -4131 1042 -4097
rect 806 -4199 840 -4165
rect 902 -4199 936 -4165
rect 1008 -4199 1042 -4165
rect 806 -4267 840 -4233
rect 902 -4267 936 -4233
rect 1008 -4267 1042 -4233
rect 806 -4335 840 -4301
rect 902 -4335 936 -4301
rect 1008 -4335 1042 -4301
rect 806 -4403 840 -4369
rect 902 -4403 936 -4369
rect 1008 -4403 1042 -4369
rect 806 -4471 840 -4437
rect 902 -4471 936 -4437
rect 1008 -4471 1042 -4437
rect 806 -4539 840 -4505
rect 902 -4539 936 -4505
rect 1008 -4539 1042 -4505
rect 806 -4607 840 -4573
rect 902 -4607 936 -4573
rect 1008 -4607 1042 -4573
rect 806 -4675 840 -4641
rect 902 -4675 936 -4641
rect 1008 -4675 1042 -4641
rect 806 -4743 840 -4709
rect 902 -4743 936 -4709
rect 1008 -4743 1042 -4709
rect 806 -4811 840 -4777
rect 902 -4811 936 -4777
rect 1008 -4811 1042 -4777
rect 806 -4879 840 -4845
rect 902 -4879 936 -4845
rect 1008 -4879 1042 -4845
rect 806 -4947 840 -4913
rect 902 -4947 936 -4913
rect 1008 -4947 1042 -4913
rect 806 -5015 840 -4981
rect 902 -5015 936 -4981
rect 1008 -5015 1042 -4981
rect 1422 -5015 1524 5015
rect -1351 -5124 -1317 -5090
rect -1283 -5124 -1249 -5090
rect -1215 -5124 -1181 -5090
rect -1147 -5124 -1113 -5090
rect -735 -5124 -701 -5090
rect -667 -5124 -633 -5090
rect -599 -5124 -565 -5090
rect -531 -5124 -497 -5090
rect -119 -5124 -85 -5090
rect -51 -5124 -17 -5090
rect 17 -5124 51 -5090
rect 85 -5124 119 -5090
rect 497 -5124 531 -5090
rect 565 -5124 599 -5090
rect 633 -5124 667 -5090
rect 701 -5124 735 -5090
rect 1113 -5124 1147 -5090
rect 1181 -5124 1215 -5090
rect 1249 -5124 1283 -5090
rect 1317 -5124 1351 -5090
<< mvndiode >>
rect -1332 4981 -1132 5000
rect -1332 -4981 -1317 4981
rect -1147 -4981 -1132 4981
rect -1332 -5000 -1132 -4981
rect -716 4981 -516 5000
rect -716 -4981 -701 4981
rect -531 -4981 -516 4981
rect -716 -5000 -516 -4981
rect -100 4981 100 5000
rect -100 -4981 -85 4981
rect 85 -4981 100 4981
rect -100 -5000 100 -4981
rect 516 4981 716 5000
rect 516 -4981 531 4981
rect 701 -4981 716 4981
rect 516 -5000 716 -4981
rect 1132 4981 1332 5000
rect 1132 -4981 1147 4981
rect 1317 -4981 1332 4981
rect 1132 -5000 1332 -4981
<< mvndiodec >>
rect -1317 -4981 -1147 4981
rect -701 -4981 -531 4981
rect -85 -4981 85 4981
rect 531 -4981 701 4981
rect 1147 -4981 1317 4981
<< locali >>
rect -1540 5124 1540 5188
rect -1540 5090 -1357 5124
rect -1317 5090 -1285 5124
rect -1249 5090 -1215 5124
rect -1179 5090 -1147 5124
rect -1107 5090 -741 5124
rect -701 5090 -669 5124
rect -633 5090 -599 5124
rect -563 5090 -531 5124
rect -491 5090 -125 5124
rect -85 5090 -53 5124
rect -17 5090 17 5124
rect 53 5090 85 5124
rect 125 5090 491 5124
rect 531 5090 563 5124
rect 599 5090 633 5124
rect 669 5090 701 5124
rect 741 5090 1107 5124
rect 1147 5090 1179 5124
rect 1215 5090 1249 5124
rect 1285 5090 1317 5124
rect 1357 5090 1540 5124
rect -1540 5057 -1422 5090
rect -1540 5023 -1528 5057
rect -1494 5023 -1422 5057
rect -1540 5021 -1422 5023
rect -1540 -5021 -1528 5021
rect -1042 5057 -806 5090
rect -1042 5023 -946 5057
rect -912 5023 -806 5057
rect -1042 5021 -806 5023
rect -1008 5015 -840 5021
rect -1320 4985 -1144 5004
rect -1320 4981 -1285 4985
rect -1179 4981 -1144 4985
rect -1320 -4981 -1317 4981
rect -1147 -4981 -1144 4981
rect -1320 -4985 -1285 -4981
rect -1179 -4985 -1144 -4981
rect -1320 -5004 -1144 -4985
rect -1008 4981 -946 5015
rect -912 4981 -840 5015
rect -426 5057 -190 5090
rect -426 5023 -330 5057
rect -296 5023 -190 5057
rect -426 5021 -190 5023
rect -392 5015 -224 5021
rect -1042 4951 -946 4981
rect -912 4951 -806 4981
rect -1042 4949 -806 4951
rect -1008 4947 -840 4949
rect -1008 4913 -946 4947
rect -912 4913 -840 4947
rect -1042 4879 -946 4913
rect -912 4879 -806 4913
rect -1008 4845 -946 4879
rect -912 4845 -840 4879
rect -1008 4843 -840 4845
rect -1042 4841 -806 4843
rect -1042 4811 -946 4841
rect -912 4811 -806 4841
rect -1008 4777 -946 4811
rect -912 4777 -840 4811
rect -1008 4771 -840 4777
rect -1042 4769 -806 4771
rect -1042 4743 -946 4769
rect -912 4743 -806 4769
rect -1008 4709 -946 4743
rect -912 4709 -840 4743
rect -1008 4699 -840 4709
rect -1042 4697 -806 4699
rect -1042 4675 -946 4697
rect -912 4675 -806 4697
rect -1008 4641 -946 4675
rect -912 4641 -840 4675
rect -1008 4627 -840 4641
rect -1042 4625 -806 4627
rect -1042 4607 -946 4625
rect -912 4607 -806 4625
rect -1008 4573 -946 4607
rect -912 4573 -840 4607
rect -1008 4555 -840 4573
rect -1042 4553 -806 4555
rect -1042 4539 -946 4553
rect -912 4539 -806 4553
rect -1008 4505 -946 4539
rect -912 4505 -840 4539
rect -1008 4483 -840 4505
rect -1042 4481 -806 4483
rect -1042 4471 -946 4481
rect -912 4471 -806 4481
rect -1008 4437 -946 4471
rect -912 4437 -840 4471
rect -1008 4411 -840 4437
rect -1042 4409 -806 4411
rect -1042 4403 -946 4409
rect -912 4403 -806 4409
rect -1008 4369 -946 4403
rect -912 4369 -840 4403
rect -1008 4339 -840 4369
rect -1042 4337 -806 4339
rect -1042 4335 -946 4337
rect -912 4335 -806 4337
rect -1008 4301 -946 4335
rect -912 4301 -840 4335
rect -1008 4267 -840 4301
rect -1008 4233 -946 4267
rect -912 4233 -840 4267
rect -1042 4231 -946 4233
rect -912 4231 -806 4233
rect -1042 4229 -806 4231
rect -1008 4199 -840 4229
rect -1008 4165 -946 4199
rect -912 4165 -840 4199
rect -1042 4159 -946 4165
rect -912 4159 -806 4165
rect -1042 4157 -806 4159
rect -1008 4131 -840 4157
rect -1008 4097 -946 4131
rect -912 4097 -840 4131
rect -1042 4087 -946 4097
rect -912 4087 -806 4097
rect -1042 4085 -806 4087
rect -1008 4063 -840 4085
rect -1008 4029 -946 4063
rect -912 4029 -840 4063
rect -1042 4015 -946 4029
rect -912 4015 -806 4029
rect -1042 4013 -806 4015
rect -1008 3995 -840 4013
rect -1008 3961 -946 3995
rect -912 3961 -840 3995
rect -1042 3943 -946 3961
rect -912 3943 -806 3961
rect -1042 3941 -806 3943
rect -1008 3927 -840 3941
rect -1008 3893 -946 3927
rect -912 3893 -840 3927
rect -1042 3871 -946 3893
rect -912 3871 -806 3893
rect -1042 3869 -806 3871
rect -1008 3859 -840 3869
rect -1008 3825 -946 3859
rect -912 3825 -840 3859
rect -1042 3799 -946 3825
rect -912 3799 -806 3825
rect -1042 3797 -806 3799
rect -1008 3791 -840 3797
rect -1008 3757 -946 3791
rect -912 3757 -840 3791
rect -1042 3727 -946 3757
rect -912 3727 -806 3757
rect -1042 3725 -806 3727
rect -1008 3723 -840 3725
rect -1008 3689 -946 3723
rect -912 3689 -840 3723
rect -1042 3655 -946 3689
rect -912 3655 -806 3689
rect -1008 3621 -946 3655
rect -912 3621 -840 3655
rect -1008 3619 -840 3621
rect -1042 3617 -806 3619
rect -1042 3587 -946 3617
rect -912 3587 -806 3617
rect -1008 3553 -946 3587
rect -912 3553 -840 3587
rect -1008 3547 -840 3553
rect -1042 3545 -806 3547
rect -1042 3519 -946 3545
rect -912 3519 -806 3545
rect -1008 3485 -946 3519
rect -912 3485 -840 3519
rect -1008 3475 -840 3485
rect -1042 3473 -806 3475
rect -1042 3451 -946 3473
rect -912 3451 -806 3473
rect -1008 3417 -946 3451
rect -912 3417 -840 3451
rect -1008 3403 -840 3417
rect -1042 3401 -806 3403
rect -1042 3383 -946 3401
rect -912 3383 -806 3401
rect -1008 3349 -946 3383
rect -912 3349 -840 3383
rect -1008 3331 -840 3349
rect -1042 3329 -806 3331
rect -1042 3315 -946 3329
rect -912 3315 -806 3329
rect -1008 3281 -946 3315
rect -912 3281 -840 3315
rect -1008 3259 -840 3281
rect -1042 3257 -806 3259
rect -1042 3247 -946 3257
rect -912 3247 -806 3257
rect -1008 3213 -946 3247
rect -912 3213 -840 3247
rect -1008 3187 -840 3213
rect -1042 3185 -806 3187
rect -1042 3179 -946 3185
rect -912 3179 -806 3185
rect -1008 3145 -946 3179
rect -912 3145 -840 3179
rect -1008 3115 -840 3145
rect -1042 3113 -806 3115
rect -1042 3111 -946 3113
rect -912 3111 -806 3113
rect -1008 3077 -946 3111
rect -912 3077 -840 3111
rect -1008 3043 -840 3077
rect -1008 3009 -946 3043
rect -912 3009 -840 3043
rect -1042 3007 -946 3009
rect -912 3007 -806 3009
rect -1042 3005 -806 3007
rect -1008 2975 -840 3005
rect -1008 2941 -946 2975
rect -912 2941 -840 2975
rect -1042 2935 -946 2941
rect -912 2935 -806 2941
rect -1042 2933 -806 2935
rect -1008 2907 -840 2933
rect -1008 2873 -946 2907
rect -912 2873 -840 2907
rect -1042 2863 -946 2873
rect -912 2863 -806 2873
rect -1042 2861 -806 2863
rect -1008 2839 -840 2861
rect -1008 2805 -946 2839
rect -912 2805 -840 2839
rect -1042 2791 -946 2805
rect -912 2791 -806 2805
rect -1042 2789 -806 2791
rect -1008 2771 -840 2789
rect -1008 2737 -946 2771
rect -912 2737 -840 2771
rect -1042 2719 -946 2737
rect -912 2719 -806 2737
rect -1042 2717 -806 2719
rect -1008 2703 -840 2717
rect -1008 2669 -946 2703
rect -912 2669 -840 2703
rect -1042 2647 -946 2669
rect -912 2647 -806 2669
rect -1042 2645 -806 2647
rect -1008 2635 -840 2645
rect -1008 2601 -946 2635
rect -912 2601 -840 2635
rect -1042 2575 -946 2601
rect -912 2575 -806 2601
rect -1042 2573 -806 2575
rect -1008 2567 -840 2573
rect -1008 2533 -946 2567
rect -912 2533 -840 2567
rect -1042 2503 -946 2533
rect -912 2503 -806 2533
rect -1042 2501 -806 2503
rect -1008 2499 -840 2501
rect -1008 2465 -946 2499
rect -912 2465 -840 2499
rect -1042 2431 -946 2465
rect -912 2431 -806 2465
rect -1008 2397 -946 2431
rect -912 2397 -840 2431
rect -1008 2395 -840 2397
rect -1042 2393 -806 2395
rect -1042 2363 -946 2393
rect -912 2363 -806 2393
rect -1008 2329 -946 2363
rect -912 2329 -840 2363
rect -1008 2323 -840 2329
rect -1042 2321 -806 2323
rect -1042 2295 -946 2321
rect -912 2295 -806 2321
rect -1008 2261 -946 2295
rect -912 2261 -840 2295
rect -1008 2251 -840 2261
rect -1042 2249 -806 2251
rect -1042 2227 -946 2249
rect -912 2227 -806 2249
rect -1008 2193 -946 2227
rect -912 2193 -840 2227
rect -1008 2179 -840 2193
rect -1042 2177 -806 2179
rect -1042 2159 -946 2177
rect -912 2159 -806 2177
rect -1008 2125 -946 2159
rect -912 2125 -840 2159
rect -1008 2107 -840 2125
rect -1042 2105 -806 2107
rect -1042 2091 -946 2105
rect -912 2091 -806 2105
rect -1008 2057 -946 2091
rect -912 2057 -840 2091
rect -1008 2035 -840 2057
rect -1042 2033 -806 2035
rect -1042 2023 -946 2033
rect -912 2023 -806 2033
rect -1008 1989 -946 2023
rect -912 1989 -840 2023
rect -1008 1963 -840 1989
rect -1042 1961 -806 1963
rect -1042 1955 -946 1961
rect -912 1955 -806 1961
rect -1008 1921 -946 1955
rect -912 1921 -840 1955
rect -1008 1891 -840 1921
rect -1042 1889 -806 1891
rect -1042 1887 -946 1889
rect -912 1887 -806 1889
rect -1008 1853 -946 1887
rect -912 1853 -840 1887
rect -1008 1819 -840 1853
rect -1008 1785 -946 1819
rect -912 1785 -840 1819
rect -1042 1783 -946 1785
rect -912 1783 -806 1785
rect -1042 1781 -806 1783
rect -1008 1751 -840 1781
rect -1008 1717 -946 1751
rect -912 1717 -840 1751
rect -1042 1711 -946 1717
rect -912 1711 -806 1717
rect -1042 1709 -806 1711
rect -1008 1683 -840 1709
rect -1008 1649 -946 1683
rect -912 1649 -840 1683
rect -1042 1639 -946 1649
rect -912 1639 -806 1649
rect -1042 1637 -806 1639
rect -1008 1615 -840 1637
rect -1008 1581 -946 1615
rect -912 1581 -840 1615
rect -1042 1567 -946 1581
rect -912 1567 -806 1581
rect -1042 1565 -806 1567
rect -1008 1547 -840 1565
rect -1008 1513 -946 1547
rect -912 1513 -840 1547
rect -1042 1495 -946 1513
rect -912 1495 -806 1513
rect -1042 1493 -806 1495
rect -1008 1479 -840 1493
rect -1008 1445 -946 1479
rect -912 1445 -840 1479
rect -1042 1423 -946 1445
rect -912 1423 -806 1445
rect -1042 1421 -806 1423
rect -1008 1411 -840 1421
rect -1008 1377 -946 1411
rect -912 1377 -840 1411
rect -1042 1351 -946 1377
rect -912 1351 -806 1377
rect -1042 1349 -806 1351
rect -1008 1343 -840 1349
rect -1008 1309 -946 1343
rect -912 1309 -840 1343
rect -1042 1279 -946 1309
rect -912 1279 -806 1309
rect -1042 1277 -806 1279
rect -1008 1275 -840 1277
rect -1008 1241 -946 1275
rect -912 1241 -840 1275
rect -1042 1207 -946 1241
rect -912 1207 -806 1241
rect -1008 1173 -946 1207
rect -912 1173 -840 1207
rect -1008 1171 -840 1173
rect -1042 1169 -806 1171
rect -1042 1139 -946 1169
rect -912 1139 -806 1169
rect -1008 1105 -946 1139
rect -912 1105 -840 1139
rect -1008 1099 -840 1105
rect -1042 1097 -806 1099
rect -1042 1071 -946 1097
rect -912 1071 -806 1097
rect -1008 1037 -946 1071
rect -912 1037 -840 1071
rect -1008 1027 -840 1037
rect -1042 1025 -806 1027
rect -1042 1003 -946 1025
rect -912 1003 -806 1025
rect -1008 969 -946 1003
rect -912 969 -840 1003
rect -1008 955 -840 969
rect -1042 953 -806 955
rect -1042 935 -946 953
rect -912 935 -806 953
rect -1008 901 -946 935
rect -912 901 -840 935
rect -1008 883 -840 901
rect -1042 881 -806 883
rect -1042 867 -946 881
rect -912 867 -806 881
rect -1008 833 -946 867
rect -912 833 -840 867
rect -1008 811 -840 833
rect -1042 809 -806 811
rect -1042 799 -946 809
rect -912 799 -806 809
rect -1008 765 -946 799
rect -912 765 -840 799
rect -1008 739 -840 765
rect -1042 737 -806 739
rect -1042 731 -946 737
rect -912 731 -806 737
rect -1008 697 -946 731
rect -912 697 -840 731
rect -1008 667 -840 697
rect -1042 665 -806 667
rect -1042 663 -946 665
rect -912 663 -806 665
rect -1008 629 -946 663
rect -912 629 -840 663
rect -1008 595 -840 629
rect -1008 561 -946 595
rect -912 561 -840 595
rect -1042 559 -946 561
rect -912 559 -806 561
rect -1042 557 -806 559
rect -1008 527 -840 557
rect -1008 493 -946 527
rect -912 493 -840 527
rect -1042 487 -946 493
rect -912 487 -806 493
rect -1042 485 -806 487
rect -1008 459 -840 485
rect -1008 425 -946 459
rect -912 425 -840 459
rect -1042 415 -946 425
rect -912 415 -806 425
rect -1042 413 -806 415
rect -1008 391 -840 413
rect -1008 357 -946 391
rect -912 357 -840 391
rect -1042 343 -946 357
rect -912 343 -806 357
rect -1042 341 -806 343
rect -1008 323 -840 341
rect -1008 289 -946 323
rect -912 289 -840 323
rect -1042 271 -946 289
rect -912 271 -806 289
rect -1042 269 -806 271
rect -1008 255 -840 269
rect -1008 221 -946 255
rect -912 221 -840 255
rect -1042 199 -946 221
rect -912 199 -806 221
rect -1042 197 -806 199
rect -1008 187 -840 197
rect -1008 153 -946 187
rect -912 153 -840 187
rect -1042 127 -946 153
rect -912 127 -806 153
rect -1042 125 -806 127
rect -1008 119 -840 125
rect -1008 85 -946 119
rect -912 85 -840 119
rect -1042 55 -946 85
rect -912 55 -806 85
rect -1042 53 -806 55
rect -1008 51 -840 53
rect -1008 17 -946 51
rect -912 17 -840 51
rect -1042 -17 -946 17
rect -912 -17 -806 17
rect -1008 -51 -946 -17
rect -912 -51 -840 -17
rect -1008 -53 -840 -51
rect -1042 -55 -806 -53
rect -1042 -85 -946 -55
rect -912 -85 -806 -55
rect -1008 -119 -946 -85
rect -912 -119 -840 -85
rect -1008 -125 -840 -119
rect -1042 -127 -806 -125
rect -1042 -153 -946 -127
rect -912 -153 -806 -127
rect -1008 -187 -946 -153
rect -912 -187 -840 -153
rect -1008 -197 -840 -187
rect -1042 -199 -806 -197
rect -1042 -221 -946 -199
rect -912 -221 -806 -199
rect -1008 -255 -946 -221
rect -912 -255 -840 -221
rect -1008 -269 -840 -255
rect -1042 -271 -806 -269
rect -1042 -289 -946 -271
rect -912 -289 -806 -271
rect -1008 -323 -946 -289
rect -912 -323 -840 -289
rect -1008 -341 -840 -323
rect -1042 -343 -806 -341
rect -1042 -357 -946 -343
rect -912 -357 -806 -343
rect -1008 -391 -946 -357
rect -912 -391 -840 -357
rect -1008 -413 -840 -391
rect -1042 -415 -806 -413
rect -1042 -425 -946 -415
rect -912 -425 -806 -415
rect -1008 -459 -946 -425
rect -912 -459 -840 -425
rect -1008 -485 -840 -459
rect -1042 -487 -806 -485
rect -1042 -493 -946 -487
rect -912 -493 -806 -487
rect -1008 -527 -946 -493
rect -912 -527 -840 -493
rect -1008 -557 -840 -527
rect -1042 -559 -806 -557
rect -1042 -561 -946 -559
rect -912 -561 -806 -559
rect -1008 -595 -946 -561
rect -912 -595 -840 -561
rect -1008 -629 -840 -595
rect -1008 -663 -946 -629
rect -912 -663 -840 -629
rect -1042 -665 -946 -663
rect -912 -665 -806 -663
rect -1042 -667 -806 -665
rect -1008 -697 -840 -667
rect -1008 -731 -946 -697
rect -912 -731 -840 -697
rect -1042 -737 -946 -731
rect -912 -737 -806 -731
rect -1042 -739 -806 -737
rect -1008 -765 -840 -739
rect -1008 -799 -946 -765
rect -912 -799 -840 -765
rect -1042 -809 -946 -799
rect -912 -809 -806 -799
rect -1042 -811 -806 -809
rect -1008 -833 -840 -811
rect -1008 -867 -946 -833
rect -912 -867 -840 -833
rect -1042 -881 -946 -867
rect -912 -881 -806 -867
rect -1042 -883 -806 -881
rect -1008 -901 -840 -883
rect -1008 -935 -946 -901
rect -912 -935 -840 -901
rect -1042 -953 -946 -935
rect -912 -953 -806 -935
rect -1042 -955 -806 -953
rect -1008 -969 -840 -955
rect -1008 -1003 -946 -969
rect -912 -1003 -840 -969
rect -1042 -1025 -946 -1003
rect -912 -1025 -806 -1003
rect -1042 -1027 -806 -1025
rect -1008 -1037 -840 -1027
rect -1008 -1071 -946 -1037
rect -912 -1071 -840 -1037
rect -1042 -1097 -946 -1071
rect -912 -1097 -806 -1071
rect -1042 -1099 -806 -1097
rect -1008 -1105 -840 -1099
rect -1008 -1139 -946 -1105
rect -912 -1139 -840 -1105
rect -1042 -1169 -946 -1139
rect -912 -1169 -806 -1139
rect -1042 -1171 -806 -1169
rect -1008 -1173 -840 -1171
rect -1008 -1207 -946 -1173
rect -912 -1207 -840 -1173
rect -1042 -1241 -946 -1207
rect -912 -1241 -806 -1207
rect -1008 -1275 -946 -1241
rect -912 -1275 -840 -1241
rect -1008 -1277 -840 -1275
rect -1042 -1279 -806 -1277
rect -1042 -1309 -946 -1279
rect -912 -1309 -806 -1279
rect -1008 -1343 -946 -1309
rect -912 -1343 -840 -1309
rect -1008 -1349 -840 -1343
rect -1042 -1351 -806 -1349
rect -1042 -1377 -946 -1351
rect -912 -1377 -806 -1351
rect -1008 -1411 -946 -1377
rect -912 -1411 -840 -1377
rect -1008 -1421 -840 -1411
rect -1042 -1423 -806 -1421
rect -1042 -1445 -946 -1423
rect -912 -1445 -806 -1423
rect -1008 -1479 -946 -1445
rect -912 -1479 -840 -1445
rect -1008 -1493 -840 -1479
rect -1042 -1495 -806 -1493
rect -1042 -1513 -946 -1495
rect -912 -1513 -806 -1495
rect -1008 -1547 -946 -1513
rect -912 -1547 -840 -1513
rect -1008 -1565 -840 -1547
rect -1042 -1567 -806 -1565
rect -1042 -1581 -946 -1567
rect -912 -1581 -806 -1567
rect -1008 -1615 -946 -1581
rect -912 -1615 -840 -1581
rect -1008 -1637 -840 -1615
rect -1042 -1639 -806 -1637
rect -1042 -1649 -946 -1639
rect -912 -1649 -806 -1639
rect -1008 -1683 -946 -1649
rect -912 -1683 -840 -1649
rect -1008 -1709 -840 -1683
rect -1042 -1711 -806 -1709
rect -1042 -1717 -946 -1711
rect -912 -1717 -806 -1711
rect -1008 -1751 -946 -1717
rect -912 -1751 -840 -1717
rect -1008 -1781 -840 -1751
rect -1042 -1783 -806 -1781
rect -1042 -1785 -946 -1783
rect -912 -1785 -806 -1783
rect -1008 -1819 -946 -1785
rect -912 -1819 -840 -1785
rect -1008 -1853 -840 -1819
rect -1008 -1887 -946 -1853
rect -912 -1887 -840 -1853
rect -1042 -1889 -946 -1887
rect -912 -1889 -806 -1887
rect -1042 -1891 -806 -1889
rect -1008 -1921 -840 -1891
rect -1008 -1955 -946 -1921
rect -912 -1955 -840 -1921
rect -1042 -1961 -946 -1955
rect -912 -1961 -806 -1955
rect -1042 -1963 -806 -1961
rect -1008 -1989 -840 -1963
rect -1008 -2023 -946 -1989
rect -912 -2023 -840 -1989
rect -1042 -2033 -946 -2023
rect -912 -2033 -806 -2023
rect -1042 -2035 -806 -2033
rect -1008 -2057 -840 -2035
rect -1008 -2091 -946 -2057
rect -912 -2091 -840 -2057
rect -1042 -2105 -946 -2091
rect -912 -2105 -806 -2091
rect -1042 -2107 -806 -2105
rect -1008 -2125 -840 -2107
rect -1008 -2159 -946 -2125
rect -912 -2159 -840 -2125
rect -1042 -2177 -946 -2159
rect -912 -2177 -806 -2159
rect -1042 -2179 -806 -2177
rect -1008 -2193 -840 -2179
rect -1008 -2227 -946 -2193
rect -912 -2227 -840 -2193
rect -1042 -2249 -946 -2227
rect -912 -2249 -806 -2227
rect -1042 -2251 -806 -2249
rect -1008 -2261 -840 -2251
rect -1008 -2295 -946 -2261
rect -912 -2295 -840 -2261
rect -1042 -2321 -946 -2295
rect -912 -2321 -806 -2295
rect -1042 -2323 -806 -2321
rect -1008 -2329 -840 -2323
rect -1008 -2363 -946 -2329
rect -912 -2363 -840 -2329
rect -1042 -2393 -946 -2363
rect -912 -2393 -806 -2363
rect -1042 -2395 -806 -2393
rect -1008 -2397 -840 -2395
rect -1008 -2431 -946 -2397
rect -912 -2431 -840 -2397
rect -1042 -2465 -946 -2431
rect -912 -2465 -806 -2431
rect -1008 -2499 -946 -2465
rect -912 -2499 -840 -2465
rect -1008 -2501 -840 -2499
rect -1042 -2503 -806 -2501
rect -1042 -2533 -946 -2503
rect -912 -2533 -806 -2503
rect -1008 -2567 -946 -2533
rect -912 -2567 -840 -2533
rect -1008 -2573 -840 -2567
rect -1042 -2575 -806 -2573
rect -1042 -2601 -946 -2575
rect -912 -2601 -806 -2575
rect -1008 -2635 -946 -2601
rect -912 -2635 -840 -2601
rect -1008 -2645 -840 -2635
rect -1042 -2647 -806 -2645
rect -1042 -2669 -946 -2647
rect -912 -2669 -806 -2647
rect -1008 -2703 -946 -2669
rect -912 -2703 -840 -2669
rect -1008 -2717 -840 -2703
rect -1042 -2719 -806 -2717
rect -1042 -2737 -946 -2719
rect -912 -2737 -806 -2719
rect -1008 -2771 -946 -2737
rect -912 -2771 -840 -2737
rect -1008 -2789 -840 -2771
rect -1042 -2791 -806 -2789
rect -1042 -2805 -946 -2791
rect -912 -2805 -806 -2791
rect -1008 -2839 -946 -2805
rect -912 -2839 -840 -2805
rect -1008 -2861 -840 -2839
rect -1042 -2863 -806 -2861
rect -1042 -2873 -946 -2863
rect -912 -2873 -806 -2863
rect -1008 -2907 -946 -2873
rect -912 -2907 -840 -2873
rect -1008 -2933 -840 -2907
rect -1042 -2935 -806 -2933
rect -1042 -2941 -946 -2935
rect -912 -2941 -806 -2935
rect -1008 -2975 -946 -2941
rect -912 -2975 -840 -2941
rect -1008 -3005 -840 -2975
rect -1042 -3007 -806 -3005
rect -1042 -3009 -946 -3007
rect -912 -3009 -806 -3007
rect -1008 -3043 -946 -3009
rect -912 -3043 -840 -3009
rect -1008 -3077 -840 -3043
rect -1008 -3111 -946 -3077
rect -912 -3111 -840 -3077
rect -1042 -3113 -946 -3111
rect -912 -3113 -806 -3111
rect -1042 -3115 -806 -3113
rect -1008 -3145 -840 -3115
rect -1008 -3179 -946 -3145
rect -912 -3179 -840 -3145
rect -1042 -3185 -946 -3179
rect -912 -3185 -806 -3179
rect -1042 -3187 -806 -3185
rect -1008 -3213 -840 -3187
rect -1008 -3247 -946 -3213
rect -912 -3247 -840 -3213
rect -1042 -3257 -946 -3247
rect -912 -3257 -806 -3247
rect -1042 -3259 -806 -3257
rect -1008 -3281 -840 -3259
rect -1008 -3315 -946 -3281
rect -912 -3315 -840 -3281
rect -1042 -3329 -946 -3315
rect -912 -3329 -806 -3315
rect -1042 -3331 -806 -3329
rect -1008 -3349 -840 -3331
rect -1008 -3383 -946 -3349
rect -912 -3383 -840 -3349
rect -1042 -3401 -946 -3383
rect -912 -3401 -806 -3383
rect -1042 -3403 -806 -3401
rect -1008 -3417 -840 -3403
rect -1008 -3451 -946 -3417
rect -912 -3451 -840 -3417
rect -1042 -3473 -946 -3451
rect -912 -3473 -806 -3451
rect -1042 -3475 -806 -3473
rect -1008 -3485 -840 -3475
rect -1008 -3519 -946 -3485
rect -912 -3519 -840 -3485
rect -1042 -3545 -946 -3519
rect -912 -3545 -806 -3519
rect -1042 -3547 -806 -3545
rect -1008 -3553 -840 -3547
rect -1008 -3587 -946 -3553
rect -912 -3587 -840 -3553
rect -1042 -3617 -946 -3587
rect -912 -3617 -806 -3587
rect -1042 -3619 -806 -3617
rect -1008 -3621 -840 -3619
rect -1008 -3655 -946 -3621
rect -912 -3655 -840 -3621
rect -1042 -3689 -946 -3655
rect -912 -3689 -806 -3655
rect -1008 -3723 -946 -3689
rect -912 -3723 -840 -3689
rect -1008 -3725 -840 -3723
rect -1042 -3727 -806 -3725
rect -1042 -3757 -946 -3727
rect -912 -3757 -806 -3727
rect -1008 -3791 -946 -3757
rect -912 -3791 -840 -3757
rect -1008 -3797 -840 -3791
rect -1042 -3799 -806 -3797
rect -1042 -3825 -946 -3799
rect -912 -3825 -806 -3799
rect -1008 -3859 -946 -3825
rect -912 -3859 -840 -3825
rect -1008 -3869 -840 -3859
rect -1042 -3871 -806 -3869
rect -1042 -3893 -946 -3871
rect -912 -3893 -806 -3871
rect -1008 -3927 -946 -3893
rect -912 -3927 -840 -3893
rect -1008 -3941 -840 -3927
rect -1042 -3943 -806 -3941
rect -1042 -3961 -946 -3943
rect -912 -3961 -806 -3943
rect -1008 -3995 -946 -3961
rect -912 -3995 -840 -3961
rect -1008 -4013 -840 -3995
rect -1042 -4015 -806 -4013
rect -1042 -4029 -946 -4015
rect -912 -4029 -806 -4015
rect -1008 -4063 -946 -4029
rect -912 -4063 -840 -4029
rect -1008 -4085 -840 -4063
rect -1042 -4087 -806 -4085
rect -1042 -4097 -946 -4087
rect -912 -4097 -806 -4087
rect -1008 -4131 -946 -4097
rect -912 -4131 -840 -4097
rect -1008 -4157 -840 -4131
rect -1042 -4159 -806 -4157
rect -1042 -4165 -946 -4159
rect -912 -4165 -806 -4159
rect -1008 -4199 -946 -4165
rect -912 -4199 -840 -4165
rect -1008 -4229 -840 -4199
rect -1042 -4231 -806 -4229
rect -1042 -4233 -946 -4231
rect -912 -4233 -806 -4231
rect -1008 -4267 -946 -4233
rect -912 -4267 -840 -4233
rect -1008 -4301 -840 -4267
rect -1008 -4335 -946 -4301
rect -912 -4335 -840 -4301
rect -1042 -4337 -946 -4335
rect -912 -4337 -806 -4335
rect -1042 -4339 -806 -4337
rect -1008 -4369 -840 -4339
rect -1008 -4403 -946 -4369
rect -912 -4403 -840 -4369
rect -1042 -4409 -946 -4403
rect -912 -4409 -806 -4403
rect -1042 -4411 -806 -4409
rect -1008 -4437 -840 -4411
rect -1008 -4471 -946 -4437
rect -912 -4471 -840 -4437
rect -1042 -4481 -946 -4471
rect -912 -4481 -806 -4471
rect -1042 -4483 -806 -4481
rect -1008 -4505 -840 -4483
rect -1008 -4539 -946 -4505
rect -912 -4539 -840 -4505
rect -1042 -4553 -946 -4539
rect -912 -4553 -806 -4539
rect -1042 -4555 -806 -4553
rect -1008 -4573 -840 -4555
rect -1008 -4607 -946 -4573
rect -912 -4607 -840 -4573
rect -1042 -4625 -946 -4607
rect -912 -4625 -806 -4607
rect -1042 -4627 -806 -4625
rect -1008 -4641 -840 -4627
rect -1008 -4675 -946 -4641
rect -912 -4675 -840 -4641
rect -1042 -4697 -946 -4675
rect -912 -4697 -806 -4675
rect -1042 -4699 -806 -4697
rect -1008 -4709 -840 -4699
rect -1008 -4743 -946 -4709
rect -912 -4743 -840 -4709
rect -1042 -4769 -946 -4743
rect -912 -4769 -806 -4743
rect -1042 -4771 -806 -4769
rect -1008 -4777 -840 -4771
rect -1008 -4811 -946 -4777
rect -912 -4811 -840 -4777
rect -1042 -4841 -946 -4811
rect -912 -4841 -806 -4811
rect -1042 -4843 -806 -4841
rect -1008 -4845 -840 -4843
rect -1008 -4879 -946 -4845
rect -912 -4879 -840 -4845
rect -1042 -4913 -946 -4879
rect -912 -4913 -806 -4879
rect -1008 -4947 -946 -4913
rect -912 -4947 -840 -4913
rect -1008 -4949 -840 -4947
rect -1042 -4951 -806 -4949
rect -1042 -4981 -946 -4951
rect -912 -4981 -806 -4951
rect -1540 -5023 -1422 -5021
rect -1540 -5057 -1528 -5023
rect -1494 -5057 -1422 -5023
rect -1540 -5090 -1422 -5057
rect -1008 -5015 -946 -4981
rect -912 -5015 -840 -4981
rect -704 4985 -528 5004
rect -704 4981 -669 4985
rect -563 4981 -528 4985
rect -704 -4981 -701 4981
rect -531 -4981 -528 4981
rect -704 -4985 -669 -4981
rect -563 -4985 -528 -4981
rect -704 -5004 -528 -4985
rect -392 4981 -330 5015
rect -296 4981 -224 5015
rect 190 5057 426 5090
rect 190 5023 286 5057
rect 320 5023 426 5057
rect 190 5021 426 5023
rect 224 5015 392 5021
rect -426 4951 -330 4981
rect -296 4951 -190 4981
rect -426 4949 -190 4951
rect -392 4947 -224 4949
rect -392 4913 -330 4947
rect -296 4913 -224 4947
rect -426 4879 -330 4913
rect -296 4879 -190 4913
rect -392 4845 -330 4879
rect -296 4845 -224 4879
rect -392 4843 -224 4845
rect -426 4841 -190 4843
rect -426 4811 -330 4841
rect -296 4811 -190 4841
rect -392 4777 -330 4811
rect -296 4777 -224 4811
rect -392 4771 -224 4777
rect -426 4769 -190 4771
rect -426 4743 -330 4769
rect -296 4743 -190 4769
rect -392 4709 -330 4743
rect -296 4709 -224 4743
rect -392 4699 -224 4709
rect -426 4697 -190 4699
rect -426 4675 -330 4697
rect -296 4675 -190 4697
rect -392 4641 -330 4675
rect -296 4641 -224 4675
rect -392 4627 -224 4641
rect -426 4625 -190 4627
rect -426 4607 -330 4625
rect -296 4607 -190 4625
rect -392 4573 -330 4607
rect -296 4573 -224 4607
rect -392 4555 -224 4573
rect -426 4553 -190 4555
rect -426 4539 -330 4553
rect -296 4539 -190 4553
rect -392 4505 -330 4539
rect -296 4505 -224 4539
rect -392 4483 -224 4505
rect -426 4481 -190 4483
rect -426 4471 -330 4481
rect -296 4471 -190 4481
rect -392 4437 -330 4471
rect -296 4437 -224 4471
rect -392 4411 -224 4437
rect -426 4409 -190 4411
rect -426 4403 -330 4409
rect -296 4403 -190 4409
rect -392 4369 -330 4403
rect -296 4369 -224 4403
rect -392 4339 -224 4369
rect -426 4337 -190 4339
rect -426 4335 -330 4337
rect -296 4335 -190 4337
rect -392 4301 -330 4335
rect -296 4301 -224 4335
rect -392 4267 -224 4301
rect -392 4233 -330 4267
rect -296 4233 -224 4267
rect -426 4231 -330 4233
rect -296 4231 -190 4233
rect -426 4229 -190 4231
rect -392 4199 -224 4229
rect -392 4165 -330 4199
rect -296 4165 -224 4199
rect -426 4159 -330 4165
rect -296 4159 -190 4165
rect -426 4157 -190 4159
rect -392 4131 -224 4157
rect -392 4097 -330 4131
rect -296 4097 -224 4131
rect -426 4087 -330 4097
rect -296 4087 -190 4097
rect -426 4085 -190 4087
rect -392 4063 -224 4085
rect -392 4029 -330 4063
rect -296 4029 -224 4063
rect -426 4015 -330 4029
rect -296 4015 -190 4029
rect -426 4013 -190 4015
rect -392 3995 -224 4013
rect -392 3961 -330 3995
rect -296 3961 -224 3995
rect -426 3943 -330 3961
rect -296 3943 -190 3961
rect -426 3941 -190 3943
rect -392 3927 -224 3941
rect -392 3893 -330 3927
rect -296 3893 -224 3927
rect -426 3871 -330 3893
rect -296 3871 -190 3893
rect -426 3869 -190 3871
rect -392 3859 -224 3869
rect -392 3825 -330 3859
rect -296 3825 -224 3859
rect -426 3799 -330 3825
rect -296 3799 -190 3825
rect -426 3797 -190 3799
rect -392 3791 -224 3797
rect -392 3757 -330 3791
rect -296 3757 -224 3791
rect -426 3727 -330 3757
rect -296 3727 -190 3757
rect -426 3725 -190 3727
rect -392 3723 -224 3725
rect -392 3689 -330 3723
rect -296 3689 -224 3723
rect -426 3655 -330 3689
rect -296 3655 -190 3689
rect -392 3621 -330 3655
rect -296 3621 -224 3655
rect -392 3619 -224 3621
rect -426 3617 -190 3619
rect -426 3587 -330 3617
rect -296 3587 -190 3617
rect -392 3553 -330 3587
rect -296 3553 -224 3587
rect -392 3547 -224 3553
rect -426 3545 -190 3547
rect -426 3519 -330 3545
rect -296 3519 -190 3545
rect -392 3485 -330 3519
rect -296 3485 -224 3519
rect -392 3475 -224 3485
rect -426 3473 -190 3475
rect -426 3451 -330 3473
rect -296 3451 -190 3473
rect -392 3417 -330 3451
rect -296 3417 -224 3451
rect -392 3403 -224 3417
rect -426 3401 -190 3403
rect -426 3383 -330 3401
rect -296 3383 -190 3401
rect -392 3349 -330 3383
rect -296 3349 -224 3383
rect -392 3331 -224 3349
rect -426 3329 -190 3331
rect -426 3315 -330 3329
rect -296 3315 -190 3329
rect -392 3281 -330 3315
rect -296 3281 -224 3315
rect -392 3259 -224 3281
rect -426 3257 -190 3259
rect -426 3247 -330 3257
rect -296 3247 -190 3257
rect -392 3213 -330 3247
rect -296 3213 -224 3247
rect -392 3187 -224 3213
rect -426 3185 -190 3187
rect -426 3179 -330 3185
rect -296 3179 -190 3185
rect -392 3145 -330 3179
rect -296 3145 -224 3179
rect -392 3115 -224 3145
rect -426 3113 -190 3115
rect -426 3111 -330 3113
rect -296 3111 -190 3113
rect -392 3077 -330 3111
rect -296 3077 -224 3111
rect -392 3043 -224 3077
rect -392 3009 -330 3043
rect -296 3009 -224 3043
rect -426 3007 -330 3009
rect -296 3007 -190 3009
rect -426 3005 -190 3007
rect -392 2975 -224 3005
rect -392 2941 -330 2975
rect -296 2941 -224 2975
rect -426 2935 -330 2941
rect -296 2935 -190 2941
rect -426 2933 -190 2935
rect -392 2907 -224 2933
rect -392 2873 -330 2907
rect -296 2873 -224 2907
rect -426 2863 -330 2873
rect -296 2863 -190 2873
rect -426 2861 -190 2863
rect -392 2839 -224 2861
rect -392 2805 -330 2839
rect -296 2805 -224 2839
rect -426 2791 -330 2805
rect -296 2791 -190 2805
rect -426 2789 -190 2791
rect -392 2771 -224 2789
rect -392 2737 -330 2771
rect -296 2737 -224 2771
rect -426 2719 -330 2737
rect -296 2719 -190 2737
rect -426 2717 -190 2719
rect -392 2703 -224 2717
rect -392 2669 -330 2703
rect -296 2669 -224 2703
rect -426 2647 -330 2669
rect -296 2647 -190 2669
rect -426 2645 -190 2647
rect -392 2635 -224 2645
rect -392 2601 -330 2635
rect -296 2601 -224 2635
rect -426 2575 -330 2601
rect -296 2575 -190 2601
rect -426 2573 -190 2575
rect -392 2567 -224 2573
rect -392 2533 -330 2567
rect -296 2533 -224 2567
rect -426 2503 -330 2533
rect -296 2503 -190 2533
rect -426 2501 -190 2503
rect -392 2499 -224 2501
rect -392 2465 -330 2499
rect -296 2465 -224 2499
rect -426 2431 -330 2465
rect -296 2431 -190 2465
rect -392 2397 -330 2431
rect -296 2397 -224 2431
rect -392 2395 -224 2397
rect -426 2393 -190 2395
rect -426 2363 -330 2393
rect -296 2363 -190 2393
rect -392 2329 -330 2363
rect -296 2329 -224 2363
rect -392 2323 -224 2329
rect -426 2321 -190 2323
rect -426 2295 -330 2321
rect -296 2295 -190 2321
rect -392 2261 -330 2295
rect -296 2261 -224 2295
rect -392 2251 -224 2261
rect -426 2249 -190 2251
rect -426 2227 -330 2249
rect -296 2227 -190 2249
rect -392 2193 -330 2227
rect -296 2193 -224 2227
rect -392 2179 -224 2193
rect -426 2177 -190 2179
rect -426 2159 -330 2177
rect -296 2159 -190 2177
rect -392 2125 -330 2159
rect -296 2125 -224 2159
rect -392 2107 -224 2125
rect -426 2105 -190 2107
rect -426 2091 -330 2105
rect -296 2091 -190 2105
rect -392 2057 -330 2091
rect -296 2057 -224 2091
rect -392 2035 -224 2057
rect -426 2033 -190 2035
rect -426 2023 -330 2033
rect -296 2023 -190 2033
rect -392 1989 -330 2023
rect -296 1989 -224 2023
rect -392 1963 -224 1989
rect -426 1961 -190 1963
rect -426 1955 -330 1961
rect -296 1955 -190 1961
rect -392 1921 -330 1955
rect -296 1921 -224 1955
rect -392 1891 -224 1921
rect -426 1889 -190 1891
rect -426 1887 -330 1889
rect -296 1887 -190 1889
rect -392 1853 -330 1887
rect -296 1853 -224 1887
rect -392 1819 -224 1853
rect -392 1785 -330 1819
rect -296 1785 -224 1819
rect -426 1783 -330 1785
rect -296 1783 -190 1785
rect -426 1781 -190 1783
rect -392 1751 -224 1781
rect -392 1717 -330 1751
rect -296 1717 -224 1751
rect -426 1711 -330 1717
rect -296 1711 -190 1717
rect -426 1709 -190 1711
rect -392 1683 -224 1709
rect -392 1649 -330 1683
rect -296 1649 -224 1683
rect -426 1639 -330 1649
rect -296 1639 -190 1649
rect -426 1637 -190 1639
rect -392 1615 -224 1637
rect -392 1581 -330 1615
rect -296 1581 -224 1615
rect -426 1567 -330 1581
rect -296 1567 -190 1581
rect -426 1565 -190 1567
rect -392 1547 -224 1565
rect -392 1513 -330 1547
rect -296 1513 -224 1547
rect -426 1495 -330 1513
rect -296 1495 -190 1513
rect -426 1493 -190 1495
rect -392 1479 -224 1493
rect -392 1445 -330 1479
rect -296 1445 -224 1479
rect -426 1423 -330 1445
rect -296 1423 -190 1445
rect -426 1421 -190 1423
rect -392 1411 -224 1421
rect -392 1377 -330 1411
rect -296 1377 -224 1411
rect -426 1351 -330 1377
rect -296 1351 -190 1377
rect -426 1349 -190 1351
rect -392 1343 -224 1349
rect -392 1309 -330 1343
rect -296 1309 -224 1343
rect -426 1279 -330 1309
rect -296 1279 -190 1309
rect -426 1277 -190 1279
rect -392 1275 -224 1277
rect -392 1241 -330 1275
rect -296 1241 -224 1275
rect -426 1207 -330 1241
rect -296 1207 -190 1241
rect -392 1173 -330 1207
rect -296 1173 -224 1207
rect -392 1171 -224 1173
rect -426 1169 -190 1171
rect -426 1139 -330 1169
rect -296 1139 -190 1169
rect -392 1105 -330 1139
rect -296 1105 -224 1139
rect -392 1099 -224 1105
rect -426 1097 -190 1099
rect -426 1071 -330 1097
rect -296 1071 -190 1097
rect -392 1037 -330 1071
rect -296 1037 -224 1071
rect -392 1027 -224 1037
rect -426 1025 -190 1027
rect -426 1003 -330 1025
rect -296 1003 -190 1025
rect -392 969 -330 1003
rect -296 969 -224 1003
rect -392 955 -224 969
rect -426 953 -190 955
rect -426 935 -330 953
rect -296 935 -190 953
rect -392 901 -330 935
rect -296 901 -224 935
rect -392 883 -224 901
rect -426 881 -190 883
rect -426 867 -330 881
rect -296 867 -190 881
rect -392 833 -330 867
rect -296 833 -224 867
rect -392 811 -224 833
rect -426 809 -190 811
rect -426 799 -330 809
rect -296 799 -190 809
rect -392 765 -330 799
rect -296 765 -224 799
rect -392 739 -224 765
rect -426 737 -190 739
rect -426 731 -330 737
rect -296 731 -190 737
rect -392 697 -330 731
rect -296 697 -224 731
rect -392 667 -224 697
rect -426 665 -190 667
rect -426 663 -330 665
rect -296 663 -190 665
rect -392 629 -330 663
rect -296 629 -224 663
rect -392 595 -224 629
rect -392 561 -330 595
rect -296 561 -224 595
rect -426 559 -330 561
rect -296 559 -190 561
rect -426 557 -190 559
rect -392 527 -224 557
rect -392 493 -330 527
rect -296 493 -224 527
rect -426 487 -330 493
rect -296 487 -190 493
rect -426 485 -190 487
rect -392 459 -224 485
rect -392 425 -330 459
rect -296 425 -224 459
rect -426 415 -330 425
rect -296 415 -190 425
rect -426 413 -190 415
rect -392 391 -224 413
rect -392 357 -330 391
rect -296 357 -224 391
rect -426 343 -330 357
rect -296 343 -190 357
rect -426 341 -190 343
rect -392 323 -224 341
rect -392 289 -330 323
rect -296 289 -224 323
rect -426 271 -330 289
rect -296 271 -190 289
rect -426 269 -190 271
rect -392 255 -224 269
rect -392 221 -330 255
rect -296 221 -224 255
rect -426 199 -330 221
rect -296 199 -190 221
rect -426 197 -190 199
rect -392 187 -224 197
rect -392 153 -330 187
rect -296 153 -224 187
rect -426 127 -330 153
rect -296 127 -190 153
rect -426 125 -190 127
rect -392 119 -224 125
rect -392 85 -330 119
rect -296 85 -224 119
rect -426 55 -330 85
rect -296 55 -190 85
rect -426 53 -190 55
rect -392 51 -224 53
rect -392 17 -330 51
rect -296 17 -224 51
rect -426 -17 -330 17
rect -296 -17 -190 17
rect -392 -51 -330 -17
rect -296 -51 -224 -17
rect -392 -53 -224 -51
rect -426 -55 -190 -53
rect -426 -85 -330 -55
rect -296 -85 -190 -55
rect -392 -119 -330 -85
rect -296 -119 -224 -85
rect -392 -125 -224 -119
rect -426 -127 -190 -125
rect -426 -153 -330 -127
rect -296 -153 -190 -127
rect -392 -187 -330 -153
rect -296 -187 -224 -153
rect -392 -197 -224 -187
rect -426 -199 -190 -197
rect -426 -221 -330 -199
rect -296 -221 -190 -199
rect -392 -255 -330 -221
rect -296 -255 -224 -221
rect -392 -269 -224 -255
rect -426 -271 -190 -269
rect -426 -289 -330 -271
rect -296 -289 -190 -271
rect -392 -323 -330 -289
rect -296 -323 -224 -289
rect -392 -341 -224 -323
rect -426 -343 -190 -341
rect -426 -357 -330 -343
rect -296 -357 -190 -343
rect -392 -391 -330 -357
rect -296 -391 -224 -357
rect -392 -413 -224 -391
rect -426 -415 -190 -413
rect -426 -425 -330 -415
rect -296 -425 -190 -415
rect -392 -459 -330 -425
rect -296 -459 -224 -425
rect -392 -485 -224 -459
rect -426 -487 -190 -485
rect -426 -493 -330 -487
rect -296 -493 -190 -487
rect -392 -527 -330 -493
rect -296 -527 -224 -493
rect -392 -557 -224 -527
rect -426 -559 -190 -557
rect -426 -561 -330 -559
rect -296 -561 -190 -559
rect -392 -595 -330 -561
rect -296 -595 -224 -561
rect -392 -629 -224 -595
rect -392 -663 -330 -629
rect -296 -663 -224 -629
rect -426 -665 -330 -663
rect -296 -665 -190 -663
rect -426 -667 -190 -665
rect -392 -697 -224 -667
rect -392 -731 -330 -697
rect -296 -731 -224 -697
rect -426 -737 -330 -731
rect -296 -737 -190 -731
rect -426 -739 -190 -737
rect -392 -765 -224 -739
rect -392 -799 -330 -765
rect -296 -799 -224 -765
rect -426 -809 -330 -799
rect -296 -809 -190 -799
rect -426 -811 -190 -809
rect -392 -833 -224 -811
rect -392 -867 -330 -833
rect -296 -867 -224 -833
rect -426 -881 -330 -867
rect -296 -881 -190 -867
rect -426 -883 -190 -881
rect -392 -901 -224 -883
rect -392 -935 -330 -901
rect -296 -935 -224 -901
rect -426 -953 -330 -935
rect -296 -953 -190 -935
rect -426 -955 -190 -953
rect -392 -969 -224 -955
rect -392 -1003 -330 -969
rect -296 -1003 -224 -969
rect -426 -1025 -330 -1003
rect -296 -1025 -190 -1003
rect -426 -1027 -190 -1025
rect -392 -1037 -224 -1027
rect -392 -1071 -330 -1037
rect -296 -1071 -224 -1037
rect -426 -1097 -330 -1071
rect -296 -1097 -190 -1071
rect -426 -1099 -190 -1097
rect -392 -1105 -224 -1099
rect -392 -1139 -330 -1105
rect -296 -1139 -224 -1105
rect -426 -1169 -330 -1139
rect -296 -1169 -190 -1139
rect -426 -1171 -190 -1169
rect -392 -1173 -224 -1171
rect -392 -1207 -330 -1173
rect -296 -1207 -224 -1173
rect -426 -1241 -330 -1207
rect -296 -1241 -190 -1207
rect -392 -1275 -330 -1241
rect -296 -1275 -224 -1241
rect -392 -1277 -224 -1275
rect -426 -1279 -190 -1277
rect -426 -1309 -330 -1279
rect -296 -1309 -190 -1279
rect -392 -1343 -330 -1309
rect -296 -1343 -224 -1309
rect -392 -1349 -224 -1343
rect -426 -1351 -190 -1349
rect -426 -1377 -330 -1351
rect -296 -1377 -190 -1351
rect -392 -1411 -330 -1377
rect -296 -1411 -224 -1377
rect -392 -1421 -224 -1411
rect -426 -1423 -190 -1421
rect -426 -1445 -330 -1423
rect -296 -1445 -190 -1423
rect -392 -1479 -330 -1445
rect -296 -1479 -224 -1445
rect -392 -1493 -224 -1479
rect -426 -1495 -190 -1493
rect -426 -1513 -330 -1495
rect -296 -1513 -190 -1495
rect -392 -1547 -330 -1513
rect -296 -1547 -224 -1513
rect -392 -1565 -224 -1547
rect -426 -1567 -190 -1565
rect -426 -1581 -330 -1567
rect -296 -1581 -190 -1567
rect -392 -1615 -330 -1581
rect -296 -1615 -224 -1581
rect -392 -1637 -224 -1615
rect -426 -1639 -190 -1637
rect -426 -1649 -330 -1639
rect -296 -1649 -190 -1639
rect -392 -1683 -330 -1649
rect -296 -1683 -224 -1649
rect -392 -1709 -224 -1683
rect -426 -1711 -190 -1709
rect -426 -1717 -330 -1711
rect -296 -1717 -190 -1711
rect -392 -1751 -330 -1717
rect -296 -1751 -224 -1717
rect -392 -1781 -224 -1751
rect -426 -1783 -190 -1781
rect -426 -1785 -330 -1783
rect -296 -1785 -190 -1783
rect -392 -1819 -330 -1785
rect -296 -1819 -224 -1785
rect -392 -1853 -224 -1819
rect -392 -1887 -330 -1853
rect -296 -1887 -224 -1853
rect -426 -1889 -330 -1887
rect -296 -1889 -190 -1887
rect -426 -1891 -190 -1889
rect -392 -1921 -224 -1891
rect -392 -1955 -330 -1921
rect -296 -1955 -224 -1921
rect -426 -1961 -330 -1955
rect -296 -1961 -190 -1955
rect -426 -1963 -190 -1961
rect -392 -1989 -224 -1963
rect -392 -2023 -330 -1989
rect -296 -2023 -224 -1989
rect -426 -2033 -330 -2023
rect -296 -2033 -190 -2023
rect -426 -2035 -190 -2033
rect -392 -2057 -224 -2035
rect -392 -2091 -330 -2057
rect -296 -2091 -224 -2057
rect -426 -2105 -330 -2091
rect -296 -2105 -190 -2091
rect -426 -2107 -190 -2105
rect -392 -2125 -224 -2107
rect -392 -2159 -330 -2125
rect -296 -2159 -224 -2125
rect -426 -2177 -330 -2159
rect -296 -2177 -190 -2159
rect -426 -2179 -190 -2177
rect -392 -2193 -224 -2179
rect -392 -2227 -330 -2193
rect -296 -2227 -224 -2193
rect -426 -2249 -330 -2227
rect -296 -2249 -190 -2227
rect -426 -2251 -190 -2249
rect -392 -2261 -224 -2251
rect -392 -2295 -330 -2261
rect -296 -2295 -224 -2261
rect -426 -2321 -330 -2295
rect -296 -2321 -190 -2295
rect -426 -2323 -190 -2321
rect -392 -2329 -224 -2323
rect -392 -2363 -330 -2329
rect -296 -2363 -224 -2329
rect -426 -2393 -330 -2363
rect -296 -2393 -190 -2363
rect -426 -2395 -190 -2393
rect -392 -2397 -224 -2395
rect -392 -2431 -330 -2397
rect -296 -2431 -224 -2397
rect -426 -2465 -330 -2431
rect -296 -2465 -190 -2431
rect -392 -2499 -330 -2465
rect -296 -2499 -224 -2465
rect -392 -2501 -224 -2499
rect -426 -2503 -190 -2501
rect -426 -2533 -330 -2503
rect -296 -2533 -190 -2503
rect -392 -2567 -330 -2533
rect -296 -2567 -224 -2533
rect -392 -2573 -224 -2567
rect -426 -2575 -190 -2573
rect -426 -2601 -330 -2575
rect -296 -2601 -190 -2575
rect -392 -2635 -330 -2601
rect -296 -2635 -224 -2601
rect -392 -2645 -224 -2635
rect -426 -2647 -190 -2645
rect -426 -2669 -330 -2647
rect -296 -2669 -190 -2647
rect -392 -2703 -330 -2669
rect -296 -2703 -224 -2669
rect -392 -2717 -224 -2703
rect -426 -2719 -190 -2717
rect -426 -2737 -330 -2719
rect -296 -2737 -190 -2719
rect -392 -2771 -330 -2737
rect -296 -2771 -224 -2737
rect -392 -2789 -224 -2771
rect -426 -2791 -190 -2789
rect -426 -2805 -330 -2791
rect -296 -2805 -190 -2791
rect -392 -2839 -330 -2805
rect -296 -2839 -224 -2805
rect -392 -2861 -224 -2839
rect -426 -2863 -190 -2861
rect -426 -2873 -330 -2863
rect -296 -2873 -190 -2863
rect -392 -2907 -330 -2873
rect -296 -2907 -224 -2873
rect -392 -2933 -224 -2907
rect -426 -2935 -190 -2933
rect -426 -2941 -330 -2935
rect -296 -2941 -190 -2935
rect -392 -2975 -330 -2941
rect -296 -2975 -224 -2941
rect -392 -3005 -224 -2975
rect -426 -3007 -190 -3005
rect -426 -3009 -330 -3007
rect -296 -3009 -190 -3007
rect -392 -3043 -330 -3009
rect -296 -3043 -224 -3009
rect -392 -3077 -224 -3043
rect -392 -3111 -330 -3077
rect -296 -3111 -224 -3077
rect -426 -3113 -330 -3111
rect -296 -3113 -190 -3111
rect -426 -3115 -190 -3113
rect -392 -3145 -224 -3115
rect -392 -3179 -330 -3145
rect -296 -3179 -224 -3145
rect -426 -3185 -330 -3179
rect -296 -3185 -190 -3179
rect -426 -3187 -190 -3185
rect -392 -3213 -224 -3187
rect -392 -3247 -330 -3213
rect -296 -3247 -224 -3213
rect -426 -3257 -330 -3247
rect -296 -3257 -190 -3247
rect -426 -3259 -190 -3257
rect -392 -3281 -224 -3259
rect -392 -3315 -330 -3281
rect -296 -3315 -224 -3281
rect -426 -3329 -330 -3315
rect -296 -3329 -190 -3315
rect -426 -3331 -190 -3329
rect -392 -3349 -224 -3331
rect -392 -3383 -330 -3349
rect -296 -3383 -224 -3349
rect -426 -3401 -330 -3383
rect -296 -3401 -190 -3383
rect -426 -3403 -190 -3401
rect -392 -3417 -224 -3403
rect -392 -3451 -330 -3417
rect -296 -3451 -224 -3417
rect -426 -3473 -330 -3451
rect -296 -3473 -190 -3451
rect -426 -3475 -190 -3473
rect -392 -3485 -224 -3475
rect -392 -3519 -330 -3485
rect -296 -3519 -224 -3485
rect -426 -3545 -330 -3519
rect -296 -3545 -190 -3519
rect -426 -3547 -190 -3545
rect -392 -3553 -224 -3547
rect -392 -3587 -330 -3553
rect -296 -3587 -224 -3553
rect -426 -3617 -330 -3587
rect -296 -3617 -190 -3587
rect -426 -3619 -190 -3617
rect -392 -3621 -224 -3619
rect -392 -3655 -330 -3621
rect -296 -3655 -224 -3621
rect -426 -3689 -330 -3655
rect -296 -3689 -190 -3655
rect -392 -3723 -330 -3689
rect -296 -3723 -224 -3689
rect -392 -3725 -224 -3723
rect -426 -3727 -190 -3725
rect -426 -3757 -330 -3727
rect -296 -3757 -190 -3727
rect -392 -3791 -330 -3757
rect -296 -3791 -224 -3757
rect -392 -3797 -224 -3791
rect -426 -3799 -190 -3797
rect -426 -3825 -330 -3799
rect -296 -3825 -190 -3799
rect -392 -3859 -330 -3825
rect -296 -3859 -224 -3825
rect -392 -3869 -224 -3859
rect -426 -3871 -190 -3869
rect -426 -3893 -330 -3871
rect -296 -3893 -190 -3871
rect -392 -3927 -330 -3893
rect -296 -3927 -224 -3893
rect -392 -3941 -224 -3927
rect -426 -3943 -190 -3941
rect -426 -3961 -330 -3943
rect -296 -3961 -190 -3943
rect -392 -3995 -330 -3961
rect -296 -3995 -224 -3961
rect -392 -4013 -224 -3995
rect -426 -4015 -190 -4013
rect -426 -4029 -330 -4015
rect -296 -4029 -190 -4015
rect -392 -4063 -330 -4029
rect -296 -4063 -224 -4029
rect -392 -4085 -224 -4063
rect -426 -4087 -190 -4085
rect -426 -4097 -330 -4087
rect -296 -4097 -190 -4087
rect -392 -4131 -330 -4097
rect -296 -4131 -224 -4097
rect -392 -4157 -224 -4131
rect -426 -4159 -190 -4157
rect -426 -4165 -330 -4159
rect -296 -4165 -190 -4159
rect -392 -4199 -330 -4165
rect -296 -4199 -224 -4165
rect -392 -4229 -224 -4199
rect -426 -4231 -190 -4229
rect -426 -4233 -330 -4231
rect -296 -4233 -190 -4231
rect -392 -4267 -330 -4233
rect -296 -4267 -224 -4233
rect -392 -4301 -224 -4267
rect -392 -4335 -330 -4301
rect -296 -4335 -224 -4301
rect -426 -4337 -330 -4335
rect -296 -4337 -190 -4335
rect -426 -4339 -190 -4337
rect -392 -4369 -224 -4339
rect -392 -4403 -330 -4369
rect -296 -4403 -224 -4369
rect -426 -4409 -330 -4403
rect -296 -4409 -190 -4403
rect -426 -4411 -190 -4409
rect -392 -4437 -224 -4411
rect -392 -4471 -330 -4437
rect -296 -4471 -224 -4437
rect -426 -4481 -330 -4471
rect -296 -4481 -190 -4471
rect -426 -4483 -190 -4481
rect -392 -4505 -224 -4483
rect -392 -4539 -330 -4505
rect -296 -4539 -224 -4505
rect -426 -4553 -330 -4539
rect -296 -4553 -190 -4539
rect -426 -4555 -190 -4553
rect -392 -4573 -224 -4555
rect -392 -4607 -330 -4573
rect -296 -4607 -224 -4573
rect -426 -4625 -330 -4607
rect -296 -4625 -190 -4607
rect -426 -4627 -190 -4625
rect -392 -4641 -224 -4627
rect -392 -4675 -330 -4641
rect -296 -4675 -224 -4641
rect -426 -4697 -330 -4675
rect -296 -4697 -190 -4675
rect -426 -4699 -190 -4697
rect -392 -4709 -224 -4699
rect -392 -4743 -330 -4709
rect -296 -4743 -224 -4709
rect -426 -4769 -330 -4743
rect -296 -4769 -190 -4743
rect -426 -4771 -190 -4769
rect -392 -4777 -224 -4771
rect -392 -4811 -330 -4777
rect -296 -4811 -224 -4777
rect -426 -4841 -330 -4811
rect -296 -4841 -190 -4811
rect -426 -4843 -190 -4841
rect -392 -4845 -224 -4843
rect -392 -4879 -330 -4845
rect -296 -4879 -224 -4845
rect -426 -4913 -330 -4879
rect -296 -4913 -190 -4879
rect -392 -4947 -330 -4913
rect -296 -4947 -224 -4913
rect -392 -4949 -224 -4947
rect -426 -4951 -190 -4949
rect -426 -4981 -330 -4951
rect -296 -4981 -190 -4951
rect -1008 -5021 -840 -5015
rect -1042 -5023 -806 -5021
rect -1042 -5057 -946 -5023
rect -912 -5057 -806 -5023
rect -1042 -5090 -806 -5057
rect -392 -5015 -330 -4981
rect -296 -5015 -224 -4981
rect -88 4985 88 5004
rect -88 4981 -53 4985
rect 53 4981 88 4985
rect -88 -4981 -85 4981
rect 85 -4981 88 4981
rect -88 -4985 -53 -4981
rect 53 -4985 88 -4981
rect -88 -5004 88 -4985
rect 224 4981 286 5015
rect 320 4981 392 5015
rect 806 5057 1042 5090
rect 806 5023 902 5057
rect 936 5023 1042 5057
rect 806 5021 1042 5023
rect 840 5015 1008 5021
rect 190 4951 286 4981
rect 320 4951 426 4981
rect 190 4949 426 4951
rect 224 4947 392 4949
rect 224 4913 286 4947
rect 320 4913 392 4947
rect 190 4879 286 4913
rect 320 4879 426 4913
rect 224 4845 286 4879
rect 320 4845 392 4879
rect 224 4843 392 4845
rect 190 4841 426 4843
rect 190 4811 286 4841
rect 320 4811 426 4841
rect 224 4777 286 4811
rect 320 4777 392 4811
rect 224 4771 392 4777
rect 190 4769 426 4771
rect 190 4743 286 4769
rect 320 4743 426 4769
rect 224 4709 286 4743
rect 320 4709 392 4743
rect 224 4699 392 4709
rect 190 4697 426 4699
rect 190 4675 286 4697
rect 320 4675 426 4697
rect 224 4641 286 4675
rect 320 4641 392 4675
rect 224 4627 392 4641
rect 190 4625 426 4627
rect 190 4607 286 4625
rect 320 4607 426 4625
rect 224 4573 286 4607
rect 320 4573 392 4607
rect 224 4555 392 4573
rect 190 4553 426 4555
rect 190 4539 286 4553
rect 320 4539 426 4553
rect 224 4505 286 4539
rect 320 4505 392 4539
rect 224 4483 392 4505
rect 190 4481 426 4483
rect 190 4471 286 4481
rect 320 4471 426 4481
rect 224 4437 286 4471
rect 320 4437 392 4471
rect 224 4411 392 4437
rect 190 4409 426 4411
rect 190 4403 286 4409
rect 320 4403 426 4409
rect 224 4369 286 4403
rect 320 4369 392 4403
rect 224 4339 392 4369
rect 190 4337 426 4339
rect 190 4335 286 4337
rect 320 4335 426 4337
rect 224 4301 286 4335
rect 320 4301 392 4335
rect 224 4267 392 4301
rect 224 4233 286 4267
rect 320 4233 392 4267
rect 190 4231 286 4233
rect 320 4231 426 4233
rect 190 4229 426 4231
rect 224 4199 392 4229
rect 224 4165 286 4199
rect 320 4165 392 4199
rect 190 4159 286 4165
rect 320 4159 426 4165
rect 190 4157 426 4159
rect 224 4131 392 4157
rect 224 4097 286 4131
rect 320 4097 392 4131
rect 190 4087 286 4097
rect 320 4087 426 4097
rect 190 4085 426 4087
rect 224 4063 392 4085
rect 224 4029 286 4063
rect 320 4029 392 4063
rect 190 4015 286 4029
rect 320 4015 426 4029
rect 190 4013 426 4015
rect 224 3995 392 4013
rect 224 3961 286 3995
rect 320 3961 392 3995
rect 190 3943 286 3961
rect 320 3943 426 3961
rect 190 3941 426 3943
rect 224 3927 392 3941
rect 224 3893 286 3927
rect 320 3893 392 3927
rect 190 3871 286 3893
rect 320 3871 426 3893
rect 190 3869 426 3871
rect 224 3859 392 3869
rect 224 3825 286 3859
rect 320 3825 392 3859
rect 190 3799 286 3825
rect 320 3799 426 3825
rect 190 3797 426 3799
rect 224 3791 392 3797
rect 224 3757 286 3791
rect 320 3757 392 3791
rect 190 3727 286 3757
rect 320 3727 426 3757
rect 190 3725 426 3727
rect 224 3723 392 3725
rect 224 3689 286 3723
rect 320 3689 392 3723
rect 190 3655 286 3689
rect 320 3655 426 3689
rect 224 3621 286 3655
rect 320 3621 392 3655
rect 224 3619 392 3621
rect 190 3617 426 3619
rect 190 3587 286 3617
rect 320 3587 426 3617
rect 224 3553 286 3587
rect 320 3553 392 3587
rect 224 3547 392 3553
rect 190 3545 426 3547
rect 190 3519 286 3545
rect 320 3519 426 3545
rect 224 3485 286 3519
rect 320 3485 392 3519
rect 224 3475 392 3485
rect 190 3473 426 3475
rect 190 3451 286 3473
rect 320 3451 426 3473
rect 224 3417 286 3451
rect 320 3417 392 3451
rect 224 3403 392 3417
rect 190 3401 426 3403
rect 190 3383 286 3401
rect 320 3383 426 3401
rect 224 3349 286 3383
rect 320 3349 392 3383
rect 224 3331 392 3349
rect 190 3329 426 3331
rect 190 3315 286 3329
rect 320 3315 426 3329
rect 224 3281 286 3315
rect 320 3281 392 3315
rect 224 3259 392 3281
rect 190 3257 426 3259
rect 190 3247 286 3257
rect 320 3247 426 3257
rect 224 3213 286 3247
rect 320 3213 392 3247
rect 224 3187 392 3213
rect 190 3185 426 3187
rect 190 3179 286 3185
rect 320 3179 426 3185
rect 224 3145 286 3179
rect 320 3145 392 3179
rect 224 3115 392 3145
rect 190 3113 426 3115
rect 190 3111 286 3113
rect 320 3111 426 3113
rect 224 3077 286 3111
rect 320 3077 392 3111
rect 224 3043 392 3077
rect 224 3009 286 3043
rect 320 3009 392 3043
rect 190 3007 286 3009
rect 320 3007 426 3009
rect 190 3005 426 3007
rect 224 2975 392 3005
rect 224 2941 286 2975
rect 320 2941 392 2975
rect 190 2935 286 2941
rect 320 2935 426 2941
rect 190 2933 426 2935
rect 224 2907 392 2933
rect 224 2873 286 2907
rect 320 2873 392 2907
rect 190 2863 286 2873
rect 320 2863 426 2873
rect 190 2861 426 2863
rect 224 2839 392 2861
rect 224 2805 286 2839
rect 320 2805 392 2839
rect 190 2791 286 2805
rect 320 2791 426 2805
rect 190 2789 426 2791
rect 224 2771 392 2789
rect 224 2737 286 2771
rect 320 2737 392 2771
rect 190 2719 286 2737
rect 320 2719 426 2737
rect 190 2717 426 2719
rect 224 2703 392 2717
rect 224 2669 286 2703
rect 320 2669 392 2703
rect 190 2647 286 2669
rect 320 2647 426 2669
rect 190 2645 426 2647
rect 224 2635 392 2645
rect 224 2601 286 2635
rect 320 2601 392 2635
rect 190 2575 286 2601
rect 320 2575 426 2601
rect 190 2573 426 2575
rect 224 2567 392 2573
rect 224 2533 286 2567
rect 320 2533 392 2567
rect 190 2503 286 2533
rect 320 2503 426 2533
rect 190 2501 426 2503
rect 224 2499 392 2501
rect 224 2465 286 2499
rect 320 2465 392 2499
rect 190 2431 286 2465
rect 320 2431 426 2465
rect 224 2397 286 2431
rect 320 2397 392 2431
rect 224 2395 392 2397
rect 190 2393 426 2395
rect 190 2363 286 2393
rect 320 2363 426 2393
rect 224 2329 286 2363
rect 320 2329 392 2363
rect 224 2323 392 2329
rect 190 2321 426 2323
rect 190 2295 286 2321
rect 320 2295 426 2321
rect 224 2261 286 2295
rect 320 2261 392 2295
rect 224 2251 392 2261
rect 190 2249 426 2251
rect 190 2227 286 2249
rect 320 2227 426 2249
rect 224 2193 286 2227
rect 320 2193 392 2227
rect 224 2179 392 2193
rect 190 2177 426 2179
rect 190 2159 286 2177
rect 320 2159 426 2177
rect 224 2125 286 2159
rect 320 2125 392 2159
rect 224 2107 392 2125
rect 190 2105 426 2107
rect 190 2091 286 2105
rect 320 2091 426 2105
rect 224 2057 286 2091
rect 320 2057 392 2091
rect 224 2035 392 2057
rect 190 2033 426 2035
rect 190 2023 286 2033
rect 320 2023 426 2033
rect 224 1989 286 2023
rect 320 1989 392 2023
rect 224 1963 392 1989
rect 190 1961 426 1963
rect 190 1955 286 1961
rect 320 1955 426 1961
rect 224 1921 286 1955
rect 320 1921 392 1955
rect 224 1891 392 1921
rect 190 1889 426 1891
rect 190 1887 286 1889
rect 320 1887 426 1889
rect 224 1853 286 1887
rect 320 1853 392 1887
rect 224 1819 392 1853
rect 224 1785 286 1819
rect 320 1785 392 1819
rect 190 1783 286 1785
rect 320 1783 426 1785
rect 190 1781 426 1783
rect 224 1751 392 1781
rect 224 1717 286 1751
rect 320 1717 392 1751
rect 190 1711 286 1717
rect 320 1711 426 1717
rect 190 1709 426 1711
rect 224 1683 392 1709
rect 224 1649 286 1683
rect 320 1649 392 1683
rect 190 1639 286 1649
rect 320 1639 426 1649
rect 190 1637 426 1639
rect 224 1615 392 1637
rect 224 1581 286 1615
rect 320 1581 392 1615
rect 190 1567 286 1581
rect 320 1567 426 1581
rect 190 1565 426 1567
rect 224 1547 392 1565
rect 224 1513 286 1547
rect 320 1513 392 1547
rect 190 1495 286 1513
rect 320 1495 426 1513
rect 190 1493 426 1495
rect 224 1479 392 1493
rect 224 1445 286 1479
rect 320 1445 392 1479
rect 190 1423 286 1445
rect 320 1423 426 1445
rect 190 1421 426 1423
rect 224 1411 392 1421
rect 224 1377 286 1411
rect 320 1377 392 1411
rect 190 1351 286 1377
rect 320 1351 426 1377
rect 190 1349 426 1351
rect 224 1343 392 1349
rect 224 1309 286 1343
rect 320 1309 392 1343
rect 190 1279 286 1309
rect 320 1279 426 1309
rect 190 1277 426 1279
rect 224 1275 392 1277
rect 224 1241 286 1275
rect 320 1241 392 1275
rect 190 1207 286 1241
rect 320 1207 426 1241
rect 224 1173 286 1207
rect 320 1173 392 1207
rect 224 1171 392 1173
rect 190 1169 426 1171
rect 190 1139 286 1169
rect 320 1139 426 1169
rect 224 1105 286 1139
rect 320 1105 392 1139
rect 224 1099 392 1105
rect 190 1097 426 1099
rect 190 1071 286 1097
rect 320 1071 426 1097
rect 224 1037 286 1071
rect 320 1037 392 1071
rect 224 1027 392 1037
rect 190 1025 426 1027
rect 190 1003 286 1025
rect 320 1003 426 1025
rect 224 969 286 1003
rect 320 969 392 1003
rect 224 955 392 969
rect 190 953 426 955
rect 190 935 286 953
rect 320 935 426 953
rect 224 901 286 935
rect 320 901 392 935
rect 224 883 392 901
rect 190 881 426 883
rect 190 867 286 881
rect 320 867 426 881
rect 224 833 286 867
rect 320 833 392 867
rect 224 811 392 833
rect 190 809 426 811
rect 190 799 286 809
rect 320 799 426 809
rect 224 765 286 799
rect 320 765 392 799
rect 224 739 392 765
rect 190 737 426 739
rect 190 731 286 737
rect 320 731 426 737
rect 224 697 286 731
rect 320 697 392 731
rect 224 667 392 697
rect 190 665 426 667
rect 190 663 286 665
rect 320 663 426 665
rect 224 629 286 663
rect 320 629 392 663
rect 224 595 392 629
rect 224 561 286 595
rect 320 561 392 595
rect 190 559 286 561
rect 320 559 426 561
rect 190 557 426 559
rect 224 527 392 557
rect 224 493 286 527
rect 320 493 392 527
rect 190 487 286 493
rect 320 487 426 493
rect 190 485 426 487
rect 224 459 392 485
rect 224 425 286 459
rect 320 425 392 459
rect 190 415 286 425
rect 320 415 426 425
rect 190 413 426 415
rect 224 391 392 413
rect 224 357 286 391
rect 320 357 392 391
rect 190 343 286 357
rect 320 343 426 357
rect 190 341 426 343
rect 224 323 392 341
rect 224 289 286 323
rect 320 289 392 323
rect 190 271 286 289
rect 320 271 426 289
rect 190 269 426 271
rect 224 255 392 269
rect 224 221 286 255
rect 320 221 392 255
rect 190 199 286 221
rect 320 199 426 221
rect 190 197 426 199
rect 224 187 392 197
rect 224 153 286 187
rect 320 153 392 187
rect 190 127 286 153
rect 320 127 426 153
rect 190 125 426 127
rect 224 119 392 125
rect 224 85 286 119
rect 320 85 392 119
rect 190 55 286 85
rect 320 55 426 85
rect 190 53 426 55
rect 224 51 392 53
rect 224 17 286 51
rect 320 17 392 51
rect 190 -17 286 17
rect 320 -17 426 17
rect 224 -51 286 -17
rect 320 -51 392 -17
rect 224 -53 392 -51
rect 190 -55 426 -53
rect 190 -85 286 -55
rect 320 -85 426 -55
rect 224 -119 286 -85
rect 320 -119 392 -85
rect 224 -125 392 -119
rect 190 -127 426 -125
rect 190 -153 286 -127
rect 320 -153 426 -127
rect 224 -187 286 -153
rect 320 -187 392 -153
rect 224 -197 392 -187
rect 190 -199 426 -197
rect 190 -221 286 -199
rect 320 -221 426 -199
rect 224 -255 286 -221
rect 320 -255 392 -221
rect 224 -269 392 -255
rect 190 -271 426 -269
rect 190 -289 286 -271
rect 320 -289 426 -271
rect 224 -323 286 -289
rect 320 -323 392 -289
rect 224 -341 392 -323
rect 190 -343 426 -341
rect 190 -357 286 -343
rect 320 -357 426 -343
rect 224 -391 286 -357
rect 320 -391 392 -357
rect 224 -413 392 -391
rect 190 -415 426 -413
rect 190 -425 286 -415
rect 320 -425 426 -415
rect 224 -459 286 -425
rect 320 -459 392 -425
rect 224 -485 392 -459
rect 190 -487 426 -485
rect 190 -493 286 -487
rect 320 -493 426 -487
rect 224 -527 286 -493
rect 320 -527 392 -493
rect 224 -557 392 -527
rect 190 -559 426 -557
rect 190 -561 286 -559
rect 320 -561 426 -559
rect 224 -595 286 -561
rect 320 -595 392 -561
rect 224 -629 392 -595
rect 224 -663 286 -629
rect 320 -663 392 -629
rect 190 -665 286 -663
rect 320 -665 426 -663
rect 190 -667 426 -665
rect 224 -697 392 -667
rect 224 -731 286 -697
rect 320 -731 392 -697
rect 190 -737 286 -731
rect 320 -737 426 -731
rect 190 -739 426 -737
rect 224 -765 392 -739
rect 224 -799 286 -765
rect 320 -799 392 -765
rect 190 -809 286 -799
rect 320 -809 426 -799
rect 190 -811 426 -809
rect 224 -833 392 -811
rect 224 -867 286 -833
rect 320 -867 392 -833
rect 190 -881 286 -867
rect 320 -881 426 -867
rect 190 -883 426 -881
rect 224 -901 392 -883
rect 224 -935 286 -901
rect 320 -935 392 -901
rect 190 -953 286 -935
rect 320 -953 426 -935
rect 190 -955 426 -953
rect 224 -969 392 -955
rect 224 -1003 286 -969
rect 320 -1003 392 -969
rect 190 -1025 286 -1003
rect 320 -1025 426 -1003
rect 190 -1027 426 -1025
rect 224 -1037 392 -1027
rect 224 -1071 286 -1037
rect 320 -1071 392 -1037
rect 190 -1097 286 -1071
rect 320 -1097 426 -1071
rect 190 -1099 426 -1097
rect 224 -1105 392 -1099
rect 224 -1139 286 -1105
rect 320 -1139 392 -1105
rect 190 -1169 286 -1139
rect 320 -1169 426 -1139
rect 190 -1171 426 -1169
rect 224 -1173 392 -1171
rect 224 -1207 286 -1173
rect 320 -1207 392 -1173
rect 190 -1241 286 -1207
rect 320 -1241 426 -1207
rect 224 -1275 286 -1241
rect 320 -1275 392 -1241
rect 224 -1277 392 -1275
rect 190 -1279 426 -1277
rect 190 -1309 286 -1279
rect 320 -1309 426 -1279
rect 224 -1343 286 -1309
rect 320 -1343 392 -1309
rect 224 -1349 392 -1343
rect 190 -1351 426 -1349
rect 190 -1377 286 -1351
rect 320 -1377 426 -1351
rect 224 -1411 286 -1377
rect 320 -1411 392 -1377
rect 224 -1421 392 -1411
rect 190 -1423 426 -1421
rect 190 -1445 286 -1423
rect 320 -1445 426 -1423
rect 224 -1479 286 -1445
rect 320 -1479 392 -1445
rect 224 -1493 392 -1479
rect 190 -1495 426 -1493
rect 190 -1513 286 -1495
rect 320 -1513 426 -1495
rect 224 -1547 286 -1513
rect 320 -1547 392 -1513
rect 224 -1565 392 -1547
rect 190 -1567 426 -1565
rect 190 -1581 286 -1567
rect 320 -1581 426 -1567
rect 224 -1615 286 -1581
rect 320 -1615 392 -1581
rect 224 -1637 392 -1615
rect 190 -1639 426 -1637
rect 190 -1649 286 -1639
rect 320 -1649 426 -1639
rect 224 -1683 286 -1649
rect 320 -1683 392 -1649
rect 224 -1709 392 -1683
rect 190 -1711 426 -1709
rect 190 -1717 286 -1711
rect 320 -1717 426 -1711
rect 224 -1751 286 -1717
rect 320 -1751 392 -1717
rect 224 -1781 392 -1751
rect 190 -1783 426 -1781
rect 190 -1785 286 -1783
rect 320 -1785 426 -1783
rect 224 -1819 286 -1785
rect 320 -1819 392 -1785
rect 224 -1853 392 -1819
rect 224 -1887 286 -1853
rect 320 -1887 392 -1853
rect 190 -1889 286 -1887
rect 320 -1889 426 -1887
rect 190 -1891 426 -1889
rect 224 -1921 392 -1891
rect 224 -1955 286 -1921
rect 320 -1955 392 -1921
rect 190 -1961 286 -1955
rect 320 -1961 426 -1955
rect 190 -1963 426 -1961
rect 224 -1989 392 -1963
rect 224 -2023 286 -1989
rect 320 -2023 392 -1989
rect 190 -2033 286 -2023
rect 320 -2033 426 -2023
rect 190 -2035 426 -2033
rect 224 -2057 392 -2035
rect 224 -2091 286 -2057
rect 320 -2091 392 -2057
rect 190 -2105 286 -2091
rect 320 -2105 426 -2091
rect 190 -2107 426 -2105
rect 224 -2125 392 -2107
rect 224 -2159 286 -2125
rect 320 -2159 392 -2125
rect 190 -2177 286 -2159
rect 320 -2177 426 -2159
rect 190 -2179 426 -2177
rect 224 -2193 392 -2179
rect 224 -2227 286 -2193
rect 320 -2227 392 -2193
rect 190 -2249 286 -2227
rect 320 -2249 426 -2227
rect 190 -2251 426 -2249
rect 224 -2261 392 -2251
rect 224 -2295 286 -2261
rect 320 -2295 392 -2261
rect 190 -2321 286 -2295
rect 320 -2321 426 -2295
rect 190 -2323 426 -2321
rect 224 -2329 392 -2323
rect 224 -2363 286 -2329
rect 320 -2363 392 -2329
rect 190 -2393 286 -2363
rect 320 -2393 426 -2363
rect 190 -2395 426 -2393
rect 224 -2397 392 -2395
rect 224 -2431 286 -2397
rect 320 -2431 392 -2397
rect 190 -2465 286 -2431
rect 320 -2465 426 -2431
rect 224 -2499 286 -2465
rect 320 -2499 392 -2465
rect 224 -2501 392 -2499
rect 190 -2503 426 -2501
rect 190 -2533 286 -2503
rect 320 -2533 426 -2503
rect 224 -2567 286 -2533
rect 320 -2567 392 -2533
rect 224 -2573 392 -2567
rect 190 -2575 426 -2573
rect 190 -2601 286 -2575
rect 320 -2601 426 -2575
rect 224 -2635 286 -2601
rect 320 -2635 392 -2601
rect 224 -2645 392 -2635
rect 190 -2647 426 -2645
rect 190 -2669 286 -2647
rect 320 -2669 426 -2647
rect 224 -2703 286 -2669
rect 320 -2703 392 -2669
rect 224 -2717 392 -2703
rect 190 -2719 426 -2717
rect 190 -2737 286 -2719
rect 320 -2737 426 -2719
rect 224 -2771 286 -2737
rect 320 -2771 392 -2737
rect 224 -2789 392 -2771
rect 190 -2791 426 -2789
rect 190 -2805 286 -2791
rect 320 -2805 426 -2791
rect 224 -2839 286 -2805
rect 320 -2839 392 -2805
rect 224 -2861 392 -2839
rect 190 -2863 426 -2861
rect 190 -2873 286 -2863
rect 320 -2873 426 -2863
rect 224 -2907 286 -2873
rect 320 -2907 392 -2873
rect 224 -2933 392 -2907
rect 190 -2935 426 -2933
rect 190 -2941 286 -2935
rect 320 -2941 426 -2935
rect 224 -2975 286 -2941
rect 320 -2975 392 -2941
rect 224 -3005 392 -2975
rect 190 -3007 426 -3005
rect 190 -3009 286 -3007
rect 320 -3009 426 -3007
rect 224 -3043 286 -3009
rect 320 -3043 392 -3009
rect 224 -3077 392 -3043
rect 224 -3111 286 -3077
rect 320 -3111 392 -3077
rect 190 -3113 286 -3111
rect 320 -3113 426 -3111
rect 190 -3115 426 -3113
rect 224 -3145 392 -3115
rect 224 -3179 286 -3145
rect 320 -3179 392 -3145
rect 190 -3185 286 -3179
rect 320 -3185 426 -3179
rect 190 -3187 426 -3185
rect 224 -3213 392 -3187
rect 224 -3247 286 -3213
rect 320 -3247 392 -3213
rect 190 -3257 286 -3247
rect 320 -3257 426 -3247
rect 190 -3259 426 -3257
rect 224 -3281 392 -3259
rect 224 -3315 286 -3281
rect 320 -3315 392 -3281
rect 190 -3329 286 -3315
rect 320 -3329 426 -3315
rect 190 -3331 426 -3329
rect 224 -3349 392 -3331
rect 224 -3383 286 -3349
rect 320 -3383 392 -3349
rect 190 -3401 286 -3383
rect 320 -3401 426 -3383
rect 190 -3403 426 -3401
rect 224 -3417 392 -3403
rect 224 -3451 286 -3417
rect 320 -3451 392 -3417
rect 190 -3473 286 -3451
rect 320 -3473 426 -3451
rect 190 -3475 426 -3473
rect 224 -3485 392 -3475
rect 224 -3519 286 -3485
rect 320 -3519 392 -3485
rect 190 -3545 286 -3519
rect 320 -3545 426 -3519
rect 190 -3547 426 -3545
rect 224 -3553 392 -3547
rect 224 -3587 286 -3553
rect 320 -3587 392 -3553
rect 190 -3617 286 -3587
rect 320 -3617 426 -3587
rect 190 -3619 426 -3617
rect 224 -3621 392 -3619
rect 224 -3655 286 -3621
rect 320 -3655 392 -3621
rect 190 -3689 286 -3655
rect 320 -3689 426 -3655
rect 224 -3723 286 -3689
rect 320 -3723 392 -3689
rect 224 -3725 392 -3723
rect 190 -3727 426 -3725
rect 190 -3757 286 -3727
rect 320 -3757 426 -3727
rect 224 -3791 286 -3757
rect 320 -3791 392 -3757
rect 224 -3797 392 -3791
rect 190 -3799 426 -3797
rect 190 -3825 286 -3799
rect 320 -3825 426 -3799
rect 224 -3859 286 -3825
rect 320 -3859 392 -3825
rect 224 -3869 392 -3859
rect 190 -3871 426 -3869
rect 190 -3893 286 -3871
rect 320 -3893 426 -3871
rect 224 -3927 286 -3893
rect 320 -3927 392 -3893
rect 224 -3941 392 -3927
rect 190 -3943 426 -3941
rect 190 -3961 286 -3943
rect 320 -3961 426 -3943
rect 224 -3995 286 -3961
rect 320 -3995 392 -3961
rect 224 -4013 392 -3995
rect 190 -4015 426 -4013
rect 190 -4029 286 -4015
rect 320 -4029 426 -4015
rect 224 -4063 286 -4029
rect 320 -4063 392 -4029
rect 224 -4085 392 -4063
rect 190 -4087 426 -4085
rect 190 -4097 286 -4087
rect 320 -4097 426 -4087
rect 224 -4131 286 -4097
rect 320 -4131 392 -4097
rect 224 -4157 392 -4131
rect 190 -4159 426 -4157
rect 190 -4165 286 -4159
rect 320 -4165 426 -4159
rect 224 -4199 286 -4165
rect 320 -4199 392 -4165
rect 224 -4229 392 -4199
rect 190 -4231 426 -4229
rect 190 -4233 286 -4231
rect 320 -4233 426 -4231
rect 224 -4267 286 -4233
rect 320 -4267 392 -4233
rect 224 -4301 392 -4267
rect 224 -4335 286 -4301
rect 320 -4335 392 -4301
rect 190 -4337 286 -4335
rect 320 -4337 426 -4335
rect 190 -4339 426 -4337
rect 224 -4369 392 -4339
rect 224 -4403 286 -4369
rect 320 -4403 392 -4369
rect 190 -4409 286 -4403
rect 320 -4409 426 -4403
rect 190 -4411 426 -4409
rect 224 -4437 392 -4411
rect 224 -4471 286 -4437
rect 320 -4471 392 -4437
rect 190 -4481 286 -4471
rect 320 -4481 426 -4471
rect 190 -4483 426 -4481
rect 224 -4505 392 -4483
rect 224 -4539 286 -4505
rect 320 -4539 392 -4505
rect 190 -4553 286 -4539
rect 320 -4553 426 -4539
rect 190 -4555 426 -4553
rect 224 -4573 392 -4555
rect 224 -4607 286 -4573
rect 320 -4607 392 -4573
rect 190 -4625 286 -4607
rect 320 -4625 426 -4607
rect 190 -4627 426 -4625
rect 224 -4641 392 -4627
rect 224 -4675 286 -4641
rect 320 -4675 392 -4641
rect 190 -4697 286 -4675
rect 320 -4697 426 -4675
rect 190 -4699 426 -4697
rect 224 -4709 392 -4699
rect 224 -4743 286 -4709
rect 320 -4743 392 -4709
rect 190 -4769 286 -4743
rect 320 -4769 426 -4743
rect 190 -4771 426 -4769
rect 224 -4777 392 -4771
rect 224 -4811 286 -4777
rect 320 -4811 392 -4777
rect 190 -4841 286 -4811
rect 320 -4841 426 -4811
rect 190 -4843 426 -4841
rect 224 -4845 392 -4843
rect 224 -4879 286 -4845
rect 320 -4879 392 -4845
rect 190 -4913 286 -4879
rect 320 -4913 426 -4879
rect 224 -4947 286 -4913
rect 320 -4947 392 -4913
rect 224 -4949 392 -4947
rect 190 -4951 426 -4949
rect 190 -4981 286 -4951
rect 320 -4981 426 -4951
rect -392 -5021 -224 -5015
rect -426 -5023 -190 -5021
rect -426 -5057 -330 -5023
rect -296 -5057 -190 -5023
rect -426 -5090 -190 -5057
rect 224 -5015 286 -4981
rect 320 -5015 392 -4981
rect 528 4985 704 5004
rect 528 4981 563 4985
rect 669 4981 704 4985
rect 528 -4981 531 4981
rect 701 -4981 704 4981
rect 528 -4985 563 -4981
rect 669 -4985 704 -4981
rect 528 -5004 704 -4985
rect 840 4981 902 5015
rect 936 4981 1008 5015
rect 1422 5057 1540 5090
rect 1422 5023 1494 5057
rect 1528 5023 1540 5057
rect 1422 5021 1540 5023
rect 806 4951 902 4981
rect 936 4951 1042 4981
rect 806 4949 1042 4951
rect 840 4947 1008 4949
rect 840 4913 902 4947
rect 936 4913 1008 4947
rect 806 4879 902 4913
rect 936 4879 1042 4913
rect 840 4845 902 4879
rect 936 4845 1008 4879
rect 840 4843 1008 4845
rect 806 4841 1042 4843
rect 806 4811 902 4841
rect 936 4811 1042 4841
rect 840 4777 902 4811
rect 936 4777 1008 4811
rect 840 4771 1008 4777
rect 806 4769 1042 4771
rect 806 4743 902 4769
rect 936 4743 1042 4769
rect 840 4709 902 4743
rect 936 4709 1008 4743
rect 840 4699 1008 4709
rect 806 4697 1042 4699
rect 806 4675 902 4697
rect 936 4675 1042 4697
rect 840 4641 902 4675
rect 936 4641 1008 4675
rect 840 4627 1008 4641
rect 806 4625 1042 4627
rect 806 4607 902 4625
rect 936 4607 1042 4625
rect 840 4573 902 4607
rect 936 4573 1008 4607
rect 840 4555 1008 4573
rect 806 4553 1042 4555
rect 806 4539 902 4553
rect 936 4539 1042 4553
rect 840 4505 902 4539
rect 936 4505 1008 4539
rect 840 4483 1008 4505
rect 806 4481 1042 4483
rect 806 4471 902 4481
rect 936 4471 1042 4481
rect 840 4437 902 4471
rect 936 4437 1008 4471
rect 840 4411 1008 4437
rect 806 4409 1042 4411
rect 806 4403 902 4409
rect 936 4403 1042 4409
rect 840 4369 902 4403
rect 936 4369 1008 4403
rect 840 4339 1008 4369
rect 806 4337 1042 4339
rect 806 4335 902 4337
rect 936 4335 1042 4337
rect 840 4301 902 4335
rect 936 4301 1008 4335
rect 840 4267 1008 4301
rect 840 4233 902 4267
rect 936 4233 1008 4267
rect 806 4231 902 4233
rect 936 4231 1042 4233
rect 806 4229 1042 4231
rect 840 4199 1008 4229
rect 840 4165 902 4199
rect 936 4165 1008 4199
rect 806 4159 902 4165
rect 936 4159 1042 4165
rect 806 4157 1042 4159
rect 840 4131 1008 4157
rect 840 4097 902 4131
rect 936 4097 1008 4131
rect 806 4087 902 4097
rect 936 4087 1042 4097
rect 806 4085 1042 4087
rect 840 4063 1008 4085
rect 840 4029 902 4063
rect 936 4029 1008 4063
rect 806 4015 902 4029
rect 936 4015 1042 4029
rect 806 4013 1042 4015
rect 840 3995 1008 4013
rect 840 3961 902 3995
rect 936 3961 1008 3995
rect 806 3943 902 3961
rect 936 3943 1042 3961
rect 806 3941 1042 3943
rect 840 3927 1008 3941
rect 840 3893 902 3927
rect 936 3893 1008 3927
rect 806 3871 902 3893
rect 936 3871 1042 3893
rect 806 3869 1042 3871
rect 840 3859 1008 3869
rect 840 3825 902 3859
rect 936 3825 1008 3859
rect 806 3799 902 3825
rect 936 3799 1042 3825
rect 806 3797 1042 3799
rect 840 3791 1008 3797
rect 840 3757 902 3791
rect 936 3757 1008 3791
rect 806 3727 902 3757
rect 936 3727 1042 3757
rect 806 3725 1042 3727
rect 840 3723 1008 3725
rect 840 3689 902 3723
rect 936 3689 1008 3723
rect 806 3655 902 3689
rect 936 3655 1042 3689
rect 840 3621 902 3655
rect 936 3621 1008 3655
rect 840 3619 1008 3621
rect 806 3617 1042 3619
rect 806 3587 902 3617
rect 936 3587 1042 3617
rect 840 3553 902 3587
rect 936 3553 1008 3587
rect 840 3547 1008 3553
rect 806 3545 1042 3547
rect 806 3519 902 3545
rect 936 3519 1042 3545
rect 840 3485 902 3519
rect 936 3485 1008 3519
rect 840 3475 1008 3485
rect 806 3473 1042 3475
rect 806 3451 902 3473
rect 936 3451 1042 3473
rect 840 3417 902 3451
rect 936 3417 1008 3451
rect 840 3403 1008 3417
rect 806 3401 1042 3403
rect 806 3383 902 3401
rect 936 3383 1042 3401
rect 840 3349 902 3383
rect 936 3349 1008 3383
rect 840 3331 1008 3349
rect 806 3329 1042 3331
rect 806 3315 902 3329
rect 936 3315 1042 3329
rect 840 3281 902 3315
rect 936 3281 1008 3315
rect 840 3259 1008 3281
rect 806 3257 1042 3259
rect 806 3247 902 3257
rect 936 3247 1042 3257
rect 840 3213 902 3247
rect 936 3213 1008 3247
rect 840 3187 1008 3213
rect 806 3185 1042 3187
rect 806 3179 902 3185
rect 936 3179 1042 3185
rect 840 3145 902 3179
rect 936 3145 1008 3179
rect 840 3115 1008 3145
rect 806 3113 1042 3115
rect 806 3111 902 3113
rect 936 3111 1042 3113
rect 840 3077 902 3111
rect 936 3077 1008 3111
rect 840 3043 1008 3077
rect 840 3009 902 3043
rect 936 3009 1008 3043
rect 806 3007 902 3009
rect 936 3007 1042 3009
rect 806 3005 1042 3007
rect 840 2975 1008 3005
rect 840 2941 902 2975
rect 936 2941 1008 2975
rect 806 2935 902 2941
rect 936 2935 1042 2941
rect 806 2933 1042 2935
rect 840 2907 1008 2933
rect 840 2873 902 2907
rect 936 2873 1008 2907
rect 806 2863 902 2873
rect 936 2863 1042 2873
rect 806 2861 1042 2863
rect 840 2839 1008 2861
rect 840 2805 902 2839
rect 936 2805 1008 2839
rect 806 2791 902 2805
rect 936 2791 1042 2805
rect 806 2789 1042 2791
rect 840 2771 1008 2789
rect 840 2737 902 2771
rect 936 2737 1008 2771
rect 806 2719 902 2737
rect 936 2719 1042 2737
rect 806 2717 1042 2719
rect 840 2703 1008 2717
rect 840 2669 902 2703
rect 936 2669 1008 2703
rect 806 2647 902 2669
rect 936 2647 1042 2669
rect 806 2645 1042 2647
rect 840 2635 1008 2645
rect 840 2601 902 2635
rect 936 2601 1008 2635
rect 806 2575 902 2601
rect 936 2575 1042 2601
rect 806 2573 1042 2575
rect 840 2567 1008 2573
rect 840 2533 902 2567
rect 936 2533 1008 2567
rect 806 2503 902 2533
rect 936 2503 1042 2533
rect 806 2501 1042 2503
rect 840 2499 1008 2501
rect 840 2465 902 2499
rect 936 2465 1008 2499
rect 806 2431 902 2465
rect 936 2431 1042 2465
rect 840 2397 902 2431
rect 936 2397 1008 2431
rect 840 2395 1008 2397
rect 806 2393 1042 2395
rect 806 2363 902 2393
rect 936 2363 1042 2393
rect 840 2329 902 2363
rect 936 2329 1008 2363
rect 840 2323 1008 2329
rect 806 2321 1042 2323
rect 806 2295 902 2321
rect 936 2295 1042 2321
rect 840 2261 902 2295
rect 936 2261 1008 2295
rect 840 2251 1008 2261
rect 806 2249 1042 2251
rect 806 2227 902 2249
rect 936 2227 1042 2249
rect 840 2193 902 2227
rect 936 2193 1008 2227
rect 840 2179 1008 2193
rect 806 2177 1042 2179
rect 806 2159 902 2177
rect 936 2159 1042 2177
rect 840 2125 902 2159
rect 936 2125 1008 2159
rect 840 2107 1008 2125
rect 806 2105 1042 2107
rect 806 2091 902 2105
rect 936 2091 1042 2105
rect 840 2057 902 2091
rect 936 2057 1008 2091
rect 840 2035 1008 2057
rect 806 2033 1042 2035
rect 806 2023 902 2033
rect 936 2023 1042 2033
rect 840 1989 902 2023
rect 936 1989 1008 2023
rect 840 1963 1008 1989
rect 806 1961 1042 1963
rect 806 1955 902 1961
rect 936 1955 1042 1961
rect 840 1921 902 1955
rect 936 1921 1008 1955
rect 840 1891 1008 1921
rect 806 1889 1042 1891
rect 806 1887 902 1889
rect 936 1887 1042 1889
rect 840 1853 902 1887
rect 936 1853 1008 1887
rect 840 1819 1008 1853
rect 840 1785 902 1819
rect 936 1785 1008 1819
rect 806 1783 902 1785
rect 936 1783 1042 1785
rect 806 1781 1042 1783
rect 840 1751 1008 1781
rect 840 1717 902 1751
rect 936 1717 1008 1751
rect 806 1711 902 1717
rect 936 1711 1042 1717
rect 806 1709 1042 1711
rect 840 1683 1008 1709
rect 840 1649 902 1683
rect 936 1649 1008 1683
rect 806 1639 902 1649
rect 936 1639 1042 1649
rect 806 1637 1042 1639
rect 840 1615 1008 1637
rect 840 1581 902 1615
rect 936 1581 1008 1615
rect 806 1567 902 1581
rect 936 1567 1042 1581
rect 806 1565 1042 1567
rect 840 1547 1008 1565
rect 840 1513 902 1547
rect 936 1513 1008 1547
rect 806 1495 902 1513
rect 936 1495 1042 1513
rect 806 1493 1042 1495
rect 840 1479 1008 1493
rect 840 1445 902 1479
rect 936 1445 1008 1479
rect 806 1423 902 1445
rect 936 1423 1042 1445
rect 806 1421 1042 1423
rect 840 1411 1008 1421
rect 840 1377 902 1411
rect 936 1377 1008 1411
rect 806 1351 902 1377
rect 936 1351 1042 1377
rect 806 1349 1042 1351
rect 840 1343 1008 1349
rect 840 1309 902 1343
rect 936 1309 1008 1343
rect 806 1279 902 1309
rect 936 1279 1042 1309
rect 806 1277 1042 1279
rect 840 1275 1008 1277
rect 840 1241 902 1275
rect 936 1241 1008 1275
rect 806 1207 902 1241
rect 936 1207 1042 1241
rect 840 1173 902 1207
rect 936 1173 1008 1207
rect 840 1171 1008 1173
rect 806 1169 1042 1171
rect 806 1139 902 1169
rect 936 1139 1042 1169
rect 840 1105 902 1139
rect 936 1105 1008 1139
rect 840 1099 1008 1105
rect 806 1097 1042 1099
rect 806 1071 902 1097
rect 936 1071 1042 1097
rect 840 1037 902 1071
rect 936 1037 1008 1071
rect 840 1027 1008 1037
rect 806 1025 1042 1027
rect 806 1003 902 1025
rect 936 1003 1042 1025
rect 840 969 902 1003
rect 936 969 1008 1003
rect 840 955 1008 969
rect 806 953 1042 955
rect 806 935 902 953
rect 936 935 1042 953
rect 840 901 902 935
rect 936 901 1008 935
rect 840 883 1008 901
rect 806 881 1042 883
rect 806 867 902 881
rect 936 867 1042 881
rect 840 833 902 867
rect 936 833 1008 867
rect 840 811 1008 833
rect 806 809 1042 811
rect 806 799 902 809
rect 936 799 1042 809
rect 840 765 902 799
rect 936 765 1008 799
rect 840 739 1008 765
rect 806 737 1042 739
rect 806 731 902 737
rect 936 731 1042 737
rect 840 697 902 731
rect 936 697 1008 731
rect 840 667 1008 697
rect 806 665 1042 667
rect 806 663 902 665
rect 936 663 1042 665
rect 840 629 902 663
rect 936 629 1008 663
rect 840 595 1008 629
rect 840 561 902 595
rect 936 561 1008 595
rect 806 559 902 561
rect 936 559 1042 561
rect 806 557 1042 559
rect 840 527 1008 557
rect 840 493 902 527
rect 936 493 1008 527
rect 806 487 902 493
rect 936 487 1042 493
rect 806 485 1042 487
rect 840 459 1008 485
rect 840 425 902 459
rect 936 425 1008 459
rect 806 415 902 425
rect 936 415 1042 425
rect 806 413 1042 415
rect 840 391 1008 413
rect 840 357 902 391
rect 936 357 1008 391
rect 806 343 902 357
rect 936 343 1042 357
rect 806 341 1042 343
rect 840 323 1008 341
rect 840 289 902 323
rect 936 289 1008 323
rect 806 271 902 289
rect 936 271 1042 289
rect 806 269 1042 271
rect 840 255 1008 269
rect 840 221 902 255
rect 936 221 1008 255
rect 806 199 902 221
rect 936 199 1042 221
rect 806 197 1042 199
rect 840 187 1008 197
rect 840 153 902 187
rect 936 153 1008 187
rect 806 127 902 153
rect 936 127 1042 153
rect 806 125 1042 127
rect 840 119 1008 125
rect 840 85 902 119
rect 936 85 1008 119
rect 806 55 902 85
rect 936 55 1042 85
rect 806 53 1042 55
rect 840 51 1008 53
rect 840 17 902 51
rect 936 17 1008 51
rect 806 -17 902 17
rect 936 -17 1042 17
rect 840 -51 902 -17
rect 936 -51 1008 -17
rect 840 -53 1008 -51
rect 806 -55 1042 -53
rect 806 -85 902 -55
rect 936 -85 1042 -55
rect 840 -119 902 -85
rect 936 -119 1008 -85
rect 840 -125 1008 -119
rect 806 -127 1042 -125
rect 806 -153 902 -127
rect 936 -153 1042 -127
rect 840 -187 902 -153
rect 936 -187 1008 -153
rect 840 -197 1008 -187
rect 806 -199 1042 -197
rect 806 -221 902 -199
rect 936 -221 1042 -199
rect 840 -255 902 -221
rect 936 -255 1008 -221
rect 840 -269 1008 -255
rect 806 -271 1042 -269
rect 806 -289 902 -271
rect 936 -289 1042 -271
rect 840 -323 902 -289
rect 936 -323 1008 -289
rect 840 -341 1008 -323
rect 806 -343 1042 -341
rect 806 -357 902 -343
rect 936 -357 1042 -343
rect 840 -391 902 -357
rect 936 -391 1008 -357
rect 840 -413 1008 -391
rect 806 -415 1042 -413
rect 806 -425 902 -415
rect 936 -425 1042 -415
rect 840 -459 902 -425
rect 936 -459 1008 -425
rect 840 -485 1008 -459
rect 806 -487 1042 -485
rect 806 -493 902 -487
rect 936 -493 1042 -487
rect 840 -527 902 -493
rect 936 -527 1008 -493
rect 840 -557 1008 -527
rect 806 -559 1042 -557
rect 806 -561 902 -559
rect 936 -561 1042 -559
rect 840 -595 902 -561
rect 936 -595 1008 -561
rect 840 -629 1008 -595
rect 840 -663 902 -629
rect 936 -663 1008 -629
rect 806 -665 902 -663
rect 936 -665 1042 -663
rect 806 -667 1042 -665
rect 840 -697 1008 -667
rect 840 -731 902 -697
rect 936 -731 1008 -697
rect 806 -737 902 -731
rect 936 -737 1042 -731
rect 806 -739 1042 -737
rect 840 -765 1008 -739
rect 840 -799 902 -765
rect 936 -799 1008 -765
rect 806 -809 902 -799
rect 936 -809 1042 -799
rect 806 -811 1042 -809
rect 840 -833 1008 -811
rect 840 -867 902 -833
rect 936 -867 1008 -833
rect 806 -881 902 -867
rect 936 -881 1042 -867
rect 806 -883 1042 -881
rect 840 -901 1008 -883
rect 840 -935 902 -901
rect 936 -935 1008 -901
rect 806 -953 902 -935
rect 936 -953 1042 -935
rect 806 -955 1042 -953
rect 840 -969 1008 -955
rect 840 -1003 902 -969
rect 936 -1003 1008 -969
rect 806 -1025 902 -1003
rect 936 -1025 1042 -1003
rect 806 -1027 1042 -1025
rect 840 -1037 1008 -1027
rect 840 -1071 902 -1037
rect 936 -1071 1008 -1037
rect 806 -1097 902 -1071
rect 936 -1097 1042 -1071
rect 806 -1099 1042 -1097
rect 840 -1105 1008 -1099
rect 840 -1139 902 -1105
rect 936 -1139 1008 -1105
rect 806 -1169 902 -1139
rect 936 -1169 1042 -1139
rect 806 -1171 1042 -1169
rect 840 -1173 1008 -1171
rect 840 -1207 902 -1173
rect 936 -1207 1008 -1173
rect 806 -1241 902 -1207
rect 936 -1241 1042 -1207
rect 840 -1275 902 -1241
rect 936 -1275 1008 -1241
rect 840 -1277 1008 -1275
rect 806 -1279 1042 -1277
rect 806 -1309 902 -1279
rect 936 -1309 1042 -1279
rect 840 -1343 902 -1309
rect 936 -1343 1008 -1309
rect 840 -1349 1008 -1343
rect 806 -1351 1042 -1349
rect 806 -1377 902 -1351
rect 936 -1377 1042 -1351
rect 840 -1411 902 -1377
rect 936 -1411 1008 -1377
rect 840 -1421 1008 -1411
rect 806 -1423 1042 -1421
rect 806 -1445 902 -1423
rect 936 -1445 1042 -1423
rect 840 -1479 902 -1445
rect 936 -1479 1008 -1445
rect 840 -1493 1008 -1479
rect 806 -1495 1042 -1493
rect 806 -1513 902 -1495
rect 936 -1513 1042 -1495
rect 840 -1547 902 -1513
rect 936 -1547 1008 -1513
rect 840 -1565 1008 -1547
rect 806 -1567 1042 -1565
rect 806 -1581 902 -1567
rect 936 -1581 1042 -1567
rect 840 -1615 902 -1581
rect 936 -1615 1008 -1581
rect 840 -1637 1008 -1615
rect 806 -1639 1042 -1637
rect 806 -1649 902 -1639
rect 936 -1649 1042 -1639
rect 840 -1683 902 -1649
rect 936 -1683 1008 -1649
rect 840 -1709 1008 -1683
rect 806 -1711 1042 -1709
rect 806 -1717 902 -1711
rect 936 -1717 1042 -1711
rect 840 -1751 902 -1717
rect 936 -1751 1008 -1717
rect 840 -1781 1008 -1751
rect 806 -1783 1042 -1781
rect 806 -1785 902 -1783
rect 936 -1785 1042 -1783
rect 840 -1819 902 -1785
rect 936 -1819 1008 -1785
rect 840 -1853 1008 -1819
rect 840 -1887 902 -1853
rect 936 -1887 1008 -1853
rect 806 -1889 902 -1887
rect 936 -1889 1042 -1887
rect 806 -1891 1042 -1889
rect 840 -1921 1008 -1891
rect 840 -1955 902 -1921
rect 936 -1955 1008 -1921
rect 806 -1961 902 -1955
rect 936 -1961 1042 -1955
rect 806 -1963 1042 -1961
rect 840 -1989 1008 -1963
rect 840 -2023 902 -1989
rect 936 -2023 1008 -1989
rect 806 -2033 902 -2023
rect 936 -2033 1042 -2023
rect 806 -2035 1042 -2033
rect 840 -2057 1008 -2035
rect 840 -2091 902 -2057
rect 936 -2091 1008 -2057
rect 806 -2105 902 -2091
rect 936 -2105 1042 -2091
rect 806 -2107 1042 -2105
rect 840 -2125 1008 -2107
rect 840 -2159 902 -2125
rect 936 -2159 1008 -2125
rect 806 -2177 902 -2159
rect 936 -2177 1042 -2159
rect 806 -2179 1042 -2177
rect 840 -2193 1008 -2179
rect 840 -2227 902 -2193
rect 936 -2227 1008 -2193
rect 806 -2249 902 -2227
rect 936 -2249 1042 -2227
rect 806 -2251 1042 -2249
rect 840 -2261 1008 -2251
rect 840 -2295 902 -2261
rect 936 -2295 1008 -2261
rect 806 -2321 902 -2295
rect 936 -2321 1042 -2295
rect 806 -2323 1042 -2321
rect 840 -2329 1008 -2323
rect 840 -2363 902 -2329
rect 936 -2363 1008 -2329
rect 806 -2393 902 -2363
rect 936 -2393 1042 -2363
rect 806 -2395 1042 -2393
rect 840 -2397 1008 -2395
rect 840 -2431 902 -2397
rect 936 -2431 1008 -2397
rect 806 -2465 902 -2431
rect 936 -2465 1042 -2431
rect 840 -2499 902 -2465
rect 936 -2499 1008 -2465
rect 840 -2501 1008 -2499
rect 806 -2503 1042 -2501
rect 806 -2533 902 -2503
rect 936 -2533 1042 -2503
rect 840 -2567 902 -2533
rect 936 -2567 1008 -2533
rect 840 -2573 1008 -2567
rect 806 -2575 1042 -2573
rect 806 -2601 902 -2575
rect 936 -2601 1042 -2575
rect 840 -2635 902 -2601
rect 936 -2635 1008 -2601
rect 840 -2645 1008 -2635
rect 806 -2647 1042 -2645
rect 806 -2669 902 -2647
rect 936 -2669 1042 -2647
rect 840 -2703 902 -2669
rect 936 -2703 1008 -2669
rect 840 -2717 1008 -2703
rect 806 -2719 1042 -2717
rect 806 -2737 902 -2719
rect 936 -2737 1042 -2719
rect 840 -2771 902 -2737
rect 936 -2771 1008 -2737
rect 840 -2789 1008 -2771
rect 806 -2791 1042 -2789
rect 806 -2805 902 -2791
rect 936 -2805 1042 -2791
rect 840 -2839 902 -2805
rect 936 -2839 1008 -2805
rect 840 -2861 1008 -2839
rect 806 -2863 1042 -2861
rect 806 -2873 902 -2863
rect 936 -2873 1042 -2863
rect 840 -2907 902 -2873
rect 936 -2907 1008 -2873
rect 840 -2933 1008 -2907
rect 806 -2935 1042 -2933
rect 806 -2941 902 -2935
rect 936 -2941 1042 -2935
rect 840 -2975 902 -2941
rect 936 -2975 1008 -2941
rect 840 -3005 1008 -2975
rect 806 -3007 1042 -3005
rect 806 -3009 902 -3007
rect 936 -3009 1042 -3007
rect 840 -3043 902 -3009
rect 936 -3043 1008 -3009
rect 840 -3077 1008 -3043
rect 840 -3111 902 -3077
rect 936 -3111 1008 -3077
rect 806 -3113 902 -3111
rect 936 -3113 1042 -3111
rect 806 -3115 1042 -3113
rect 840 -3145 1008 -3115
rect 840 -3179 902 -3145
rect 936 -3179 1008 -3145
rect 806 -3185 902 -3179
rect 936 -3185 1042 -3179
rect 806 -3187 1042 -3185
rect 840 -3213 1008 -3187
rect 840 -3247 902 -3213
rect 936 -3247 1008 -3213
rect 806 -3257 902 -3247
rect 936 -3257 1042 -3247
rect 806 -3259 1042 -3257
rect 840 -3281 1008 -3259
rect 840 -3315 902 -3281
rect 936 -3315 1008 -3281
rect 806 -3329 902 -3315
rect 936 -3329 1042 -3315
rect 806 -3331 1042 -3329
rect 840 -3349 1008 -3331
rect 840 -3383 902 -3349
rect 936 -3383 1008 -3349
rect 806 -3401 902 -3383
rect 936 -3401 1042 -3383
rect 806 -3403 1042 -3401
rect 840 -3417 1008 -3403
rect 840 -3451 902 -3417
rect 936 -3451 1008 -3417
rect 806 -3473 902 -3451
rect 936 -3473 1042 -3451
rect 806 -3475 1042 -3473
rect 840 -3485 1008 -3475
rect 840 -3519 902 -3485
rect 936 -3519 1008 -3485
rect 806 -3545 902 -3519
rect 936 -3545 1042 -3519
rect 806 -3547 1042 -3545
rect 840 -3553 1008 -3547
rect 840 -3587 902 -3553
rect 936 -3587 1008 -3553
rect 806 -3617 902 -3587
rect 936 -3617 1042 -3587
rect 806 -3619 1042 -3617
rect 840 -3621 1008 -3619
rect 840 -3655 902 -3621
rect 936 -3655 1008 -3621
rect 806 -3689 902 -3655
rect 936 -3689 1042 -3655
rect 840 -3723 902 -3689
rect 936 -3723 1008 -3689
rect 840 -3725 1008 -3723
rect 806 -3727 1042 -3725
rect 806 -3757 902 -3727
rect 936 -3757 1042 -3727
rect 840 -3791 902 -3757
rect 936 -3791 1008 -3757
rect 840 -3797 1008 -3791
rect 806 -3799 1042 -3797
rect 806 -3825 902 -3799
rect 936 -3825 1042 -3799
rect 840 -3859 902 -3825
rect 936 -3859 1008 -3825
rect 840 -3869 1008 -3859
rect 806 -3871 1042 -3869
rect 806 -3893 902 -3871
rect 936 -3893 1042 -3871
rect 840 -3927 902 -3893
rect 936 -3927 1008 -3893
rect 840 -3941 1008 -3927
rect 806 -3943 1042 -3941
rect 806 -3961 902 -3943
rect 936 -3961 1042 -3943
rect 840 -3995 902 -3961
rect 936 -3995 1008 -3961
rect 840 -4013 1008 -3995
rect 806 -4015 1042 -4013
rect 806 -4029 902 -4015
rect 936 -4029 1042 -4015
rect 840 -4063 902 -4029
rect 936 -4063 1008 -4029
rect 840 -4085 1008 -4063
rect 806 -4087 1042 -4085
rect 806 -4097 902 -4087
rect 936 -4097 1042 -4087
rect 840 -4131 902 -4097
rect 936 -4131 1008 -4097
rect 840 -4157 1008 -4131
rect 806 -4159 1042 -4157
rect 806 -4165 902 -4159
rect 936 -4165 1042 -4159
rect 840 -4199 902 -4165
rect 936 -4199 1008 -4165
rect 840 -4229 1008 -4199
rect 806 -4231 1042 -4229
rect 806 -4233 902 -4231
rect 936 -4233 1042 -4231
rect 840 -4267 902 -4233
rect 936 -4267 1008 -4233
rect 840 -4301 1008 -4267
rect 840 -4335 902 -4301
rect 936 -4335 1008 -4301
rect 806 -4337 902 -4335
rect 936 -4337 1042 -4335
rect 806 -4339 1042 -4337
rect 840 -4369 1008 -4339
rect 840 -4403 902 -4369
rect 936 -4403 1008 -4369
rect 806 -4409 902 -4403
rect 936 -4409 1042 -4403
rect 806 -4411 1042 -4409
rect 840 -4437 1008 -4411
rect 840 -4471 902 -4437
rect 936 -4471 1008 -4437
rect 806 -4481 902 -4471
rect 936 -4481 1042 -4471
rect 806 -4483 1042 -4481
rect 840 -4505 1008 -4483
rect 840 -4539 902 -4505
rect 936 -4539 1008 -4505
rect 806 -4553 902 -4539
rect 936 -4553 1042 -4539
rect 806 -4555 1042 -4553
rect 840 -4573 1008 -4555
rect 840 -4607 902 -4573
rect 936 -4607 1008 -4573
rect 806 -4625 902 -4607
rect 936 -4625 1042 -4607
rect 806 -4627 1042 -4625
rect 840 -4641 1008 -4627
rect 840 -4675 902 -4641
rect 936 -4675 1008 -4641
rect 806 -4697 902 -4675
rect 936 -4697 1042 -4675
rect 806 -4699 1042 -4697
rect 840 -4709 1008 -4699
rect 840 -4743 902 -4709
rect 936 -4743 1008 -4709
rect 806 -4769 902 -4743
rect 936 -4769 1042 -4743
rect 806 -4771 1042 -4769
rect 840 -4777 1008 -4771
rect 840 -4811 902 -4777
rect 936 -4811 1008 -4777
rect 806 -4841 902 -4811
rect 936 -4841 1042 -4811
rect 806 -4843 1042 -4841
rect 840 -4845 1008 -4843
rect 840 -4879 902 -4845
rect 936 -4879 1008 -4845
rect 806 -4913 902 -4879
rect 936 -4913 1042 -4879
rect 840 -4947 902 -4913
rect 936 -4947 1008 -4913
rect 840 -4949 1008 -4947
rect 806 -4951 1042 -4949
rect 806 -4981 902 -4951
rect 936 -4981 1042 -4951
rect 224 -5021 392 -5015
rect 190 -5023 426 -5021
rect 190 -5057 286 -5023
rect 320 -5057 426 -5023
rect 190 -5090 426 -5057
rect 840 -5015 902 -4981
rect 936 -5015 1008 -4981
rect 1144 4985 1320 5004
rect 1144 4981 1179 4985
rect 1285 4981 1320 4985
rect 1144 -4981 1147 4981
rect 1317 -4981 1320 4981
rect 1144 -4985 1179 -4981
rect 1285 -4985 1320 -4981
rect 1144 -5004 1320 -4985
rect 840 -5021 1008 -5015
rect 806 -5023 1042 -5021
rect 806 -5057 902 -5023
rect 936 -5057 1042 -5023
rect 806 -5090 1042 -5057
rect 1528 -5021 1540 5021
rect 1422 -5023 1540 -5021
rect 1422 -5057 1494 -5023
rect 1528 -5057 1540 -5023
rect 1422 -5090 1540 -5057
rect -1540 -5124 -1357 -5090
rect -1317 -5124 -1285 -5090
rect -1249 -5124 -1215 -5090
rect -1179 -5124 -1147 -5090
rect -1107 -5124 -741 -5090
rect -701 -5124 -669 -5090
rect -633 -5124 -599 -5090
rect -563 -5124 -531 -5090
rect -491 -5124 -125 -5090
rect -85 -5124 -53 -5090
rect -17 -5124 17 -5090
rect 53 -5124 85 -5090
rect 125 -5124 491 -5090
rect 531 -5124 563 -5090
rect 599 -5124 633 -5090
rect 669 -5124 701 -5090
rect 741 -5124 1107 -5090
rect 1147 -5124 1179 -5090
rect 1215 -5124 1249 -5090
rect 1285 -5124 1317 -5090
rect 1357 -5124 1540 -5090
rect -1540 -5188 1540 -5124
<< viali >>
rect -1357 5090 -1351 5124
rect -1351 5090 -1323 5124
rect -1285 5090 -1283 5124
rect -1283 5090 -1251 5124
rect -1213 5090 -1181 5124
rect -1181 5090 -1179 5124
rect -1141 5090 -1113 5124
rect -1113 5090 -1107 5124
rect -741 5090 -735 5124
rect -735 5090 -707 5124
rect -669 5090 -667 5124
rect -667 5090 -635 5124
rect -597 5090 -565 5124
rect -565 5090 -563 5124
rect -525 5090 -497 5124
rect -497 5090 -491 5124
rect -125 5090 -119 5124
rect -119 5090 -91 5124
rect -53 5090 -51 5124
rect -51 5090 -19 5124
rect 19 5090 51 5124
rect 51 5090 53 5124
rect 91 5090 119 5124
rect 119 5090 125 5124
rect 491 5090 497 5124
rect 497 5090 525 5124
rect 563 5090 565 5124
rect 565 5090 597 5124
rect 635 5090 667 5124
rect 667 5090 669 5124
rect 707 5090 735 5124
rect 735 5090 741 5124
rect 1107 5090 1113 5124
rect 1113 5090 1141 5124
rect 1179 5090 1181 5124
rect 1181 5090 1213 5124
rect 1251 5090 1283 5124
rect 1283 5090 1285 5124
rect 1323 5090 1351 5124
rect 1351 5090 1357 5124
rect -1528 5023 -1494 5057
rect -1528 5015 -1422 5021
rect -1528 -5015 -1524 5015
rect -1524 -5015 -1422 5015
rect -946 5023 -912 5057
rect -1042 5015 -1008 5021
rect -840 5015 -806 5021
rect -1285 4981 -1179 4985
rect -1285 -4981 -1179 4981
rect -1285 -4985 -1179 -4981
rect -1042 4987 -1008 5015
rect -946 4981 -912 4985
rect -840 4987 -806 5015
rect -330 5023 -296 5057
rect -426 5015 -392 5021
rect -224 5015 -190 5021
rect -946 4951 -912 4981
rect -1042 4947 -1008 4949
rect -840 4947 -806 4949
rect -1042 4915 -1008 4947
rect -840 4915 -806 4947
rect -946 4879 -912 4913
rect -1042 4845 -1008 4877
rect -840 4845 -806 4877
rect -1042 4843 -1008 4845
rect -840 4843 -806 4845
rect -946 4811 -912 4841
rect -1042 4777 -1008 4805
rect -946 4807 -912 4811
rect -840 4777 -806 4805
rect -1042 4771 -1008 4777
rect -840 4771 -806 4777
rect -946 4743 -912 4769
rect -1042 4709 -1008 4733
rect -946 4735 -912 4743
rect -840 4709 -806 4733
rect -1042 4699 -1008 4709
rect -840 4699 -806 4709
rect -946 4675 -912 4697
rect -1042 4641 -1008 4661
rect -946 4663 -912 4675
rect -840 4641 -806 4661
rect -1042 4627 -1008 4641
rect -840 4627 -806 4641
rect -946 4607 -912 4625
rect -1042 4573 -1008 4589
rect -946 4591 -912 4607
rect -840 4573 -806 4589
rect -1042 4555 -1008 4573
rect -840 4555 -806 4573
rect -946 4539 -912 4553
rect -1042 4505 -1008 4517
rect -946 4519 -912 4539
rect -840 4505 -806 4517
rect -1042 4483 -1008 4505
rect -840 4483 -806 4505
rect -946 4471 -912 4481
rect -1042 4437 -1008 4445
rect -946 4447 -912 4471
rect -840 4437 -806 4445
rect -1042 4411 -1008 4437
rect -840 4411 -806 4437
rect -946 4403 -912 4409
rect -1042 4369 -1008 4373
rect -946 4375 -912 4403
rect -840 4369 -806 4373
rect -1042 4339 -1008 4369
rect -840 4339 -806 4369
rect -946 4335 -912 4337
rect -946 4303 -912 4335
rect -1042 4267 -1008 4301
rect -840 4267 -806 4301
rect -946 4233 -912 4265
rect -946 4231 -912 4233
rect -1042 4199 -1008 4229
rect -840 4199 -806 4229
rect -1042 4195 -1008 4199
rect -946 4165 -912 4193
rect -840 4195 -806 4199
rect -946 4159 -912 4165
rect -1042 4131 -1008 4157
rect -840 4131 -806 4157
rect -1042 4123 -1008 4131
rect -946 4097 -912 4121
rect -840 4123 -806 4131
rect -946 4087 -912 4097
rect -1042 4063 -1008 4085
rect -840 4063 -806 4085
rect -1042 4051 -1008 4063
rect -946 4029 -912 4049
rect -840 4051 -806 4063
rect -946 4015 -912 4029
rect -1042 3995 -1008 4013
rect -840 3995 -806 4013
rect -1042 3979 -1008 3995
rect -946 3961 -912 3977
rect -840 3979 -806 3995
rect -946 3943 -912 3961
rect -1042 3927 -1008 3941
rect -840 3927 -806 3941
rect -1042 3907 -1008 3927
rect -946 3893 -912 3905
rect -840 3907 -806 3927
rect -946 3871 -912 3893
rect -1042 3859 -1008 3869
rect -840 3859 -806 3869
rect -1042 3835 -1008 3859
rect -946 3825 -912 3833
rect -840 3835 -806 3859
rect -946 3799 -912 3825
rect -1042 3791 -1008 3797
rect -840 3791 -806 3797
rect -1042 3763 -1008 3791
rect -946 3757 -912 3761
rect -840 3763 -806 3791
rect -946 3727 -912 3757
rect -1042 3723 -1008 3725
rect -840 3723 -806 3725
rect -1042 3691 -1008 3723
rect -840 3691 -806 3723
rect -946 3655 -912 3689
rect -1042 3621 -1008 3653
rect -840 3621 -806 3653
rect -1042 3619 -1008 3621
rect -840 3619 -806 3621
rect -946 3587 -912 3617
rect -1042 3553 -1008 3581
rect -946 3583 -912 3587
rect -840 3553 -806 3581
rect -1042 3547 -1008 3553
rect -840 3547 -806 3553
rect -946 3519 -912 3545
rect -1042 3485 -1008 3509
rect -946 3511 -912 3519
rect -840 3485 -806 3509
rect -1042 3475 -1008 3485
rect -840 3475 -806 3485
rect -946 3451 -912 3473
rect -1042 3417 -1008 3437
rect -946 3439 -912 3451
rect -840 3417 -806 3437
rect -1042 3403 -1008 3417
rect -840 3403 -806 3417
rect -946 3383 -912 3401
rect -1042 3349 -1008 3365
rect -946 3367 -912 3383
rect -840 3349 -806 3365
rect -1042 3331 -1008 3349
rect -840 3331 -806 3349
rect -946 3315 -912 3329
rect -1042 3281 -1008 3293
rect -946 3295 -912 3315
rect -840 3281 -806 3293
rect -1042 3259 -1008 3281
rect -840 3259 -806 3281
rect -946 3247 -912 3257
rect -1042 3213 -1008 3221
rect -946 3223 -912 3247
rect -840 3213 -806 3221
rect -1042 3187 -1008 3213
rect -840 3187 -806 3213
rect -946 3179 -912 3185
rect -1042 3145 -1008 3149
rect -946 3151 -912 3179
rect -840 3145 -806 3149
rect -1042 3115 -1008 3145
rect -840 3115 -806 3145
rect -946 3111 -912 3113
rect -946 3079 -912 3111
rect -1042 3043 -1008 3077
rect -840 3043 -806 3077
rect -946 3009 -912 3041
rect -946 3007 -912 3009
rect -1042 2975 -1008 3005
rect -840 2975 -806 3005
rect -1042 2971 -1008 2975
rect -946 2941 -912 2969
rect -840 2971 -806 2975
rect -946 2935 -912 2941
rect -1042 2907 -1008 2933
rect -840 2907 -806 2933
rect -1042 2899 -1008 2907
rect -946 2873 -912 2897
rect -840 2899 -806 2907
rect -946 2863 -912 2873
rect -1042 2839 -1008 2861
rect -840 2839 -806 2861
rect -1042 2827 -1008 2839
rect -946 2805 -912 2825
rect -840 2827 -806 2839
rect -946 2791 -912 2805
rect -1042 2771 -1008 2789
rect -840 2771 -806 2789
rect -1042 2755 -1008 2771
rect -946 2737 -912 2753
rect -840 2755 -806 2771
rect -946 2719 -912 2737
rect -1042 2703 -1008 2717
rect -840 2703 -806 2717
rect -1042 2683 -1008 2703
rect -946 2669 -912 2681
rect -840 2683 -806 2703
rect -946 2647 -912 2669
rect -1042 2635 -1008 2645
rect -840 2635 -806 2645
rect -1042 2611 -1008 2635
rect -946 2601 -912 2609
rect -840 2611 -806 2635
rect -946 2575 -912 2601
rect -1042 2567 -1008 2573
rect -840 2567 -806 2573
rect -1042 2539 -1008 2567
rect -946 2533 -912 2537
rect -840 2539 -806 2567
rect -946 2503 -912 2533
rect -1042 2499 -1008 2501
rect -840 2499 -806 2501
rect -1042 2467 -1008 2499
rect -840 2467 -806 2499
rect -946 2431 -912 2465
rect -1042 2397 -1008 2429
rect -840 2397 -806 2429
rect -1042 2395 -1008 2397
rect -840 2395 -806 2397
rect -946 2363 -912 2393
rect -1042 2329 -1008 2357
rect -946 2359 -912 2363
rect -840 2329 -806 2357
rect -1042 2323 -1008 2329
rect -840 2323 -806 2329
rect -946 2295 -912 2321
rect -1042 2261 -1008 2285
rect -946 2287 -912 2295
rect -840 2261 -806 2285
rect -1042 2251 -1008 2261
rect -840 2251 -806 2261
rect -946 2227 -912 2249
rect -1042 2193 -1008 2213
rect -946 2215 -912 2227
rect -840 2193 -806 2213
rect -1042 2179 -1008 2193
rect -840 2179 -806 2193
rect -946 2159 -912 2177
rect -1042 2125 -1008 2141
rect -946 2143 -912 2159
rect -840 2125 -806 2141
rect -1042 2107 -1008 2125
rect -840 2107 -806 2125
rect -946 2091 -912 2105
rect -1042 2057 -1008 2069
rect -946 2071 -912 2091
rect -840 2057 -806 2069
rect -1042 2035 -1008 2057
rect -840 2035 -806 2057
rect -946 2023 -912 2033
rect -1042 1989 -1008 1997
rect -946 1999 -912 2023
rect -840 1989 -806 1997
rect -1042 1963 -1008 1989
rect -840 1963 -806 1989
rect -946 1955 -912 1961
rect -1042 1921 -1008 1925
rect -946 1927 -912 1955
rect -840 1921 -806 1925
rect -1042 1891 -1008 1921
rect -840 1891 -806 1921
rect -946 1887 -912 1889
rect -946 1855 -912 1887
rect -1042 1819 -1008 1853
rect -840 1819 -806 1853
rect -946 1785 -912 1817
rect -946 1783 -912 1785
rect -1042 1751 -1008 1781
rect -840 1751 -806 1781
rect -1042 1747 -1008 1751
rect -946 1717 -912 1745
rect -840 1747 -806 1751
rect -946 1711 -912 1717
rect -1042 1683 -1008 1709
rect -840 1683 -806 1709
rect -1042 1675 -1008 1683
rect -946 1649 -912 1673
rect -840 1675 -806 1683
rect -946 1639 -912 1649
rect -1042 1615 -1008 1637
rect -840 1615 -806 1637
rect -1042 1603 -1008 1615
rect -946 1581 -912 1601
rect -840 1603 -806 1615
rect -946 1567 -912 1581
rect -1042 1547 -1008 1565
rect -840 1547 -806 1565
rect -1042 1531 -1008 1547
rect -946 1513 -912 1529
rect -840 1531 -806 1547
rect -946 1495 -912 1513
rect -1042 1479 -1008 1493
rect -840 1479 -806 1493
rect -1042 1459 -1008 1479
rect -946 1445 -912 1457
rect -840 1459 -806 1479
rect -946 1423 -912 1445
rect -1042 1411 -1008 1421
rect -840 1411 -806 1421
rect -1042 1387 -1008 1411
rect -946 1377 -912 1385
rect -840 1387 -806 1411
rect -946 1351 -912 1377
rect -1042 1343 -1008 1349
rect -840 1343 -806 1349
rect -1042 1315 -1008 1343
rect -946 1309 -912 1313
rect -840 1315 -806 1343
rect -946 1279 -912 1309
rect -1042 1275 -1008 1277
rect -840 1275 -806 1277
rect -1042 1243 -1008 1275
rect -840 1243 -806 1275
rect -946 1207 -912 1241
rect -1042 1173 -1008 1205
rect -840 1173 -806 1205
rect -1042 1171 -1008 1173
rect -840 1171 -806 1173
rect -946 1139 -912 1169
rect -1042 1105 -1008 1133
rect -946 1135 -912 1139
rect -840 1105 -806 1133
rect -1042 1099 -1008 1105
rect -840 1099 -806 1105
rect -946 1071 -912 1097
rect -1042 1037 -1008 1061
rect -946 1063 -912 1071
rect -840 1037 -806 1061
rect -1042 1027 -1008 1037
rect -840 1027 -806 1037
rect -946 1003 -912 1025
rect -1042 969 -1008 989
rect -946 991 -912 1003
rect -840 969 -806 989
rect -1042 955 -1008 969
rect -840 955 -806 969
rect -946 935 -912 953
rect -1042 901 -1008 917
rect -946 919 -912 935
rect -840 901 -806 917
rect -1042 883 -1008 901
rect -840 883 -806 901
rect -946 867 -912 881
rect -1042 833 -1008 845
rect -946 847 -912 867
rect -840 833 -806 845
rect -1042 811 -1008 833
rect -840 811 -806 833
rect -946 799 -912 809
rect -1042 765 -1008 773
rect -946 775 -912 799
rect -840 765 -806 773
rect -1042 739 -1008 765
rect -840 739 -806 765
rect -946 731 -912 737
rect -1042 697 -1008 701
rect -946 703 -912 731
rect -840 697 -806 701
rect -1042 667 -1008 697
rect -840 667 -806 697
rect -946 663 -912 665
rect -946 631 -912 663
rect -1042 595 -1008 629
rect -840 595 -806 629
rect -946 561 -912 593
rect -946 559 -912 561
rect -1042 527 -1008 557
rect -840 527 -806 557
rect -1042 523 -1008 527
rect -946 493 -912 521
rect -840 523 -806 527
rect -946 487 -912 493
rect -1042 459 -1008 485
rect -840 459 -806 485
rect -1042 451 -1008 459
rect -946 425 -912 449
rect -840 451 -806 459
rect -946 415 -912 425
rect -1042 391 -1008 413
rect -840 391 -806 413
rect -1042 379 -1008 391
rect -946 357 -912 377
rect -840 379 -806 391
rect -946 343 -912 357
rect -1042 323 -1008 341
rect -840 323 -806 341
rect -1042 307 -1008 323
rect -946 289 -912 305
rect -840 307 -806 323
rect -946 271 -912 289
rect -1042 255 -1008 269
rect -840 255 -806 269
rect -1042 235 -1008 255
rect -946 221 -912 233
rect -840 235 -806 255
rect -946 199 -912 221
rect -1042 187 -1008 197
rect -840 187 -806 197
rect -1042 163 -1008 187
rect -946 153 -912 161
rect -840 163 -806 187
rect -946 127 -912 153
rect -1042 119 -1008 125
rect -840 119 -806 125
rect -1042 91 -1008 119
rect -946 85 -912 89
rect -840 91 -806 119
rect -946 55 -912 85
rect -1042 51 -1008 53
rect -840 51 -806 53
rect -1042 19 -1008 51
rect -840 19 -806 51
rect -946 -17 -912 17
rect -1042 -51 -1008 -19
rect -840 -51 -806 -19
rect -1042 -53 -1008 -51
rect -840 -53 -806 -51
rect -946 -85 -912 -55
rect -1042 -119 -1008 -91
rect -946 -89 -912 -85
rect -840 -119 -806 -91
rect -1042 -125 -1008 -119
rect -840 -125 -806 -119
rect -946 -153 -912 -127
rect -1042 -187 -1008 -163
rect -946 -161 -912 -153
rect -840 -187 -806 -163
rect -1042 -197 -1008 -187
rect -840 -197 -806 -187
rect -946 -221 -912 -199
rect -1042 -255 -1008 -235
rect -946 -233 -912 -221
rect -840 -255 -806 -235
rect -1042 -269 -1008 -255
rect -840 -269 -806 -255
rect -946 -289 -912 -271
rect -1042 -323 -1008 -307
rect -946 -305 -912 -289
rect -840 -323 -806 -307
rect -1042 -341 -1008 -323
rect -840 -341 -806 -323
rect -946 -357 -912 -343
rect -1042 -391 -1008 -379
rect -946 -377 -912 -357
rect -840 -391 -806 -379
rect -1042 -413 -1008 -391
rect -840 -413 -806 -391
rect -946 -425 -912 -415
rect -1042 -459 -1008 -451
rect -946 -449 -912 -425
rect -840 -459 -806 -451
rect -1042 -485 -1008 -459
rect -840 -485 -806 -459
rect -946 -493 -912 -487
rect -1042 -527 -1008 -523
rect -946 -521 -912 -493
rect -840 -527 -806 -523
rect -1042 -557 -1008 -527
rect -840 -557 -806 -527
rect -946 -561 -912 -559
rect -946 -593 -912 -561
rect -1042 -629 -1008 -595
rect -840 -629 -806 -595
rect -946 -663 -912 -631
rect -946 -665 -912 -663
rect -1042 -697 -1008 -667
rect -840 -697 -806 -667
rect -1042 -701 -1008 -697
rect -946 -731 -912 -703
rect -840 -701 -806 -697
rect -946 -737 -912 -731
rect -1042 -765 -1008 -739
rect -840 -765 -806 -739
rect -1042 -773 -1008 -765
rect -946 -799 -912 -775
rect -840 -773 -806 -765
rect -946 -809 -912 -799
rect -1042 -833 -1008 -811
rect -840 -833 -806 -811
rect -1042 -845 -1008 -833
rect -946 -867 -912 -847
rect -840 -845 -806 -833
rect -946 -881 -912 -867
rect -1042 -901 -1008 -883
rect -840 -901 -806 -883
rect -1042 -917 -1008 -901
rect -946 -935 -912 -919
rect -840 -917 -806 -901
rect -946 -953 -912 -935
rect -1042 -969 -1008 -955
rect -840 -969 -806 -955
rect -1042 -989 -1008 -969
rect -946 -1003 -912 -991
rect -840 -989 -806 -969
rect -946 -1025 -912 -1003
rect -1042 -1037 -1008 -1027
rect -840 -1037 -806 -1027
rect -1042 -1061 -1008 -1037
rect -946 -1071 -912 -1063
rect -840 -1061 -806 -1037
rect -946 -1097 -912 -1071
rect -1042 -1105 -1008 -1099
rect -840 -1105 -806 -1099
rect -1042 -1133 -1008 -1105
rect -946 -1139 -912 -1135
rect -840 -1133 -806 -1105
rect -946 -1169 -912 -1139
rect -1042 -1173 -1008 -1171
rect -840 -1173 -806 -1171
rect -1042 -1205 -1008 -1173
rect -840 -1205 -806 -1173
rect -946 -1241 -912 -1207
rect -1042 -1275 -1008 -1243
rect -840 -1275 -806 -1243
rect -1042 -1277 -1008 -1275
rect -840 -1277 -806 -1275
rect -946 -1309 -912 -1279
rect -1042 -1343 -1008 -1315
rect -946 -1313 -912 -1309
rect -840 -1343 -806 -1315
rect -1042 -1349 -1008 -1343
rect -840 -1349 -806 -1343
rect -946 -1377 -912 -1351
rect -1042 -1411 -1008 -1387
rect -946 -1385 -912 -1377
rect -840 -1411 -806 -1387
rect -1042 -1421 -1008 -1411
rect -840 -1421 -806 -1411
rect -946 -1445 -912 -1423
rect -1042 -1479 -1008 -1459
rect -946 -1457 -912 -1445
rect -840 -1479 -806 -1459
rect -1042 -1493 -1008 -1479
rect -840 -1493 -806 -1479
rect -946 -1513 -912 -1495
rect -1042 -1547 -1008 -1531
rect -946 -1529 -912 -1513
rect -840 -1547 -806 -1531
rect -1042 -1565 -1008 -1547
rect -840 -1565 -806 -1547
rect -946 -1581 -912 -1567
rect -1042 -1615 -1008 -1603
rect -946 -1601 -912 -1581
rect -840 -1615 -806 -1603
rect -1042 -1637 -1008 -1615
rect -840 -1637 -806 -1615
rect -946 -1649 -912 -1639
rect -1042 -1683 -1008 -1675
rect -946 -1673 -912 -1649
rect -840 -1683 -806 -1675
rect -1042 -1709 -1008 -1683
rect -840 -1709 -806 -1683
rect -946 -1717 -912 -1711
rect -1042 -1751 -1008 -1747
rect -946 -1745 -912 -1717
rect -840 -1751 -806 -1747
rect -1042 -1781 -1008 -1751
rect -840 -1781 -806 -1751
rect -946 -1785 -912 -1783
rect -946 -1817 -912 -1785
rect -1042 -1853 -1008 -1819
rect -840 -1853 -806 -1819
rect -946 -1887 -912 -1855
rect -946 -1889 -912 -1887
rect -1042 -1921 -1008 -1891
rect -840 -1921 -806 -1891
rect -1042 -1925 -1008 -1921
rect -946 -1955 -912 -1927
rect -840 -1925 -806 -1921
rect -946 -1961 -912 -1955
rect -1042 -1989 -1008 -1963
rect -840 -1989 -806 -1963
rect -1042 -1997 -1008 -1989
rect -946 -2023 -912 -1999
rect -840 -1997 -806 -1989
rect -946 -2033 -912 -2023
rect -1042 -2057 -1008 -2035
rect -840 -2057 -806 -2035
rect -1042 -2069 -1008 -2057
rect -946 -2091 -912 -2071
rect -840 -2069 -806 -2057
rect -946 -2105 -912 -2091
rect -1042 -2125 -1008 -2107
rect -840 -2125 -806 -2107
rect -1042 -2141 -1008 -2125
rect -946 -2159 -912 -2143
rect -840 -2141 -806 -2125
rect -946 -2177 -912 -2159
rect -1042 -2193 -1008 -2179
rect -840 -2193 -806 -2179
rect -1042 -2213 -1008 -2193
rect -946 -2227 -912 -2215
rect -840 -2213 -806 -2193
rect -946 -2249 -912 -2227
rect -1042 -2261 -1008 -2251
rect -840 -2261 -806 -2251
rect -1042 -2285 -1008 -2261
rect -946 -2295 -912 -2287
rect -840 -2285 -806 -2261
rect -946 -2321 -912 -2295
rect -1042 -2329 -1008 -2323
rect -840 -2329 -806 -2323
rect -1042 -2357 -1008 -2329
rect -946 -2363 -912 -2359
rect -840 -2357 -806 -2329
rect -946 -2393 -912 -2363
rect -1042 -2397 -1008 -2395
rect -840 -2397 -806 -2395
rect -1042 -2429 -1008 -2397
rect -840 -2429 -806 -2397
rect -946 -2465 -912 -2431
rect -1042 -2499 -1008 -2467
rect -840 -2499 -806 -2467
rect -1042 -2501 -1008 -2499
rect -840 -2501 -806 -2499
rect -946 -2533 -912 -2503
rect -1042 -2567 -1008 -2539
rect -946 -2537 -912 -2533
rect -840 -2567 -806 -2539
rect -1042 -2573 -1008 -2567
rect -840 -2573 -806 -2567
rect -946 -2601 -912 -2575
rect -1042 -2635 -1008 -2611
rect -946 -2609 -912 -2601
rect -840 -2635 -806 -2611
rect -1042 -2645 -1008 -2635
rect -840 -2645 -806 -2635
rect -946 -2669 -912 -2647
rect -1042 -2703 -1008 -2683
rect -946 -2681 -912 -2669
rect -840 -2703 -806 -2683
rect -1042 -2717 -1008 -2703
rect -840 -2717 -806 -2703
rect -946 -2737 -912 -2719
rect -1042 -2771 -1008 -2755
rect -946 -2753 -912 -2737
rect -840 -2771 -806 -2755
rect -1042 -2789 -1008 -2771
rect -840 -2789 -806 -2771
rect -946 -2805 -912 -2791
rect -1042 -2839 -1008 -2827
rect -946 -2825 -912 -2805
rect -840 -2839 -806 -2827
rect -1042 -2861 -1008 -2839
rect -840 -2861 -806 -2839
rect -946 -2873 -912 -2863
rect -1042 -2907 -1008 -2899
rect -946 -2897 -912 -2873
rect -840 -2907 -806 -2899
rect -1042 -2933 -1008 -2907
rect -840 -2933 -806 -2907
rect -946 -2941 -912 -2935
rect -1042 -2975 -1008 -2971
rect -946 -2969 -912 -2941
rect -840 -2975 -806 -2971
rect -1042 -3005 -1008 -2975
rect -840 -3005 -806 -2975
rect -946 -3009 -912 -3007
rect -946 -3041 -912 -3009
rect -1042 -3077 -1008 -3043
rect -840 -3077 -806 -3043
rect -946 -3111 -912 -3079
rect -946 -3113 -912 -3111
rect -1042 -3145 -1008 -3115
rect -840 -3145 -806 -3115
rect -1042 -3149 -1008 -3145
rect -946 -3179 -912 -3151
rect -840 -3149 -806 -3145
rect -946 -3185 -912 -3179
rect -1042 -3213 -1008 -3187
rect -840 -3213 -806 -3187
rect -1042 -3221 -1008 -3213
rect -946 -3247 -912 -3223
rect -840 -3221 -806 -3213
rect -946 -3257 -912 -3247
rect -1042 -3281 -1008 -3259
rect -840 -3281 -806 -3259
rect -1042 -3293 -1008 -3281
rect -946 -3315 -912 -3295
rect -840 -3293 -806 -3281
rect -946 -3329 -912 -3315
rect -1042 -3349 -1008 -3331
rect -840 -3349 -806 -3331
rect -1042 -3365 -1008 -3349
rect -946 -3383 -912 -3367
rect -840 -3365 -806 -3349
rect -946 -3401 -912 -3383
rect -1042 -3417 -1008 -3403
rect -840 -3417 -806 -3403
rect -1042 -3437 -1008 -3417
rect -946 -3451 -912 -3439
rect -840 -3437 -806 -3417
rect -946 -3473 -912 -3451
rect -1042 -3485 -1008 -3475
rect -840 -3485 -806 -3475
rect -1042 -3509 -1008 -3485
rect -946 -3519 -912 -3511
rect -840 -3509 -806 -3485
rect -946 -3545 -912 -3519
rect -1042 -3553 -1008 -3547
rect -840 -3553 -806 -3547
rect -1042 -3581 -1008 -3553
rect -946 -3587 -912 -3583
rect -840 -3581 -806 -3553
rect -946 -3617 -912 -3587
rect -1042 -3621 -1008 -3619
rect -840 -3621 -806 -3619
rect -1042 -3653 -1008 -3621
rect -840 -3653 -806 -3621
rect -946 -3689 -912 -3655
rect -1042 -3723 -1008 -3691
rect -840 -3723 -806 -3691
rect -1042 -3725 -1008 -3723
rect -840 -3725 -806 -3723
rect -946 -3757 -912 -3727
rect -1042 -3791 -1008 -3763
rect -946 -3761 -912 -3757
rect -840 -3791 -806 -3763
rect -1042 -3797 -1008 -3791
rect -840 -3797 -806 -3791
rect -946 -3825 -912 -3799
rect -1042 -3859 -1008 -3835
rect -946 -3833 -912 -3825
rect -840 -3859 -806 -3835
rect -1042 -3869 -1008 -3859
rect -840 -3869 -806 -3859
rect -946 -3893 -912 -3871
rect -1042 -3927 -1008 -3907
rect -946 -3905 -912 -3893
rect -840 -3927 -806 -3907
rect -1042 -3941 -1008 -3927
rect -840 -3941 -806 -3927
rect -946 -3961 -912 -3943
rect -1042 -3995 -1008 -3979
rect -946 -3977 -912 -3961
rect -840 -3995 -806 -3979
rect -1042 -4013 -1008 -3995
rect -840 -4013 -806 -3995
rect -946 -4029 -912 -4015
rect -1042 -4063 -1008 -4051
rect -946 -4049 -912 -4029
rect -840 -4063 -806 -4051
rect -1042 -4085 -1008 -4063
rect -840 -4085 -806 -4063
rect -946 -4097 -912 -4087
rect -1042 -4131 -1008 -4123
rect -946 -4121 -912 -4097
rect -840 -4131 -806 -4123
rect -1042 -4157 -1008 -4131
rect -840 -4157 -806 -4131
rect -946 -4165 -912 -4159
rect -1042 -4199 -1008 -4195
rect -946 -4193 -912 -4165
rect -840 -4199 -806 -4195
rect -1042 -4229 -1008 -4199
rect -840 -4229 -806 -4199
rect -946 -4233 -912 -4231
rect -946 -4265 -912 -4233
rect -1042 -4301 -1008 -4267
rect -840 -4301 -806 -4267
rect -946 -4335 -912 -4303
rect -946 -4337 -912 -4335
rect -1042 -4369 -1008 -4339
rect -840 -4369 -806 -4339
rect -1042 -4373 -1008 -4369
rect -946 -4403 -912 -4375
rect -840 -4373 -806 -4369
rect -946 -4409 -912 -4403
rect -1042 -4437 -1008 -4411
rect -840 -4437 -806 -4411
rect -1042 -4445 -1008 -4437
rect -946 -4471 -912 -4447
rect -840 -4445 -806 -4437
rect -946 -4481 -912 -4471
rect -1042 -4505 -1008 -4483
rect -840 -4505 -806 -4483
rect -1042 -4517 -1008 -4505
rect -946 -4539 -912 -4519
rect -840 -4517 -806 -4505
rect -946 -4553 -912 -4539
rect -1042 -4573 -1008 -4555
rect -840 -4573 -806 -4555
rect -1042 -4589 -1008 -4573
rect -946 -4607 -912 -4591
rect -840 -4589 -806 -4573
rect -946 -4625 -912 -4607
rect -1042 -4641 -1008 -4627
rect -840 -4641 -806 -4627
rect -1042 -4661 -1008 -4641
rect -946 -4675 -912 -4663
rect -840 -4661 -806 -4641
rect -946 -4697 -912 -4675
rect -1042 -4709 -1008 -4699
rect -840 -4709 -806 -4699
rect -1042 -4733 -1008 -4709
rect -946 -4743 -912 -4735
rect -840 -4733 -806 -4709
rect -946 -4769 -912 -4743
rect -1042 -4777 -1008 -4771
rect -840 -4777 -806 -4771
rect -1042 -4805 -1008 -4777
rect -946 -4811 -912 -4807
rect -840 -4805 -806 -4777
rect -946 -4841 -912 -4811
rect -1042 -4845 -1008 -4843
rect -840 -4845 -806 -4843
rect -1042 -4877 -1008 -4845
rect -840 -4877 -806 -4845
rect -946 -4913 -912 -4879
rect -1042 -4947 -1008 -4915
rect -840 -4947 -806 -4915
rect -1042 -4949 -1008 -4947
rect -840 -4949 -806 -4947
rect -946 -4981 -912 -4951
rect -1528 -5021 -1422 -5015
rect -1528 -5057 -1494 -5023
rect -1042 -5015 -1008 -4987
rect -946 -4985 -912 -4981
rect -840 -5015 -806 -4987
rect -669 4981 -563 4985
rect -669 -4981 -563 4981
rect -669 -4985 -563 -4981
rect -426 4987 -392 5015
rect -330 4981 -296 4985
rect -224 4987 -190 5015
rect 286 5023 320 5057
rect 190 5015 224 5021
rect 392 5015 426 5021
rect -330 4951 -296 4981
rect -426 4947 -392 4949
rect -224 4947 -190 4949
rect -426 4915 -392 4947
rect -224 4915 -190 4947
rect -330 4879 -296 4913
rect -426 4845 -392 4877
rect -224 4845 -190 4877
rect -426 4843 -392 4845
rect -224 4843 -190 4845
rect -330 4811 -296 4841
rect -426 4777 -392 4805
rect -330 4807 -296 4811
rect -224 4777 -190 4805
rect -426 4771 -392 4777
rect -224 4771 -190 4777
rect -330 4743 -296 4769
rect -426 4709 -392 4733
rect -330 4735 -296 4743
rect -224 4709 -190 4733
rect -426 4699 -392 4709
rect -224 4699 -190 4709
rect -330 4675 -296 4697
rect -426 4641 -392 4661
rect -330 4663 -296 4675
rect -224 4641 -190 4661
rect -426 4627 -392 4641
rect -224 4627 -190 4641
rect -330 4607 -296 4625
rect -426 4573 -392 4589
rect -330 4591 -296 4607
rect -224 4573 -190 4589
rect -426 4555 -392 4573
rect -224 4555 -190 4573
rect -330 4539 -296 4553
rect -426 4505 -392 4517
rect -330 4519 -296 4539
rect -224 4505 -190 4517
rect -426 4483 -392 4505
rect -224 4483 -190 4505
rect -330 4471 -296 4481
rect -426 4437 -392 4445
rect -330 4447 -296 4471
rect -224 4437 -190 4445
rect -426 4411 -392 4437
rect -224 4411 -190 4437
rect -330 4403 -296 4409
rect -426 4369 -392 4373
rect -330 4375 -296 4403
rect -224 4369 -190 4373
rect -426 4339 -392 4369
rect -224 4339 -190 4369
rect -330 4335 -296 4337
rect -330 4303 -296 4335
rect -426 4267 -392 4301
rect -224 4267 -190 4301
rect -330 4233 -296 4265
rect -330 4231 -296 4233
rect -426 4199 -392 4229
rect -224 4199 -190 4229
rect -426 4195 -392 4199
rect -330 4165 -296 4193
rect -224 4195 -190 4199
rect -330 4159 -296 4165
rect -426 4131 -392 4157
rect -224 4131 -190 4157
rect -426 4123 -392 4131
rect -330 4097 -296 4121
rect -224 4123 -190 4131
rect -330 4087 -296 4097
rect -426 4063 -392 4085
rect -224 4063 -190 4085
rect -426 4051 -392 4063
rect -330 4029 -296 4049
rect -224 4051 -190 4063
rect -330 4015 -296 4029
rect -426 3995 -392 4013
rect -224 3995 -190 4013
rect -426 3979 -392 3995
rect -330 3961 -296 3977
rect -224 3979 -190 3995
rect -330 3943 -296 3961
rect -426 3927 -392 3941
rect -224 3927 -190 3941
rect -426 3907 -392 3927
rect -330 3893 -296 3905
rect -224 3907 -190 3927
rect -330 3871 -296 3893
rect -426 3859 -392 3869
rect -224 3859 -190 3869
rect -426 3835 -392 3859
rect -330 3825 -296 3833
rect -224 3835 -190 3859
rect -330 3799 -296 3825
rect -426 3791 -392 3797
rect -224 3791 -190 3797
rect -426 3763 -392 3791
rect -330 3757 -296 3761
rect -224 3763 -190 3791
rect -330 3727 -296 3757
rect -426 3723 -392 3725
rect -224 3723 -190 3725
rect -426 3691 -392 3723
rect -224 3691 -190 3723
rect -330 3655 -296 3689
rect -426 3621 -392 3653
rect -224 3621 -190 3653
rect -426 3619 -392 3621
rect -224 3619 -190 3621
rect -330 3587 -296 3617
rect -426 3553 -392 3581
rect -330 3583 -296 3587
rect -224 3553 -190 3581
rect -426 3547 -392 3553
rect -224 3547 -190 3553
rect -330 3519 -296 3545
rect -426 3485 -392 3509
rect -330 3511 -296 3519
rect -224 3485 -190 3509
rect -426 3475 -392 3485
rect -224 3475 -190 3485
rect -330 3451 -296 3473
rect -426 3417 -392 3437
rect -330 3439 -296 3451
rect -224 3417 -190 3437
rect -426 3403 -392 3417
rect -224 3403 -190 3417
rect -330 3383 -296 3401
rect -426 3349 -392 3365
rect -330 3367 -296 3383
rect -224 3349 -190 3365
rect -426 3331 -392 3349
rect -224 3331 -190 3349
rect -330 3315 -296 3329
rect -426 3281 -392 3293
rect -330 3295 -296 3315
rect -224 3281 -190 3293
rect -426 3259 -392 3281
rect -224 3259 -190 3281
rect -330 3247 -296 3257
rect -426 3213 -392 3221
rect -330 3223 -296 3247
rect -224 3213 -190 3221
rect -426 3187 -392 3213
rect -224 3187 -190 3213
rect -330 3179 -296 3185
rect -426 3145 -392 3149
rect -330 3151 -296 3179
rect -224 3145 -190 3149
rect -426 3115 -392 3145
rect -224 3115 -190 3145
rect -330 3111 -296 3113
rect -330 3079 -296 3111
rect -426 3043 -392 3077
rect -224 3043 -190 3077
rect -330 3009 -296 3041
rect -330 3007 -296 3009
rect -426 2975 -392 3005
rect -224 2975 -190 3005
rect -426 2971 -392 2975
rect -330 2941 -296 2969
rect -224 2971 -190 2975
rect -330 2935 -296 2941
rect -426 2907 -392 2933
rect -224 2907 -190 2933
rect -426 2899 -392 2907
rect -330 2873 -296 2897
rect -224 2899 -190 2907
rect -330 2863 -296 2873
rect -426 2839 -392 2861
rect -224 2839 -190 2861
rect -426 2827 -392 2839
rect -330 2805 -296 2825
rect -224 2827 -190 2839
rect -330 2791 -296 2805
rect -426 2771 -392 2789
rect -224 2771 -190 2789
rect -426 2755 -392 2771
rect -330 2737 -296 2753
rect -224 2755 -190 2771
rect -330 2719 -296 2737
rect -426 2703 -392 2717
rect -224 2703 -190 2717
rect -426 2683 -392 2703
rect -330 2669 -296 2681
rect -224 2683 -190 2703
rect -330 2647 -296 2669
rect -426 2635 -392 2645
rect -224 2635 -190 2645
rect -426 2611 -392 2635
rect -330 2601 -296 2609
rect -224 2611 -190 2635
rect -330 2575 -296 2601
rect -426 2567 -392 2573
rect -224 2567 -190 2573
rect -426 2539 -392 2567
rect -330 2533 -296 2537
rect -224 2539 -190 2567
rect -330 2503 -296 2533
rect -426 2499 -392 2501
rect -224 2499 -190 2501
rect -426 2467 -392 2499
rect -224 2467 -190 2499
rect -330 2431 -296 2465
rect -426 2397 -392 2429
rect -224 2397 -190 2429
rect -426 2395 -392 2397
rect -224 2395 -190 2397
rect -330 2363 -296 2393
rect -426 2329 -392 2357
rect -330 2359 -296 2363
rect -224 2329 -190 2357
rect -426 2323 -392 2329
rect -224 2323 -190 2329
rect -330 2295 -296 2321
rect -426 2261 -392 2285
rect -330 2287 -296 2295
rect -224 2261 -190 2285
rect -426 2251 -392 2261
rect -224 2251 -190 2261
rect -330 2227 -296 2249
rect -426 2193 -392 2213
rect -330 2215 -296 2227
rect -224 2193 -190 2213
rect -426 2179 -392 2193
rect -224 2179 -190 2193
rect -330 2159 -296 2177
rect -426 2125 -392 2141
rect -330 2143 -296 2159
rect -224 2125 -190 2141
rect -426 2107 -392 2125
rect -224 2107 -190 2125
rect -330 2091 -296 2105
rect -426 2057 -392 2069
rect -330 2071 -296 2091
rect -224 2057 -190 2069
rect -426 2035 -392 2057
rect -224 2035 -190 2057
rect -330 2023 -296 2033
rect -426 1989 -392 1997
rect -330 1999 -296 2023
rect -224 1989 -190 1997
rect -426 1963 -392 1989
rect -224 1963 -190 1989
rect -330 1955 -296 1961
rect -426 1921 -392 1925
rect -330 1927 -296 1955
rect -224 1921 -190 1925
rect -426 1891 -392 1921
rect -224 1891 -190 1921
rect -330 1887 -296 1889
rect -330 1855 -296 1887
rect -426 1819 -392 1853
rect -224 1819 -190 1853
rect -330 1785 -296 1817
rect -330 1783 -296 1785
rect -426 1751 -392 1781
rect -224 1751 -190 1781
rect -426 1747 -392 1751
rect -330 1717 -296 1745
rect -224 1747 -190 1751
rect -330 1711 -296 1717
rect -426 1683 -392 1709
rect -224 1683 -190 1709
rect -426 1675 -392 1683
rect -330 1649 -296 1673
rect -224 1675 -190 1683
rect -330 1639 -296 1649
rect -426 1615 -392 1637
rect -224 1615 -190 1637
rect -426 1603 -392 1615
rect -330 1581 -296 1601
rect -224 1603 -190 1615
rect -330 1567 -296 1581
rect -426 1547 -392 1565
rect -224 1547 -190 1565
rect -426 1531 -392 1547
rect -330 1513 -296 1529
rect -224 1531 -190 1547
rect -330 1495 -296 1513
rect -426 1479 -392 1493
rect -224 1479 -190 1493
rect -426 1459 -392 1479
rect -330 1445 -296 1457
rect -224 1459 -190 1479
rect -330 1423 -296 1445
rect -426 1411 -392 1421
rect -224 1411 -190 1421
rect -426 1387 -392 1411
rect -330 1377 -296 1385
rect -224 1387 -190 1411
rect -330 1351 -296 1377
rect -426 1343 -392 1349
rect -224 1343 -190 1349
rect -426 1315 -392 1343
rect -330 1309 -296 1313
rect -224 1315 -190 1343
rect -330 1279 -296 1309
rect -426 1275 -392 1277
rect -224 1275 -190 1277
rect -426 1243 -392 1275
rect -224 1243 -190 1275
rect -330 1207 -296 1241
rect -426 1173 -392 1205
rect -224 1173 -190 1205
rect -426 1171 -392 1173
rect -224 1171 -190 1173
rect -330 1139 -296 1169
rect -426 1105 -392 1133
rect -330 1135 -296 1139
rect -224 1105 -190 1133
rect -426 1099 -392 1105
rect -224 1099 -190 1105
rect -330 1071 -296 1097
rect -426 1037 -392 1061
rect -330 1063 -296 1071
rect -224 1037 -190 1061
rect -426 1027 -392 1037
rect -224 1027 -190 1037
rect -330 1003 -296 1025
rect -426 969 -392 989
rect -330 991 -296 1003
rect -224 969 -190 989
rect -426 955 -392 969
rect -224 955 -190 969
rect -330 935 -296 953
rect -426 901 -392 917
rect -330 919 -296 935
rect -224 901 -190 917
rect -426 883 -392 901
rect -224 883 -190 901
rect -330 867 -296 881
rect -426 833 -392 845
rect -330 847 -296 867
rect -224 833 -190 845
rect -426 811 -392 833
rect -224 811 -190 833
rect -330 799 -296 809
rect -426 765 -392 773
rect -330 775 -296 799
rect -224 765 -190 773
rect -426 739 -392 765
rect -224 739 -190 765
rect -330 731 -296 737
rect -426 697 -392 701
rect -330 703 -296 731
rect -224 697 -190 701
rect -426 667 -392 697
rect -224 667 -190 697
rect -330 663 -296 665
rect -330 631 -296 663
rect -426 595 -392 629
rect -224 595 -190 629
rect -330 561 -296 593
rect -330 559 -296 561
rect -426 527 -392 557
rect -224 527 -190 557
rect -426 523 -392 527
rect -330 493 -296 521
rect -224 523 -190 527
rect -330 487 -296 493
rect -426 459 -392 485
rect -224 459 -190 485
rect -426 451 -392 459
rect -330 425 -296 449
rect -224 451 -190 459
rect -330 415 -296 425
rect -426 391 -392 413
rect -224 391 -190 413
rect -426 379 -392 391
rect -330 357 -296 377
rect -224 379 -190 391
rect -330 343 -296 357
rect -426 323 -392 341
rect -224 323 -190 341
rect -426 307 -392 323
rect -330 289 -296 305
rect -224 307 -190 323
rect -330 271 -296 289
rect -426 255 -392 269
rect -224 255 -190 269
rect -426 235 -392 255
rect -330 221 -296 233
rect -224 235 -190 255
rect -330 199 -296 221
rect -426 187 -392 197
rect -224 187 -190 197
rect -426 163 -392 187
rect -330 153 -296 161
rect -224 163 -190 187
rect -330 127 -296 153
rect -426 119 -392 125
rect -224 119 -190 125
rect -426 91 -392 119
rect -330 85 -296 89
rect -224 91 -190 119
rect -330 55 -296 85
rect -426 51 -392 53
rect -224 51 -190 53
rect -426 19 -392 51
rect -224 19 -190 51
rect -330 -17 -296 17
rect -426 -51 -392 -19
rect -224 -51 -190 -19
rect -426 -53 -392 -51
rect -224 -53 -190 -51
rect -330 -85 -296 -55
rect -426 -119 -392 -91
rect -330 -89 -296 -85
rect -224 -119 -190 -91
rect -426 -125 -392 -119
rect -224 -125 -190 -119
rect -330 -153 -296 -127
rect -426 -187 -392 -163
rect -330 -161 -296 -153
rect -224 -187 -190 -163
rect -426 -197 -392 -187
rect -224 -197 -190 -187
rect -330 -221 -296 -199
rect -426 -255 -392 -235
rect -330 -233 -296 -221
rect -224 -255 -190 -235
rect -426 -269 -392 -255
rect -224 -269 -190 -255
rect -330 -289 -296 -271
rect -426 -323 -392 -307
rect -330 -305 -296 -289
rect -224 -323 -190 -307
rect -426 -341 -392 -323
rect -224 -341 -190 -323
rect -330 -357 -296 -343
rect -426 -391 -392 -379
rect -330 -377 -296 -357
rect -224 -391 -190 -379
rect -426 -413 -392 -391
rect -224 -413 -190 -391
rect -330 -425 -296 -415
rect -426 -459 -392 -451
rect -330 -449 -296 -425
rect -224 -459 -190 -451
rect -426 -485 -392 -459
rect -224 -485 -190 -459
rect -330 -493 -296 -487
rect -426 -527 -392 -523
rect -330 -521 -296 -493
rect -224 -527 -190 -523
rect -426 -557 -392 -527
rect -224 -557 -190 -527
rect -330 -561 -296 -559
rect -330 -593 -296 -561
rect -426 -629 -392 -595
rect -224 -629 -190 -595
rect -330 -663 -296 -631
rect -330 -665 -296 -663
rect -426 -697 -392 -667
rect -224 -697 -190 -667
rect -426 -701 -392 -697
rect -330 -731 -296 -703
rect -224 -701 -190 -697
rect -330 -737 -296 -731
rect -426 -765 -392 -739
rect -224 -765 -190 -739
rect -426 -773 -392 -765
rect -330 -799 -296 -775
rect -224 -773 -190 -765
rect -330 -809 -296 -799
rect -426 -833 -392 -811
rect -224 -833 -190 -811
rect -426 -845 -392 -833
rect -330 -867 -296 -847
rect -224 -845 -190 -833
rect -330 -881 -296 -867
rect -426 -901 -392 -883
rect -224 -901 -190 -883
rect -426 -917 -392 -901
rect -330 -935 -296 -919
rect -224 -917 -190 -901
rect -330 -953 -296 -935
rect -426 -969 -392 -955
rect -224 -969 -190 -955
rect -426 -989 -392 -969
rect -330 -1003 -296 -991
rect -224 -989 -190 -969
rect -330 -1025 -296 -1003
rect -426 -1037 -392 -1027
rect -224 -1037 -190 -1027
rect -426 -1061 -392 -1037
rect -330 -1071 -296 -1063
rect -224 -1061 -190 -1037
rect -330 -1097 -296 -1071
rect -426 -1105 -392 -1099
rect -224 -1105 -190 -1099
rect -426 -1133 -392 -1105
rect -330 -1139 -296 -1135
rect -224 -1133 -190 -1105
rect -330 -1169 -296 -1139
rect -426 -1173 -392 -1171
rect -224 -1173 -190 -1171
rect -426 -1205 -392 -1173
rect -224 -1205 -190 -1173
rect -330 -1241 -296 -1207
rect -426 -1275 -392 -1243
rect -224 -1275 -190 -1243
rect -426 -1277 -392 -1275
rect -224 -1277 -190 -1275
rect -330 -1309 -296 -1279
rect -426 -1343 -392 -1315
rect -330 -1313 -296 -1309
rect -224 -1343 -190 -1315
rect -426 -1349 -392 -1343
rect -224 -1349 -190 -1343
rect -330 -1377 -296 -1351
rect -426 -1411 -392 -1387
rect -330 -1385 -296 -1377
rect -224 -1411 -190 -1387
rect -426 -1421 -392 -1411
rect -224 -1421 -190 -1411
rect -330 -1445 -296 -1423
rect -426 -1479 -392 -1459
rect -330 -1457 -296 -1445
rect -224 -1479 -190 -1459
rect -426 -1493 -392 -1479
rect -224 -1493 -190 -1479
rect -330 -1513 -296 -1495
rect -426 -1547 -392 -1531
rect -330 -1529 -296 -1513
rect -224 -1547 -190 -1531
rect -426 -1565 -392 -1547
rect -224 -1565 -190 -1547
rect -330 -1581 -296 -1567
rect -426 -1615 -392 -1603
rect -330 -1601 -296 -1581
rect -224 -1615 -190 -1603
rect -426 -1637 -392 -1615
rect -224 -1637 -190 -1615
rect -330 -1649 -296 -1639
rect -426 -1683 -392 -1675
rect -330 -1673 -296 -1649
rect -224 -1683 -190 -1675
rect -426 -1709 -392 -1683
rect -224 -1709 -190 -1683
rect -330 -1717 -296 -1711
rect -426 -1751 -392 -1747
rect -330 -1745 -296 -1717
rect -224 -1751 -190 -1747
rect -426 -1781 -392 -1751
rect -224 -1781 -190 -1751
rect -330 -1785 -296 -1783
rect -330 -1817 -296 -1785
rect -426 -1853 -392 -1819
rect -224 -1853 -190 -1819
rect -330 -1887 -296 -1855
rect -330 -1889 -296 -1887
rect -426 -1921 -392 -1891
rect -224 -1921 -190 -1891
rect -426 -1925 -392 -1921
rect -330 -1955 -296 -1927
rect -224 -1925 -190 -1921
rect -330 -1961 -296 -1955
rect -426 -1989 -392 -1963
rect -224 -1989 -190 -1963
rect -426 -1997 -392 -1989
rect -330 -2023 -296 -1999
rect -224 -1997 -190 -1989
rect -330 -2033 -296 -2023
rect -426 -2057 -392 -2035
rect -224 -2057 -190 -2035
rect -426 -2069 -392 -2057
rect -330 -2091 -296 -2071
rect -224 -2069 -190 -2057
rect -330 -2105 -296 -2091
rect -426 -2125 -392 -2107
rect -224 -2125 -190 -2107
rect -426 -2141 -392 -2125
rect -330 -2159 -296 -2143
rect -224 -2141 -190 -2125
rect -330 -2177 -296 -2159
rect -426 -2193 -392 -2179
rect -224 -2193 -190 -2179
rect -426 -2213 -392 -2193
rect -330 -2227 -296 -2215
rect -224 -2213 -190 -2193
rect -330 -2249 -296 -2227
rect -426 -2261 -392 -2251
rect -224 -2261 -190 -2251
rect -426 -2285 -392 -2261
rect -330 -2295 -296 -2287
rect -224 -2285 -190 -2261
rect -330 -2321 -296 -2295
rect -426 -2329 -392 -2323
rect -224 -2329 -190 -2323
rect -426 -2357 -392 -2329
rect -330 -2363 -296 -2359
rect -224 -2357 -190 -2329
rect -330 -2393 -296 -2363
rect -426 -2397 -392 -2395
rect -224 -2397 -190 -2395
rect -426 -2429 -392 -2397
rect -224 -2429 -190 -2397
rect -330 -2465 -296 -2431
rect -426 -2499 -392 -2467
rect -224 -2499 -190 -2467
rect -426 -2501 -392 -2499
rect -224 -2501 -190 -2499
rect -330 -2533 -296 -2503
rect -426 -2567 -392 -2539
rect -330 -2537 -296 -2533
rect -224 -2567 -190 -2539
rect -426 -2573 -392 -2567
rect -224 -2573 -190 -2567
rect -330 -2601 -296 -2575
rect -426 -2635 -392 -2611
rect -330 -2609 -296 -2601
rect -224 -2635 -190 -2611
rect -426 -2645 -392 -2635
rect -224 -2645 -190 -2635
rect -330 -2669 -296 -2647
rect -426 -2703 -392 -2683
rect -330 -2681 -296 -2669
rect -224 -2703 -190 -2683
rect -426 -2717 -392 -2703
rect -224 -2717 -190 -2703
rect -330 -2737 -296 -2719
rect -426 -2771 -392 -2755
rect -330 -2753 -296 -2737
rect -224 -2771 -190 -2755
rect -426 -2789 -392 -2771
rect -224 -2789 -190 -2771
rect -330 -2805 -296 -2791
rect -426 -2839 -392 -2827
rect -330 -2825 -296 -2805
rect -224 -2839 -190 -2827
rect -426 -2861 -392 -2839
rect -224 -2861 -190 -2839
rect -330 -2873 -296 -2863
rect -426 -2907 -392 -2899
rect -330 -2897 -296 -2873
rect -224 -2907 -190 -2899
rect -426 -2933 -392 -2907
rect -224 -2933 -190 -2907
rect -330 -2941 -296 -2935
rect -426 -2975 -392 -2971
rect -330 -2969 -296 -2941
rect -224 -2975 -190 -2971
rect -426 -3005 -392 -2975
rect -224 -3005 -190 -2975
rect -330 -3009 -296 -3007
rect -330 -3041 -296 -3009
rect -426 -3077 -392 -3043
rect -224 -3077 -190 -3043
rect -330 -3111 -296 -3079
rect -330 -3113 -296 -3111
rect -426 -3145 -392 -3115
rect -224 -3145 -190 -3115
rect -426 -3149 -392 -3145
rect -330 -3179 -296 -3151
rect -224 -3149 -190 -3145
rect -330 -3185 -296 -3179
rect -426 -3213 -392 -3187
rect -224 -3213 -190 -3187
rect -426 -3221 -392 -3213
rect -330 -3247 -296 -3223
rect -224 -3221 -190 -3213
rect -330 -3257 -296 -3247
rect -426 -3281 -392 -3259
rect -224 -3281 -190 -3259
rect -426 -3293 -392 -3281
rect -330 -3315 -296 -3295
rect -224 -3293 -190 -3281
rect -330 -3329 -296 -3315
rect -426 -3349 -392 -3331
rect -224 -3349 -190 -3331
rect -426 -3365 -392 -3349
rect -330 -3383 -296 -3367
rect -224 -3365 -190 -3349
rect -330 -3401 -296 -3383
rect -426 -3417 -392 -3403
rect -224 -3417 -190 -3403
rect -426 -3437 -392 -3417
rect -330 -3451 -296 -3439
rect -224 -3437 -190 -3417
rect -330 -3473 -296 -3451
rect -426 -3485 -392 -3475
rect -224 -3485 -190 -3475
rect -426 -3509 -392 -3485
rect -330 -3519 -296 -3511
rect -224 -3509 -190 -3485
rect -330 -3545 -296 -3519
rect -426 -3553 -392 -3547
rect -224 -3553 -190 -3547
rect -426 -3581 -392 -3553
rect -330 -3587 -296 -3583
rect -224 -3581 -190 -3553
rect -330 -3617 -296 -3587
rect -426 -3621 -392 -3619
rect -224 -3621 -190 -3619
rect -426 -3653 -392 -3621
rect -224 -3653 -190 -3621
rect -330 -3689 -296 -3655
rect -426 -3723 -392 -3691
rect -224 -3723 -190 -3691
rect -426 -3725 -392 -3723
rect -224 -3725 -190 -3723
rect -330 -3757 -296 -3727
rect -426 -3791 -392 -3763
rect -330 -3761 -296 -3757
rect -224 -3791 -190 -3763
rect -426 -3797 -392 -3791
rect -224 -3797 -190 -3791
rect -330 -3825 -296 -3799
rect -426 -3859 -392 -3835
rect -330 -3833 -296 -3825
rect -224 -3859 -190 -3835
rect -426 -3869 -392 -3859
rect -224 -3869 -190 -3859
rect -330 -3893 -296 -3871
rect -426 -3927 -392 -3907
rect -330 -3905 -296 -3893
rect -224 -3927 -190 -3907
rect -426 -3941 -392 -3927
rect -224 -3941 -190 -3927
rect -330 -3961 -296 -3943
rect -426 -3995 -392 -3979
rect -330 -3977 -296 -3961
rect -224 -3995 -190 -3979
rect -426 -4013 -392 -3995
rect -224 -4013 -190 -3995
rect -330 -4029 -296 -4015
rect -426 -4063 -392 -4051
rect -330 -4049 -296 -4029
rect -224 -4063 -190 -4051
rect -426 -4085 -392 -4063
rect -224 -4085 -190 -4063
rect -330 -4097 -296 -4087
rect -426 -4131 -392 -4123
rect -330 -4121 -296 -4097
rect -224 -4131 -190 -4123
rect -426 -4157 -392 -4131
rect -224 -4157 -190 -4131
rect -330 -4165 -296 -4159
rect -426 -4199 -392 -4195
rect -330 -4193 -296 -4165
rect -224 -4199 -190 -4195
rect -426 -4229 -392 -4199
rect -224 -4229 -190 -4199
rect -330 -4233 -296 -4231
rect -330 -4265 -296 -4233
rect -426 -4301 -392 -4267
rect -224 -4301 -190 -4267
rect -330 -4335 -296 -4303
rect -330 -4337 -296 -4335
rect -426 -4369 -392 -4339
rect -224 -4369 -190 -4339
rect -426 -4373 -392 -4369
rect -330 -4403 -296 -4375
rect -224 -4373 -190 -4369
rect -330 -4409 -296 -4403
rect -426 -4437 -392 -4411
rect -224 -4437 -190 -4411
rect -426 -4445 -392 -4437
rect -330 -4471 -296 -4447
rect -224 -4445 -190 -4437
rect -330 -4481 -296 -4471
rect -426 -4505 -392 -4483
rect -224 -4505 -190 -4483
rect -426 -4517 -392 -4505
rect -330 -4539 -296 -4519
rect -224 -4517 -190 -4505
rect -330 -4553 -296 -4539
rect -426 -4573 -392 -4555
rect -224 -4573 -190 -4555
rect -426 -4589 -392 -4573
rect -330 -4607 -296 -4591
rect -224 -4589 -190 -4573
rect -330 -4625 -296 -4607
rect -426 -4641 -392 -4627
rect -224 -4641 -190 -4627
rect -426 -4661 -392 -4641
rect -330 -4675 -296 -4663
rect -224 -4661 -190 -4641
rect -330 -4697 -296 -4675
rect -426 -4709 -392 -4699
rect -224 -4709 -190 -4699
rect -426 -4733 -392 -4709
rect -330 -4743 -296 -4735
rect -224 -4733 -190 -4709
rect -330 -4769 -296 -4743
rect -426 -4777 -392 -4771
rect -224 -4777 -190 -4771
rect -426 -4805 -392 -4777
rect -330 -4811 -296 -4807
rect -224 -4805 -190 -4777
rect -330 -4841 -296 -4811
rect -426 -4845 -392 -4843
rect -224 -4845 -190 -4843
rect -426 -4877 -392 -4845
rect -224 -4877 -190 -4845
rect -330 -4913 -296 -4879
rect -426 -4947 -392 -4915
rect -224 -4947 -190 -4915
rect -426 -4949 -392 -4947
rect -224 -4949 -190 -4947
rect -330 -4981 -296 -4951
rect -1042 -5021 -1008 -5015
rect -840 -5021 -806 -5015
rect -946 -5057 -912 -5023
rect -426 -5015 -392 -4987
rect -330 -4985 -296 -4981
rect -224 -5015 -190 -4987
rect -53 4981 53 4985
rect -53 -4981 53 4981
rect -53 -4985 53 -4981
rect 190 4987 224 5015
rect 286 4981 320 4985
rect 392 4987 426 5015
rect 902 5023 936 5057
rect 806 5015 840 5021
rect 1008 5015 1042 5021
rect 286 4951 320 4981
rect 190 4947 224 4949
rect 392 4947 426 4949
rect 190 4915 224 4947
rect 392 4915 426 4947
rect 286 4879 320 4913
rect 190 4845 224 4877
rect 392 4845 426 4877
rect 190 4843 224 4845
rect 392 4843 426 4845
rect 286 4811 320 4841
rect 190 4777 224 4805
rect 286 4807 320 4811
rect 392 4777 426 4805
rect 190 4771 224 4777
rect 392 4771 426 4777
rect 286 4743 320 4769
rect 190 4709 224 4733
rect 286 4735 320 4743
rect 392 4709 426 4733
rect 190 4699 224 4709
rect 392 4699 426 4709
rect 286 4675 320 4697
rect 190 4641 224 4661
rect 286 4663 320 4675
rect 392 4641 426 4661
rect 190 4627 224 4641
rect 392 4627 426 4641
rect 286 4607 320 4625
rect 190 4573 224 4589
rect 286 4591 320 4607
rect 392 4573 426 4589
rect 190 4555 224 4573
rect 392 4555 426 4573
rect 286 4539 320 4553
rect 190 4505 224 4517
rect 286 4519 320 4539
rect 392 4505 426 4517
rect 190 4483 224 4505
rect 392 4483 426 4505
rect 286 4471 320 4481
rect 190 4437 224 4445
rect 286 4447 320 4471
rect 392 4437 426 4445
rect 190 4411 224 4437
rect 392 4411 426 4437
rect 286 4403 320 4409
rect 190 4369 224 4373
rect 286 4375 320 4403
rect 392 4369 426 4373
rect 190 4339 224 4369
rect 392 4339 426 4369
rect 286 4335 320 4337
rect 286 4303 320 4335
rect 190 4267 224 4301
rect 392 4267 426 4301
rect 286 4233 320 4265
rect 286 4231 320 4233
rect 190 4199 224 4229
rect 392 4199 426 4229
rect 190 4195 224 4199
rect 286 4165 320 4193
rect 392 4195 426 4199
rect 286 4159 320 4165
rect 190 4131 224 4157
rect 392 4131 426 4157
rect 190 4123 224 4131
rect 286 4097 320 4121
rect 392 4123 426 4131
rect 286 4087 320 4097
rect 190 4063 224 4085
rect 392 4063 426 4085
rect 190 4051 224 4063
rect 286 4029 320 4049
rect 392 4051 426 4063
rect 286 4015 320 4029
rect 190 3995 224 4013
rect 392 3995 426 4013
rect 190 3979 224 3995
rect 286 3961 320 3977
rect 392 3979 426 3995
rect 286 3943 320 3961
rect 190 3927 224 3941
rect 392 3927 426 3941
rect 190 3907 224 3927
rect 286 3893 320 3905
rect 392 3907 426 3927
rect 286 3871 320 3893
rect 190 3859 224 3869
rect 392 3859 426 3869
rect 190 3835 224 3859
rect 286 3825 320 3833
rect 392 3835 426 3859
rect 286 3799 320 3825
rect 190 3791 224 3797
rect 392 3791 426 3797
rect 190 3763 224 3791
rect 286 3757 320 3761
rect 392 3763 426 3791
rect 286 3727 320 3757
rect 190 3723 224 3725
rect 392 3723 426 3725
rect 190 3691 224 3723
rect 392 3691 426 3723
rect 286 3655 320 3689
rect 190 3621 224 3653
rect 392 3621 426 3653
rect 190 3619 224 3621
rect 392 3619 426 3621
rect 286 3587 320 3617
rect 190 3553 224 3581
rect 286 3583 320 3587
rect 392 3553 426 3581
rect 190 3547 224 3553
rect 392 3547 426 3553
rect 286 3519 320 3545
rect 190 3485 224 3509
rect 286 3511 320 3519
rect 392 3485 426 3509
rect 190 3475 224 3485
rect 392 3475 426 3485
rect 286 3451 320 3473
rect 190 3417 224 3437
rect 286 3439 320 3451
rect 392 3417 426 3437
rect 190 3403 224 3417
rect 392 3403 426 3417
rect 286 3383 320 3401
rect 190 3349 224 3365
rect 286 3367 320 3383
rect 392 3349 426 3365
rect 190 3331 224 3349
rect 392 3331 426 3349
rect 286 3315 320 3329
rect 190 3281 224 3293
rect 286 3295 320 3315
rect 392 3281 426 3293
rect 190 3259 224 3281
rect 392 3259 426 3281
rect 286 3247 320 3257
rect 190 3213 224 3221
rect 286 3223 320 3247
rect 392 3213 426 3221
rect 190 3187 224 3213
rect 392 3187 426 3213
rect 286 3179 320 3185
rect 190 3145 224 3149
rect 286 3151 320 3179
rect 392 3145 426 3149
rect 190 3115 224 3145
rect 392 3115 426 3145
rect 286 3111 320 3113
rect 286 3079 320 3111
rect 190 3043 224 3077
rect 392 3043 426 3077
rect 286 3009 320 3041
rect 286 3007 320 3009
rect 190 2975 224 3005
rect 392 2975 426 3005
rect 190 2971 224 2975
rect 286 2941 320 2969
rect 392 2971 426 2975
rect 286 2935 320 2941
rect 190 2907 224 2933
rect 392 2907 426 2933
rect 190 2899 224 2907
rect 286 2873 320 2897
rect 392 2899 426 2907
rect 286 2863 320 2873
rect 190 2839 224 2861
rect 392 2839 426 2861
rect 190 2827 224 2839
rect 286 2805 320 2825
rect 392 2827 426 2839
rect 286 2791 320 2805
rect 190 2771 224 2789
rect 392 2771 426 2789
rect 190 2755 224 2771
rect 286 2737 320 2753
rect 392 2755 426 2771
rect 286 2719 320 2737
rect 190 2703 224 2717
rect 392 2703 426 2717
rect 190 2683 224 2703
rect 286 2669 320 2681
rect 392 2683 426 2703
rect 286 2647 320 2669
rect 190 2635 224 2645
rect 392 2635 426 2645
rect 190 2611 224 2635
rect 286 2601 320 2609
rect 392 2611 426 2635
rect 286 2575 320 2601
rect 190 2567 224 2573
rect 392 2567 426 2573
rect 190 2539 224 2567
rect 286 2533 320 2537
rect 392 2539 426 2567
rect 286 2503 320 2533
rect 190 2499 224 2501
rect 392 2499 426 2501
rect 190 2467 224 2499
rect 392 2467 426 2499
rect 286 2431 320 2465
rect 190 2397 224 2429
rect 392 2397 426 2429
rect 190 2395 224 2397
rect 392 2395 426 2397
rect 286 2363 320 2393
rect 190 2329 224 2357
rect 286 2359 320 2363
rect 392 2329 426 2357
rect 190 2323 224 2329
rect 392 2323 426 2329
rect 286 2295 320 2321
rect 190 2261 224 2285
rect 286 2287 320 2295
rect 392 2261 426 2285
rect 190 2251 224 2261
rect 392 2251 426 2261
rect 286 2227 320 2249
rect 190 2193 224 2213
rect 286 2215 320 2227
rect 392 2193 426 2213
rect 190 2179 224 2193
rect 392 2179 426 2193
rect 286 2159 320 2177
rect 190 2125 224 2141
rect 286 2143 320 2159
rect 392 2125 426 2141
rect 190 2107 224 2125
rect 392 2107 426 2125
rect 286 2091 320 2105
rect 190 2057 224 2069
rect 286 2071 320 2091
rect 392 2057 426 2069
rect 190 2035 224 2057
rect 392 2035 426 2057
rect 286 2023 320 2033
rect 190 1989 224 1997
rect 286 1999 320 2023
rect 392 1989 426 1997
rect 190 1963 224 1989
rect 392 1963 426 1989
rect 286 1955 320 1961
rect 190 1921 224 1925
rect 286 1927 320 1955
rect 392 1921 426 1925
rect 190 1891 224 1921
rect 392 1891 426 1921
rect 286 1887 320 1889
rect 286 1855 320 1887
rect 190 1819 224 1853
rect 392 1819 426 1853
rect 286 1785 320 1817
rect 286 1783 320 1785
rect 190 1751 224 1781
rect 392 1751 426 1781
rect 190 1747 224 1751
rect 286 1717 320 1745
rect 392 1747 426 1751
rect 286 1711 320 1717
rect 190 1683 224 1709
rect 392 1683 426 1709
rect 190 1675 224 1683
rect 286 1649 320 1673
rect 392 1675 426 1683
rect 286 1639 320 1649
rect 190 1615 224 1637
rect 392 1615 426 1637
rect 190 1603 224 1615
rect 286 1581 320 1601
rect 392 1603 426 1615
rect 286 1567 320 1581
rect 190 1547 224 1565
rect 392 1547 426 1565
rect 190 1531 224 1547
rect 286 1513 320 1529
rect 392 1531 426 1547
rect 286 1495 320 1513
rect 190 1479 224 1493
rect 392 1479 426 1493
rect 190 1459 224 1479
rect 286 1445 320 1457
rect 392 1459 426 1479
rect 286 1423 320 1445
rect 190 1411 224 1421
rect 392 1411 426 1421
rect 190 1387 224 1411
rect 286 1377 320 1385
rect 392 1387 426 1411
rect 286 1351 320 1377
rect 190 1343 224 1349
rect 392 1343 426 1349
rect 190 1315 224 1343
rect 286 1309 320 1313
rect 392 1315 426 1343
rect 286 1279 320 1309
rect 190 1275 224 1277
rect 392 1275 426 1277
rect 190 1243 224 1275
rect 392 1243 426 1275
rect 286 1207 320 1241
rect 190 1173 224 1205
rect 392 1173 426 1205
rect 190 1171 224 1173
rect 392 1171 426 1173
rect 286 1139 320 1169
rect 190 1105 224 1133
rect 286 1135 320 1139
rect 392 1105 426 1133
rect 190 1099 224 1105
rect 392 1099 426 1105
rect 286 1071 320 1097
rect 190 1037 224 1061
rect 286 1063 320 1071
rect 392 1037 426 1061
rect 190 1027 224 1037
rect 392 1027 426 1037
rect 286 1003 320 1025
rect 190 969 224 989
rect 286 991 320 1003
rect 392 969 426 989
rect 190 955 224 969
rect 392 955 426 969
rect 286 935 320 953
rect 190 901 224 917
rect 286 919 320 935
rect 392 901 426 917
rect 190 883 224 901
rect 392 883 426 901
rect 286 867 320 881
rect 190 833 224 845
rect 286 847 320 867
rect 392 833 426 845
rect 190 811 224 833
rect 392 811 426 833
rect 286 799 320 809
rect 190 765 224 773
rect 286 775 320 799
rect 392 765 426 773
rect 190 739 224 765
rect 392 739 426 765
rect 286 731 320 737
rect 190 697 224 701
rect 286 703 320 731
rect 392 697 426 701
rect 190 667 224 697
rect 392 667 426 697
rect 286 663 320 665
rect 286 631 320 663
rect 190 595 224 629
rect 392 595 426 629
rect 286 561 320 593
rect 286 559 320 561
rect 190 527 224 557
rect 392 527 426 557
rect 190 523 224 527
rect 286 493 320 521
rect 392 523 426 527
rect 286 487 320 493
rect 190 459 224 485
rect 392 459 426 485
rect 190 451 224 459
rect 286 425 320 449
rect 392 451 426 459
rect 286 415 320 425
rect 190 391 224 413
rect 392 391 426 413
rect 190 379 224 391
rect 286 357 320 377
rect 392 379 426 391
rect 286 343 320 357
rect 190 323 224 341
rect 392 323 426 341
rect 190 307 224 323
rect 286 289 320 305
rect 392 307 426 323
rect 286 271 320 289
rect 190 255 224 269
rect 392 255 426 269
rect 190 235 224 255
rect 286 221 320 233
rect 392 235 426 255
rect 286 199 320 221
rect 190 187 224 197
rect 392 187 426 197
rect 190 163 224 187
rect 286 153 320 161
rect 392 163 426 187
rect 286 127 320 153
rect 190 119 224 125
rect 392 119 426 125
rect 190 91 224 119
rect 286 85 320 89
rect 392 91 426 119
rect 286 55 320 85
rect 190 51 224 53
rect 392 51 426 53
rect 190 19 224 51
rect 392 19 426 51
rect 286 -17 320 17
rect 190 -51 224 -19
rect 392 -51 426 -19
rect 190 -53 224 -51
rect 392 -53 426 -51
rect 286 -85 320 -55
rect 190 -119 224 -91
rect 286 -89 320 -85
rect 392 -119 426 -91
rect 190 -125 224 -119
rect 392 -125 426 -119
rect 286 -153 320 -127
rect 190 -187 224 -163
rect 286 -161 320 -153
rect 392 -187 426 -163
rect 190 -197 224 -187
rect 392 -197 426 -187
rect 286 -221 320 -199
rect 190 -255 224 -235
rect 286 -233 320 -221
rect 392 -255 426 -235
rect 190 -269 224 -255
rect 392 -269 426 -255
rect 286 -289 320 -271
rect 190 -323 224 -307
rect 286 -305 320 -289
rect 392 -323 426 -307
rect 190 -341 224 -323
rect 392 -341 426 -323
rect 286 -357 320 -343
rect 190 -391 224 -379
rect 286 -377 320 -357
rect 392 -391 426 -379
rect 190 -413 224 -391
rect 392 -413 426 -391
rect 286 -425 320 -415
rect 190 -459 224 -451
rect 286 -449 320 -425
rect 392 -459 426 -451
rect 190 -485 224 -459
rect 392 -485 426 -459
rect 286 -493 320 -487
rect 190 -527 224 -523
rect 286 -521 320 -493
rect 392 -527 426 -523
rect 190 -557 224 -527
rect 392 -557 426 -527
rect 286 -561 320 -559
rect 286 -593 320 -561
rect 190 -629 224 -595
rect 392 -629 426 -595
rect 286 -663 320 -631
rect 286 -665 320 -663
rect 190 -697 224 -667
rect 392 -697 426 -667
rect 190 -701 224 -697
rect 286 -731 320 -703
rect 392 -701 426 -697
rect 286 -737 320 -731
rect 190 -765 224 -739
rect 392 -765 426 -739
rect 190 -773 224 -765
rect 286 -799 320 -775
rect 392 -773 426 -765
rect 286 -809 320 -799
rect 190 -833 224 -811
rect 392 -833 426 -811
rect 190 -845 224 -833
rect 286 -867 320 -847
rect 392 -845 426 -833
rect 286 -881 320 -867
rect 190 -901 224 -883
rect 392 -901 426 -883
rect 190 -917 224 -901
rect 286 -935 320 -919
rect 392 -917 426 -901
rect 286 -953 320 -935
rect 190 -969 224 -955
rect 392 -969 426 -955
rect 190 -989 224 -969
rect 286 -1003 320 -991
rect 392 -989 426 -969
rect 286 -1025 320 -1003
rect 190 -1037 224 -1027
rect 392 -1037 426 -1027
rect 190 -1061 224 -1037
rect 286 -1071 320 -1063
rect 392 -1061 426 -1037
rect 286 -1097 320 -1071
rect 190 -1105 224 -1099
rect 392 -1105 426 -1099
rect 190 -1133 224 -1105
rect 286 -1139 320 -1135
rect 392 -1133 426 -1105
rect 286 -1169 320 -1139
rect 190 -1173 224 -1171
rect 392 -1173 426 -1171
rect 190 -1205 224 -1173
rect 392 -1205 426 -1173
rect 286 -1241 320 -1207
rect 190 -1275 224 -1243
rect 392 -1275 426 -1243
rect 190 -1277 224 -1275
rect 392 -1277 426 -1275
rect 286 -1309 320 -1279
rect 190 -1343 224 -1315
rect 286 -1313 320 -1309
rect 392 -1343 426 -1315
rect 190 -1349 224 -1343
rect 392 -1349 426 -1343
rect 286 -1377 320 -1351
rect 190 -1411 224 -1387
rect 286 -1385 320 -1377
rect 392 -1411 426 -1387
rect 190 -1421 224 -1411
rect 392 -1421 426 -1411
rect 286 -1445 320 -1423
rect 190 -1479 224 -1459
rect 286 -1457 320 -1445
rect 392 -1479 426 -1459
rect 190 -1493 224 -1479
rect 392 -1493 426 -1479
rect 286 -1513 320 -1495
rect 190 -1547 224 -1531
rect 286 -1529 320 -1513
rect 392 -1547 426 -1531
rect 190 -1565 224 -1547
rect 392 -1565 426 -1547
rect 286 -1581 320 -1567
rect 190 -1615 224 -1603
rect 286 -1601 320 -1581
rect 392 -1615 426 -1603
rect 190 -1637 224 -1615
rect 392 -1637 426 -1615
rect 286 -1649 320 -1639
rect 190 -1683 224 -1675
rect 286 -1673 320 -1649
rect 392 -1683 426 -1675
rect 190 -1709 224 -1683
rect 392 -1709 426 -1683
rect 286 -1717 320 -1711
rect 190 -1751 224 -1747
rect 286 -1745 320 -1717
rect 392 -1751 426 -1747
rect 190 -1781 224 -1751
rect 392 -1781 426 -1751
rect 286 -1785 320 -1783
rect 286 -1817 320 -1785
rect 190 -1853 224 -1819
rect 392 -1853 426 -1819
rect 286 -1887 320 -1855
rect 286 -1889 320 -1887
rect 190 -1921 224 -1891
rect 392 -1921 426 -1891
rect 190 -1925 224 -1921
rect 286 -1955 320 -1927
rect 392 -1925 426 -1921
rect 286 -1961 320 -1955
rect 190 -1989 224 -1963
rect 392 -1989 426 -1963
rect 190 -1997 224 -1989
rect 286 -2023 320 -1999
rect 392 -1997 426 -1989
rect 286 -2033 320 -2023
rect 190 -2057 224 -2035
rect 392 -2057 426 -2035
rect 190 -2069 224 -2057
rect 286 -2091 320 -2071
rect 392 -2069 426 -2057
rect 286 -2105 320 -2091
rect 190 -2125 224 -2107
rect 392 -2125 426 -2107
rect 190 -2141 224 -2125
rect 286 -2159 320 -2143
rect 392 -2141 426 -2125
rect 286 -2177 320 -2159
rect 190 -2193 224 -2179
rect 392 -2193 426 -2179
rect 190 -2213 224 -2193
rect 286 -2227 320 -2215
rect 392 -2213 426 -2193
rect 286 -2249 320 -2227
rect 190 -2261 224 -2251
rect 392 -2261 426 -2251
rect 190 -2285 224 -2261
rect 286 -2295 320 -2287
rect 392 -2285 426 -2261
rect 286 -2321 320 -2295
rect 190 -2329 224 -2323
rect 392 -2329 426 -2323
rect 190 -2357 224 -2329
rect 286 -2363 320 -2359
rect 392 -2357 426 -2329
rect 286 -2393 320 -2363
rect 190 -2397 224 -2395
rect 392 -2397 426 -2395
rect 190 -2429 224 -2397
rect 392 -2429 426 -2397
rect 286 -2465 320 -2431
rect 190 -2499 224 -2467
rect 392 -2499 426 -2467
rect 190 -2501 224 -2499
rect 392 -2501 426 -2499
rect 286 -2533 320 -2503
rect 190 -2567 224 -2539
rect 286 -2537 320 -2533
rect 392 -2567 426 -2539
rect 190 -2573 224 -2567
rect 392 -2573 426 -2567
rect 286 -2601 320 -2575
rect 190 -2635 224 -2611
rect 286 -2609 320 -2601
rect 392 -2635 426 -2611
rect 190 -2645 224 -2635
rect 392 -2645 426 -2635
rect 286 -2669 320 -2647
rect 190 -2703 224 -2683
rect 286 -2681 320 -2669
rect 392 -2703 426 -2683
rect 190 -2717 224 -2703
rect 392 -2717 426 -2703
rect 286 -2737 320 -2719
rect 190 -2771 224 -2755
rect 286 -2753 320 -2737
rect 392 -2771 426 -2755
rect 190 -2789 224 -2771
rect 392 -2789 426 -2771
rect 286 -2805 320 -2791
rect 190 -2839 224 -2827
rect 286 -2825 320 -2805
rect 392 -2839 426 -2827
rect 190 -2861 224 -2839
rect 392 -2861 426 -2839
rect 286 -2873 320 -2863
rect 190 -2907 224 -2899
rect 286 -2897 320 -2873
rect 392 -2907 426 -2899
rect 190 -2933 224 -2907
rect 392 -2933 426 -2907
rect 286 -2941 320 -2935
rect 190 -2975 224 -2971
rect 286 -2969 320 -2941
rect 392 -2975 426 -2971
rect 190 -3005 224 -2975
rect 392 -3005 426 -2975
rect 286 -3009 320 -3007
rect 286 -3041 320 -3009
rect 190 -3077 224 -3043
rect 392 -3077 426 -3043
rect 286 -3111 320 -3079
rect 286 -3113 320 -3111
rect 190 -3145 224 -3115
rect 392 -3145 426 -3115
rect 190 -3149 224 -3145
rect 286 -3179 320 -3151
rect 392 -3149 426 -3145
rect 286 -3185 320 -3179
rect 190 -3213 224 -3187
rect 392 -3213 426 -3187
rect 190 -3221 224 -3213
rect 286 -3247 320 -3223
rect 392 -3221 426 -3213
rect 286 -3257 320 -3247
rect 190 -3281 224 -3259
rect 392 -3281 426 -3259
rect 190 -3293 224 -3281
rect 286 -3315 320 -3295
rect 392 -3293 426 -3281
rect 286 -3329 320 -3315
rect 190 -3349 224 -3331
rect 392 -3349 426 -3331
rect 190 -3365 224 -3349
rect 286 -3383 320 -3367
rect 392 -3365 426 -3349
rect 286 -3401 320 -3383
rect 190 -3417 224 -3403
rect 392 -3417 426 -3403
rect 190 -3437 224 -3417
rect 286 -3451 320 -3439
rect 392 -3437 426 -3417
rect 286 -3473 320 -3451
rect 190 -3485 224 -3475
rect 392 -3485 426 -3475
rect 190 -3509 224 -3485
rect 286 -3519 320 -3511
rect 392 -3509 426 -3485
rect 286 -3545 320 -3519
rect 190 -3553 224 -3547
rect 392 -3553 426 -3547
rect 190 -3581 224 -3553
rect 286 -3587 320 -3583
rect 392 -3581 426 -3553
rect 286 -3617 320 -3587
rect 190 -3621 224 -3619
rect 392 -3621 426 -3619
rect 190 -3653 224 -3621
rect 392 -3653 426 -3621
rect 286 -3689 320 -3655
rect 190 -3723 224 -3691
rect 392 -3723 426 -3691
rect 190 -3725 224 -3723
rect 392 -3725 426 -3723
rect 286 -3757 320 -3727
rect 190 -3791 224 -3763
rect 286 -3761 320 -3757
rect 392 -3791 426 -3763
rect 190 -3797 224 -3791
rect 392 -3797 426 -3791
rect 286 -3825 320 -3799
rect 190 -3859 224 -3835
rect 286 -3833 320 -3825
rect 392 -3859 426 -3835
rect 190 -3869 224 -3859
rect 392 -3869 426 -3859
rect 286 -3893 320 -3871
rect 190 -3927 224 -3907
rect 286 -3905 320 -3893
rect 392 -3927 426 -3907
rect 190 -3941 224 -3927
rect 392 -3941 426 -3927
rect 286 -3961 320 -3943
rect 190 -3995 224 -3979
rect 286 -3977 320 -3961
rect 392 -3995 426 -3979
rect 190 -4013 224 -3995
rect 392 -4013 426 -3995
rect 286 -4029 320 -4015
rect 190 -4063 224 -4051
rect 286 -4049 320 -4029
rect 392 -4063 426 -4051
rect 190 -4085 224 -4063
rect 392 -4085 426 -4063
rect 286 -4097 320 -4087
rect 190 -4131 224 -4123
rect 286 -4121 320 -4097
rect 392 -4131 426 -4123
rect 190 -4157 224 -4131
rect 392 -4157 426 -4131
rect 286 -4165 320 -4159
rect 190 -4199 224 -4195
rect 286 -4193 320 -4165
rect 392 -4199 426 -4195
rect 190 -4229 224 -4199
rect 392 -4229 426 -4199
rect 286 -4233 320 -4231
rect 286 -4265 320 -4233
rect 190 -4301 224 -4267
rect 392 -4301 426 -4267
rect 286 -4335 320 -4303
rect 286 -4337 320 -4335
rect 190 -4369 224 -4339
rect 392 -4369 426 -4339
rect 190 -4373 224 -4369
rect 286 -4403 320 -4375
rect 392 -4373 426 -4369
rect 286 -4409 320 -4403
rect 190 -4437 224 -4411
rect 392 -4437 426 -4411
rect 190 -4445 224 -4437
rect 286 -4471 320 -4447
rect 392 -4445 426 -4437
rect 286 -4481 320 -4471
rect 190 -4505 224 -4483
rect 392 -4505 426 -4483
rect 190 -4517 224 -4505
rect 286 -4539 320 -4519
rect 392 -4517 426 -4505
rect 286 -4553 320 -4539
rect 190 -4573 224 -4555
rect 392 -4573 426 -4555
rect 190 -4589 224 -4573
rect 286 -4607 320 -4591
rect 392 -4589 426 -4573
rect 286 -4625 320 -4607
rect 190 -4641 224 -4627
rect 392 -4641 426 -4627
rect 190 -4661 224 -4641
rect 286 -4675 320 -4663
rect 392 -4661 426 -4641
rect 286 -4697 320 -4675
rect 190 -4709 224 -4699
rect 392 -4709 426 -4699
rect 190 -4733 224 -4709
rect 286 -4743 320 -4735
rect 392 -4733 426 -4709
rect 286 -4769 320 -4743
rect 190 -4777 224 -4771
rect 392 -4777 426 -4771
rect 190 -4805 224 -4777
rect 286 -4811 320 -4807
rect 392 -4805 426 -4777
rect 286 -4841 320 -4811
rect 190 -4845 224 -4843
rect 392 -4845 426 -4843
rect 190 -4877 224 -4845
rect 392 -4877 426 -4845
rect 286 -4913 320 -4879
rect 190 -4947 224 -4915
rect 392 -4947 426 -4915
rect 190 -4949 224 -4947
rect 392 -4949 426 -4947
rect 286 -4981 320 -4951
rect -426 -5021 -392 -5015
rect -224 -5021 -190 -5015
rect -330 -5057 -296 -5023
rect 190 -5015 224 -4987
rect 286 -4985 320 -4981
rect 392 -5015 426 -4987
rect 563 4981 669 4985
rect 563 -4981 669 4981
rect 563 -4985 669 -4981
rect 806 4987 840 5015
rect 902 4981 936 4985
rect 1008 4987 1042 5015
rect 1494 5023 1528 5057
rect 1422 5015 1528 5021
rect 902 4951 936 4981
rect 806 4947 840 4949
rect 1008 4947 1042 4949
rect 806 4915 840 4947
rect 1008 4915 1042 4947
rect 902 4879 936 4913
rect 806 4845 840 4877
rect 1008 4845 1042 4877
rect 806 4843 840 4845
rect 1008 4843 1042 4845
rect 902 4811 936 4841
rect 806 4777 840 4805
rect 902 4807 936 4811
rect 1008 4777 1042 4805
rect 806 4771 840 4777
rect 1008 4771 1042 4777
rect 902 4743 936 4769
rect 806 4709 840 4733
rect 902 4735 936 4743
rect 1008 4709 1042 4733
rect 806 4699 840 4709
rect 1008 4699 1042 4709
rect 902 4675 936 4697
rect 806 4641 840 4661
rect 902 4663 936 4675
rect 1008 4641 1042 4661
rect 806 4627 840 4641
rect 1008 4627 1042 4641
rect 902 4607 936 4625
rect 806 4573 840 4589
rect 902 4591 936 4607
rect 1008 4573 1042 4589
rect 806 4555 840 4573
rect 1008 4555 1042 4573
rect 902 4539 936 4553
rect 806 4505 840 4517
rect 902 4519 936 4539
rect 1008 4505 1042 4517
rect 806 4483 840 4505
rect 1008 4483 1042 4505
rect 902 4471 936 4481
rect 806 4437 840 4445
rect 902 4447 936 4471
rect 1008 4437 1042 4445
rect 806 4411 840 4437
rect 1008 4411 1042 4437
rect 902 4403 936 4409
rect 806 4369 840 4373
rect 902 4375 936 4403
rect 1008 4369 1042 4373
rect 806 4339 840 4369
rect 1008 4339 1042 4369
rect 902 4335 936 4337
rect 902 4303 936 4335
rect 806 4267 840 4301
rect 1008 4267 1042 4301
rect 902 4233 936 4265
rect 902 4231 936 4233
rect 806 4199 840 4229
rect 1008 4199 1042 4229
rect 806 4195 840 4199
rect 902 4165 936 4193
rect 1008 4195 1042 4199
rect 902 4159 936 4165
rect 806 4131 840 4157
rect 1008 4131 1042 4157
rect 806 4123 840 4131
rect 902 4097 936 4121
rect 1008 4123 1042 4131
rect 902 4087 936 4097
rect 806 4063 840 4085
rect 1008 4063 1042 4085
rect 806 4051 840 4063
rect 902 4029 936 4049
rect 1008 4051 1042 4063
rect 902 4015 936 4029
rect 806 3995 840 4013
rect 1008 3995 1042 4013
rect 806 3979 840 3995
rect 902 3961 936 3977
rect 1008 3979 1042 3995
rect 902 3943 936 3961
rect 806 3927 840 3941
rect 1008 3927 1042 3941
rect 806 3907 840 3927
rect 902 3893 936 3905
rect 1008 3907 1042 3927
rect 902 3871 936 3893
rect 806 3859 840 3869
rect 1008 3859 1042 3869
rect 806 3835 840 3859
rect 902 3825 936 3833
rect 1008 3835 1042 3859
rect 902 3799 936 3825
rect 806 3791 840 3797
rect 1008 3791 1042 3797
rect 806 3763 840 3791
rect 902 3757 936 3761
rect 1008 3763 1042 3791
rect 902 3727 936 3757
rect 806 3723 840 3725
rect 1008 3723 1042 3725
rect 806 3691 840 3723
rect 1008 3691 1042 3723
rect 902 3655 936 3689
rect 806 3621 840 3653
rect 1008 3621 1042 3653
rect 806 3619 840 3621
rect 1008 3619 1042 3621
rect 902 3587 936 3617
rect 806 3553 840 3581
rect 902 3583 936 3587
rect 1008 3553 1042 3581
rect 806 3547 840 3553
rect 1008 3547 1042 3553
rect 902 3519 936 3545
rect 806 3485 840 3509
rect 902 3511 936 3519
rect 1008 3485 1042 3509
rect 806 3475 840 3485
rect 1008 3475 1042 3485
rect 902 3451 936 3473
rect 806 3417 840 3437
rect 902 3439 936 3451
rect 1008 3417 1042 3437
rect 806 3403 840 3417
rect 1008 3403 1042 3417
rect 902 3383 936 3401
rect 806 3349 840 3365
rect 902 3367 936 3383
rect 1008 3349 1042 3365
rect 806 3331 840 3349
rect 1008 3331 1042 3349
rect 902 3315 936 3329
rect 806 3281 840 3293
rect 902 3295 936 3315
rect 1008 3281 1042 3293
rect 806 3259 840 3281
rect 1008 3259 1042 3281
rect 902 3247 936 3257
rect 806 3213 840 3221
rect 902 3223 936 3247
rect 1008 3213 1042 3221
rect 806 3187 840 3213
rect 1008 3187 1042 3213
rect 902 3179 936 3185
rect 806 3145 840 3149
rect 902 3151 936 3179
rect 1008 3145 1042 3149
rect 806 3115 840 3145
rect 1008 3115 1042 3145
rect 902 3111 936 3113
rect 902 3079 936 3111
rect 806 3043 840 3077
rect 1008 3043 1042 3077
rect 902 3009 936 3041
rect 902 3007 936 3009
rect 806 2975 840 3005
rect 1008 2975 1042 3005
rect 806 2971 840 2975
rect 902 2941 936 2969
rect 1008 2971 1042 2975
rect 902 2935 936 2941
rect 806 2907 840 2933
rect 1008 2907 1042 2933
rect 806 2899 840 2907
rect 902 2873 936 2897
rect 1008 2899 1042 2907
rect 902 2863 936 2873
rect 806 2839 840 2861
rect 1008 2839 1042 2861
rect 806 2827 840 2839
rect 902 2805 936 2825
rect 1008 2827 1042 2839
rect 902 2791 936 2805
rect 806 2771 840 2789
rect 1008 2771 1042 2789
rect 806 2755 840 2771
rect 902 2737 936 2753
rect 1008 2755 1042 2771
rect 902 2719 936 2737
rect 806 2703 840 2717
rect 1008 2703 1042 2717
rect 806 2683 840 2703
rect 902 2669 936 2681
rect 1008 2683 1042 2703
rect 902 2647 936 2669
rect 806 2635 840 2645
rect 1008 2635 1042 2645
rect 806 2611 840 2635
rect 902 2601 936 2609
rect 1008 2611 1042 2635
rect 902 2575 936 2601
rect 806 2567 840 2573
rect 1008 2567 1042 2573
rect 806 2539 840 2567
rect 902 2533 936 2537
rect 1008 2539 1042 2567
rect 902 2503 936 2533
rect 806 2499 840 2501
rect 1008 2499 1042 2501
rect 806 2467 840 2499
rect 1008 2467 1042 2499
rect 902 2431 936 2465
rect 806 2397 840 2429
rect 1008 2397 1042 2429
rect 806 2395 840 2397
rect 1008 2395 1042 2397
rect 902 2363 936 2393
rect 806 2329 840 2357
rect 902 2359 936 2363
rect 1008 2329 1042 2357
rect 806 2323 840 2329
rect 1008 2323 1042 2329
rect 902 2295 936 2321
rect 806 2261 840 2285
rect 902 2287 936 2295
rect 1008 2261 1042 2285
rect 806 2251 840 2261
rect 1008 2251 1042 2261
rect 902 2227 936 2249
rect 806 2193 840 2213
rect 902 2215 936 2227
rect 1008 2193 1042 2213
rect 806 2179 840 2193
rect 1008 2179 1042 2193
rect 902 2159 936 2177
rect 806 2125 840 2141
rect 902 2143 936 2159
rect 1008 2125 1042 2141
rect 806 2107 840 2125
rect 1008 2107 1042 2125
rect 902 2091 936 2105
rect 806 2057 840 2069
rect 902 2071 936 2091
rect 1008 2057 1042 2069
rect 806 2035 840 2057
rect 1008 2035 1042 2057
rect 902 2023 936 2033
rect 806 1989 840 1997
rect 902 1999 936 2023
rect 1008 1989 1042 1997
rect 806 1963 840 1989
rect 1008 1963 1042 1989
rect 902 1955 936 1961
rect 806 1921 840 1925
rect 902 1927 936 1955
rect 1008 1921 1042 1925
rect 806 1891 840 1921
rect 1008 1891 1042 1921
rect 902 1887 936 1889
rect 902 1855 936 1887
rect 806 1819 840 1853
rect 1008 1819 1042 1853
rect 902 1785 936 1817
rect 902 1783 936 1785
rect 806 1751 840 1781
rect 1008 1751 1042 1781
rect 806 1747 840 1751
rect 902 1717 936 1745
rect 1008 1747 1042 1751
rect 902 1711 936 1717
rect 806 1683 840 1709
rect 1008 1683 1042 1709
rect 806 1675 840 1683
rect 902 1649 936 1673
rect 1008 1675 1042 1683
rect 902 1639 936 1649
rect 806 1615 840 1637
rect 1008 1615 1042 1637
rect 806 1603 840 1615
rect 902 1581 936 1601
rect 1008 1603 1042 1615
rect 902 1567 936 1581
rect 806 1547 840 1565
rect 1008 1547 1042 1565
rect 806 1531 840 1547
rect 902 1513 936 1529
rect 1008 1531 1042 1547
rect 902 1495 936 1513
rect 806 1479 840 1493
rect 1008 1479 1042 1493
rect 806 1459 840 1479
rect 902 1445 936 1457
rect 1008 1459 1042 1479
rect 902 1423 936 1445
rect 806 1411 840 1421
rect 1008 1411 1042 1421
rect 806 1387 840 1411
rect 902 1377 936 1385
rect 1008 1387 1042 1411
rect 902 1351 936 1377
rect 806 1343 840 1349
rect 1008 1343 1042 1349
rect 806 1315 840 1343
rect 902 1309 936 1313
rect 1008 1315 1042 1343
rect 902 1279 936 1309
rect 806 1275 840 1277
rect 1008 1275 1042 1277
rect 806 1243 840 1275
rect 1008 1243 1042 1275
rect 902 1207 936 1241
rect 806 1173 840 1205
rect 1008 1173 1042 1205
rect 806 1171 840 1173
rect 1008 1171 1042 1173
rect 902 1139 936 1169
rect 806 1105 840 1133
rect 902 1135 936 1139
rect 1008 1105 1042 1133
rect 806 1099 840 1105
rect 1008 1099 1042 1105
rect 902 1071 936 1097
rect 806 1037 840 1061
rect 902 1063 936 1071
rect 1008 1037 1042 1061
rect 806 1027 840 1037
rect 1008 1027 1042 1037
rect 902 1003 936 1025
rect 806 969 840 989
rect 902 991 936 1003
rect 1008 969 1042 989
rect 806 955 840 969
rect 1008 955 1042 969
rect 902 935 936 953
rect 806 901 840 917
rect 902 919 936 935
rect 1008 901 1042 917
rect 806 883 840 901
rect 1008 883 1042 901
rect 902 867 936 881
rect 806 833 840 845
rect 902 847 936 867
rect 1008 833 1042 845
rect 806 811 840 833
rect 1008 811 1042 833
rect 902 799 936 809
rect 806 765 840 773
rect 902 775 936 799
rect 1008 765 1042 773
rect 806 739 840 765
rect 1008 739 1042 765
rect 902 731 936 737
rect 806 697 840 701
rect 902 703 936 731
rect 1008 697 1042 701
rect 806 667 840 697
rect 1008 667 1042 697
rect 902 663 936 665
rect 902 631 936 663
rect 806 595 840 629
rect 1008 595 1042 629
rect 902 561 936 593
rect 902 559 936 561
rect 806 527 840 557
rect 1008 527 1042 557
rect 806 523 840 527
rect 902 493 936 521
rect 1008 523 1042 527
rect 902 487 936 493
rect 806 459 840 485
rect 1008 459 1042 485
rect 806 451 840 459
rect 902 425 936 449
rect 1008 451 1042 459
rect 902 415 936 425
rect 806 391 840 413
rect 1008 391 1042 413
rect 806 379 840 391
rect 902 357 936 377
rect 1008 379 1042 391
rect 902 343 936 357
rect 806 323 840 341
rect 1008 323 1042 341
rect 806 307 840 323
rect 902 289 936 305
rect 1008 307 1042 323
rect 902 271 936 289
rect 806 255 840 269
rect 1008 255 1042 269
rect 806 235 840 255
rect 902 221 936 233
rect 1008 235 1042 255
rect 902 199 936 221
rect 806 187 840 197
rect 1008 187 1042 197
rect 806 163 840 187
rect 902 153 936 161
rect 1008 163 1042 187
rect 902 127 936 153
rect 806 119 840 125
rect 1008 119 1042 125
rect 806 91 840 119
rect 902 85 936 89
rect 1008 91 1042 119
rect 902 55 936 85
rect 806 51 840 53
rect 1008 51 1042 53
rect 806 19 840 51
rect 1008 19 1042 51
rect 902 -17 936 17
rect 806 -51 840 -19
rect 1008 -51 1042 -19
rect 806 -53 840 -51
rect 1008 -53 1042 -51
rect 902 -85 936 -55
rect 806 -119 840 -91
rect 902 -89 936 -85
rect 1008 -119 1042 -91
rect 806 -125 840 -119
rect 1008 -125 1042 -119
rect 902 -153 936 -127
rect 806 -187 840 -163
rect 902 -161 936 -153
rect 1008 -187 1042 -163
rect 806 -197 840 -187
rect 1008 -197 1042 -187
rect 902 -221 936 -199
rect 806 -255 840 -235
rect 902 -233 936 -221
rect 1008 -255 1042 -235
rect 806 -269 840 -255
rect 1008 -269 1042 -255
rect 902 -289 936 -271
rect 806 -323 840 -307
rect 902 -305 936 -289
rect 1008 -323 1042 -307
rect 806 -341 840 -323
rect 1008 -341 1042 -323
rect 902 -357 936 -343
rect 806 -391 840 -379
rect 902 -377 936 -357
rect 1008 -391 1042 -379
rect 806 -413 840 -391
rect 1008 -413 1042 -391
rect 902 -425 936 -415
rect 806 -459 840 -451
rect 902 -449 936 -425
rect 1008 -459 1042 -451
rect 806 -485 840 -459
rect 1008 -485 1042 -459
rect 902 -493 936 -487
rect 806 -527 840 -523
rect 902 -521 936 -493
rect 1008 -527 1042 -523
rect 806 -557 840 -527
rect 1008 -557 1042 -527
rect 902 -561 936 -559
rect 902 -593 936 -561
rect 806 -629 840 -595
rect 1008 -629 1042 -595
rect 902 -663 936 -631
rect 902 -665 936 -663
rect 806 -697 840 -667
rect 1008 -697 1042 -667
rect 806 -701 840 -697
rect 902 -731 936 -703
rect 1008 -701 1042 -697
rect 902 -737 936 -731
rect 806 -765 840 -739
rect 1008 -765 1042 -739
rect 806 -773 840 -765
rect 902 -799 936 -775
rect 1008 -773 1042 -765
rect 902 -809 936 -799
rect 806 -833 840 -811
rect 1008 -833 1042 -811
rect 806 -845 840 -833
rect 902 -867 936 -847
rect 1008 -845 1042 -833
rect 902 -881 936 -867
rect 806 -901 840 -883
rect 1008 -901 1042 -883
rect 806 -917 840 -901
rect 902 -935 936 -919
rect 1008 -917 1042 -901
rect 902 -953 936 -935
rect 806 -969 840 -955
rect 1008 -969 1042 -955
rect 806 -989 840 -969
rect 902 -1003 936 -991
rect 1008 -989 1042 -969
rect 902 -1025 936 -1003
rect 806 -1037 840 -1027
rect 1008 -1037 1042 -1027
rect 806 -1061 840 -1037
rect 902 -1071 936 -1063
rect 1008 -1061 1042 -1037
rect 902 -1097 936 -1071
rect 806 -1105 840 -1099
rect 1008 -1105 1042 -1099
rect 806 -1133 840 -1105
rect 902 -1139 936 -1135
rect 1008 -1133 1042 -1105
rect 902 -1169 936 -1139
rect 806 -1173 840 -1171
rect 1008 -1173 1042 -1171
rect 806 -1205 840 -1173
rect 1008 -1205 1042 -1173
rect 902 -1241 936 -1207
rect 806 -1275 840 -1243
rect 1008 -1275 1042 -1243
rect 806 -1277 840 -1275
rect 1008 -1277 1042 -1275
rect 902 -1309 936 -1279
rect 806 -1343 840 -1315
rect 902 -1313 936 -1309
rect 1008 -1343 1042 -1315
rect 806 -1349 840 -1343
rect 1008 -1349 1042 -1343
rect 902 -1377 936 -1351
rect 806 -1411 840 -1387
rect 902 -1385 936 -1377
rect 1008 -1411 1042 -1387
rect 806 -1421 840 -1411
rect 1008 -1421 1042 -1411
rect 902 -1445 936 -1423
rect 806 -1479 840 -1459
rect 902 -1457 936 -1445
rect 1008 -1479 1042 -1459
rect 806 -1493 840 -1479
rect 1008 -1493 1042 -1479
rect 902 -1513 936 -1495
rect 806 -1547 840 -1531
rect 902 -1529 936 -1513
rect 1008 -1547 1042 -1531
rect 806 -1565 840 -1547
rect 1008 -1565 1042 -1547
rect 902 -1581 936 -1567
rect 806 -1615 840 -1603
rect 902 -1601 936 -1581
rect 1008 -1615 1042 -1603
rect 806 -1637 840 -1615
rect 1008 -1637 1042 -1615
rect 902 -1649 936 -1639
rect 806 -1683 840 -1675
rect 902 -1673 936 -1649
rect 1008 -1683 1042 -1675
rect 806 -1709 840 -1683
rect 1008 -1709 1042 -1683
rect 902 -1717 936 -1711
rect 806 -1751 840 -1747
rect 902 -1745 936 -1717
rect 1008 -1751 1042 -1747
rect 806 -1781 840 -1751
rect 1008 -1781 1042 -1751
rect 902 -1785 936 -1783
rect 902 -1817 936 -1785
rect 806 -1853 840 -1819
rect 1008 -1853 1042 -1819
rect 902 -1887 936 -1855
rect 902 -1889 936 -1887
rect 806 -1921 840 -1891
rect 1008 -1921 1042 -1891
rect 806 -1925 840 -1921
rect 902 -1955 936 -1927
rect 1008 -1925 1042 -1921
rect 902 -1961 936 -1955
rect 806 -1989 840 -1963
rect 1008 -1989 1042 -1963
rect 806 -1997 840 -1989
rect 902 -2023 936 -1999
rect 1008 -1997 1042 -1989
rect 902 -2033 936 -2023
rect 806 -2057 840 -2035
rect 1008 -2057 1042 -2035
rect 806 -2069 840 -2057
rect 902 -2091 936 -2071
rect 1008 -2069 1042 -2057
rect 902 -2105 936 -2091
rect 806 -2125 840 -2107
rect 1008 -2125 1042 -2107
rect 806 -2141 840 -2125
rect 902 -2159 936 -2143
rect 1008 -2141 1042 -2125
rect 902 -2177 936 -2159
rect 806 -2193 840 -2179
rect 1008 -2193 1042 -2179
rect 806 -2213 840 -2193
rect 902 -2227 936 -2215
rect 1008 -2213 1042 -2193
rect 902 -2249 936 -2227
rect 806 -2261 840 -2251
rect 1008 -2261 1042 -2251
rect 806 -2285 840 -2261
rect 902 -2295 936 -2287
rect 1008 -2285 1042 -2261
rect 902 -2321 936 -2295
rect 806 -2329 840 -2323
rect 1008 -2329 1042 -2323
rect 806 -2357 840 -2329
rect 902 -2363 936 -2359
rect 1008 -2357 1042 -2329
rect 902 -2393 936 -2363
rect 806 -2397 840 -2395
rect 1008 -2397 1042 -2395
rect 806 -2429 840 -2397
rect 1008 -2429 1042 -2397
rect 902 -2465 936 -2431
rect 806 -2499 840 -2467
rect 1008 -2499 1042 -2467
rect 806 -2501 840 -2499
rect 1008 -2501 1042 -2499
rect 902 -2533 936 -2503
rect 806 -2567 840 -2539
rect 902 -2537 936 -2533
rect 1008 -2567 1042 -2539
rect 806 -2573 840 -2567
rect 1008 -2573 1042 -2567
rect 902 -2601 936 -2575
rect 806 -2635 840 -2611
rect 902 -2609 936 -2601
rect 1008 -2635 1042 -2611
rect 806 -2645 840 -2635
rect 1008 -2645 1042 -2635
rect 902 -2669 936 -2647
rect 806 -2703 840 -2683
rect 902 -2681 936 -2669
rect 1008 -2703 1042 -2683
rect 806 -2717 840 -2703
rect 1008 -2717 1042 -2703
rect 902 -2737 936 -2719
rect 806 -2771 840 -2755
rect 902 -2753 936 -2737
rect 1008 -2771 1042 -2755
rect 806 -2789 840 -2771
rect 1008 -2789 1042 -2771
rect 902 -2805 936 -2791
rect 806 -2839 840 -2827
rect 902 -2825 936 -2805
rect 1008 -2839 1042 -2827
rect 806 -2861 840 -2839
rect 1008 -2861 1042 -2839
rect 902 -2873 936 -2863
rect 806 -2907 840 -2899
rect 902 -2897 936 -2873
rect 1008 -2907 1042 -2899
rect 806 -2933 840 -2907
rect 1008 -2933 1042 -2907
rect 902 -2941 936 -2935
rect 806 -2975 840 -2971
rect 902 -2969 936 -2941
rect 1008 -2975 1042 -2971
rect 806 -3005 840 -2975
rect 1008 -3005 1042 -2975
rect 902 -3009 936 -3007
rect 902 -3041 936 -3009
rect 806 -3077 840 -3043
rect 1008 -3077 1042 -3043
rect 902 -3111 936 -3079
rect 902 -3113 936 -3111
rect 806 -3145 840 -3115
rect 1008 -3145 1042 -3115
rect 806 -3149 840 -3145
rect 902 -3179 936 -3151
rect 1008 -3149 1042 -3145
rect 902 -3185 936 -3179
rect 806 -3213 840 -3187
rect 1008 -3213 1042 -3187
rect 806 -3221 840 -3213
rect 902 -3247 936 -3223
rect 1008 -3221 1042 -3213
rect 902 -3257 936 -3247
rect 806 -3281 840 -3259
rect 1008 -3281 1042 -3259
rect 806 -3293 840 -3281
rect 902 -3315 936 -3295
rect 1008 -3293 1042 -3281
rect 902 -3329 936 -3315
rect 806 -3349 840 -3331
rect 1008 -3349 1042 -3331
rect 806 -3365 840 -3349
rect 902 -3383 936 -3367
rect 1008 -3365 1042 -3349
rect 902 -3401 936 -3383
rect 806 -3417 840 -3403
rect 1008 -3417 1042 -3403
rect 806 -3437 840 -3417
rect 902 -3451 936 -3439
rect 1008 -3437 1042 -3417
rect 902 -3473 936 -3451
rect 806 -3485 840 -3475
rect 1008 -3485 1042 -3475
rect 806 -3509 840 -3485
rect 902 -3519 936 -3511
rect 1008 -3509 1042 -3485
rect 902 -3545 936 -3519
rect 806 -3553 840 -3547
rect 1008 -3553 1042 -3547
rect 806 -3581 840 -3553
rect 902 -3587 936 -3583
rect 1008 -3581 1042 -3553
rect 902 -3617 936 -3587
rect 806 -3621 840 -3619
rect 1008 -3621 1042 -3619
rect 806 -3653 840 -3621
rect 1008 -3653 1042 -3621
rect 902 -3689 936 -3655
rect 806 -3723 840 -3691
rect 1008 -3723 1042 -3691
rect 806 -3725 840 -3723
rect 1008 -3725 1042 -3723
rect 902 -3757 936 -3727
rect 806 -3791 840 -3763
rect 902 -3761 936 -3757
rect 1008 -3791 1042 -3763
rect 806 -3797 840 -3791
rect 1008 -3797 1042 -3791
rect 902 -3825 936 -3799
rect 806 -3859 840 -3835
rect 902 -3833 936 -3825
rect 1008 -3859 1042 -3835
rect 806 -3869 840 -3859
rect 1008 -3869 1042 -3859
rect 902 -3893 936 -3871
rect 806 -3927 840 -3907
rect 902 -3905 936 -3893
rect 1008 -3927 1042 -3907
rect 806 -3941 840 -3927
rect 1008 -3941 1042 -3927
rect 902 -3961 936 -3943
rect 806 -3995 840 -3979
rect 902 -3977 936 -3961
rect 1008 -3995 1042 -3979
rect 806 -4013 840 -3995
rect 1008 -4013 1042 -3995
rect 902 -4029 936 -4015
rect 806 -4063 840 -4051
rect 902 -4049 936 -4029
rect 1008 -4063 1042 -4051
rect 806 -4085 840 -4063
rect 1008 -4085 1042 -4063
rect 902 -4097 936 -4087
rect 806 -4131 840 -4123
rect 902 -4121 936 -4097
rect 1008 -4131 1042 -4123
rect 806 -4157 840 -4131
rect 1008 -4157 1042 -4131
rect 902 -4165 936 -4159
rect 806 -4199 840 -4195
rect 902 -4193 936 -4165
rect 1008 -4199 1042 -4195
rect 806 -4229 840 -4199
rect 1008 -4229 1042 -4199
rect 902 -4233 936 -4231
rect 902 -4265 936 -4233
rect 806 -4301 840 -4267
rect 1008 -4301 1042 -4267
rect 902 -4335 936 -4303
rect 902 -4337 936 -4335
rect 806 -4369 840 -4339
rect 1008 -4369 1042 -4339
rect 806 -4373 840 -4369
rect 902 -4403 936 -4375
rect 1008 -4373 1042 -4369
rect 902 -4409 936 -4403
rect 806 -4437 840 -4411
rect 1008 -4437 1042 -4411
rect 806 -4445 840 -4437
rect 902 -4471 936 -4447
rect 1008 -4445 1042 -4437
rect 902 -4481 936 -4471
rect 806 -4505 840 -4483
rect 1008 -4505 1042 -4483
rect 806 -4517 840 -4505
rect 902 -4539 936 -4519
rect 1008 -4517 1042 -4505
rect 902 -4553 936 -4539
rect 806 -4573 840 -4555
rect 1008 -4573 1042 -4555
rect 806 -4589 840 -4573
rect 902 -4607 936 -4591
rect 1008 -4589 1042 -4573
rect 902 -4625 936 -4607
rect 806 -4641 840 -4627
rect 1008 -4641 1042 -4627
rect 806 -4661 840 -4641
rect 902 -4675 936 -4663
rect 1008 -4661 1042 -4641
rect 902 -4697 936 -4675
rect 806 -4709 840 -4699
rect 1008 -4709 1042 -4699
rect 806 -4733 840 -4709
rect 902 -4743 936 -4735
rect 1008 -4733 1042 -4709
rect 902 -4769 936 -4743
rect 806 -4777 840 -4771
rect 1008 -4777 1042 -4771
rect 806 -4805 840 -4777
rect 902 -4811 936 -4807
rect 1008 -4805 1042 -4777
rect 902 -4841 936 -4811
rect 806 -4845 840 -4843
rect 1008 -4845 1042 -4843
rect 806 -4877 840 -4845
rect 1008 -4877 1042 -4845
rect 902 -4913 936 -4879
rect 806 -4947 840 -4915
rect 1008 -4947 1042 -4915
rect 806 -4949 840 -4947
rect 1008 -4949 1042 -4947
rect 902 -4981 936 -4951
rect 190 -5021 224 -5015
rect 392 -5021 426 -5015
rect 286 -5057 320 -5023
rect 806 -5015 840 -4987
rect 902 -4985 936 -4981
rect 1008 -5015 1042 -4987
rect 1179 4981 1285 4985
rect 1179 -4981 1285 4981
rect 1179 -4985 1285 -4981
rect 806 -5021 840 -5015
rect 1008 -5021 1042 -5015
rect 902 -5057 936 -5023
rect 1422 -5015 1524 5015
rect 1524 -5015 1528 5015
rect 1422 -5021 1528 -5015
rect 1494 -5057 1528 -5023
rect -1357 -5124 -1351 -5090
rect -1351 -5124 -1323 -5090
rect -1285 -5124 -1283 -5090
rect -1283 -5124 -1251 -5090
rect -1213 -5124 -1181 -5090
rect -1181 -5124 -1179 -5090
rect -1141 -5124 -1113 -5090
rect -1113 -5124 -1107 -5090
rect -741 -5124 -735 -5090
rect -735 -5124 -707 -5090
rect -669 -5124 -667 -5090
rect -667 -5124 -635 -5090
rect -597 -5124 -565 -5090
rect -565 -5124 -563 -5090
rect -525 -5124 -497 -5090
rect -497 -5124 -491 -5090
rect -125 -5124 -119 -5090
rect -119 -5124 -91 -5090
rect -53 -5124 -51 -5090
rect -51 -5124 -19 -5090
rect 19 -5124 51 -5090
rect 51 -5124 53 -5090
rect 91 -5124 119 -5090
rect 119 -5124 125 -5090
rect 491 -5124 497 -5090
rect 497 -5124 525 -5090
rect 563 -5124 565 -5090
rect 565 -5124 597 -5090
rect 635 -5124 667 -5090
rect 667 -5124 669 -5090
rect 707 -5124 735 -5090
rect 735 -5124 741 -5090
rect 1107 -5124 1113 -5090
rect 1113 -5124 1141 -5090
rect 1179 -5124 1181 -5090
rect 1181 -5124 1213 -5090
rect 1251 -5124 1283 -5090
rect 1283 -5124 1285 -5090
rect 1323 -5124 1351 -5090
rect 1351 -5124 1357 -5090
<< metal1 >>
rect -1540 5124 1540 5188
rect -1540 5090 -1357 5124
rect -1323 5090 -1285 5124
rect -1251 5090 -1213 5124
rect -1179 5090 -1141 5124
rect -1107 5090 -741 5124
rect -707 5090 -669 5124
rect -635 5090 -597 5124
rect -563 5090 -525 5124
rect -491 5090 -125 5124
rect -91 5090 -53 5124
rect -19 5090 19 5124
rect 53 5090 91 5124
rect 125 5090 491 5124
rect 525 5090 563 5124
rect 597 5090 635 5124
rect 669 5090 707 5124
rect 741 5090 1107 5124
rect 1141 5090 1179 5124
rect 1213 5090 1251 5124
rect 1285 5090 1323 5124
rect 1357 5090 1540 5124
rect -1540 5084 1540 5090
rect -1540 5062 -1398 5084
tri -1398 5062 -1376 5084 nw
tri -1088 5062 -1066 5084 ne
rect -1066 5062 -782 5084
tri -782 5062 -760 5084 nw
tri -472 5062 -450 5084 ne
rect -450 5062 -166 5084
tri -166 5062 -144 5084 nw
tri 144 5062 166 5084 ne
rect 166 5062 450 5084
tri 450 5062 472 5084 nw
tri 760 5062 782 5084 ne
rect 782 5062 1066 5084
tri 1066 5062 1088 5084 nw
tri 1376 5062 1398 5084 ne
rect 1398 5062 1540 5084
rect -1540 5057 -1403 5062
tri -1403 5057 -1398 5062 nw
tri -1066 5057 -1061 5062 ne
rect -1061 5057 -787 5062
tri -787 5057 -782 5062 nw
tri -450 5057 -445 5062 ne
rect -445 5057 -171 5062
tri -171 5057 -166 5062 nw
tri 166 5057 171 5062 ne
rect 171 5057 445 5062
tri 445 5057 450 5062 nw
tri 782 5057 787 5062 ne
rect 787 5057 1061 5062
tri 1061 5057 1066 5062 nw
tri 1398 5057 1403 5062 ne
rect 1403 5057 1540 5062
rect -1540 5023 -1528 5057
rect -1494 5023 -1416 5057
tri -1416 5044 -1403 5057 nw
tri -1061 5044 -1048 5057 ne
rect -1540 5021 -1416 5023
rect -1540 -5021 -1528 5021
rect -1422 -5021 -1416 5021
rect -1048 5023 -946 5057
rect -912 5023 -800 5057
tri -800 5044 -787 5057 nw
tri -445 5044 -432 5057 ne
rect -1048 5021 -800 5023
tri -1326 5000 -1306 5020 se
rect -1306 5000 -1158 5020
tri -1158 5000 -1138 5020 sw
rect -1326 4985 -1138 5000
rect -1326 -4985 -1285 4985
rect -1179 -4985 -1138 4985
rect -1326 -5000 -1138 -4985
tri -1326 -5020 -1306 -5000 ne
rect -1306 -5020 -1158 -5000
tri -1158 -5020 -1138 -5000 nw
rect -1048 4987 -1042 5021
rect -1008 4987 -840 5021
rect -806 4987 -800 5021
rect -432 5023 -330 5057
rect -296 5023 -184 5057
tri -184 5044 -171 5057 nw
tri 171 5044 184 5057 ne
rect -432 5021 -184 5023
rect -1048 4985 -800 4987
rect -1048 4951 -946 4985
rect -912 4951 -800 4985
rect -1048 4949 -800 4951
rect -1048 4915 -1042 4949
rect -1008 4915 -840 4949
rect -806 4915 -800 4949
rect -1048 4913 -800 4915
rect -1048 4879 -946 4913
rect -912 4879 -800 4913
rect -1048 4877 -800 4879
rect -1048 4843 -1042 4877
rect -1008 4843 -840 4877
rect -806 4843 -800 4877
rect -1048 4841 -800 4843
rect -1048 4807 -946 4841
rect -912 4807 -800 4841
rect -1048 4805 -800 4807
rect -1048 4771 -1042 4805
rect -1008 4771 -840 4805
rect -806 4771 -800 4805
rect -1048 4769 -800 4771
rect -1048 4735 -946 4769
rect -912 4735 -800 4769
rect -1048 4733 -800 4735
rect -1048 4699 -1042 4733
rect -1008 4699 -840 4733
rect -806 4699 -800 4733
rect -1048 4697 -800 4699
rect -1048 4663 -946 4697
rect -912 4663 -800 4697
rect -1048 4661 -800 4663
rect -1048 4627 -1042 4661
rect -1008 4627 -840 4661
rect -806 4627 -800 4661
rect -1048 4625 -800 4627
rect -1048 4591 -946 4625
rect -912 4591 -800 4625
rect -1048 4589 -800 4591
rect -1048 4555 -1042 4589
rect -1008 4555 -840 4589
rect -806 4555 -800 4589
rect -1048 4553 -800 4555
rect -1048 4519 -946 4553
rect -912 4519 -800 4553
rect -1048 4517 -800 4519
rect -1048 4483 -1042 4517
rect -1008 4483 -840 4517
rect -806 4483 -800 4517
rect -1048 4481 -800 4483
rect -1048 4447 -946 4481
rect -912 4447 -800 4481
rect -1048 4445 -800 4447
rect -1048 4411 -1042 4445
rect -1008 4411 -840 4445
rect -806 4411 -800 4445
rect -1048 4409 -800 4411
rect -1048 4375 -946 4409
rect -912 4375 -800 4409
rect -1048 4373 -800 4375
rect -1048 4339 -1042 4373
rect -1008 4339 -840 4373
rect -806 4339 -800 4373
rect -1048 4337 -800 4339
rect -1048 4303 -946 4337
rect -912 4303 -800 4337
rect -1048 4301 -800 4303
rect -1048 4267 -1042 4301
rect -1008 4267 -840 4301
rect -806 4267 -800 4301
rect -1048 4265 -800 4267
rect -1048 4231 -946 4265
rect -912 4231 -800 4265
rect -1048 4229 -800 4231
rect -1048 4195 -1042 4229
rect -1008 4195 -840 4229
rect -806 4195 -800 4229
rect -1048 4193 -800 4195
rect -1048 4159 -946 4193
rect -912 4159 -800 4193
rect -1048 4157 -800 4159
rect -1048 4123 -1042 4157
rect -1008 4123 -840 4157
rect -806 4123 -800 4157
rect -1048 4121 -800 4123
rect -1048 4087 -946 4121
rect -912 4087 -800 4121
rect -1048 4085 -800 4087
rect -1048 4051 -1042 4085
rect -1008 4051 -840 4085
rect -806 4051 -800 4085
rect -1048 4049 -800 4051
rect -1048 4015 -946 4049
rect -912 4015 -800 4049
rect -1048 4013 -800 4015
rect -1048 3979 -1042 4013
rect -1008 3979 -840 4013
rect -806 3979 -800 4013
rect -1048 3977 -800 3979
rect -1048 3943 -946 3977
rect -912 3943 -800 3977
rect -1048 3941 -800 3943
rect -1048 3907 -1042 3941
rect -1008 3907 -840 3941
rect -806 3907 -800 3941
rect -1048 3905 -800 3907
rect -1048 3871 -946 3905
rect -912 3871 -800 3905
rect -1048 3869 -800 3871
rect -1048 3835 -1042 3869
rect -1008 3835 -840 3869
rect -806 3835 -800 3869
rect -1048 3833 -800 3835
rect -1048 3799 -946 3833
rect -912 3799 -800 3833
rect -1048 3797 -800 3799
rect -1048 3763 -1042 3797
rect -1008 3763 -840 3797
rect -806 3763 -800 3797
rect -1048 3761 -800 3763
rect -1048 3727 -946 3761
rect -912 3727 -800 3761
rect -1048 3725 -800 3727
rect -1048 3691 -1042 3725
rect -1008 3691 -840 3725
rect -806 3691 -800 3725
rect -1048 3689 -800 3691
rect -1048 3655 -946 3689
rect -912 3655 -800 3689
rect -1048 3653 -800 3655
rect -1048 3619 -1042 3653
rect -1008 3619 -840 3653
rect -806 3619 -800 3653
rect -1048 3617 -800 3619
rect -1048 3583 -946 3617
rect -912 3583 -800 3617
rect -1048 3581 -800 3583
rect -1048 3547 -1042 3581
rect -1008 3547 -840 3581
rect -806 3547 -800 3581
rect -1048 3545 -800 3547
rect -1048 3511 -946 3545
rect -912 3511 -800 3545
rect -1048 3509 -800 3511
rect -1048 3475 -1042 3509
rect -1008 3475 -840 3509
rect -806 3475 -800 3509
rect -1048 3473 -800 3475
rect -1048 3439 -946 3473
rect -912 3439 -800 3473
rect -1048 3437 -800 3439
rect -1048 3403 -1042 3437
rect -1008 3403 -840 3437
rect -806 3403 -800 3437
rect -1048 3401 -800 3403
rect -1048 3367 -946 3401
rect -912 3367 -800 3401
rect -1048 3365 -800 3367
rect -1048 3331 -1042 3365
rect -1008 3331 -840 3365
rect -806 3331 -800 3365
rect -1048 3329 -800 3331
rect -1048 3295 -946 3329
rect -912 3295 -800 3329
rect -1048 3293 -800 3295
rect -1048 3259 -1042 3293
rect -1008 3259 -840 3293
rect -806 3259 -800 3293
rect -1048 3257 -800 3259
rect -1048 3223 -946 3257
rect -912 3223 -800 3257
rect -1048 3221 -800 3223
rect -1048 3187 -1042 3221
rect -1008 3187 -840 3221
rect -806 3187 -800 3221
rect -1048 3185 -800 3187
rect -1048 3151 -946 3185
rect -912 3151 -800 3185
rect -1048 3149 -800 3151
rect -1048 3115 -1042 3149
rect -1008 3115 -840 3149
rect -806 3115 -800 3149
rect -1048 3113 -800 3115
rect -1048 3079 -946 3113
rect -912 3079 -800 3113
rect -1048 3077 -800 3079
rect -1048 3043 -1042 3077
rect -1008 3043 -840 3077
rect -806 3043 -800 3077
rect -1048 3041 -800 3043
rect -1048 3007 -946 3041
rect -912 3007 -800 3041
rect -1048 3005 -800 3007
rect -1048 2971 -1042 3005
rect -1008 2971 -840 3005
rect -806 2971 -800 3005
rect -1048 2969 -800 2971
rect -1048 2935 -946 2969
rect -912 2935 -800 2969
rect -1048 2933 -800 2935
rect -1048 2899 -1042 2933
rect -1008 2899 -840 2933
rect -806 2899 -800 2933
rect -1048 2897 -800 2899
rect -1048 2863 -946 2897
rect -912 2863 -800 2897
rect -1048 2861 -800 2863
rect -1048 2827 -1042 2861
rect -1008 2827 -840 2861
rect -806 2827 -800 2861
rect -1048 2825 -800 2827
rect -1048 2791 -946 2825
rect -912 2791 -800 2825
rect -1048 2789 -800 2791
rect -1048 2755 -1042 2789
rect -1008 2755 -840 2789
rect -806 2755 -800 2789
rect -1048 2753 -800 2755
rect -1048 2719 -946 2753
rect -912 2719 -800 2753
rect -1048 2717 -800 2719
rect -1048 2683 -1042 2717
rect -1008 2683 -840 2717
rect -806 2683 -800 2717
rect -1048 2681 -800 2683
rect -1048 2647 -946 2681
rect -912 2647 -800 2681
rect -1048 2645 -800 2647
rect -1048 2611 -1042 2645
rect -1008 2611 -840 2645
rect -806 2611 -800 2645
rect -1048 2609 -800 2611
rect -1048 2575 -946 2609
rect -912 2575 -800 2609
rect -1048 2573 -800 2575
rect -1048 2539 -1042 2573
rect -1008 2539 -840 2573
rect -806 2539 -800 2573
rect -1048 2537 -800 2539
rect -1048 2503 -946 2537
rect -912 2503 -800 2537
rect -1048 2501 -800 2503
rect -1048 2467 -1042 2501
rect -1008 2467 -840 2501
rect -806 2467 -800 2501
rect -1048 2465 -800 2467
rect -1048 2431 -946 2465
rect -912 2431 -800 2465
rect -1048 2429 -800 2431
rect -1048 2395 -1042 2429
rect -1008 2395 -840 2429
rect -806 2395 -800 2429
rect -1048 2393 -800 2395
rect -1048 2359 -946 2393
rect -912 2359 -800 2393
rect -1048 2357 -800 2359
rect -1048 2323 -1042 2357
rect -1008 2323 -840 2357
rect -806 2323 -800 2357
rect -1048 2321 -800 2323
rect -1048 2287 -946 2321
rect -912 2287 -800 2321
rect -1048 2285 -800 2287
rect -1048 2251 -1042 2285
rect -1008 2251 -840 2285
rect -806 2251 -800 2285
rect -1048 2249 -800 2251
rect -1048 2215 -946 2249
rect -912 2215 -800 2249
rect -1048 2213 -800 2215
rect -1048 2179 -1042 2213
rect -1008 2179 -840 2213
rect -806 2179 -800 2213
rect -1048 2177 -800 2179
rect -1048 2143 -946 2177
rect -912 2143 -800 2177
rect -1048 2141 -800 2143
rect -1048 2107 -1042 2141
rect -1008 2107 -840 2141
rect -806 2107 -800 2141
rect -1048 2105 -800 2107
rect -1048 2071 -946 2105
rect -912 2071 -800 2105
rect -1048 2069 -800 2071
rect -1048 2035 -1042 2069
rect -1008 2035 -840 2069
rect -806 2035 -800 2069
rect -1048 2033 -800 2035
rect -1048 1999 -946 2033
rect -912 1999 -800 2033
rect -1048 1997 -800 1999
rect -1048 1963 -1042 1997
rect -1008 1963 -840 1997
rect -806 1963 -800 1997
rect -1048 1961 -800 1963
rect -1048 1927 -946 1961
rect -912 1927 -800 1961
rect -1048 1925 -800 1927
rect -1048 1891 -1042 1925
rect -1008 1891 -840 1925
rect -806 1891 -800 1925
rect -1048 1889 -800 1891
rect -1048 1855 -946 1889
rect -912 1855 -800 1889
rect -1048 1853 -800 1855
rect -1048 1819 -1042 1853
rect -1008 1819 -840 1853
rect -806 1819 -800 1853
rect -1048 1817 -800 1819
rect -1048 1783 -946 1817
rect -912 1783 -800 1817
rect -1048 1781 -800 1783
rect -1048 1747 -1042 1781
rect -1008 1747 -840 1781
rect -806 1747 -800 1781
rect -1048 1745 -800 1747
rect -1048 1711 -946 1745
rect -912 1711 -800 1745
rect -1048 1709 -800 1711
rect -1048 1675 -1042 1709
rect -1008 1675 -840 1709
rect -806 1675 -800 1709
rect -1048 1673 -800 1675
rect -1048 1639 -946 1673
rect -912 1639 -800 1673
rect -1048 1637 -800 1639
rect -1048 1603 -1042 1637
rect -1008 1603 -840 1637
rect -806 1603 -800 1637
rect -1048 1601 -800 1603
rect -1048 1567 -946 1601
rect -912 1567 -800 1601
rect -1048 1565 -800 1567
rect -1048 1531 -1042 1565
rect -1008 1531 -840 1565
rect -806 1531 -800 1565
rect -1048 1529 -800 1531
rect -1048 1495 -946 1529
rect -912 1495 -800 1529
rect -1048 1493 -800 1495
rect -1048 1459 -1042 1493
rect -1008 1459 -840 1493
rect -806 1459 -800 1493
rect -1048 1457 -800 1459
rect -1048 1423 -946 1457
rect -912 1423 -800 1457
rect -1048 1421 -800 1423
rect -1048 1387 -1042 1421
rect -1008 1387 -840 1421
rect -806 1387 -800 1421
rect -1048 1385 -800 1387
rect -1048 1351 -946 1385
rect -912 1351 -800 1385
rect -1048 1349 -800 1351
rect -1048 1315 -1042 1349
rect -1008 1315 -840 1349
rect -806 1315 -800 1349
rect -1048 1313 -800 1315
rect -1048 1279 -946 1313
rect -912 1279 -800 1313
rect -1048 1277 -800 1279
rect -1048 1243 -1042 1277
rect -1008 1243 -840 1277
rect -806 1243 -800 1277
rect -1048 1241 -800 1243
rect -1048 1207 -946 1241
rect -912 1207 -800 1241
rect -1048 1205 -800 1207
rect -1048 1171 -1042 1205
rect -1008 1171 -840 1205
rect -806 1171 -800 1205
rect -1048 1169 -800 1171
rect -1048 1135 -946 1169
rect -912 1135 -800 1169
rect -1048 1133 -800 1135
rect -1048 1099 -1042 1133
rect -1008 1099 -840 1133
rect -806 1099 -800 1133
rect -1048 1097 -800 1099
rect -1048 1063 -946 1097
rect -912 1063 -800 1097
rect -1048 1061 -800 1063
rect -1048 1027 -1042 1061
rect -1008 1027 -840 1061
rect -806 1027 -800 1061
rect -1048 1025 -800 1027
rect -1048 991 -946 1025
rect -912 991 -800 1025
rect -1048 989 -800 991
rect -1048 955 -1042 989
rect -1008 955 -840 989
rect -806 955 -800 989
rect -1048 953 -800 955
rect -1048 919 -946 953
rect -912 919 -800 953
rect -1048 917 -800 919
rect -1048 883 -1042 917
rect -1008 883 -840 917
rect -806 883 -800 917
rect -1048 881 -800 883
rect -1048 847 -946 881
rect -912 847 -800 881
rect -1048 845 -800 847
rect -1048 811 -1042 845
rect -1008 811 -840 845
rect -806 811 -800 845
rect -1048 809 -800 811
rect -1048 775 -946 809
rect -912 775 -800 809
rect -1048 773 -800 775
rect -1048 739 -1042 773
rect -1008 739 -840 773
rect -806 739 -800 773
rect -1048 737 -800 739
rect -1048 703 -946 737
rect -912 703 -800 737
rect -1048 701 -800 703
rect -1048 667 -1042 701
rect -1008 667 -840 701
rect -806 667 -800 701
rect -1048 665 -800 667
rect -1048 631 -946 665
rect -912 631 -800 665
rect -1048 629 -800 631
rect -1048 595 -1042 629
rect -1008 595 -840 629
rect -806 595 -800 629
rect -1048 593 -800 595
rect -1048 559 -946 593
rect -912 559 -800 593
rect -1048 557 -800 559
rect -1048 523 -1042 557
rect -1008 523 -840 557
rect -806 523 -800 557
rect -1048 521 -800 523
rect -1048 487 -946 521
rect -912 487 -800 521
rect -1048 485 -800 487
rect -1048 451 -1042 485
rect -1008 451 -840 485
rect -806 451 -800 485
rect -1048 449 -800 451
rect -1048 415 -946 449
rect -912 415 -800 449
rect -1048 413 -800 415
rect -1048 379 -1042 413
rect -1008 379 -840 413
rect -806 379 -800 413
rect -1048 377 -800 379
rect -1048 343 -946 377
rect -912 343 -800 377
rect -1048 341 -800 343
rect -1048 307 -1042 341
rect -1008 307 -840 341
rect -806 307 -800 341
rect -1048 305 -800 307
rect -1048 271 -946 305
rect -912 271 -800 305
rect -1048 269 -800 271
rect -1048 235 -1042 269
rect -1008 235 -840 269
rect -806 235 -800 269
rect -1048 233 -800 235
rect -1048 199 -946 233
rect -912 199 -800 233
rect -1048 197 -800 199
rect -1048 163 -1042 197
rect -1008 163 -840 197
rect -806 163 -800 197
rect -1048 161 -800 163
rect -1048 127 -946 161
rect -912 127 -800 161
rect -1048 125 -800 127
rect -1048 91 -1042 125
rect -1008 91 -840 125
rect -806 91 -800 125
rect -1048 89 -800 91
rect -1048 55 -946 89
rect -912 55 -800 89
rect -1048 53 -800 55
rect -1048 19 -1042 53
rect -1008 19 -840 53
rect -806 19 -800 53
rect -1048 17 -800 19
rect -1048 -17 -946 17
rect -912 -17 -800 17
rect -1048 -19 -800 -17
rect -1048 -53 -1042 -19
rect -1008 -53 -840 -19
rect -806 -53 -800 -19
rect -1048 -55 -800 -53
rect -1048 -89 -946 -55
rect -912 -89 -800 -55
rect -1048 -91 -800 -89
rect -1048 -125 -1042 -91
rect -1008 -125 -840 -91
rect -806 -125 -800 -91
rect -1048 -127 -800 -125
rect -1048 -161 -946 -127
rect -912 -161 -800 -127
rect -1048 -163 -800 -161
rect -1048 -197 -1042 -163
rect -1008 -197 -840 -163
rect -806 -197 -800 -163
rect -1048 -199 -800 -197
rect -1048 -233 -946 -199
rect -912 -233 -800 -199
rect -1048 -235 -800 -233
rect -1048 -269 -1042 -235
rect -1008 -269 -840 -235
rect -806 -269 -800 -235
rect -1048 -271 -800 -269
rect -1048 -305 -946 -271
rect -912 -305 -800 -271
rect -1048 -307 -800 -305
rect -1048 -341 -1042 -307
rect -1008 -341 -840 -307
rect -806 -341 -800 -307
rect -1048 -343 -800 -341
rect -1048 -377 -946 -343
rect -912 -377 -800 -343
rect -1048 -379 -800 -377
rect -1048 -413 -1042 -379
rect -1008 -413 -840 -379
rect -806 -413 -800 -379
rect -1048 -415 -800 -413
rect -1048 -449 -946 -415
rect -912 -449 -800 -415
rect -1048 -451 -800 -449
rect -1048 -485 -1042 -451
rect -1008 -485 -840 -451
rect -806 -485 -800 -451
rect -1048 -487 -800 -485
rect -1048 -521 -946 -487
rect -912 -521 -800 -487
rect -1048 -523 -800 -521
rect -1048 -557 -1042 -523
rect -1008 -557 -840 -523
rect -806 -557 -800 -523
rect -1048 -559 -800 -557
rect -1048 -593 -946 -559
rect -912 -593 -800 -559
rect -1048 -595 -800 -593
rect -1048 -629 -1042 -595
rect -1008 -629 -840 -595
rect -806 -629 -800 -595
rect -1048 -631 -800 -629
rect -1048 -665 -946 -631
rect -912 -665 -800 -631
rect -1048 -667 -800 -665
rect -1048 -701 -1042 -667
rect -1008 -701 -840 -667
rect -806 -701 -800 -667
rect -1048 -703 -800 -701
rect -1048 -737 -946 -703
rect -912 -737 -800 -703
rect -1048 -739 -800 -737
rect -1048 -773 -1042 -739
rect -1008 -773 -840 -739
rect -806 -773 -800 -739
rect -1048 -775 -800 -773
rect -1048 -809 -946 -775
rect -912 -809 -800 -775
rect -1048 -811 -800 -809
rect -1048 -845 -1042 -811
rect -1008 -845 -840 -811
rect -806 -845 -800 -811
rect -1048 -847 -800 -845
rect -1048 -881 -946 -847
rect -912 -881 -800 -847
rect -1048 -883 -800 -881
rect -1048 -917 -1042 -883
rect -1008 -917 -840 -883
rect -806 -917 -800 -883
rect -1048 -919 -800 -917
rect -1048 -953 -946 -919
rect -912 -953 -800 -919
rect -1048 -955 -800 -953
rect -1048 -989 -1042 -955
rect -1008 -989 -840 -955
rect -806 -989 -800 -955
rect -1048 -991 -800 -989
rect -1048 -1025 -946 -991
rect -912 -1025 -800 -991
rect -1048 -1027 -800 -1025
rect -1048 -1061 -1042 -1027
rect -1008 -1061 -840 -1027
rect -806 -1061 -800 -1027
rect -1048 -1063 -800 -1061
rect -1048 -1097 -946 -1063
rect -912 -1097 -800 -1063
rect -1048 -1099 -800 -1097
rect -1048 -1133 -1042 -1099
rect -1008 -1133 -840 -1099
rect -806 -1133 -800 -1099
rect -1048 -1135 -800 -1133
rect -1048 -1169 -946 -1135
rect -912 -1169 -800 -1135
rect -1048 -1171 -800 -1169
rect -1048 -1205 -1042 -1171
rect -1008 -1205 -840 -1171
rect -806 -1205 -800 -1171
rect -1048 -1207 -800 -1205
rect -1048 -1241 -946 -1207
rect -912 -1241 -800 -1207
rect -1048 -1243 -800 -1241
rect -1048 -1277 -1042 -1243
rect -1008 -1277 -840 -1243
rect -806 -1277 -800 -1243
rect -1048 -1279 -800 -1277
rect -1048 -1313 -946 -1279
rect -912 -1313 -800 -1279
rect -1048 -1315 -800 -1313
rect -1048 -1349 -1042 -1315
rect -1008 -1349 -840 -1315
rect -806 -1349 -800 -1315
rect -1048 -1351 -800 -1349
rect -1048 -1385 -946 -1351
rect -912 -1385 -800 -1351
rect -1048 -1387 -800 -1385
rect -1048 -1421 -1042 -1387
rect -1008 -1421 -840 -1387
rect -806 -1421 -800 -1387
rect -1048 -1423 -800 -1421
rect -1048 -1457 -946 -1423
rect -912 -1457 -800 -1423
rect -1048 -1459 -800 -1457
rect -1048 -1493 -1042 -1459
rect -1008 -1493 -840 -1459
rect -806 -1493 -800 -1459
rect -1048 -1495 -800 -1493
rect -1048 -1529 -946 -1495
rect -912 -1529 -800 -1495
rect -1048 -1531 -800 -1529
rect -1048 -1565 -1042 -1531
rect -1008 -1565 -840 -1531
rect -806 -1565 -800 -1531
rect -1048 -1567 -800 -1565
rect -1048 -1601 -946 -1567
rect -912 -1601 -800 -1567
rect -1048 -1603 -800 -1601
rect -1048 -1637 -1042 -1603
rect -1008 -1637 -840 -1603
rect -806 -1637 -800 -1603
rect -1048 -1639 -800 -1637
rect -1048 -1673 -946 -1639
rect -912 -1673 -800 -1639
rect -1048 -1675 -800 -1673
rect -1048 -1709 -1042 -1675
rect -1008 -1709 -840 -1675
rect -806 -1709 -800 -1675
rect -1048 -1711 -800 -1709
rect -1048 -1745 -946 -1711
rect -912 -1745 -800 -1711
rect -1048 -1747 -800 -1745
rect -1048 -1781 -1042 -1747
rect -1008 -1781 -840 -1747
rect -806 -1781 -800 -1747
rect -1048 -1783 -800 -1781
rect -1048 -1817 -946 -1783
rect -912 -1817 -800 -1783
rect -1048 -1819 -800 -1817
rect -1048 -1853 -1042 -1819
rect -1008 -1853 -840 -1819
rect -806 -1853 -800 -1819
rect -1048 -1855 -800 -1853
rect -1048 -1889 -946 -1855
rect -912 -1889 -800 -1855
rect -1048 -1891 -800 -1889
rect -1048 -1925 -1042 -1891
rect -1008 -1925 -840 -1891
rect -806 -1925 -800 -1891
rect -1048 -1927 -800 -1925
rect -1048 -1961 -946 -1927
rect -912 -1961 -800 -1927
rect -1048 -1963 -800 -1961
rect -1048 -1997 -1042 -1963
rect -1008 -1997 -840 -1963
rect -806 -1997 -800 -1963
rect -1048 -1999 -800 -1997
rect -1048 -2033 -946 -1999
rect -912 -2033 -800 -1999
rect -1048 -2035 -800 -2033
rect -1048 -2069 -1042 -2035
rect -1008 -2069 -840 -2035
rect -806 -2069 -800 -2035
rect -1048 -2071 -800 -2069
rect -1048 -2105 -946 -2071
rect -912 -2105 -800 -2071
rect -1048 -2107 -800 -2105
rect -1048 -2141 -1042 -2107
rect -1008 -2141 -840 -2107
rect -806 -2141 -800 -2107
rect -1048 -2143 -800 -2141
rect -1048 -2177 -946 -2143
rect -912 -2177 -800 -2143
rect -1048 -2179 -800 -2177
rect -1048 -2213 -1042 -2179
rect -1008 -2213 -840 -2179
rect -806 -2213 -800 -2179
rect -1048 -2215 -800 -2213
rect -1048 -2249 -946 -2215
rect -912 -2249 -800 -2215
rect -1048 -2251 -800 -2249
rect -1048 -2285 -1042 -2251
rect -1008 -2285 -840 -2251
rect -806 -2285 -800 -2251
rect -1048 -2287 -800 -2285
rect -1048 -2321 -946 -2287
rect -912 -2321 -800 -2287
rect -1048 -2323 -800 -2321
rect -1048 -2357 -1042 -2323
rect -1008 -2357 -840 -2323
rect -806 -2357 -800 -2323
rect -1048 -2359 -800 -2357
rect -1048 -2393 -946 -2359
rect -912 -2393 -800 -2359
rect -1048 -2395 -800 -2393
rect -1048 -2429 -1042 -2395
rect -1008 -2429 -840 -2395
rect -806 -2429 -800 -2395
rect -1048 -2431 -800 -2429
rect -1048 -2465 -946 -2431
rect -912 -2465 -800 -2431
rect -1048 -2467 -800 -2465
rect -1048 -2501 -1042 -2467
rect -1008 -2501 -840 -2467
rect -806 -2501 -800 -2467
rect -1048 -2503 -800 -2501
rect -1048 -2537 -946 -2503
rect -912 -2537 -800 -2503
rect -1048 -2539 -800 -2537
rect -1048 -2573 -1042 -2539
rect -1008 -2573 -840 -2539
rect -806 -2573 -800 -2539
rect -1048 -2575 -800 -2573
rect -1048 -2609 -946 -2575
rect -912 -2609 -800 -2575
rect -1048 -2611 -800 -2609
rect -1048 -2645 -1042 -2611
rect -1008 -2645 -840 -2611
rect -806 -2645 -800 -2611
rect -1048 -2647 -800 -2645
rect -1048 -2681 -946 -2647
rect -912 -2681 -800 -2647
rect -1048 -2683 -800 -2681
rect -1048 -2717 -1042 -2683
rect -1008 -2717 -840 -2683
rect -806 -2717 -800 -2683
rect -1048 -2719 -800 -2717
rect -1048 -2753 -946 -2719
rect -912 -2753 -800 -2719
rect -1048 -2755 -800 -2753
rect -1048 -2789 -1042 -2755
rect -1008 -2789 -840 -2755
rect -806 -2789 -800 -2755
rect -1048 -2791 -800 -2789
rect -1048 -2825 -946 -2791
rect -912 -2825 -800 -2791
rect -1048 -2827 -800 -2825
rect -1048 -2861 -1042 -2827
rect -1008 -2861 -840 -2827
rect -806 -2861 -800 -2827
rect -1048 -2863 -800 -2861
rect -1048 -2897 -946 -2863
rect -912 -2897 -800 -2863
rect -1048 -2899 -800 -2897
rect -1048 -2933 -1042 -2899
rect -1008 -2933 -840 -2899
rect -806 -2933 -800 -2899
rect -1048 -2935 -800 -2933
rect -1048 -2969 -946 -2935
rect -912 -2969 -800 -2935
rect -1048 -2971 -800 -2969
rect -1048 -3005 -1042 -2971
rect -1008 -3005 -840 -2971
rect -806 -3005 -800 -2971
rect -1048 -3007 -800 -3005
rect -1048 -3041 -946 -3007
rect -912 -3041 -800 -3007
rect -1048 -3043 -800 -3041
rect -1048 -3077 -1042 -3043
rect -1008 -3077 -840 -3043
rect -806 -3077 -800 -3043
rect -1048 -3079 -800 -3077
rect -1048 -3113 -946 -3079
rect -912 -3113 -800 -3079
rect -1048 -3115 -800 -3113
rect -1048 -3149 -1042 -3115
rect -1008 -3149 -840 -3115
rect -806 -3149 -800 -3115
rect -1048 -3151 -800 -3149
rect -1048 -3185 -946 -3151
rect -912 -3185 -800 -3151
rect -1048 -3187 -800 -3185
rect -1048 -3221 -1042 -3187
rect -1008 -3221 -840 -3187
rect -806 -3221 -800 -3187
rect -1048 -3223 -800 -3221
rect -1048 -3257 -946 -3223
rect -912 -3257 -800 -3223
rect -1048 -3259 -800 -3257
rect -1048 -3293 -1042 -3259
rect -1008 -3293 -840 -3259
rect -806 -3293 -800 -3259
rect -1048 -3295 -800 -3293
rect -1048 -3329 -946 -3295
rect -912 -3329 -800 -3295
rect -1048 -3331 -800 -3329
rect -1048 -3365 -1042 -3331
rect -1008 -3365 -840 -3331
rect -806 -3365 -800 -3331
rect -1048 -3367 -800 -3365
rect -1048 -3401 -946 -3367
rect -912 -3401 -800 -3367
rect -1048 -3403 -800 -3401
rect -1048 -3437 -1042 -3403
rect -1008 -3437 -840 -3403
rect -806 -3437 -800 -3403
rect -1048 -3439 -800 -3437
rect -1048 -3473 -946 -3439
rect -912 -3473 -800 -3439
rect -1048 -3475 -800 -3473
rect -1048 -3509 -1042 -3475
rect -1008 -3509 -840 -3475
rect -806 -3509 -800 -3475
rect -1048 -3511 -800 -3509
rect -1048 -3545 -946 -3511
rect -912 -3545 -800 -3511
rect -1048 -3547 -800 -3545
rect -1048 -3581 -1042 -3547
rect -1008 -3581 -840 -3547
rect -806 -3581 -800 -3547
rect -1048 -3583 -800 -3581
rect -1048 -3617 -946 -3583
rect -912 -3617 -800 -3583
rect -1048 -3619 -800 -3617
rect -1048 -3653 -1042 -3619
rect -1008 -3653 -840 -3619
rect -806 -3653 -800 -3619
rect -1048 -3655 -800 -3653
rect -1048 -3689 -946 -3655
rect -912 -3689 -800 -3655
rect -1048 -3691 -800 -3689
rect -1048 -3725 -1042 -3691
rect -1008 -3725 -840 -3691
rect -806 -3725 -800 -3691
rect -1048 -3727 -800 -3725
rect -1048 -3761 -946 -3727
rect -912 -3761 -800 -3727
rect -1048 -3763 -800 -3761
rect -1048 -3797 -1042 -3763
rect -1008 -3797 -840 -3763
rect -806 -3797 -800 -3763
rect -1048 -3799 -800 -3797
rect -1048 -3833 -946 -3799
rect -912 -3833 -800 -3799
rect -1048 -3835 -800 -3833
rect -1048 -3869 -1042 -3835
rect -1008 -3869 -840 -3835
rect -806 -3869 -800 -3835
rect -1048 -3871 -800 -3869
rect -1048 -3905 -946 -3871
rect -912 -3905 -800 -3871
rect -1048 -3907 -800 -3905
rect -1048 -3941 -1042 -3907
rect -1008 -3941 -840 -3907
rect -806 -3941 -800 -3907
rect -1048 -3943 -800 -3941
rect -1048 -3977 -946 -3943
rect -912 -3977 -800 -3943
rect -1048 -3979 -800 -3977
rect -1048 -4013 -1042 -3979
rect -1008 -4013 -840 -3979
rect -806 -4013 -800 -3979
rect -1048 -4015 -800 -4013
rect -1048 -4049 -946 -4015
rect -912 -4049 -800 -4015
rect -1048 -4051 -800 -4049
rect -1048 -4085 -1042 -4051
rect -1008 -4085 -840 -4051
rect -806 -4085 -800 -4051
rect -1048 -4087 -800 -4085
rect -1048 -4121 -946 -4087
rect -912 -4121 -800 -4087
rect -1048 -4123 -800 -4121
rect -1048 -4157 -1042 -4123
rect -1008 -4157 -840 -4123
rect -806 -4157 -800 -4123
rect -1048 -4159 -800 -4157
rect -1048 -4193 -946 -4159
rect -912 -4193 -800 -4159
rect -1048 -4195 -800 -4193
rect -1048 -4229 -1042 -4195
rect -1008 -4229 -840 -4195
rect -806 -4229 -800 -4195
rect -1048 -4231 -800 -4229
rect -1048 -4265 -946 -4231
rect -912 -4265 -800 -4231
rect -1048 -4267 -800 -4265
rect -1048 -4301 -1042 -4267
rect -1008 -4301 -840 -4267
rect -806 -4301 -800 -4267
rect -1048 -4303 -800 -4301
rect -1048 -4337 -946 -4303
rect -912 -4337 -800 -4303
rect -1048 -4339 -800 -4337
rect -1048 -4373 -1042 -4339
rect -1008 -4373 -840 -4339
rect -806 -4373 -800 -4339
rect -1048 -4375 -800 -4373
rect -1048 -4409 -946 -4375
rect -912 -4409 -800 -4375
rect -1048 -4411 -800 -4409
rect -1048 -4445 -1042 -4411
rect -1008 -4445 -840 -4411
rect -806 -4445 -800 -4411
rect -1048 -4447 -800 -4445
rect -1048 -4481 -946 -4447
rect -912 -4481 -800 -4447
rect -1048 -4483 -800 -4481
rect -1048 -4517 -1042 -4483
rect -1008 -4517 -840 -4483
rect -806 -4517 -800 -4483
rect -1048 -4519 -800 -4517
rect -1048 -4553 -946 -4519
rect -912 -4553 -800 -4519
rect -1048 -4555 -800 -4553
rect -1048 -4589 -1042 -4555
rect -1008 -4589 -840 -4555
rect -806 -4589 -800 -4555
rect -1048 -4591 -800 -4589
rect -1048 -4625 -946 -4591
rect -912 -4625 -800 -4591
rect -1048 -4627 -800 -4625
rect -1048 -4661 -1042 -4627
rect -1008 -4661 -840 -4627
rect -806 -4661 -800 -4627
rect -1048 -4663 -800 -4661
rect -1048 -4697 -946 -4663
rect -912 -4697 -800 -4663
rect -1048 -4699 -800 -4697
rect -1048 -4733 -1042 -4699
rect -1008 -4733 -840 -4699
rect -806 -4733 -800 -4699
rect -1048 -4735 -800 -4733
rect -1048 -4769 -946 -4735
rect -912 -4769 -800 -4735
rect -1048 -4771 -800 -4769
rect -1048 -4805 -1042 -4771
rect -1008 -4805 -840 -4771
rect -806 -4805 -800 -4771
rect -1048 -4807 -800 -4805
rect -1048 -4841 -946 -4807
rect -912 -4841 -800 -4807
rect -1048 -4843 -800 -4841
rect -1048 -4877 -1042 -4843
rect -1008 -4877 -840 -4843
rect -806 -4877 -800 -4843
rect -1048 -4879 -800 -4877
rect -1048 -4913 -946 -4879
rect -912 -4913 -800 -4879
rect -1048 -4915 -800 -4913
rect -1048 -4949 -1042 -4915
rect -1008 -4949 -840 -4915
rect -806 -4949 -800 -4915
rect -1048 -4951 -800 -4949
rect -1048 -4985 -946 -4951
rect -912 -4985 -800 -4951
rect -1048 -4987 -800 -4985
rect -1540 -5023 -1416 -5021
rect -1540 -5057 -1528 -5023
rect -1494 -5057 -1416 -5023
rect -1048 -5021 -1042 -4987
rect -1008 -5021 -840 -4987
rect -806 -5021 -800 -4987
tri -710 5000 -690 5020 se
rect -690 5000 -542 5020
tri -542 5000 -522 5020 sw
rect -710 4985 -522 5000
rect -710 -4985 -669 4985
rect -563 -4985 -522 4985
rect -710 -5000 -522 -4985
tri -710 -5020 -690 -5000 ne
rect -690 -5020 -542 -5000
tri -542 -5020 -522 -5000 nw
rect -432 4987 -426 5021
rect -392 4987 -224 5021
rect -190 4987 -184 5021
rect 184 5023 286 5057
rect 320 5023 432 5057
tri 432 5044 445 5057 nw
tri 787 5044 800 5057 ne
rect 184 5021 432 5023
rect -432 4985 -184 4987
rect -432 4951 -330 4985
rect -296 4951 -184 4985
rect -432 4949 -184 4951
rect -432 4915 -426 4949
rect -392 4915 -224 4949
rect -190 4915 -184 4949
rect -432 4913 -184 4915
rect -432 4879 -330 4913
rect -296 4879 -184 4913
rect -432 4877 -184 4879
rect -432 4843 -426 4877
rect -392 4843 -224 4877
rect -190 4843 -184 4877
rect -432 4841 -184 4843
rect -432 4807 -330 4841
rect -296 4807 -184 4841
rect -432 4805 -184 4807
rect -432 4771 -426 4805
rect -392 4771 -224 4805
rect -190 4771 -184 4805
rect -432 4769 -184 4771
rect -432 4735 -330 4769
rect -296 4735 -184 4769
rect -432 4733 -184 4735
rect -432 4699 -426 4733
rect -392 4699 -224 4733
rect -190 4699 -184 4733
rect -432 4697 -184 4699
rect -432 4663 -330 4697
rect -296 4663 -184 4697
rect -432 4661 -184 4663
rect -432 4627 -426 4661
rect -392 4627 -224 4661
rect -190 4627 -184 4661
rect -432 4625 -184 4627
rect -432 4591 -330 4625
rect -296 4591 -184 4625
rect -432 4589 -184 4591
rect -432 4555 -426 4589
rect -392 4555 -224 4589
rect -190 4555 -184 4589
rect -432 4553 -184 4555
rect -432 4519 -330 4553
rect -296 4519 -184 4553
rect -432 4517 -184 4519
rect -432 4483 -426 4517
rect -392 4483 -224 4517
rect -190 4483 -184 4517
rect -432 4481 -184 4483
rect -432 4447 -330 4481
rect -296 4447 -184 4481
rect -432 4445 -184 4447
rect -432 4411 -426 4445
rect -392 4411 -224 4445
rect -190 4411 -184 4445
rect -432 4409 -184 4411
rect -432 4375 -330 4409
rect -296 4375 -184 4409
rect -432 4373 -184 4375
rect -432 4339 -426 4373
rect -392 4339 -224 4373
rect -190 4339 -184 4373
rect -432 4337 -184 4339
rect -432 4303 -330 4337
rect -296 4303 -184 4337
rect -432 4301 -184 4303
rect -432 4267 -426 4301
rect -392 4267 -224 4301
rect -190 4267 -184 4301
rect -432 4265 -184 4267
rect -432 4231 -330 4265
rect -296 4231 -184 4265
rect -432 4229 -184 4231
rect -432 4195 -426 4229
rect -392 4195 -224 4229
rect -190 4195 -184 4229
rect -432 4193 -184 4195
rect -432 4159 -330 4193
rect -296 4159 -184 4193
rect -432 4157 -184 4159
rect -432 4123 -426 4157
rect -392 4123 -224 4157
rect -190 4123 -184 4157
rect -432 4121 -184 4123
rect -432 4087 -330 4121
rect -296 4087 -184 4121
rect -432 4085 -184 4087
rect -432 4051 -426 4085
rect -392 4051 -224 4085
rect -190 4051 -184 4085
rect -432 4049 -184 4051
rect -432 4015 -330 4049
rect -296 4015 -184 4049
rect -432 4013 -184 4015
rect -432 3979 -426 4013
rect -392 3979 -224 4013
rect -190 3979 -184 4013
rect -432 3977 -184 3979
rect -432 3943 -330 3977
rect -296 3943 -184 3977
rect -432 3941 -184 3943
rect -432 3907 -426 3941
rect -392 3907 -224 3941
rect -190 3907 -184 3941
rect -432 3905 -184 3907
rect -432 3871 -330 3905
rect -296 3871 -184 3905
rect -432 3869 -184 3871
rect -432 3835 -426 3869
rect -392 3835 -224 3869
rect -190 3835 -184 3869
rect -432 3833 -184 3835
rect -432 3799 -330 3833
rect -296 3799 -184 3833
rect -432 3797 -184 3799
rect -432 3763 -426 3797
rect -392 3763 -224 3797
rect -190 3763 -184 3797
rect -432 3761 -184 3763
rect -432 3727 -330 3761
rect -296 3727 -184 3761
rect -432 3725 -184 3727
rect -432 3691 -426 3725
rect -392 3691 -224 3725
rect -190 3691 -184 3725
rect -432 3689 -184 3691
rect -432 3655 -330 3689
rect -296 3655 -184 3689
rect -432 3653 -184 3655
rect -432 3619 -426 3653
rect -392 3619 -224 3653
rect -190 3619 -184 3653
rect -432 3617 -184 3619
rect -432 3583 -330 3617
rect -296 3583 -184 3617
rect -432 3581 -184 3583
rect -432 3547 -426 3581
rect -392 3547 -224 3581
rect -190 3547 -184 3581
rect -432 3545 -184 3547
rect -432 3511 -330 3545
rect -296 3511 -184 3545
rect -432 3509 -184 3511
rect -432 3475 -426 3509
rect -392 3475 -224 3509
rect -190 3475 -184 3509
rect -432 3473 -184 3475
rect -432 3439 -330 3473
rect -296 3439 -184 3473
rect -432 3437 -184 3439
rect -432 3403 -426 3437
rect -392 3403 -224 3437
rect -190 3403 -184 3437
rect -432 3401 -184 3403
rect -432 3367 -330 3401
rect -296 3367 -184 3401
rect -432 3365 -184 3367
rect -432 3331 -426 3365
rect -392 3331 -224 3365
rect -190 3331 -184 3365
rect -432 3329 -184 3331
rect -432 3295 -330 3329
rect -296 3295 -184 3329
rect -432 3293 -184 3295
rect -432 3259 -426 3293
rect -392 3259 -224 3293
rect -190 3259 -184 3293
rect -432 3257 -184 3259
rect -432 3223 -330 3257
rect -296 3223 -184 3257
rect -432 3221 -184 3223
rect -432 3187 -426 3221
rect -392 3187 -224 3221
rect -190 3187 -184 3221
rect -432 3185 -184 3187
rect -432 3151 -330 3185
rect -296 3151 -184 3185
rect -432 3149 -184 3151
rect -432 3115 -426 3149
rect -392 3115 -224 3149
rect -190 3115 -184 3149
rect -432 3113 -184 3115
rect -432 3079 -330 3113
rect -296 3079 -184 3113
rect -432 3077 -184 3079
rect -432 3043 -426 3077
rect -392 3043 -224 3077
rect -190 3043 -184 3077
rect -432 3041 -184 3043
rect -432 3007 -330 3041
rect -296 3007 -184 3041
rect -432 3005 -184 3007
rect -432 2971 -426 3005
rect -392 2971 -224 3005
rect -190 2971 -184 3005
rect -432 2969 -184 2971
rect -432 2935 -330 2969
rect -296 2935 -184 2969
rect -432 2933 -184 2935
rect -432 2899 -426 2933
rect -392 2899 -224 2933
rect -190 2899 -184 2933
rect -432 2897 -184 2899
rect -432 2863 -330 2897
rect -296 2863 -184 2897
rect -432 2861 -184 2863
rect -432 2827 -426 2861
rect -392 2827 -224 2861
rect -190 2827 -184 2861
rect -432 2825 -184 2827
rect -432 2791 -330 2825
rect -296 2791 -184 2825
rect -432 2789 -184 2791
rect -432 2755 -426 2789
rect -392 2755 -224 2789
rect -190 2755 -184 2789
rect -432 2753 -184 2755
rect -432 2719 -330 2753
rect -296 2719 -184 2753
rect -432 2717 -184 2719
rect -432 2683 -426 2717
rect -392 2683 -224 2717
rect -190 2683 -184 2717
rect -432 2681 -184 2683
rect -432 2647 -330 2681
rect -296 2647 -184 2681
rect -432 2645 -184 2647
rect -432 2611 -426 2645
rect -392 2611 -224 2645
rect -190 2611 -184 2645
rect -432 2609 -184 2611
rect -432 2575 -330 2609
rect -296 2575 -184 2609
rect -432 2573 -184 2575
rect -432 2539 -426 2573
rect -392 2539 -224 2573
rect -190 2539 -184 2573
rect -432 2537 -184 2539
rect -432 2503 -330 2537
rect -296 2503 -184 2537
rect -432 2501 -184 2503
rect -432 2467 -426 2501
rect -392 2467 -224 2501
rect -190 2467 -184 2501
rect -432 2465 -184 2467
rect -432 2431 -330 2465
rect -296 2431 -184 2465
rect -432 2429 -184 2431
rect -432 2395 -426 2429
rect -392 2395 -224 2429
rect -190 2395 -184 2429
rect -432 2393 -184 2395
rect -432 2359 -330 2393
rect -296 2359 -184 2393
rect -432 2357 -184 2359
rect -432 2323 -426 2357
rect -392 2323 -224 2357
rect -190 2323 -184 2357
rect -432 2321 -184 2323
rect -432 2287 -330 2321
rect -296 2287 -184 2321
rect -432 2285 -184 2287
rect -432 2251 -426 2285
rect -392 2251 -224 2285
rect -190 2251 -184 2285
rect -432 2249 -184 2251
rect -432 2215 -330 2249
rect -296 2215 -184 2249
rect -432 2213 -184 2215
rect -432 2179 -426 2213
rect -392 2179 -224 2213
rect -190 2179 -184 2213
rect -432 2177 -184 2179
rect -432 2143 -330 2177
rect -296 2143 -184 2177
rect -432 2141 -184 2143
rect -432 2107 -426 2141
rect -392 2107 -224 2141
rect -190 2107 -184 2141
rect -432 2105 -184 2107
rect -432 2071 -330 2105
rect -296 2071 -184 2105
rect -432 2069 -184 2071
rect -432 2035 -426 2069
rect -392 2035 -224 2069
rect -190 2035 -184 2069
rect -432 2033 -184 2035
rect -432 1999 -330 2033
rect -296 1999 -184 2033
rect -432 1997 -184 1999
rect -432 1963 -426 1997
rect -392 1963 -224 1997
rect -190 1963 -184 1997
rect -432 1961 -184 1963
rect -432 1927 -330 1961
rect -296 1927 -184 1961
rect -432 1925 -184 1927
rect -432 1891 -426 1925
rect -392 1891 -224 1925
rect -190 1891 -184 1925
rect -432 1889 -184 1891
rect -432 1855 -330 1889
rect -296 1855 -184 1889
rect -432 1853 -184 1855
rect -432 1819 -426 1853
rect -392 1819 -224 1853
rect -190 1819 -184 1853
rect -432 1817 -184 1819
rect -432 1783 -330 1817
rect -296 1783 -184 1817
rect -432 1781 -184 1783
rect -432 1747 -426 1781
rect -392 1747 -224 1781
rect -190 1747 -184 1781
rect -432 1745 -184 1747
rect -432 1711 -330 1745
rect -296 1711 -184 1745
rect -432 1709 -184 1711
rect -432 1675 -426 1709
rect -392 1675 -224 1709
rect -190 1675 -184 1709
rect -432 1673 -184 1675
rect -432 1639 -330 1673
rect -296 1639 -184 1673
rect -432 1637 -184 1639
rect -432 1603 -426 1637
rect -392 1603 -224 1637
rect -190 1603 -184 1637
rect -432 1601 -184 1603
rect -432 1567 -330 1601
rect -296 1567 -184 1601
rect -432 1565 -184 1567
rect -432 1531 -426 1565
rect -392 1531 -224 1565
rect -190 1531 -184 1565
rect -432 1529 -184 1531
rect -432 1495 -330 1529
rect -296 1495 -184 1529
rect -432 1493 -184 1495
rect -432 1459 -426 1493
rect -392 1459 -224 1493
rect -190 1459 -184 1493
rect -432 1457 -184 1459
rect -432 1423 -330 1457
rect -296 1423 -184 1457
rect -432 1421 -184 1423
rect -432 1387 -426 1421
rect -392 1387 -224 1421
rect -190 1387 -184 1421
rect -432 1385 -184 1387
rect -432 1351 -330 1385
rect -296 1351 -184 1385
rect -432 1349 -184 1351
rect -432 1315 -426 1349
rect -392 1315 -224 1349
rect -190 1315 -184 1349
rect -432 1313 -184 1315
rect -432 1279 -330 1313
rect -296 1279 -184 1313
rect -432 1277 -184 1279
rect -432 1243 -426 1277
rect -392 1243 -224 1277
rect -190 1243 -184 1277
rect -432 1241 -184 1243
rect -432 1207 -330 1241
rect -296 1207 -184 1241
rect -432 1205 -184 1207
rect -432 1171 -426 1205
rect -392 1171 -224 1205
rect -190 1171 -184 1205
rect -432 1169 -184 1171
rect -432 1135 -330 1169
rect -296 1135 -184 1169
rect -432 1133 -184 1135
rect -432 1099 -426 1133
rect -392 1099 -224 1133
rect -190 1099 -184 1133
rect -432 1097 -184 1099
rect -432 1063 -330 1097
rect -296 1063 -184 1097
rect -432 1061 -184 1063
rect -432 1027 -426 1061
rect -392 1027 -224 1061
rect -190 1027 -184 1061
rect -432 1025 -184 1027
rect -432 991 -330 1025
rect -296 991 -184 1025
rect -432 989 -184 991
rect -432 955 -426 989
rect -392 955 -224 989
rect -190 955 -184 989
rect -432 953 -184 955
rect -432 919 -330 953
rect -296 919 -184 953
rect -432 917 -184 919
rect -432 883 -426 917
rect -392 883 -224 917
rect -190 883 -184 917
rect -432 881 -184 883
rect -432 847 -330 881
rect -296 847 -184 881
rect -432 845 -184 847
rect -432 811 -426 845
rect -392 811 -224 845
rect -190 811 -184 845
rect -432 809 -184 811
rect -432 775 -330 809
rect -296 775 -184 809
rect -432 773 -184 775
rect -432 739 -426 773
rect -392 739 -224 773
rect -190 739 -184 773
rect -432 737 -184 739
rect -432 703 -330 737
rect -296 703 -184 737
rect -432 701 -184 703
rect -432 667 -426 701
rect -392 667 -224 701
rect -190 667 -184 701
rect -432 665 -184 667
rect -432 631 -330 665
rect -296 631 -184 665
rect -432 629 -184 631
rect -432 595 -426 629
rect -392 595 -224 629
rect -190 595 -184 629
rect -432 593 -184 595
rect -432 559 -330 593
rect -296 559 -184 593
rect -432 557 -184 559
rect -432 523 -426 557
rect -392 523 -224 557
rect -190 523 -184 557
rect -432 521 -184 523
rect -432 487 -330 521
rect -296 487 -184 521
rect -432 485 -184 487
rect -432 451 -426 485
rect -392 451 -224 485
rect -190 451 -184 485
rect -432 449 -184 451
rect -432 415 -330 449
rect -296 415 -184 449
rect -432 413 -184 415
rect -432 379 -426 413
rect -392 379 -224 413
rect -190 379 -184 413
rect -432 377 -184 379
rect -432 343 -330 377
rect -296 343 -184 377
rect -432 341 -184 343
rect -432 307 -426 341
rect -392 307 -224 341
rect -190 307 -184 341
rect -432 305 -184 307
rect -432 271 -330 305
rect -296 271 -184 305
rect -432 269 -184 271
rect -432 235 -426 269
rect -392 235 -224 269
rect -190 235 -184 269
rect -432 233 -184 235
rect -432 199 -330 233
rect -296 199 -184 233
rect -432 197 -184 199
rect -432 163 -426 197
rect -392 163 -224 197
rect -190 163 -184 197
rect -432 161 -184 163
rect -432 127 -330 161
rect -296 127 -184 161
rect -432 125 -184 127
rect -432 91 -426 125
rect -392 91 -224 125
rect -190 91 -184 125
rect -432 89 -184 91
rect -432 55 -330 89
rect -296 55 -184 89
rect -432 53 -184 55
rect -432 19 -426 53
rect -392 19 -224 53
rect -190 19 -184 53
rect -432 17 -184 19
rect -432 -17 -330 17
rect -296 -17 -184 17
rect -432 -19 -184 -17
rect -432 -53 -426 -19
rect -392 -53 -224 -19
rect -190 -53 -184 -19
rect -432 -55 -184 -53
rect -432 -89 -330 -55
rect -296 -89 -184 -55
rect -432 -91 -184 -89
rect -432 -125 -426 -91
rect -392 -125 -224 -91
rect -190 -125 -184 -91
rect -432 -127 -184 -125
rect -432 -161 -330 -127
rect -296 -161 -184 -127
rect -432 -163 -184 -161
rect -432 -197 -426 -163
rect -392 -197 -224 -163
rect -190 -197 -184 -163
rect -432 -199 -184 -197
rect -432 -233 -330 -199
rect -296 -233 -184 -199
rect -432 -235 -184 -233
rect -432 -269 -426 -235
rect -392 -269 -224 -235
rect -190 -269 -184 -235
rect -432 -271 -184 -269
rect -432 -305 -330 -271
rect -296 -305 -184 -271
rect -432 -307 -184 -305
rect -432 -341 -426 -307
rect -392 -341 -224 -307
rect -190 -341 -184 -307
rect -432 -343 -184 -341
rect -432 -377 -330 -343
rect -296 -377 -184 -343
rect -432 -379 -184 -377
rect -432 -413 -426 -379
rect -392 -413 -224 -379
rect -190 -413 -184 -379
rect -432 -415 -184 -413
rect -432 -449 -330 -415
rect -296 -449 -184 -415
rect -432 -451 -184 -449
rect -432 -485 -426 -451
rect -392 -485 -224 -451
rect -190 -485 -184 -451
rect -432 -487 -184 -485
rect -432 -521 -330 -487
rect -296 -521 -184 -487
rect -432 -523 -184 -521
rect -432 -557 -426 -523
rect -392 -557 -224 -523
rect -190 -557 -184 -523
rect -432 -559 -184 -557
rect -432 -593 -330 -559
rect -296 -593 -184 -559
rect -432 -595 -184 -593
rect -432 -629 -426 -595
rect -392 -629 -224 -595
rect -190 -629 -184 -595
rect -432 -631 -184 -629
rect -432 -665 -330 -631
rect -296 -665 -184 -631
rect -432 -667 -184 -665
rect -432 -701 -426 -667
rect -392 -701 -224 -667
rect -190 -701 -184 -667
rect -432 -703 -184 -701
rect -432 -737 -330 -703
rect -296 -737 -184 -703
rect -432 -739 -184 -737
rect -432 -773 -426 -739
rect -392 -773 -224 -739
rect -190 -773 -184 -739
rect -432 -775 -184 -773
rect -432 -809 -330 -775
rect -296 -809 -184 -775
rect -432 -811 -184 -809
rect -432 -845 -426 -811
rect -392 -845 -224 -811
rect -190 -845 -184 -811
rect -432 -847 -184 -845
rect -432 -881 -330 -847
rect -296 -881 -184 -847
rect -432 -883 -184 -881
rect -432 -917 -426 -883
rect -392 -917 -224 -883
rect -190 -917 -184 -883
rect -432 -919 -184 -917
rect -432 -953 -330 -919
rect -296 -953 -184 -919
rect -432 -955 -184 -953
rect -432 -989 -426 -955
rect -392 -989 -224 -955
rect -190 -989 -184 -955
rect -432 -991 -184 -989
rect -432 -1025 -330 -991
rect -296 -1025 -184 -991
rect -432 -1027 -184 -1025
rect -432 -1061 -426 -1027
rect -392 -1061 -224 -1027
rect -190 -1061 -184 -1027
rect -432 -1063 -184 -1061
rect -432 -1097 -330 -1063
rect -296 -1097 -184 -1063
rect -432 -1099 -184 -1097
rect -432 -1133 -426 -1099
rect -392 -1133 -224 -1099
rect -190 -1133 -184 -1099
rect -432 -1135 -184 -1133
rect -432 -1169 -330 -1135
rect -296 -1169 -184 -1135
rect -432 -1171 -184 -1169
rect -432 -1205 -426 -1171
rect -392 -1205 -224 -1171
rect -190 -1205 -184 -1171
rect -432 -1207 -184 -1205
rect -432 -1241 -330 -1207
rect -296 -1241 -184 -1207
rect -432 -1243 -184 -1241
rect -432 -1277 -426 -1243
rect -392 -1277 -224 -1243
rect -190 -1277 -184 -1243
rect -432 -1279 -184 -1277
rect -432 -1313 -330 -1279
rect -296 -1313 -184 -1279
rect -432 -1315 -184 -1313
rect -432 -1349 -426 -1315
rect -392 -1349 -224 -1315
rect -190 -1349 -184 -1315
rect -432 -1351 -184 -1349
rect -432 -1385 -330 -1351
rect -296 -1385 -184 -1351
rect -432 -1387 -184 -1385
rect -432 -1421 -426 -1387
rect -392 -1421 -224 -1387
rect -190 -1421 -184 -1387
rect -432 -1423 -184 -1421
rect -432 -1457 -330 -1423
rect -296 -1457 -184 -1423
rect -432 -1459 -184 -1457
rect -432 -1493 -426 -1459
rect -392 -1493 -224 -1459
rect -190 -1493 -184 -1459
rect -432 -1495 -184 -1493
rect -432 -1529 -330 -1495
rect -296 -1529 -184 -1495
rect -432 -1531 -184 -1529
rect -432 -1565 -426 -1531
rect -392 -1565 -224 -1531
rect -190 -1565 -184 -1531
rect -432 -1567 -184 -1565
rect -432 -1601 -330 -1567
rect -296 -1601 -184 -1567
rect -432 -1603 -184 -1601
rect -432 -1637 -426 -1603
rect -392 -1637 -224 -1603
rect -190 -1637 -184 -1603
rect -432 -1639 -184 -1637
rect -432 -1673 -330 -1639
rect -296 -1673 -184 -1639
rect -432 -1675 -184 -1673
rect -432 -1709 -426 -1675
rect -392 -1709 -224 -1675
rect -190 -1709 -184 -1675
rect -432 -1711 -184 -1709
rect -432 -1745 -330 -1711
rect -296 -1745 -184 -1711
rect -432 -1747 -184 -1745
rect -432 -1781 -426 -1747
rect -392 -1781 -224 -1747
rect -190 -1781 -184 -1747
rect -432 -1783 -184 -1781
rect -432 -1817 -330 -1783
rect -296 -1817 -184 -1783
rect -432 -1819 -184 -1817
rect -432 -1853 -426 -1819
rect -392 -1853 -224 -1819
rect -190 -1853 -184 -1819
rect -432 -1855 -184 -1853
rect -432 -1889 -330 -1855
rect -296 -1889 -184 -1855
rect -432 -1891 -184 -1889
rect -432 -1925 -426 -1891
rect -392 -1925 -224 -1891
rect -190 -1925 -184 -1891
rect -432 -1927 -184 -1925
rect -432 -1961 -330 -1927
rect -296 -1961 -184 -1927
rect -432 -1963 -184 -1961
rect -432 -1997 -426 -1963
rect -392 -1997 -224 -1963
rect -190 -1997 -184 -1963
rect -432 -1999 -184 -1997
rect -432 -2033 -330 -1999
rect -296 -2033 -184 -1999
rect -432 -2035 -184 -2033
rect -432 -2069 -426 -2035
rect -392 -2069 -224 -2035
rect -190 -2069 -184 -2035
rect -432 -2071 -184 -2069
rect -432 -2105 -330 -2071
rect -296 -2105 -184 -2071
rect -432 -2107 -184 -2105
rect -432 -2141 -426 -2107
rect -392 -2141 -224 -2107
rect -190 -2141 -184 -2107
rect -432 -2143 -184 -2141
rect -432 -2177 -330 -2143
rect -296 -2177 -184 -2143
rect -432 -2179 -184 -2177
rect -432 -2213 -426 -2179
rect -392 -2213 -224 -2179
rect -190 -2213 -184 -2179
rect -432 -2215 -184 -2213
rect -432 -2249 -330 -2215
rect -296 -2249 -184 -2215
rect -432 -2251 -184 -2249
rect -432 -2285 -426 -2251
rect -392 -2285 -224 -2251
rect -190 -2285 -184 -2251
rect -432 -2287 -184 -2285
rect -432 -2321 -330 -2287
rect -296 -2321 -184 -2287
rect -432 -2323 -184 -2321
rect -432 -2357 -426 -2323
rect -392 -2357 -224 -2323
rect -190 -2357 -184 -2323
rect -432 -2359 -184 -2357
rect -432 -2393 -330 -2359
rect -296 -2393 -184 -2359
rect -432 -2395 -184 -2393
rect -432 -2429 -426 -2395
rect -392 -2429 -224 -2395
rect -190 -2429 -184 -2395
rect -432 -2431 -184 -2429
rect -432 -2465 -330 -2431
rect -296 -2465 -184 -2431
rect -432 -2467 -184 -2465
rect -432 -2501 -426 -2467
rect -392 -2501 -224 -2467
rect -190 -2501 -184 -2467
rect -432 -2503 -184 -2501
rect -432 -2537 -330 -2503
rect -296 -2537 -184 -2503
rect -432 -2539 -184 -2537
rect -432 -2573 -426 -2539
rect -392 -2573 -224 -2539
rect -190 -2573 -184 -2539
rect -432 -2575 -184 -2573
rect -432 -2609 -330 -2575
rect -296 -2609 -184 -2575
rect -432 -2611 -184 -2609
rect -432 -2645 -426 -2611
rect -392 -2645 -224 -2611
rect -190 -2645 -184 -2611
rect -432 -2647 -184 -2645
rect -432 -2681 -330 -2647
rect -296 -2681 -184 -2647
rect -432 -2683 -184 -2681
rect -432 -2717 -426 -2683
rect -392 -2717 -224 -2683
rect -190 -2717 -184 -2683
rect -432 -2719 -184 -2717
rect -432 -2753 -330 -2719
rect -296 -2753 -184 -2719
rect -432 -2755 -184 -2753
rect -432 -2789 -426 -2755
rect -392 -2789 -224 -2755
rect -190 -2789 -184 -2755
rect -432 -2791 -184 -2789
rect -432 -2825 -330 -2791
rect -296 -2825 -184 -2791
rect -432 -2827 -184 -2825
rect -432 -2861 -426 -2827
rect -392 -2861 -224 -2827
rect -190 -2861 -184 -2827
rect -432 -2863 -184 -2861
rect -432 -2897 -330 -2863
rect -296 -2897 -184 -2863
rect -432 -2899 -184 -2897
rect -432 -2933 -426 -2899
rect -392 -2933 -224 -2899
rect -190 -2933 -184 -2899
rect -432 -2935 -184 -2933
rect -432 -2969 -330 -2935
rect -296 -2969 -184 -2935
rect -432 -2971 -184 -2969
rect -432 -3005 -426 -2971
rect -392 -3005 -224 -2971
rect -190 -3005 -184 -2971
rect -432 -3007 -184 -3005
rect -432 -3041 -330 -3007
rect -296 -3041 -184 -3007
rect -432 -3043 -184 -3041
rect -432 -3077 -426 -3043
rect -392 -3077 -224 -3043
rect -190 -3077 -184 -3043
rect -432 -3079 -184 -3077
rect -432 -3113 -330 -3079
rect -296 -3113 -184 -3079
rect -432 -3115 -184 -3113
rect -432 -3149 -426 -3115
rect -392 -3149 -224 -3115
rect -190 -3149 -184 -3115
rect -432 -3151 -184 -3149
rect -432 -3185 -330 -3151
rect -296 -3185 -184 -3151
rect -432 -3187 -184 -3185
rect -432 -3221 -426 -3187
rect -392 -3221 -224 -3187
rect -190 -3221 -184 -3187
rect -432 -3223 -184 -3221
rect -432 -3257 -330 -3223
rect -296 -3257 -184 -3223
rect -432 -3259 -184 -3257
rect -432 -3293 -426 -3259
rect -392 -3293 -224 -3259
rect -190 -3293 -184 -3259
rect -432 -3295 -184 -3293
rect -432 -3329 -330 -3295
rect -296 -3329 -184 -3295
rect -432 -3331 -184 -3329
rect -432 -3365 -426 -3331
rect -392 -3365 -224 -3331
rect -190 -3365 -184 -3331
rect -432 -3367 -184 -3365
rect -432 -3401 -330 -3367
rect -296 -3401 -184 -3367
rect -432 -3403 -184 -3401
rect -432 -3437 -426 -3403
rect -392 -3437 -224 -3403
rect -190 -3437 -184 -3403
rect -432 -3439 -184 -3437
rect -432 -3473 -330 -3439
rect -296 -3473 -184 -3439
rect -432 -3475 -184 -3473
rect -432 -3509 -426 -3475
rect -392 -3509 -224 -3475
rect -190 -3509 -184 -3475
rect -432 -3511 -184 -3509
rect -432 -3545 -330 -3511
rect -296 -3545 -184 -3511
rect -432 -3547 -184 -3545
rect -432 -3581 -426 -3547
rect -392 -3581 -224 -3547
rect -190 -3581 -184 -3547
rect -432 -3583 -184 -3581
rect -432 -3617 -330 -3583
rect -296 -3617 -184 -3583
rect -432 -3619 -184 -3617
rect -432 -3653 -426 -3619
rect -392 -3653 -224 -3619
rect -190 -3653 -184 -3619
rect -432 -3655 -184 -3653
rect -432 -3689 -330 -3655
rect -296 -3689 -184 -3655
rect -432 -3691 -184 -3689
rect -432 -3725 -426 -3691
rect -392 -3725 -224 -3691
rect -190 -3725 -184 -3691
rect -432 -3727 -184 -3725
rect -432 -3761 -330 -3727
rect -296 -3761 -184 -3727
rect -432 -3763 -184 -3761
rect -432 -3797 -426 -3763
rect -392 -3797 -224 -3763
rect -190 -3797 -184 -3763
rect -432 -3799 -184 -3797
rect -432 -3833 -330 -3799
rect -296 -3833 -184 -3799
rect -432 -3835 -184 -3833
rect -432 -3869 -426 -3835
rect -392 -3869 -224 -3835
rect -190 -3869 -184 -3835
rect -432 -3871 -184 -3869
rect -432 -3905 -330 -3871
rect -296 -3905 -184 -3871
rect -432 -3907 -184 -3905
rect -432 -3941 -426 -3907
rect -392 -3941 -224 -3907
rect -190 -3941 -184 -3907
rect -432 -3943 -184 -3941
rect -432 -3977 -330 -3943
rect -296 -3977 -184 -3943
rect -432 -3979 -184 -3977
rect -432 -4013 -426 -3979
rect -392 -4013 -224 -3979
rect -190 -4013 -184 -3979
rect -432 -4015 -184 -4013
rect -432 -4049 -330 -4015
rect -296 -4049 -184 -4015
rect -432 -4051 -184 -4049
rect -432 -4085 -426 -4051
rect -392 -4085 -224 -4051
rect -190 -4085 -184 -4051
rect -432 -4087 -184 -4085
rect -432 -4121 -330 -4087
rect -296 -4121 -184 -4087
rect -432 -4123 -184 -4121
rect -432 -4157 -426 -4123
rect -392 -4157 -224 -4123
rect -190 -4157 -184 -4123
rect -432 -4159 -184 -4157
rect -432 -4193 -330 -4159
rect -296 -4193 -184 -4159
rect -432 -4195 -184 -4193
rect -432 -4229 -426 -4195
rect -392 -4229 -224 -4195
rect -190 -4229 -184 -4195
rect -432 -4231 -184 -4229
rect -432 -4265 -330 -4231
rect -296 -4265 -184 -4231
rect -432 -4267 -184 -4265
rect -432 -4301 -426 -4267
rect -392 -4301 -224 -4267
rect -190 -4301 -184 -4267
rect -432 -4303 -184 -4301
rect -432 -4337 -330 -4303
rect -296 -4337 -184 -4303
rect -432 -4339 -184 -4337
rect -432 -4373 -426 -4339
rect -392 -4373 -224 -4339
rect -190 -4373 -184 -4339
rect -432 -4375 -184 -4373
rect -432 -4409 -330 -4375
rect -296 -4409 -184 -4375
rect -432 -4411 -184 -4409
rect -432 -4445 -426 -4411
rect -392 -4445 -224 -4411
rect -190 -4445 -184 -4411
rect -432 -4447 -184 -4445
rect -432 -4481 -330 -4447
rect -296 -4481 -184 -4447
rect -432 -4483 -184 -4481
rect -432 -4517 -426 -4483
rect -392 -4517 -224 -4483
rect -190 -4517 -184 -4483
rect -432 -4519 -184 -4517
rect -432 -4553 -330 -4519
rect -296 -4553 -184 -4519
rect -432 -4555 -184 -4553
rect -432 -4589 -426 -4555
rect -392 -4589 -224 -4555
rect -190 -4589 -184 -4555
rect -432 -4591 -184 -4589
rect -432 -4625 -330 -4591
rect -296 -4625 -184 -4591
rect -432 -4627 -184 -4625
rect -432 -4661 -426 -4627
rect -392 -4661 -224 -4627
rect -190 -4661 -184 -4627
rect -432 -4663 -184 -4661
rect -432 -4697 -330 -4663
rect -296 -4697 -184 -4663
rect -432 -4699 -184 -4697
rect -432 -4733 -426 -4699
rect -392 -4733 -224 -4699
rect -190 -4733 -184 -4699
rect -432 -4735 -184 -4733
rect -432 -4769 -330 -4735
rect -296 -4769 -184 -4735
rect -432 -4771 -184 -4769
rect -432 -4805 -426 -4771
rect -392 -4805 -224 -4771
rect -190 -4805 -184 -4771
rect -432 -4807 -184 -4805
rect -432 -4841 -330 -4807
rect -296 -4841 -184 -4807
rect -432 -4843 -184 -4841
rect -432 -4877 -426 -4843
rect -392 -4877 -224 -4843
rect -190 -4877 -184 -4843
rect -432 -4879 -184 -4877
rect -432 -4913 -330 -4879
rect -296 -4913 -184 -4879
rect -432 -4915 -184 -4913
rect -432 -4949 -426 -4915
rect -392 -4949 -224 -4915
rect -190 -4949 -184 -4915
rect -432 -4951 -184 -4949
rect -432 -4985 -330 -4951
rect -296 -4985 -184 -4951
rect -432 -4987 -184 -4985
rect -1048 -5023 -800 -5021
tri -1416 -5057 -1403 -5044 sw
tri -1061 -5057 -1048 -5044 se
rect -1048 -5057 -946 -5023
rect -912 -5057 -800 -5023
rect -432 -5021 -426 -4987
rect -392 -5021 -224 -4987
rect -190 -5021 -184 -4987
tri -94 5000 -74 5020 se
rect -74 5000 74 5020
tri 74 5000 94 5020 sw
rect -94 4985 94 5000
rect -94 -4985 -53 4985
rect 53 -4985 94 4985
rect -94 -5000 94 -4985
tri -94 -5020 -74 -5000 ne
rect -74 -5020 74 -5000
tri 74 -5020 94 -5000 nw
rect 184 4987 190 5021
rect 224 4987 392 5021
rect 426 4987 432 5021
rect 800 5023 902 5057
rect 936 5023 1048 5057
tri 1048 5044 1061 5057 nw
tri 1403 5044 1416 5057 ne
rect 800 5021 1048 5023
rect 184 4985 432 4987
rect 184 4951 286 4985
rect 320 4951 432 4985
rect 184 4949 432 4951
rect 184 4915 190 4949
rect 224 4915 392 4949
rect 426 4915 432 4949
rect 184 4913 432 4915
rect 184 4879 286 4913
rect 320 4879 432 4913
rect 184 4877 432 4879
rect 184 4843 190 4877
rect 224 4843 392 4877
rect 426 4843 432 4877
rect 184 4841 432 4843
rect 184 4807 286 4841
rect 320 4807 432 4841
rect 184 4805 432 4807
rect 184 4771 190 4805
rect 224 4771 392 4805
rect 426 4771 432 4805
rect 184 4769 432 4771
rect 184 4735 286 4769
rect 320 4735 432 4769
rect 184 4733 432 4735
rect 184 4699 190 4733
rect 224 4699 392 4733
rect 426 4699 432 4733
rect 184 4697 432 4699
rect 184 4663 286 4697
rect 320 4663 432 4697
rect 184 4661 432 4663
rect 184 4627 190 4661
rect 224 4627 392 4661
rect 426 4627 432 4661
rect 184 4625 432 4627
rect 184 4591 286 4625
rect 320 4591 432 4625
rect 184 4589 432 4591
rect 184 4555 190 4589
rect 224 4555 392 4589
rect 426 4555 432 4589
rect 184 4553 432 4555
rect 184 4519 286 4553
rect 320 4519 432 4553
rect 184 4517 432 4519
rect 184 4483 190 4517
rect 224 4483 392 4517
rect 426 4483 432 4517
rect 184 4481 432 4483
rect 184 4447 286 4481
rect 320 4447 432 4481
rect 184 4445 432 4447
rect 184 4411 190 4445
rect 224 4411 392 4445
rect 426 4411 432 4445
rect 184 4409 432 4411
rect 184 4375 286 4409
rect 320 4375 432 4409
rect 184 4373 432 4375
rect 184 4339 190 4373
rect 224 4339 392 4373
rect 426 4339 432 4373
rect 184 4337 432 4339
rect 184 4303 286 4337
rect 320 4303 432 4337
rect 184 4301 432 4303
rect 184 4267 190 4301
rect 224 4267 392 4301
rect 426 4267 432 4301
rect 184 4265 432 4267
rect 184 4231 286 4265
rect 320 4231 432 4265
rect 184 4229 432 4231
rect 184 4195 190 4229
rect 224 4195 392 4229
rect 426 4195 432 4229
rect 184 4193 432 4195
rect 184 4159 286 4193
rect 320 4159 432 4193
rect 184 4157 432 4159
rect 184 4123 190 4157
rect 224 4123 392 4157
rect 426 4123 432 4157
rect 184 4121 432 4123
rect 184 4087 286 4121
rect 320 4087 432 4121
rect 184 4085 432 4087
rect 184 4051 190 4085
rect 224 4051 392 4085
rect 426 4051 432 4085
rect 184 4049 432 4051
rect 184 4015 286 4049
rect 320 4015 432 4049
rect 184 4013 432 4015
rect 184 3979 190 4013
rect 224 3979 392 4013
rect 426 3979 432 4013
rect 184 3977 432 3979
rect 184 3943 286 3977
rect 320 3943 432 3977
rect 184 3941 432 3943
rect 184 3907 190 3941
rect 224 3907 392 3941
rect 426 3907 432 3941
rect 184 3905 432 3907
rect 184 3871 286 3905
rect 320 3871 432 3905
rect 184 3869 432 3871
rect 184 3835 190 3869
rect 224 3835 392 3869
rect 426 3835 432 3869
rect 184 3833 432 3835
rect 184 3799 286 3833
rect 320 3799 432 3833
rect 184 3797 432 3799
rect 184 3763 190 3797
rect 224 3763 392 3797
rect 426 3763 432 3797
rect 184 3761 432 3763
rect 184 3727 286 3761
rect 320 3727 432 3761
rect 184 3725 432 3727
rect 184 3691 190 3725
rect 224 3691 392 3725
rect 426 3691 432 3725
rect 184 3689 432 3691
rect 184 3655 286 3689
rect 320 3655 432 3689
rect 184 3653 432 3655
rect 184 3619 190 3653
rect 224 3619 392 3653
rect 426 3619 432 3653
rect 184 3617 432 3619
rect 184 3583 286 3617
rect 320 3583 432 3617
rect 184 3581 432 3583
rect 184 3547 190 3581
rect 224 3547 392 3581
rect 426 3547 432 3581
rect 184 3545 432 3547
rect 184 3511 286 3545
rect 320 3511 432 3545
rect 184 3509 432 3511
rect 184 3475 190 3509
rect 224 3475 392 3509
rect 426 3475 432 3509
rect 184 3473 432 3475
rect 184 3439 286 3473
rect 320 3439 432 3473
rect 184 3437 432 3439
rect 184 3403 190 3437
rect 224 3403 392 3437
rect 426 3403 432 3437
rect 184 3401 432 3403
rect 184 3367 286 3401
rect 320 3367 432 3401
rect 184 3365 432 3367
rect 184 3331 190 3365
rect 224 3331 392 3365
rect 426 3331 432 3365
rect 184 3329 432 3331
rect 184 3295 286 3329
rect 320 3295 432 3329
rect 184 3293 432 3295
rect 184 3259 190 3293
rect 224 3259 392 3293
rect 426 3259 432 3293
rect 184 3257 432 3259
rect 184 3223 286 3257
rect 320 3223 432 3257
rect 184 3221 432 3223
rect 184 3187 190 3221
rect 224 3187 392 3221
rect 426 3187 432 3221
rect 184 3185 432 3187
rect 184 3151 286 3185
rect 320 3151 432 3185
rect 184 3149 432 3151
rect 184 3115 190 3149
rect 224 3115 392 3149
rect 426 3115 432 3149
rect 184 3113 432 3115
rect 184 3079 286 3113
rect 320 3079 432 3113
rect 184 3077 432 3079
rect 184 3043 190 3077
rect 224 3043 392 3077
rect 426 3043 432 3077
rect 184 3041 432 3043
rect 184 3007 286 3041
rect 320 3007 432 3041
rect 184 3005 432 3007
rect 184 2971 190 3005
rect 224 2971 392 3005
rect 426 2971 432 3005
rect 184 2969 432 2971
rect 184 2935 286 2969
rect 320 2935 432 2969
rect 184 2933 432 2935
rect 184 2899 190 2933
rect 224 2899 392 2933
rect 426 2899 432 2933
rect 184 2897 432 2899
rect 184 2863 286 2897
rect 320 2863 432 2897
rect 184 2861 432 2863
rect 184 2827 190 2861
rect 224 2827 392 2861
rect 426 2827 432 2861
rect 184 2825 432 2827
rect 184 2791 286 2825
rect 320 2791 432 2825
rect 184 2789 432 2791
rect 184 2755 190 2789
rect 224 2755 392 2789
rect 426 2755 432 2789
rect 184 2753 432 2755
rect 184 2719 286 2753
rect 320 2719 432 2753
rect 184 2717 432 2719
rect 184 2683 190 2717
rect 224 2683 392 2717
rect 426 2683 432 2717
rect 184 2681 432 2683
rect 184 2647 286 2681
rect 320 2647 432 2681
rect 184 2645 432 2647
rect 184 2611 190 2645
rect 224 2611 392 2645
rect 426 2611 432 2645
rect 184 2609 432 2611
rect 184 2575 286 2609
rect 320 2575 432 2609
rect 184 2573 432 2575
rect 184 2539 190 2573
rect 224 2539 392 2573
rect 426 2539 432 2573
rect 184 2537 432 2539
rect 184 2503 286 2537
rect 320 2503 432 2537
rect 184 2501 432 2503
rect 184 2467 190 2501
rect 224 2467 392 2501
rect 426 2467 432 2501
rect 184 2465 432 2467
rect 184 2431 286 2465
rect 320 2431 432 2465
rect 184 2429 432 2431
rect 184 2395 190 2429
rect 224 2395 392 2429
rect 426 2395 432 2429
rect 184 2393 432 2395
rect 184 2359 286 2393
rect 320 2359 432 2393
rect 184 2357 432 2359
rect 184 2323 190 2357
rect 224 2323 392 2357
rect 426 2323 432 2357
rect 184 2321 432 2323
rect 184 2287 286 2321
rect 320 2287 432 2321
rect 184 2285 432 2287
rect 184 2251 190 2285
rect 224 2251 392 2285
rect 426 2251 432 2285
rect 184 2249 432 2251
rect 184 2215 286 2249
rect 320 2215 432 2249
rect 184 2213 432 2215
rect 184 2179 190 2213
rect 224 2179 392 2213
rect 426 2179 432 2213
rect 184 2177 432 2179
rect 184 2143 286 2177
rect 320 2143 432 2177
rect 184 2141 432 2143
rect 184 2107 190 2141
rect 224 2107 392 2141
rect 426 2107 432 2141
rect 184 2105 432 2107
rect 184 2071 286 2105
rect 320 2071 432 2105
rect 184 2069 432 2071
rect 184 2035 190 2069
rect 224 2035 392 2069
rect 426 2035 432 2069
rect 184 2033 432 2035
rect 184 1999 286 2033
rect 320 1999 432 2033
rect 184 1997 432 1999
rect 184 1963 190 1997
rect 224 1963 392 1997
rect 426 1963 432 1997
rect 184 1961 432 1963
rect 184 1927 286 1961
rect 320 1927 432 1961
rect 184 1925 432 1927
rect 184 1891 190 1925
rect 224 1891 392 1925
rect 426 1891 432 1925
rect 184 1889 432 1891
rect 184 1855 286 1889
rect 320 1855 432 1889
rect 184 1853 432 1855
rect 184 1819 190 1853
rect 224 1819 392 1853
rect 426 1819 432 1853
rect 184 1817 432 1819
rect 184 1783 286 1817
rect 320 1783 432 1817
rect 184 1781 432 1783
rect 184 1747 190 1781
rect 224 1747 392 1781
rect 426 1747 432 1781
rect 184 1745 432 1747
rect 184 1711 286 1745
rect 320 1711 432 1745
rect 184 1709 432 1711
rect 184 1675 190 1709
rect 224 1675 392 1709
rect 426 1675 432 1709
rect 184 1673 432 1675
rect 184 1639 286 1673
rect 320 1639 432 1673
rect 184 1637 432 1639
rect 184 1603 190 1637
rect 224 1603 392 1637
rect 426 1603 432 1637
rect 184 1601 432 1603
rect 184 1567 286 1601
rect 320 1567 432 1601
rect 184 1565 432 1567
rect 184 1531 190 1565
rect 224 1531 392 1565
rect 426 1531 432 1565
rect 184 1529 432 1531
rect 184 1495 286 1529
rect 320 1495 432 1529
rect 184 1493 432 1495
rect 184 1459 190 1493
rect 224 1459 392 1493
rect 426 1459 432 1493
rect 184 1457 432 1459
rect 184 1423 286 1457
rect 320 1423 432 1457
rect 184 1421 432 1423
rect 184 1387 190 1421
rect 224 1387 392 1421
rect 426 1387 432 1421
rect 184 1385 432 1387
rect 184 1351 286 1385
rect 320 1351 432 1385
rect 184 1349 432 1351
rect 184 1315 190 1349
rect 224 1315 392 1349
rect 426 1315 432 1349
rect 184 1313 432 1315
rect 184 1279 286 1313
rect 320 1279 432 1313
rect 184 1277 432 1279
rect 184 1243 190 1277
rect 224 1243 392 1277
rect 426 1243 432 1277
rect 184 1241 432 1243
rect 184 1207 286 1241
rect 320 1207 432 1241
rect 184 1205 432 1207
rect 184 1171 190 1205
rect 224 1171 392 1205
rect 426 1171 432 1205
rect 184 1169 432 1171
rect 184 1135 286 1169
rect 320 1135 432 1169
rect 184 1133 432 1135
rect 184 1099 190 1133
rect 224 1099 392 1133
rect 426 1099 432 1133
rect 184 1097 432 1099
rect 184 1063 286 1097
rect 320 1063 432 1097
rect 184 1061 432 1063
rect 184 1027 190 1061
rect 224 1027 392 1061
rect 426 1027 432 1061
rect 184 1025 432 1027
rect 184 991 286 1025
rect 320 991 432 1025
rect 184 989 432 991
rect 184 955 190 989
rect 224 955 392 989
rect 426 955 432 989
rect 184 953 432 955
rect 184 919 286 953
rect 320 919 432 953
rect 184 917 432 919
rect 184 883 190 917
rect 224 883 392 917
rect 426 883 432 917
rect 184 881 432 883
rect 184 847 286 881
rect 320 847 432 881
rect 184 845 432 847
rect 184 811 190 845
rect 224 811 392 845
rect 426 811 432 845
rect 184 809 432 811
rect 184 775 286 809
rect 320 775 432 809
rect 184 773 432 775
rect 184 739 190 773
rect 224 739 392 773
rect 426 739 432 773
rect 184 737 432 739
rect 184 703 286 737
rect 320 703 432 737
rect 184 701 432 703
rect 184 667 190 701
rect 224 667 392 701
rect 426 667 432 701
rect 184 665 432 667
rect 184 631 286 665
rect 320 631 432 665
rect 184 629 432 631
rect 184 595 190 629
rect 224 595 392 629
rect 426 595 432 629
rect 184 593 432 595
rect 184 559 286 593
rect 320 559 432 593
rect 184 557 432 559
rect 184 523 190 557
rect 224 523 392 557
rect 426 523 432 557
rect 184 521 432 523
rect 184 487 286 521
rect 320 487 432 521
rect 184 485 432 487
rect 184 451 190 485
rect 224 451 392 485
rect 426 451 432 485
rect 184 449 432 451
rect 184 415 286 449
rect 320 415 432 449
rect 184 413 432 415
rect 184 379 190 413
rect 224 379 392 413
rect 426 379 432 413
rect 184 377 432 379
rect 184 343 286 377
rect 320 343 432 377
rect 184 341 432 343
rect 184 307 190 341
rect 224 307 392 341
rect 426 307 432 341
rect 184 305 432 307
rect 184 271 286 305
rect 320 271 432 305
rect 184 269 432 271
rect 184 235 190 269
rect 224 235 392 269
rect 426 235 432 269
rect 184 233 432 235
rect 184 199 286 233
rect 320 199 432 233
rect 184 197 432 199
rect 184 163 190 197
rect 224 163 392 197
rect 426 163 432 197
rect 184 161 432 163
rect 184 127 286 161
rect 320 127 432 161
rect 184 125 432 127
rect 184 91 190 125
rect 224 91 392 125
rect 426 91 432 125
rect 184 89 432 91
rect 184 55 286 89
rect 320 55 432 89
rect 184 53 432 55
rect 184 19 190 53
rect 224 19 392 53
rect 426 19 432 53
rect 184 17 432 19
rect 184 -17 286 17
rect 320 -17 432 17
rect 184 -19 432 -17
rect 184 -53 190 -19
rect 224 -53 392 -19
rect 426 -53 432 -19
rect 184 -55 432 -53
rect 184 -89 286 -55
rect 320 -89 432 -55
rect 184 -91 432 -89
rect 184 -125 190 -91
rect 224 -125 392 -91
rect 426 -125 432 -91
rect 184 -127 432 -125
rect 184 -161 286 -127
rect 320 -161 432 -127
rect 184 -163 432 -161
rect 184 -197 190 -163
rect 224 -197 392 -163
rect 426 -197 432 -163
rect 184 -199 432 -197
rect 184 -233 286 -199
rect 320 -233 432 -199
rect 184 -235 432 -233
rect 184 -269 190 -235
rect 224 -269 392 -235
rect 426 -269 432 -235
rect 184 -271 432 -269
rect 184 -305 286 -271
rect 320 -305 432 -271
rect 184 -307 432 -305
rect 184 -341 190 -307
rect 224 -341 392 -307
rect 426 -341 432 -307
rect 184 -343 432 -341
rect 184 -377 286 -343
rect 320 -377 432 -343
rect 184 -379 432 -377
rect 184 -413 190 -379
rect 224 -413 392 -379
rect 426 -413 432 -379
rect 184 -415 432 -413
rect 184 -449 286 -415
rect 320 -449 432 -415
rect 184 -451 432 -449
rect 184 -485 190 -451
rect 224 -485 392 -451
rect 426 -485 432 -451
rect 184 -487 432 -485
rect 184 -521 286 -487
rect 320 -521 432 -487
rect 184 -523 432 -521
rect 184 -557 190 -523
rect 224 -557 392 -523
rect 426 -557 432 -523
rect 184 -559 432 -557
rect 184 -593 286 -559
rect 320 -593 432 -559
rect 184 -595 432 -593
rect 184 -629 190 -595
rect 224 -629 392 -595
rect 426 -629 432 -595
rect 184 -631 432 -629
rect 184 -665 286 -631
rect 320 -665 432 -631
rect 184 -667 432 -665
rect 184 -701 190 -667
rect 224 -701 392 -667
rect 426 -701 432 -667
rect 184 -703 432 -701
rect 184 -737 286 -703
rect 320 -737 432 -703
rect 184 -739 432 -737
rect 184 -773 190 -739
rect 224 -773 392 -739
rect 426 -773 432 -739
rect 184 -775 432 -773
rect 184 -809 286 -775
rect 320 -809 432 -775
rect 184 -811 432 -809
rect 184 -845 190 -811
rect 224 -845 392 -811
rect 426 -845 432 -811
rect 184 -847 432 -845
rect 184 -881 286 -847
rect 320 -881 432 -847
rect 184 -883 432 -881
rect 184 -917 190 -883
rect 224 -917 392 -883
rect 426 -917 432 -883
rect 184 -919 432 -917
rect 184 -953 286 -919
rect 320 -953 432 -919
rect 184 -955 432 -953
rect 184 -989 190 -955
rect 224 -989 392 -955
rect 426 -989 432 -955
rect 184 -991 432 -989
rect 184 -1025 286 -991
rect 320 -1025 432 -991
rect 184 -1027 432 -1025
rect 184 -1061 190 -1027
rect 224 -1061 392 -1027
rect 426 -1061 432 -1027
rect 184 -1063 432 -1061
rect 184 -1097 286 -1063
rect 320 -1097 432 -1063
rect 184 -1099 432 -1097
rect 184 -1133 190 -1099
rect 224 -1133 392 -1099
rect 426 -1133 432 -1099
rect 184 -1135 432 -1133
rect 184 -1169 286 -1135
rect 320 -1169 432 -1135
rect 184 -1171 432 -1169
rect 184 -1205 190 -1171
rect 224 -1205 392 -1171
rect 426 -1205 432 -1171
rect 184 -1207 432 -1205
rect 184 -1241 286 -1207
rect 320 -1241 432 -1207
rect 184 -1243 432 -1241
rect 184 -1277 190 -1243
rect 224 -1277 392 -1243
rect 426 -1277 432 -1243
rect 184 -1279 432 -1277
rect 184 -1313 286 -1279
rect 320 -1313 432 -1279
rect 184 -1315 432 -1313
rect 184 -1349 190 -1315
rect 224 -1349 392 -1315
rect 426 -1349 432 -1315
rect 184 -1351 432 -1349
rect 184 -1385 286 -1351
rect 320 -1385 432 -1351
rect 184 -1387 432 -1385
rect 184 -1421 190 -1387
rect 224 -1421 392 -1387
rect 426 -1421 432 -1387
rect 184 -1423 432 -1421
rect 184 -1457 286 -1423
rect 320 -1457 432 -1423
rect 184 -1459 432 -1457
rect 184 -1493 190 -1459
rect 224 -1493 392 -1459
rect 426 -1493 432 -1459
rect 184 -1495 432 -1493
rect 184 -1529 286 -1495
rect 320 -1529 432 -1495
rect 184 -1531 432 -1529
rect 184 -1565 190 -1531
rect 224 -1565 392 -1531
rect 426 -1565 432 -1531
rect 184 -1567 432 -1565
rect 184 -1601 286 -1567
rect 320 -1601 432 -1567
rect 184 -1603 432 -1601
rect 184 -1637 190 -1603
rect 224 -1637 392 -1603
rect 426 -1637 432 -1603
rect 184 -1639 432 -1637
rect 184 -1673 286 -1639
rect 320 -1673 432 -1639
rect 184 -1675 432 -1673
rect 184 -1709 190 -1675
rect 224 -1709 392 -1675
rect 426 -1709 432 -1675
rect 184 -1711 432 -1709
rect 184 -1745 286 -1711
rect 320 -1745 432 -1711
rect 184 -1747 432 -1745
rect 184 -1781 190 -1747
rect 224 -1781 392 -1747
rect 426 -1781 432 -1747
rect 184 -1783 432 -1781
rect 184 -1817 286 -1783
rect 320 -1817 432 -1783
rect 184 -1819 432 -1817
rect 184 -1853 190 -1819
rect 224 -1853 392 -1819
rect 426 -1853 432 -1819
rect 184 -1855 432 -1853
rect 184 -1889 286 -1855
rect 320 -1889 432 -1855
rect 184 -1891 432 -1889
rect 184 -1925 190 -1891
rect 224 -1925 392 -1891
rect 426 -1925 432 -1891
rect 184 -1927 432 -1925
rect 184 -1961 286 -1927
rect 320 -1961 432 -1927
rect 184 -1963 432 -1961
rect 184 -1997 190 -1963
rect 224 -1997 392 -1963
rect 426 -1997 432 -1963
rect 184 -1999 432 -1997
rect 184 -2033 286 -1999
rect 320 -2033 432 -1999
rect 184 -2035 432 -2033
rect 184 -2069 190 -2035
rect 224 -2069 392 -2035
rect 426 -2069 432 -2035
rect 184 -2071 432 -2069
rect 184 -2105 286 -2071
rect 320 -2105 432 -2071
rect 184 -2107 432 -2105
rect 184 -2141 190 -2107
rect 224 -2141 392 -2107
rect 426 -2141 432 -2107
rect 184 -2143 432 -2141
rect 184 -2177 286 -2143
rect 320 -2177 432 -2143
rect 184 -2179 432 -2177
rect 184 -2213 190 -2179
rect 224 -2213 392 -2179
rect 426 -2213 432 -2179
rect 184 -2215 432 -2213
rect 184 -2249 286 -2215
rect 320 -2249 432 -2215
rect 184 -2251 432 -2249
rect 184 -2285 190 -2251
rect 224 -2285 392 -2251
rect 426 -2285 432 -2251
rect 184 -2287 432 -2285
rect 184 -2321 286 -2287
rect 320 -2321 432 -2287
rect 184 -2323 432 -2321
rect 184 -2357 190 -2323
rect 224 -2357 392 -2323
rect 426 -2357 432 -2323
rect 184 -2359 432 -2357
rect 184 -2393 286 -2359
rect 320 -2393 432 -2359
rect 184 -2395 432 -2393
rect 184 -2429 190 -2395
rect 224 -2429 392 -2395
rect 426 -2429 432 -2395
rect 184 -2431 432 -2429
rect 184 -2465 286 -2431
rect 320 -2465 432 -2431
rect 184 -2467 432 -2465
rect 184 -2501 190 -2467
rect 224 -2501 392 -2467
rect 426 -2501 432 -2467
rect 184 -2503 432 -2501
rect 184 -2537 286 -2503
rect 320 -2537 432 -2503
rect 184 -2539 432 -2537
rect 184 -2573 190 -2539
rect 224 -2573 392 -2539
rect 426 -2573 432 -2539
rect 184 -2575 432 -2573
rect 184 -2609 286 -2575
rect 320 -2609 432 -2575
rect 184 -2611 432 -2609
rect 184 -2645 190 -2611
rect 224 -2645 392 -2611
rect 426 -2645 432 -2611
rect 184 -2647 432 -2645
rect 184 -2681 286 -2647
rect 320 -2681 432 -2647
rect 184 -2683 432 -2681
rect 184 -2717 190 -2683
rect 224 -2717 392 -2683
rect 426 -2717 432 -2683
rect 184 -2719 432 -2717
rect 184 -2753 286 -2719
rect 320 -2753 432 -2719
rect 184 -2755 432 -2753
rect 184 -2789 190 -2755
rect 224 -2789 392 -2755
rect 426 -2789 432 -2755
rect 184 -2791 432 -2789
rect 184 -2825 286 -2791
rect 320 -2825 432 -2791
rect 184 -2827 432 -2825
rect 184 -2861 190 -2827
rect 224 -2861 392 -2827
rect 426 -2861 432 -2827
rect 184 -2863 432 -2861
rect 184 -2897 286 -2863
rect 320 -2897 432 -2863
rect 184 -2899 432 -2897
rect 184 -2933 190 -2899
rect 224 -2933 392 -2899
rect 426 -2933 432 -2899
rect 184 -2935 432 -2933
rect 184 -2969 286 -2935
rect 320 -2969 432 -2935
rect 184 -2971 432 -2969
rect 184 -3005 190 -2971
rect 224 -3005 392 -2971
rect 426 -3005 432 -2971
rect 184 -3007 432 -3005
rect 184 -3041 286 -3007
rect 320 -3041 432 -3007
rect 184 -3043 432 -3041
rect 184 -3077 190 -3043
rect 224 -3077 392 -3043
rect 426 -3077 432 -3043
rect 184 -3079 432 -3077
rect 184 -3113 286 -3079
rect 320 -3113 432 -3079
rect 184 -3115 432 -3113
rect 184 -3149 190 -3115
rect 224 -3149 392 -3115
rect 426 -3149 432 -3115
rect 184 -3151 432 -3149
rect 184 -3185 286 -3151
rect 320 -3185 432 -3151
rect 184 -3187 432 -3185
rect 184 -3221 190 -3187
rect 224 -3221 392 -3187
rect 426 -3221 432 -3187
rect 184 -3223 432 -3221
rect 184 -3257 286 -3223
rect 320 -3257 432 -3223
rect 184 -3259 432 -3257
rect 184 -3293 190 -3259
rect 224 -3293 392 -3259
rect 426 -3293 432 -3259
rect 184 -3295 432 -3293
rect 184 -3329 286 -3295
rect 320 -3329 432 -3295
rect 184 -3331 432 -3329
rect 184 -3365 190 -3331
rect 224 -3365 392 -3331
rect 426 -3365 432 -3331
rect 184 -3367 432 -3365
rect 184 -3401 286 -3367
rect 320 -3401 432 -3367
rect 184 -3403 432 -3401
rect 184 -3437 190 -3403
rect 224 -3437 392 -3403
rect 426 -3437 432 -3403
rect 184 -3439 432 -3437
rect 184 -3473 286 -3439
rect 320 -3473 432 -3439
rect 184 -3475 432 -3473
rect 184 -3509 190 -3475
rect 224 -3509 392 -3475
rect 426 -3509 432 -3475
rect 184 -3511 432 -3509
rect 184 -3545 286 -3511
rect 320 -3545 432 -3511
rect 184 -3547 432 -3545
rect 184 -3581 190 -3547
rect 224 -3581 392 -3547
rect 426 -3581 432 -3547
rect 184 -3583 432 -3581
rect 184 -3617 286 -3583
rect 320 -3617 432 -3583
rect 184 -3619 432 -3617
rect 184 -3653 190 -3619
rect 224 -3653 392 -3619
rect 426 -3653 432 -3619
rect 184 -3655 432 -3653
rect 184 -3689 286 -3655
rect 320 -3689 432 -3655
rect 184 -3691 432 -3689
rect 184 -3725 190 -3691
rect 224 -3725 392 -3691
rect 426 -3725 432 -3691
rect 184 -3727 432 -3725
rect 184 -3761 286 -3727
rect 320 -3761 432 -3727
rect 184 -3763 432 -3761
rect 184 -3797 190 -3763
rect 224 -3797 392 -3763
rect 426 -3797 432 -3763
rect 184 -3799 432 -3797
rect 184 -3833 286 -3799
rect 320 -3833 432 -3799
rect 184 -3835 432 -3833
rect 184 -3869 190 -3835
rect 224 -3869 392 -3835
rect 426 -3869 432 -3835
rect 184 -3871 432 -3869
rect 184 -3905 286 -3871
rect 320 -3905 432 -3871
rect 184 -3907 432 -3905
rect 184 -3941 190 -3907
rect 224 -3941 392 -3907
rect 426 -3941 432 -3907
rect 184 -3943 432 -3941
rect 184 -3977 286 -3943
rect 320 -3977 432 -3943
rect 184 -3979 432 -3977
rect 184 -4013 190 -3979
rect 224 -4013 392 -3979
rect 426 -4013 432 -3979
rect 184 -4015 432 -4013
rect 184 -4049 286 -4015
rect 320 -4049 432 -4015
rect 184 -4051 432 -4049
rect 184 -4085 190 -4051
rect 224 -4085 392 -4051
rect 426 -4085 432 -4051
rect 184 -4087 432 -4085
rect 184 -4121 286 -4087
rect 320 -4121 432 -4087
rect 184 -4123 432 -4121
rect 184 -4157 190 -4123
rect 224 -4157 392 -4123
rect 426 -4157 432 -4123
rect 184 -4159 432 -4157
rect 184 -4193 286 -4159
rect 320 -4193 432 -4159
rect 184 -4195 432 -4193
rect 184 -4229 190 -4195
rect 224 -4229 392 -4195
rect 426 -4229 432 -4195
rect 184 -4231 432 -4229
rect 184 -4265 286 -4231
rect 320 -4265 432 -4231
rect 184 -4267 432 -4265
rect 184 -4301 190 -4267
rect 224 -4301 392 -4267
rect 426 -4301 432 -4267
rect 184 -4303 432 -4301
rect 184 -4337 286 -4303
rect 320 -4337 432 -4303
rect 184 -4339 432 -4337
rect 184 -4373 190 -4339
rect 224 -4373 392 -4339
rect 426 -4373 432 -4339
rect 184 -4375 432 -4373
rect 184 -4409 286 -4375
rect 320 -4409 432 -4375
rect 184 -4411 432 -4409
rect 184 -4445 190 -4411
rect 224 -4445 392 -4411
rect 426 -4445 432 -4411
rect 184 -4447 432 -4445
rect 184 -4481 286 -4447
rect 320 -4481 432 -4447
rect 184 -4483 432 -4481
rect 184 -4517 190 -4483
rect 224 -4517 392 -4483
rect 426 -4517 432 -4483
rect 184 -4519 432 -4517
rect 184 -4553 286 -4519
rect 320 -4553 432 -4519
rect 184 -4555 432 -4553
rect 184 -4589 190 -4555
rect 224 -4589 392 -4555
rect 426 -4589 432 -4555
rect 184 -4591 432 -4589
rect 184 -4625 286 -4591
rect 320 -4625 432 -4591
rect 184 -4627 432 -4625
rect 184 -4661 190 -4627
rect 224 -4661 392 -4627
rect 426 -4661 432 -4627
rect 184 -4663 432 -4661
rect 184 -4697 286 -4663
rect 320 -4697 432 -4663
rect 184 -4699 432 -4697
rect 184 -4733 190 -4699
rect 224 -4733 392 -4699
rect 426 -4733 432 -4699
rect 184 -4735 432 -4733
rect 184 -4769 286 -4735
rect 320 -4769 432 -4735
rect 184 -4771 432 -4769
rect 184 -4805 190 -4771
rect 224 -4805 392 -4771
rect 426 -4805 432 -4771
rect 184 -4807 432 -4805
rect 184 -4841 286 -4807
rect 320 -4841 432 -4807
rect 184 -4843 432 -4841
rect 184 -4877 190 -4843
rect 224 -4877 392 -4843
rect 426 -4877 432 -4843
rect 184 -4879 432 -4877
rect 184 -4913 286 -4879
rect 320 -4913 432 -4879
rect 184 -4915 432 -4913
rect 184 -4949 190 -4915
rect 224 -4949 392 -4915
rect 426 -4949 432 -4915
rect 184 -4951 432 -4949
rect 184 -4985 286 -4951
rect 320 -4985 432 -4951
rect 184 -4987 432 -4985
rect -432 -5023 -184 -5021
tri -800 -5057 -787 -5044 sw
tri -445 -5057 -432 -5044 se
rect -432 -5057 -330 -5023
rect -296 -5057 -184 -5023
rect 184 -5021 190 -4987
rect 224 -5021 392 -4987
rect 426 -5021 432 -4987
tri 522 5000 542 5020 se
rect 542 5000 690 5020
tri 690 5000 710 5020 sw
rect 522 4985 710 5000
rect 522 -4985 563 4985
rect 669 -4985 710 4985
rect 522 -5000 710 -4985
tri 522 -5020 542 -5000 ne
rect 542 -5020 690 -5000
tri 690 -5020 710 -5000 nw
rect 800 4987 806 5021
rect 840 4987 1008 5021
rect 1042 4987 1048 5021
rect 1416 5023 1494 5057
rect 1528 5023 1540 5057
rect 1416 5021 1540 5023
rect 800 4985 1048 4987
rect 800 4951 902 4985
rect 936 4951 1048 4985
rect 800 4949 1048 4951
rect 800 4915 806 4949
rect 840 4915 1008 4949
rect 1042 4915 1048 4949
rect 800 4913 1048 4915
rect 800 4879 902 4913
rect 936 4879 1048 4913
rect 800 4877 1048 4879
rect 800 4843 806 4877
rect 840 4843 1008 4877
rect 1042 4843 1048 4877
rect 800 4841 1048 4843
rect 800 4807 902 4841
rect 936 4807 1048 4841
rect 800 4805 1048 4807
rect 800 4771 806 4805
rect 840 4771 1008 4805
rect 1042 4771 1048 4805
rect 800 4769 1048 4771
rect 800 4735 902 4769
rect 936 4735 1048 4769
rect 800 4733 1048 4735
rect 800 4699 806 4733
rect 840 4699 1008 4733
rect 1042 4699 1048 4733
rect 800 4697 1048 4699
rect 800 4663 902 4697
rect 936 4663 1048 4697
rect 800 4661 1048 4663
rect 800 4627 806 4661
rect 840 4627 1008 4661
rect 1042 4627 1048 4661
rect 800 4625 1048 4627
rect 800 4591 902 4625
rect 936 4591 1048 4625
rect 800 4589 1048 4591
rect 800 4555 806 4589
rect 840 4555 1008 4589
rect 1042 4555 1048 4589
rect 800 4553 1048 4555
rect 800 4519 902 4553
rect 936 4519 1048 4553
rect 800 4517 1048 4519
rect 800 4483 806 4517
rect 840 4483 1008 4517
rect 1042 4483 1048 4517
rect 800 4481 1048 4483
rect 800 4447 902 4481
rect 936 4447 1048 4481
rect 800 4445 1048 4447
rect 800 4411 806 4445
rect 840 4411 1008 4445
rect 1042 4411 1048 4445
rect 800 4409 1048 4411
rect 800 4375 902 4409
rect 936 4375 1048 4409
rect 800 4373 1048 4375
rect 800 4339 806 4373
rect 840 4339 1008 4373
rect 1042 4339 1048 4373
rect 800 4337 1048 4339
rect 800 4303 902 4337
rect 936 4303 1048 4337
rect 800 4301 1048 4303
rect 800 4267 806 4301
rect 840 4267 1008 4301
rect 1042 4267 1048 4301
rect 800 4265 1048 4267
rect 800 4231 902 4265
rect 936 4231 1048 4265
rect 800 4229 1048 4231
rect 800 4195 806 4229
rect 840 4195 1008 4229
rect 1042 4195 1048 4229
rect 800 4193 1048 4195
rect 800 4159 902 4193
rect 936 4159 1048 4193
rect 800 4157 1048 4159
rect 800 4123 806 4157
rect 840 4123 1008 4157
rect 1042 4123 1048 4157
rect 800 4121 1048 4123
rect 800 4087 902 4121
rect 936 4087 1048 4121
rect 800 4085 1048 4087
rect 800 4051 806 4085
rect 840 4051 1008 4085
rect 1042 4051 1048 4085
rect 800 4049 1048 4051
rect 800 4015 902 4049
rect 936 4015 1048 4049
rect 800 4013 1048 4015
rect 800 3979 806 4013
rect 840 3979 1008 4013
rect 1042 3979 1048 4013
rect 800 3977 1048 3979
rect 800 3943 902 3977
rect 936 3943 1048 3977
rect 800 3941 1048 3943
rect 800 3907 806 3941
rect 840 3907 1008 3941
rect 1042 3907 1048 3941
rect 800 3905 1048 3907
rect 800 3871 902 3905
rect 936 3871 1048 3905
rect 800 3869 1048 3871
rect 800 3835 806 3869
rect 840 3835 1008 3869
rect 1042 3835 1048 3869
rect 800 3833 1048 3835
rect 800 3799 902 3833
rect 936 3799 1048 3833
rect 800 3797 1048 3799
rect 800 3763 806 3797
rect 840 3763 1008 3797
rect 1042 3763 1048 3797
rect 800 3761 1048 3763
rect 800 3727 902 3761
rect 936 3727 1048 3761
rect 800 3725 1048 3727
rect 800 3691 806 3725
rect 840 3691 1008 3725
rect 1042 3691 1048 3725
rect 800 3689 1048 3691
rect 800 3655 902 3689
rect 936 3655 1048 3689
rect 800 3653 1048 3655
rect 800 3619 806 3653
rect 840 3619 1008 3653
rect 1042 3619 1048 3653
rect 800 3617 1048 3619
rect 800 3583 902 3617
rect 936 3583 1048 3617
rect 800 3581 1048 3583
rect 800 3547 806 3581
rect 840 3547 1008 3581
rect 1042 3547 1048 3581
rect 800 3545 1048 3547
rect 800 3511 902 3545
rect 936 3511 1048 3545
rect 800 3509 1048 3511
rect 800 3475 806 3509
rect 840 3475 1008 3509
rect 1042 3475 1048 3509
rect 800 3473 1048 3475
rect 800 3439 902 3473
rect 936 3439 1048 3473
rect 800 3437 1048 3439
rect 800 3403 806 3437
rect 840 3403 1008 3437
rect 1042 3403 1048 3437
rect 800 3401 1048 3403
rect 800 3367 902 3401
rect 936 3367 1048 3401
rect 800 3365 1048 3367
rect 800 3331 806 3365
rect 840 3331 1008 3365
rect 1042 3331 1048 3365
rect 800 3329 1048 3331
rect 800 3295 902 3329
rect 936 3295 1048 3329
rect 800 3293 1048 3295
rect 800 3259 806 3293
rect 840 3259 1008 3293
rect 1042 3259 1048 3293
rect 800 3257 1048 3259
rect 800 3223 902 3257
rect 936 3223 1048 3257
rect 800 3221 1048 3223
rect 800 3187 806 3221
rect 840 3187 1008 3221
rect 1042 3187 1048 3221
rect 800 3185 1048 3187
rect 800 3151 902 3185
rect 936 3151 1048 3185
rect 800 3149 1048 3151
rect 800 3115 806 3149
rect 840 3115 1008 3149
rect 1042 3115 1048 3149
rect 800 3113 1048 3115
rect 800 3079 902 3113
rect 936 3079 1048 3113
rect 800 3077 1048 3079
rect 800 3043 806 3077
rect 840 3043 1008 3077
rect 1042 3043 1048 3077
rect 800 3041 1048 3043
rect 800 3007 902 3041
rect 936 3007 1048 3041
rect 800 3005 1048 3007
rect 800 2971 806 3005
rect 840 2971 1008 3005
rect 1042 2971 1048 3005
rect 800 2969 1048 2971
rect 800 2935 902 2969
rect 936 2935 1048 2969
rect 800 2933 1048 2935
rect 800 2899 806 2933
rect 840 2899 1008 2933
rect 1042 2899 1048 2933
rect 800 2897 1048 2899
rect 800 2863 902 2897
rect 936 2863 1048 2897
rect 800 2861 1048 2863
rect 800 2827 806 2861
rect 840 2827 1008 2861
rect 1042 2827 1048 2861
rect 800 2825 1048 2827
rect 800 2791 902 2825
rect 936 2791 1048 2825
rect 800 2789 1048 2791
rect 800 2755 806 2789
rect 840 2755 1008 2789
rect 1042 2755 1048 2789
rect 800 2753 1048 2755
rect 800 2719 902 2753
rect 936 2719 1048 2753
rect 800 2717 1048 2719
rect 800 2683 806 2717
rect 840 2683 1008 2717
rect 1042 2683 1048 2717
rect 800 2681 1048 2683
rect 800 2647 902 2681
rect 936 2647 1048 2681
rect 800 2645 1048 2647
rect 800 2611 806 2645
rect 840 2611 1008 2645
rect 1042 2611 1048 2645
rect 800 2609 1048 2611
rect 800 2575 902 2609
rect 936 2575 1048 2609
rect 800 2573 1048 2575
rect 800 2539 806 2573
rect 840 2539 1008 2573
rect 1042 2539 1048 2573
rect 800 2537 1048 2539
rect 800 2503 902 2537
rect 936 2503 1048 2537
rect 800 2501 1048 2503
rect 800 2467 806 2501
rect 840 2467 1008 2501
rect 1042 2467 1048 2501
rect 800 2465 1048 2467
rect 800 2431 902 2465
rect 936 2431 1048 2465
rect 800 2429 1048 2431
rect 800 2395 806 2429
rect 840 2395 1008 2429
rect 1042 2395 1048 2429
rect 800 2393 1048 2395
rect 800 2359 902 2393
rect 936 2359 1048 2393
rect 800 2357 1048 2359
rect 800 2323 806 2357
rect 840 2323 1008 2357
rect 1042 2323 1048 2357
rect 800 2321 1048 2323
rect 800 2287 902 2321
rect 936 2287 1048 2321
rect 800 2285 1048 2287
rect 800 2251 806 2285
rect 840 2251 1008 2285
rect 1042 2251 1048 2285
rect 800 2249 1048 2251
rect 800 2215 902 2249
rect 936 2215 1048 2249
rect 800 2213 1048 2215
rect 800 2179 806 2213
rect 840 2179 1008 2213
rect 1042 2179 1048 2213
rect 800 2177 1048 2179
rect 800 2143 902 2177
rect 936 2143 1048 2177
rect 800 2141 1048 2143
rect 800 2107 806 2141
rect 840 2107 1008 2141
rect 1042 2107 1048 2141
rect 800 2105 1048 2107
rect 800 2071 902 2105
rect 936 2071 1048 2105
rect 800 2069 1048 2071
rect 800 2035 806 2069
rect 840 2035 1008 2069
rect 1042 2035 1048 2069
rect 800 2033 1048 2035
rect 800 1999 902 2033
rect 936 1999 1048 2033
rect 800 1997 1048 1999
rect 800 1963 806 1997
rect 840 1963 1008 1997
rect 1042 1963 1048 1997
rect 800 1961 1048 1963
rect 800 1927 902 1961
rect 936 1927 1048 1961
rect 800 1925 1048 1927
rect 800 1891 806 1925
rect 840 1891 1008 1925
rect 1042 1891 1048 1925
rect 800 1889 1048 1891
rect 800 1855 902 1889
rect 936 1855 1048 1889
rect 800 1853 1048 1855
rect 800 1819 806 1853
rect 840 1819 1008 1853
rect 1042 1819 1048 1853
rect 800 1817 1048 1819
rect 800 1783 902 1817
rect 936 1783 1048 1817
rect 800 1781 1048 1783
rect 800 1747 806 1781
rect 840 1747 1008 1781
rect 1042 1747 1048 1781
rect 800 1745 1048 1747
rect 800 1711 902 1745
rect 936 1711 1048 1745
rect 800 1709 1048 1711
rect 800 1675 806 1709
rect 840 1675 1008 1709
rect 1042 1675 1048 1709
rect 800 1673 1048 1675
rect 800 1639 902 1673
rect 936 1639 1048 1673
rect 800 1637 1048 1639
rect 800 1603 806 1637
rect 840 1603 1008 1637
rect 1042 1603 1048 1637
rect 800 1601 1048 1603
rect 800 1567 902 1601
rect 936 1567 1048 1601
rect 800 1565 1048 1567
rect 800 1531 806 1565
rect 840 1531 1008 1565
rect 1042 1531 1048 1565
rect 800 1529 1048 1531
rect 800 1495 902 1529
rect 936 1495 1048 1529
rect 800 1493 1048 1495
rect 800 1459 806 1493
rect 840 1459 1008 1493
rect 1042 1459 1048 1493
rect 800 1457 1048 1459
rect 800 1423 902 1457
rect 936 1423 1048 1457
rect 800 1421 1048 1423
rect 800 1387 806 1421
rect 840 1387 1008 1421
rect 1042 1387 1048 1421
rect 800 1385 1048 1387
rect 800 1351 902 1385
rect 936 1351 1048 1385
rect 800 1349 1048 1351
rect 800 1315 806 1349
rect 840 1315 1008 1349
rect 1042 1315 1048 1349
rect 800 1313 1048 1315
rect 800 1279 902 1313
rect 936 1279 1048 1313
rect 800 1277 1048 1279
rect 800 1243 806 1277
rect 840 1243 1008 1277
rect 1042 1243 1048 1277
rect 800 1241 1048 1243
rect 800 1207 902 1241
rect 936 1207 1048 1241
rect 800 1205 1048 1207
rect 800 1171 806 1205
rect 840 1171 1008 1205
rect 1042 1171 1048 1205
rect 800 1169 1048 1171
rect 800 1135 902 1169
rect 936 1135 1048 1169
rect 800 1133 1048 1135
rect 800 1099 806 1133
rect 840 1099 1008 1133
rect 1042 1099 1048 1133
rect 800 1097 1048 1099
rect 800 1063 902 1097
rect 936 1063 1048 1097
rect 800 1061 1048 1063
rect 800 1027 806 1061
rect 840 1027 1008 1061
rect 1042 1027 1048 1061
rect 800 1025 1048 1027
rect 800 991 902 1025
rect 936 991 1048 1025
rect 800 989 1048 991
rect 800 955 806 989
rect 840 955 1008 989
rect 1042 955 1048 989
rect 800 953 1048 955
rect 800 919 902 953
rect 936 919 1048 953
rect 800 917 1048 919
rect 800 883 806 917
rect 840 883 1008 917
rect 1042 883 1048 917
rect 800 881 1048 883
rect 800 847 902 881
rect 936 847 1048 881
rect 800 845 1048 847
rect 800 811 806 845
rect 840 811 1008 845
rect 1042 811 1048 845
rect 800 809 1048 811
rect 800 775 902 809
rect 936 775 1048 809
rect 800 773 1048 775
rect 800 739 806 773
rect 840 739 1008 773
rect 1042 739 1048 773
rect 800 737 1048 739
rect 800 703 902 737
rect 936 703 1048 737
rect 800 701 1048 703
rect 800 667 806 701
rect 840 667 1008 701
rect 1042 667 1048 701
rect 800 665 1048 667
rect 800 631 902 665
rect 936 631 1048 665
rect 800 629 1048 631
rect 800 595 806 629
rect 840 595 1008 629
rect 1042 595 1048 629
rect 800 593 1048 595
rect 800 559 902 593
rect 936 559 1048 593
rect 800 557 1048 559
rect 800 523 806 557
rect 840 523 1008 557
rect 1042 523 1048 557
rect 800 521 1048 523
rect 800 487 902 521
rect 936 487 1048 521
rect 800 485 1048 487
rect 800 451 806 485
rect 840 451 1008 485
rect 1042 451 1048 485
rect 800 449 1048 451
rect 800 415 902 449
rect 936 415 1048 449
rect 800 413 1048 415
rect 800 379 806 413
rect 840 379 1008 413
rect 1042 379 1048 413
rect 800 377 1048 379
rect 800 343 902 377
rect 936 343 1048 377
rect 800 341 1048 343
rect 800 307 806 341
rect 840 307 1008 341
rect 1042 307 1048 341
rect 800 305 1048 307
rect 800 271 902 305
rect 936 271 1048 305
rect 800 269 1048 271
rect 800 235 806 269
rect 840 235 1008 269
rect 1042 235 1048 269
rect 800 233 1048 235
rect 800 199 902 233
rect 936 199 1048 233
rect 800 197 1048 199
rect 800 163 806 197
rect 840 163 1008 197
rect 1042 163 1048 197
rect 800 161 1048 163
rect 800 127 902 161
rect 936 127 1048 161
rect 800 125 1048 127
rect 800 91 806 125
rect 840 91 1008 125
rect 1042 91 1048 125
rect 800 89 1048 91
rect 800 55 902 89
rect 936 55 1048 89
rect 800 53 1048 55
rect 800 19 806 53
rect 840 19 1008 53
rect 1042 19 1048 53
rect 800 17 1048 19
rect 800 -17 902 17
rect 936 -17 1048 17
rect 800 -19 1048 -17
rect 800 -53 806 -19
rect 840 -53 1008 -19
rect 1042 -53 1048 -19
rect 800 -55 1048 -53
rect 800 -89 902 -55
rect 936 -89 1048 -55
rect 800 -91 1048 -89
rect 800 -125 806 -91
rect 840 -125 1008 -91
rect 1042 -125 1048 -91
rect 800 -127 1048 -125
rect 800 -161 902 -127
rect 936 -161 1048 -127
rect 800 -163 1048 -161
rect 800 -197 806 -163
rect 840 -197 1008 -163
rect 1042 -197 1048 -163
rect 800 -199 1048 -197
rect 800 -233 902 -199
rect 936 -233 1048 -199
rect 800 -235 1048 -233
rect 800 -269 806 -235
rect 840 -269 1008 -235
rect 1042 -269 1048 -235
rect 800 -271 1048 -269
rect 800 -305 902 -271
rect 936 -305 1048 -271
rect 800 -307 1048 -305
rect 800 -341 806 -307
rect 840 -341 1008 -307
rect 1042 -341 1048 -307
rect 800 -343 1048 -341
rect 800 -377 902 -343
rect 936 -377 1048 -343
rect 800 -379 1048 -377
rect 800 -413 806 -379
rect 840 -413 1008 -379
rect 1042 -413 1048 -379
rect 800 -415 1048 -413
rect 800 -449 902 -415
rect 936 -449 1048 -415
rect 800 -451 1048 -449
rect 800 -485 806 -451
rect 840 -485 1008 -451
rect 1042 -485 1048 -451
rect 800 -487 1048 -485
rect 800 -521 902 -487
rect 936 -521 1048 -487
rect 800 -523 1048 -521
rect 800 -557 806 -523
rect 840 -557 1008 -523
rect 1042 -557 1048 -523
rect 800 -559 1048 -557
rect 800 -593 902 -559
rect 936 -593 1048 -559
rect 800 -595 1048 -593
rect 800 -629 806 -595
rect 840 -629 1008 -595
rect 1042 -629 1048 -595
rect 800 -631 1048 -629
rect 800 -665 902 -631
rect 936 -665 1048 -631
rect 800 -667 1048 -665
rect 800 -701 806 -667
rect 840 -701 1008 -667
rect 1042 -701 1048 -667
rect 800 -703 1048 -701
rect 800 -737 902 -703
rect 936 -737 1048 -703
rect 800 -739 1048 -737
rect 800 -773 806 -739
rect 840 -773 1008 -739
rect 1042 -773 1048 -739
rect 800 -775 1048 -773
rect 800 -809 902 -775
rect 936 -809 1048 -775
rect 800 -811 1048 -809
rect 800 -845 806 -811
rect 840 -845 1008 -811
rect 1042 -845 1048 -811
rect 800 -847 1048 -845
rect 800 -881 902 -847
rect 936 -881 1048 -847
rect 800 -883 1048 -881
rect 800 -917 806 -883
rect 840 -917 1008 -883
rect 1042 -917 1048 -883
rect 800 -919 1048 -917
rect 800 -953 902 -919
rect 936 -953 1048 -919
rect 800 -955 1048 -953
rect 800 -989 806 -955
rect 840 -989 1008 -955
rect 1042 -989 1048 -955
rect 800 -991 1048 -989
rect 800 -1025 902 -991
rect 936 -1025 1048 -991
rect 800 -1027 1048 -1025
rect 800 -1061 806 -1027
rect 840 -1061 1008 -1027
rect 1042 -1061 1048 -1027
rect 800 -1063 1048 -1061
rect 800 -1097 902 -1063
rect 936 -1097 1048 -1063
rect 800 -1099 1048 -1097
rect 800 -1133 806 -1099
rect 840 -1133 1008 -1099
rect 1042 -1133 1048 -1099
rect 800 -1135 1048 -1133
rect 800 -1169 902 -1135
rect 936 -1169 1048 -1135
rect 800 -1171 1048 -1169
rect 800 -1205 806 -1171
rect 840 -1205 1008 -1171
rect 1042 -1205 1048 -1171
rect 800 -1207 1048 -1205
rect 800 -1241 902 -1207
rect 936 -1241 1048 -1207
rect 800 -1243 1048 -1241
rect 800 -1277 806 -1243
rect 840 -1277 1008 -1243
rect 1042 -1277 1048 -1243
rect 800 -1279 1048 -1277
rect 800 -1313 902 -1279
rect 936 -1313 1048 -1279
rect 800 -1315 1048 -1313
rect 800 -1349 806 -1315
rect 840 -1349 1008 -1315
rect 1042 -1349 1048 -1315
rect 800 -1351 1048 -1349
rect 800 -1385 902 -1351
rect 936 -1385 1048 -1351
rect 800 -1387 1048 -1385
rect 800 -1421 806 -1387
rect 840 -1421 1008 -1387
rect 1042 -1421 1048 -1387
rect 800 -1423 1048 -1421
rect 800 -1457 902 -1423
rect 936 -1457 1048 -1423
rect 800 -1459 1048 -1457
rect 800 -1493 806 -1459
rect 840 -1493 1008 -1459
rect 1042 -1493 1048 -1459
rect 800 -1495 1048 -1493
rect 800 -1529 902 -1495
rect 936 -1529 1048 -1495
rect 800 -1531 1048 -1529
rect 800 -1565 806 -1531
rect 840 -1565 1008 -1531
rect 1042 -1565 1048 -1531
rect 800 -1567 1048 -1565
rect 800 -1601 902 -1567
rect 936 -1601 1048 -1567
rect 800 -1603 1048 -1601
rect 800 -1637 806 -1603
rect 840 -1637 1008 -1603
rect 1042 -1637 1048 -1603
rect 800 -1639 1048 -1637
rect 800 -1673 902 -1639
rect 936 -1673 1048 -1639
rect 800 -1675 1048 -1673
rect 800 -1709 806 -1675
rect 840 -1709 1008 -1675
rect 1042 -1709 1048 -1675
rect 800 -1711 1048 -1709
rect 800 -1745 902 -1711
rect 936 -1745 1048 -1711
rect 800 -1747 1048 -1745
rect 800 -1781 806 -1747
rect 840 -1781 1008 -1747
rect 1042 -1781 1048 -1747
rect 800 -1783 1048 -1781
rect 800 -1817 902 -1783
rect 936 -1817 1048 -1783
rect 800 -1819 1048 -1817
rect 800 -1853 806 -1819
rect 840 -1853 1008 -1819
rect 1042 -1853 1048 -1819
rect 800 -1855 1048 -1853
rect 800 -1889 902 -1855
rect 936 -1889 1048 -1855
rect 800 -1891 1048 -1889
rect 800 -1925 806 -1891
rect 840 -1925 1008 -1891
rect 1042 -1925 1048 -1891
rect 800 -1927 1048 -1925
rect 800 -1961 902 -1927
rect 936 -1961 1048 -1927
rect 800 -1963 1048 -1961
rect 800 -1997 806 -1963
rect 840 -1997 1008 -1963
rect 1042 -1997 1048 -1963
rect 800 -1999 1048 -1997
rect 800 -2033 902 -1999
rect 936 -2033 1048 -1999
rect 800 -2035 1048 -2033
rect 800 -2069 806 -2035
rect 840 -2069 1008 -2035
rect 1042 -2069 1048 -2035
rect 800 -2071 1048 -2069
rect 800 -2105 902 -2071
rect 936 -2105 1048 -2071
rect 800 -2107 1048 -2105
rect 800 -2141 806 -2107
rect 840 -2141 1008 -2107
rect 1042 -2141 1048 -2107
rect 800 -2143 1048 -2141
rect 800 -2177 902 -2143
rect 936 -2177 1048 -2143
rect 800 -2179 1048 -2177
rect 800 -2213 806 -2179
rect 840 -2213 1008 -2179
rect 1042 -2213 1048 -2179
rect 800 -2215 1048 -2213
rect 800 -2249 902 -2215
rect 936 -2249 1048 -2215
rect 800 -2251 1048 -2249
rect 800 -2285 806 -2251
rect 840 -2285 1008 -2251
rect 1042 -2285 1048 -2251
rect 800 -2287 1048 -2285
rect 800 -2321 902 -2287
rect 936 -2321 1048 -2287
rect 800 -2323 1048 -2321
rect 800 -2357 806 -2323
rect 840 -2357 1008 -2323
rect 1042 -2357 1048 -2323
rect 800 -2359 1048 -2357
rect 800 -2393 902 -2359
rect 936 -2393 1048 -2359
rect 800 -2395 1048 -2393
rect 800 -2429 806 -2395
rect 840 -2429 1008 -2395
rect 1042 -2429 1048 -2395
rect 800 -2431 1048 -2429
rect 800 -2465 902 -2431
rect 936 -2465 1048 -2431
rect 800 -2467 1048 -2465
rect 800 -2501 806 -2467
rect 840 -2501 1008 -2467
rect 1042 -2501 1048 -2467
rect 800 -2503 1048 -2501
rect 800 -2537 902 -2503
rect 936 -2537 1048 -2503
rect 800 -2539 1048 -2537
rect 800 -2573 806 -2539
rect 840 -2573 1008 -2539
rect 1042 -2573 1048 -2539
rect 800 -2575 1048 -2573
rect 800 -2609 902 -2575
rect 936 -2609 1048 -2575
rect 800 -2611 1048 -2609
rect 800 -2645 806 -2611
rect 840 -2645 1008 -2611
rect 1042 -2645 1048 -2611
rect 800 -2647 1048 -2645
rect 800 -2681 902 -2647
rect 936 -2681 1048 -2647
rect 800 -2683 1048 -2681
rect 800 -2717 806 -2683
rect 840 -2717 1008 -2683
rect 1042 -2717 1048 -2683
rect 800 -2719 1048 -2717
rect 800 -2753 902 -2719
rect 936 -2753 1048 -2719
rect 800 -2755 1048 -2753
rect 800 -2789 806 -2755
rect 840 -2789 1008 -2755
rect 1042 -2789 1048 -2755
rect 800 -2791 1048 -2789
rect 800 -2825 902 -2791
rect 936 -2825 1048 -2791
rect 800 -2827 1048 -2825
rect 800 -2861 806 -2827
rect 840 -2861 1008 -2827
rect 1042 -2861 1048 -2827
rect 800 -2863 1048 -2861
rect 800 -2897 902 -2863
rect 936 -2897 1048 -2863
rect 800 -2899 1048 -2897
rect 800 -2933 806 -2899
rect 840 -2933 1008 -2899
rect 1042 -2933 1048 -2899
rect 800 -2935 1048 -2933
rect 800 -2969 902 -2935
rect 936 -2969 1048 -2935
rect 800 -2971 1048 -2969
rect 800 -3005 806 -2971
rect 840 -3005 1008 -2971
rect 1042 -3005 1048 -2971
rect 800 -3007 1048 -3005
rect 800 -3041 902 -3007
rect 936 -3041 1048 -3007
rect 800 -3043 1048 -3041
rect 800 -3077 806 -3043
rect 840 -3077 1008 -3043
rect 1042 -3077 1048 -3043
rect 800 -3079 1048 -3077
rect 800 -3113 902 -3079
rect 936 -3113 1048 -3079
rect 800 -3115 1048 -3113
rect 800 -3149 806 -3115
rect 840 -3149 1008 -3115
rect 1042 -3149 1048 -3115
rect 800 -3151 1048 -3149
rect 800 -3185 902 -3151
rect 936 -3185 1048 -3151
rect 800 -3187 1048 -3185
rect 800 -3221 806 -3187
rect 840 -3221 1008 -3187
rect 1042 -3221 1048 -3187
rect 800 -3223 1048 -3221
rect 800 -3257 902 -3223
rect 936 -3257 1048 -3223
rect 800 -3259 1048 -3257
rect 800 -3293 806 -3259
rect 840 -3293 1008 -3259
rect 1042 -3293 1048 -3259
rect 800 -3295 1048 -3293
rect 800 -3329 902 -3295
rect 936 -3329 1048 -3295
rect 800 -3331 1048 -3329
rect 800 -3365 806 -3331
rect 840 -3365 1008 -3331
rect 1042 -3365 1048 -3331
rect 800 -3367 1048 -3365
rect 800 -3401 902 -3367
rect 936 -3401 1048 -3367
rect 800 -3403 1048 -3401
rect 800 -3437 806 -3403
rect 840 -3437 1008 -3403
rect 1042 -3437 1048 -3403
rect 800 -3439 1048 -3437
rect 800 -3473 902 -3439
rect 936 -3473 1048 -3439
rect 800 -3475 1048 -3473
rect 800 -3509 806 -3475
rect 840 -3509 1008 -3475
rect 1042 -3509 1048 -3475
rect 800 -3511 1048 -3509
rect 800 -3545 902 -3511
rect 936 -3545 1048 -3511
rect 800 -3547 1048 -3545
rect 800 -3581 806 -3547
rect 840 -3581 1008 -3547
rect 1042 -3581 1048 -3547
rect 800 -3583 1048 -3581
rect 800 -3617 902 -3583
rect 936 -3617 1048 -3583
rect 800 -3619 1048 -3617
rect 800 -3653 806 -3619
rect 840 -3653 1008 -3619
rect 1042 -3653 1048 -3619
rect 800 -3655 1048 -3653
rect 800 -3689 902 -3655
rect 936 -3689 1048 -3655
rect 800 -3691 1048 -3689
rect 800 -3725 806 -3691
rect 840 -3725 1008 -3691
rect 1042 -3725 1048 -3691
rect 800 -3727 1048 -3725
rect 800 -3761 902 -3727
rect 936 -3761 1048 -3727
rect 800 -3763 1048 -3761
rect 800 -3797 806 -3763
rect 840 -3797 1008 -3763
rect 1042 -3797 1048 -3763
rect 800 -3799 1048 -3797
rect 800 -3833 902 -3799
rect 936 -3833 1048 -3799
rect 800 -3835 1048 -3833
rect 800 -3869 806 -3835
rect 840 -3869 1008 -3835
rect 1042 -3869 1048 -3835
rect 800 -3871 1048 -3869
rect 800 -3905 902 -3871
rect 936 -3905 1048 -3871
rect 800 -3907 1048 -3905
rect 800 -3941 806 -3907
rect 840 -3941 1008 -3907
rect 1042 -3941 1048 -3907
rect 800 -3943 1048 -3941
rect 800 -3977 902 -3943
rect 936 -3977 1048 -3943
rect 800 -3979 1048 -3977
rect 800 -4013 806 -3979
rect 840 -4013 1008 -3979
rect 1042 -4013 1048 -3979
rect 800 -4015 1048 -4013
rect 800 -4049 902 -4015
rect 936 -4049 1048 -4015
rect 800 -4051 1048 -4049
rect 800 -4085 806 -4051
rect 840 -4085 1008 -4051
rect 1042 -4085 1048 -4051
rect 800 -4087 1048 -4085
rect 800 -4121 902 -4087
rect 936 -4121 1048 -4087
rect 800 -4123 1048 -4121
rect 800 -4157 806 -4123
rect 840 -4157 1008 -4123
rect 1042 -4157 1048 -4123
rect 800 -4159 1048 -4157
rect 800 -4193 902 -4159
rect 936 -4193 1048 -4159
rect 800 -4195 1048 -4193
rect 800 -4229 806 -4195
rect 840 -4229 1008 -4195
rect 1042 -4229 1048 -4195
rect 800 -4231 1048 -4229
rect 800 -4265 902 -4231
rect 936 -4265 1048 -4231
rect 800 -4267 1048 -4265
rect 800 -4301 806 -4267
rect 840 -4301 1008 -4267
rect 1042 -4301 1048 -4267
rect 800 -4303 1048 -4301
rect 800 -4337 902 -4303
rect 936 -4337 1048 -4303
rect 800 -4339 1048 -4337
rect 800 -4373 806 -4339
rect 840 -4373 1008 -4339
rect 1042 -4373 1048 -4339
rect 800 -4375 1048 -4373
rect 800 -4409 902 -4375
rect 936 -4409 1048 -4375
rect 800 -4411 1048 -4409
rect 800 -4445 806 -4411
rect 840 -4445 1008 -4411
rect 1042 -4445 1048 -4411
rect 800 -4447 1048 -4445
rect 800 -4481 902 -4447
rect 936 -4481 1048 -4447
rect 800 -4483 1048 -4481
rect 800 -4517 806 -4483
rect 840 -4517 1008 -4483
rect 1042 -4517 1048 -4483
rect 800 -4519 1048 -4517
rect 800 -4553 902 -4519
rect 936 -4553 1048 -4519
rect 800 -4555 1048 -4553
rect 800 -4589 806 -4555
rect 840 -4589 1008 -4555
rect 1042 -4589 1048 -4555
rect 800 -4591 1048 -4589
rect 800 -4625 902 -4591
rect 936 -4625 1048 -4591
rect 800 -4627 1048 -4625
rect 800 -4661 806 -4627
rect 840 -4661 1008 -4627
rect 1042 -4661 1048 -4627
rect 800 -4663 1048 -4661
rect 800 -4697 902 -4663
rect 936 -4697 1048 -4663
rect 800 -4699 1048 -4697
rect 800 -4733 806 -4699
rect 840 -4733 1008 -4699
rect 1042 -4733 1048 -4699
rect 800 -4735 1048 -4733
rect 800 -4769 902 -4735
rect 936 -4769 1048 -4735
rect 800 -4771 1048 -4769
rect 800 -4805 806 -4771
rect 840 -4805 1008 -4771
rect 1042 -4805 1048 -4771
rect 800 -4807 1048 -4805
rect 800 -4841 902 -4807
rect 936 -4841 1048 -4807
rect 800 -4843 1048 -4841
rect 800 -4877 806 -4843
rect 840 -4877 1008 -4843
rect 1042 -4877 1048 -4843
rect 800 -4879 1048 -4877
rect 800 -4913 902 -4879
rect 936 -4913 1048 -4879
rect 800 -4915 1048 -4913
rect 800 -4949 806 -4915
rect 840 -4949 1008 -4915
rect 1042 -4949 1048 -4915
rect 800 -4951 1048 -4949
rect 800 -4985 902 -4951
rect 936 -4985 1048 -4951
rect 800 -4987 1048 -4985
rect 184 -5023 432 -5021
tri -184 -5057 -171 -5044 sw
tri 171 -5057 184 -5044 se
rect 184 -5057 286 -5023
rect 320 -5057 432 -5023
rect 800 -5021 806 -4987
rect 840 -5021 1008 -4987
rect 1042 -5021 1048 -4987
tri 1138 5000 1158 5020 se
rect 1158 5000 1306 5020
tri 1306 5000 1326 5020 sw
rect 1138 4985 1326 5000
rect 1138 -4985 1179 4985
rect 1285 -4985 1326 4985
rect 1138 -5000 1326 -4985
tri 1138 -5020 1158 -5000 ne
rect 1158 -5020 1306 -5000
tri 1306 -5020 1326 -5000 nw
rect 800 -5023 1048 -5021
tri 432 -5057 445 -5044 sw
tri 787 -5057 800 -5044 se
rect 800 -5057 902 -5023
rect 936 -5057 1048 -5023
rect 1416 -5021 1422 5021
rect 1528 -5021 1540 5021
rect 1416 -5023 1540 -5021
tri 1048 -5057 1061 -5044 sw
tri 1403 -5057 1416 -5044 se
rect 1416 -5057 1494 -5023
rect 1528 -5057 1540 -5023
rect -1540 -5062 -1403 -5057
tri -1403 -5062 -1398 -5057 sw
tri -1066 -5062 -1061 -5057 se
rect -1061 -5062 -787 -5057
tri -787 -5062 -782 -5057 sw
tri -450 -5062 -445 -5057 se
rect -445 -5062 -171 -5057
tri -171 -5062 -166 -5057 sw
tri 166 -5062 171 -5057 se
rect 171 -5062 445 -5057
tri 445 -5062 450 -5057 sw
tri 782 -5062 787 -5057 se
rect 787 -5062 1061 -5057
tri 1061 -5062 1066 -5057 sw
tri 1398 -5062 1403 -5057 se
rect 1403 -5062 1540 -5057
rect -1540 -5084 -1398 -5062
tri -1398 -5084 -1376 -5062 sw
tri -1088 -5084 -1066 -5062 se
rect -1066 -5084 -782 -5062
tri -782 -5084 -760 -5062 sw
tri -472 -5084 -450 -5062 se
rect -450 -5084 -166 -5062
tri -166 -5084 -144 -5062 sw
tri 144 -5084 166 -5062 se
rect 166 -5084 450 -5062
tri 450 -5084 472 -5062 sw
tri 760 -5084 782 -5062 se
rect 782 -5084 1066 -5062
tri 1066 -5084 1088 -5062 sw
tri 1376 -5084 1398 -5062 se
rect 1398 -5084 1540 -5062
rect -1540 -5090 1540 -5084
rect -1540 -5124 -1357 -5090
rect -1323 -5124 -1285 -5090
rect -1251 -5124 -1213 -5090
rect -1179 -5124 -1141 -5090
rect -1107 -5124 -741 -5090
rect -707 -5124 -669 -5090
rect -635 -5124 -597 -5090
rect -563 -5124 -525 -5090
rect -491 -5124 -125 -5090
rect -91 -5124 -53 -5090
rect -19 -5124 19 -5090
rect 53 -5124 91 -5090
rect 125 -5124 491 -5090
rect 525 -5124 563 -5090
rect 597 -5124 635 -5090
rect 669 -5124 707 -5090
rect 741 -5124 1107 -5090
rect 1141 -5124 1179 -5090
rect 1213 -5124 1251 -5090
rect 1285 -5124 1323 -5090
rect 1357 -5124 1540 -5090
rect -1540 -5188 1540 -5124
<< properties >>
string FIXED_BBOX 1024 -5106 1438 5106
string GDS_END 1270914
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 731550
<< end >>
