// input external delay: 4 ns
// in delay: 0.011365 ns
// input delay: 0.010861 ns
// output delay: 0.175128 ns
// out delay: 0.000627 ns
// total extra delay: 4.197981 ns
// critical path time: 20.308298 ns
// total inverter delay needed: 20.308298 - 4.197981 = 16.110317 ns
// average one inverter delay: 0.03012 ns
// inverters needed: 532

module inverter(input wire a, output wire y);
    not (y, a);
endmodule

module issue_replica(input wire in, output wire out);
	wire [530:0] interconnections; // Wires to connect inverters

	// Instantiate 532 inverters and chain them
	inverter inv0(in, interconnections[0]);
	inverter inv1(interconnections[0], interconnections[1]);
	inverter inv2(interconnections[1], interconnections[2]);
	inverter inv3(interconnections[2], interconnections[3]);
	inverter inv4(interconnections[3], interconnections[4]);
	inverter inv5(interconnections[4], interconnections[5]);
	inverter inv6(interconnections[5], interconnections[6]);
	inverter inv7(interconnections[6], interconnections[7]);
	inverter inv8(interconnections[7], interconnections[8]);
	inverter inv9(interconnections[8], interconnections[9]);
	inverter inv10(interconnections[9], interconnections[10]);
	inverter inv11(interconnections[10], interconnections[11]);
	inverter inv12(interconnections[11], interconnections[12]);
	inverter inv13(interconnections[12], interconnections[13]);
	inverter inv14(interconnections[13], interconnections[14]);
	inverter inv15(interconnections[14], interconnections[15]);
	inverter inv16(interconnections[15], interconnections[16]);
	inverter inv17(interconnections[16], interconnections[17]);
	inverter inv18(interconnections[17], interconnections[18]);
	inverter inv19(interconnections[18], interconnections[19]);
	inverter inv20(interconnections[19], interconnections[20]);
	inverter inv21(interconnections[20], interconnections[21]);
	inverter inv22(interconnections[21], interconnections[22]);
	inverter inv23(interconnections[22], interconnections[23]);
	inverter inv24(interconnections[23], interconnections[24]);
	inverter inv25(interconnections[24], interconnections[25]);
	inverter inv26(interconnections[25], interconnections[26]);
	inverter inv27(interconnections[26], interconnections[27]);
	inverter inv28(interconnections[27], interconnections[28]);
	inverter inv29(interconnections[28], interconnections[29]);
	inverter inv30(interconnections[29], interconnections[30]);
	inverter inv31(interconnections[30], interconnections[31]);
	inverter inv32(interconnections[31], interconnections[32]);
	inverter inv33(interconnections[32], interconnections[33]);
	inverter inv34(interconnections[33], interconnections[34]);
	inverter inv35(interconnections[34], interconnections[35]);
	inverter inv36(interconnections[35], interconnections[36]);
	inverter inv37(interconnections[36], interconnections[37]);
	inverter inv38(interconnections[37], interconnections[38]);
	inverter inv39(interconnections[38], interconnections[39]);
	inverter inv40(interconnections[39], interconnections[40]);
	inverter inv41(interconnections[40], interconnections[41]);
	inverter inv42(interconnections[41], interconnections[42]);
	inverter inv43(interconnections[42], interconnections[43]);
	inverter inv44(interconnections[43], interconnections[44]);
	inverter inv45(interconnections[44], interconnections[45]);
	inverter inv46(interconnections[45], interconnections[46]);
	inverter inv47(interconnections[46], interconnections[47]);
	inverter inv48(interconnections[47], interconnections[48]);
	inverter inv49(interconnections[48], interconnections[49]);
	inverter inv50(interconnections[49], interconnections[50]);
	inverter inv51(interconnections[50], interconnections[51]);
	inverter inv52(interconnections[51], interconnections[52]);
	inverter inv53(interconnections[52], interconnections[53]);
	inverter inv54(interconnections[53], interconnections[54]);
	inverter inv55(interconnections[54], interconnections[55]);
	inverter inv56(interconnections[55], interconnections[56]);
	inverter inv57(interconnections[56], interconnections[57]);
	inverter inv58(interconnections[57], interconnections[58]);
	inverter inv59(interconnections[58], interconnections[59]);
	inverter inv60(interconnections[59], interconnections[60]);
	inverter inv61(interconnections[60], interconnections[61]);
	inverter inv62(interconnections[61], interconnections[62]);
	inverter inv63(interconnections[62], interconnections[63]);
	inverter inv64(interconnections[63], interconnections[64]);
	inverter inv65(interconnections[64], interconnections[65]);
	inverter inv66(interconnections[65], interconnections[66]);
	inverter inv67(interconnections[66], interconnections[67]);
	inverter inv68(interconnections[67], interconnections[68]);
	inverter inv69(interconnections[68], interconnections[69]);
	inverter inv70(interconnections[69], interconnections[70]);
	inverter inv71(interconnections[70], interconnections[71]);
	inverter inv72(interconnections[71], interconnections[72]);
	inverter inv73(interconnections[72], interconnections[73]);
	inverter inv74(interconnections[73], interconnections[74]);
	inverter inv75(interconnections[74], interconnections[75]);
	inverter inv76(interconnections[75], interconnections[76]);
	inverter inv77(interconnections[76], interconnections[77]);
	inverter inv78(interconnections[77], interconnections[78]);
	inverter inv79(interconnections[78], interconnections[79]);
	inverter inv80(interconnections[79], interconnections[80]);
	inverter inv81(interconnections[80], interconnections[81]);
	inverter inv82(interconnections[81], interconnections[82]);
	inverter inv83(interconnections[82], interconnections[83]);
	inverter inv84(interconnections[83], interconnections[84]);
	inverter inv85(interconnections[84], interconnections[85]);
	inverter inv86(interconnections[85], interconnections[86]);
	inverter inv87(interconnections[86], interconnections[87]);
	inverter inv88(interconnections[87], interconnections[88]);
	inverter inv89(interconnections[88], interconnections[89]);
	inverter inv90(interconnections[89], interconnections[90]);
	inverter inv91(interconnections[90], interconnections[91]);
	inverter inv92(interconnections[91], interconnections[92]);
	inverter inv93(interconnections[92], interconnections[93]);
	inverter inv94(interconnections[93], interconnections[94]);
	inverter inv95(interconnections[94], interconnections[95]);
	inverter inv96(interconnections[95], interconnections[96]);
	inverter inv97(interconnections[96], interconnections[97]);
	inverter inv98(interconnections[97], interconnections[98]);
	inverter inv99(interconnections[98], interconnections[99]);
	inverter inv100(interconnections[99], interconnections[100]);
	inverter inv101(interconnections[100], interconnections[101]);
	inverter inv102(interconnections[101], interconnections[102]);
	inverter inv103(interconnections[102], interconnections[103]);
	inverter inv104(interconnections[103], interconnections[104]);
	inverter inv105(interconnections[104], interconnections[105]);
	inverter inv106(interconnections[105], interconnections[106]);
	inverter inv107(interconnections[106], interconnections[107]);
	inverter inv108(interconnections[107], interconnections[108]);
	inverter inv109(interconnections[108], interconnections[109]);
	inverter inv110(interconnections[109], interconnections[110]);
	inverter inv111(interconnections[110], interconnections[111]);
	inverter inv112(interconnections[111], interconnections[112]);
	inverter inv113(interconnections[112], interconnections[113]);
	inverter inv114(interconnections[113], interconnections[114]);
	inverter inv115(interconnections[114], interconnections[115]);
	inverter inv116(interconnections[115], interconnections[116]);
	inverter inv117(interconnections[116], interconnections[117]);
	inverter inv118(interconnections[117], interconnections[118]);
	inverter inv119(interconnections[118], interconnections[119]);
	inverter inv120(interconnections[119], interconnections[120]);
	inverter inv121(interconnections[120], interconnections[121]);
	inverter inv122(interconnections[121], interconnections[122]);
	inverter inv123(interconnections[122], interconnections[123]);
	inverter inv124(interconnections[123], interconnections[124]);
	inverter inv125(interconnections[124], interconnections[125]);
	inverter inv126(interconnections[125], interconnections[126]);
	inverter inv127(interconnections[126], interconnections[127]);
	inverter inv128(interconnections[127], interconnections[128]);
	inverter inv129(interconnections[128], interconnections[129]);
	inverter inv130(interconnections[129], interconnections[130]);
    inverter inv131(interconnections[130], interconnections[131]);
	inverter inv132(interconnections[131], interconnections[132]);
	inverter inv133(interconnections[132], interconnections[133]);
	inverter inv134(interconnections[133], interconnections[134]);
	inverter inv135(interconnections[134], interconnections[135]);
	inverter inv136(interconnections[135], interconnections[136]);
	inverter inv137(interconnections[136], interconnections[137]);
	inverter inv138(interconnections[137], interconnections[138]);
	inverter inv139(interconnections[138], interconnections[139]);
	inverter inv140(interconnections[139], interconnections[140]);
    inverter inv141(interconnections[140], interconnections[141]);
	inverter inv142(interconnections[141], interconnections[142]);
	inverter inv143(interconnections[142], interconnections[143]);
	inverter inv144(interconnections[143], interconnections[144]);
	inverter inv145(interconnections[144], interconnections[145]);
	inverter inv146(interconnections[145], interconnections[146]);
	inverter inv147(interconnections[146], interconnections[147]);
	inverter inv148(interconnections[147], interconnections[148]);
	inverter inv149(interconnections[148], interconnections[149]);
	inverter inv150(interconnections[149], interconnections[150]);
    inverter inv151(interconnections[150], interconnections[151]);
	inverter inv152(interconnections[151], interconnections[152]);
	inverter inv153(interconnections[152], interconnections[153]);
	inverter inv154(interconnections[153], interconnections[154]);
	inverter inv155(interconnections[154], interconnections[155]);
	inverter inv156(interconnections[155], interconnections[156]);
	inverter inv157(interconnections[156], interconnections[157]);
	inverter inv158(interconnections[157], interconnections[158]);
	inverter inv159(interconnections[158], interconnections[159]);
	inverter inv160(interconnections[159], interconnections[160]);
    inverter inv161(interconnections[160], interconnections[161]);
	inverter inv162(interconnections[161], interconnections[162]);
	inverter inv163(interconnections[162], interconnections[163]);
	inverter inv164(interconnections[163], interconnections[164]);
	inverter inv165(interconnections[164], interconnections[165]);
	inverter inv166(interconnections[165], interconnections[166]);
	inverter inv167(interconnections[166], interconnections[167]);
	inverter inv168(interconnections[167], interconnections[168]);
	inverter inv169(interconnections[168], interconnections[169]);
	inverter inv170(interconnections[169], interconnections[170]);
	inverter inv171(interconnections[170], interconnections[171]);
	inverter inv172(interconnections[171], interconnections[172]);
	inverter inv173(interconnections[172], interconnections[173]);
	inverter inv174(interconnections[173], interconnections[174]);
	inverter inv175(interconnections[174], interconnections[175]);
	inverter inv176(interconnections[175], interconnections[176]);
	inverter inv177(interconnections[176], interconnections[177]);
	inverter inv178(interconnections[177], interconnections[178]);
	inverter inv179(interconnections[178], interconnections[179]);
	inverter inv180(interconnections[179], interconnections[180]);
	inverter inv181(interconnections[180], interconnections[181]);
	inverter inv182(interconnections[181], interconnections[182]);
	inverter inv183(interconnections[182], interconnections[183]);
	inverter inv184(interconnections[183], interconnections[184]);
	inverter inv185(interconnections[184], interconnections[185]);
	inverter inv186(interconnections[185], interconnections[186]);
	inverter inv187(interconnections[186], interconnections[187]);
	inverter inv188(interconnections[187], interconnections[188]);
	inverter inv189(interconnections[188], interconnections[189]);
	inverter inv190(interconnections[189], interconnections[190]);
	inverter inv191(interconnections[190], interconnections[191]);
	inverter inv192(interconnections[191], interconnections[192]);
	inverter inv193(interconnections[192], interconnections[193]);
	inverter inv194(interconnections[193], interconnections[194]);
	inverter inv195(interconnections[194], interconnections[195]);
	inverter inv196(interconnections[195], interconnections[196]);
	inverter inv197(interconnections[196], interconnections[197]);
	inverter inv198(interconnections[197], interconnections[198]);
	inverter inv199(interconnections[198], interconnections[199]);
	inverter inv200(interconnections[199], interconnections[200]);
	inverter inv201(interconnections[200], interconnections[201]);
	inverter inv202(interconnections[201], interconnections[202]);
	inverter inv203(interconnections[202], interconnections[203]);
	inverter inv204(interconnections[203], interconnections[204]);
	inverter inv205(interconnections[204], interconnections[205]);
	inverter inv206(interconnections[205], interconnections[206]);
	inverter inv207(interconnections[206], interconnections[207]);
	inverter inv208(interconnections[207], interconnections[208]);
	inverter inv209(interconnections[208], interconnections[209]);
	inverter inv210(interconnections[209], interconnections[210]);
	inverter inv211(interconnections[210], interconnections[211]);
	inverter inv212(interconnections[211], interconnections[212]);
	inverter inv213(interconnections[212], interconnections[213]);
	inverter inv214(interconnections[213], interconnections[214]);
	inverter inv215(interconnections[214], interconnections[215]);
	inverter inv216(interconnections[215], interconnections[216]);
	inverter inv217(interconnections[216], interconnections[217]);
	inverter inv218(interconnections[217], interconnections[218]);
	inverter inv219(interconnections[218], interconnections[219]);
	inverter inv220(interconnections[219], interconnections[220]);
	inverter inv221(interconnections[220], interconnections[221]);
	inverter inv222(interconnections[221], interconnections[222]);
	inverter inv223(interconnections[222], interconnections[223]);
	inverter inv224(interconnections[223], interconnections[224]);
	inverter inv225(interconnections[224], interconnections[225]);
	inverter inv226(interconnections[225], interconnections[226]);
	inverter inv227(interconnections[226], interconnections[227]);
	inverter inv228(interconnections[227], interconnections[228]);
	inverter inv229(interconnections[228], interconnections[229]);
	inverter inv230(interconnections[229], interconnections[230]);
	inverter inv231(interconnections[230], interconnections[231]);
	inverter inv232(interconnections[231], interconnections[232]);
	inverter inv233(interconnections[232], interconnections[233]);
	inverter inv234(interconnections[233], interconnections[234]);
	inverter inv235(interconnections[234], interconnections[235]);
	inverter inv236(interconnections[235], interconnections[236]);
	inverter inv237(interconnections[236], interconnections[237]);
	inverter inv238(interconnections[237], interconnections[238]);
	inverter inv239(interconnections[238], interconnections[239]);
	inverter inv240(interconnections[239], interconnections[240]);
	inverter inv241(interconnections[240], interconnections[241]);
	inverter inv242(interconnections[241], interconnections[242]);
	inverter inv243(interconnections[242], interconnections[243]);
	inverter inv244(interconnections[243], interconnections[244]);
	inverter inv245(interconnections[244], interconnections[245]);
	inverter inv246(interconnections[245], interconnections[246]);
	inverter inv247(interconnections[246], interconnections[247]);
	inverter inv248(interconnections[247], interconnections[248]);
	inverter inv249(interconnections[248], interconnections[249]);
	inverter inv250(interconnections[249], interconnections[250]);
	inverter inv251(interconnections[250], interconnections[251]);
	inverter inv252(interconnections[251], interconnections[252]);
	inverter inv253(interconnections[252], interconnections[253]);
	inverter inv254(interconnections[253], interconnections[254]);
	inverter inv255(interconnections[254], interconnections[255]);
	inverter inv256(interconnections[255], interconnections[256]);
	inverter inv257(interconnections[256], interconnections[257]);
	inverter inv258(interconnections[257], interconnections[258]);
	inverter inv259(interconnections[258], interconnections[259]);
	inverter inv260(interconnections[259], interconnections[260]);
	inverter inv261(interconnections[260], interconnections[261]);
	inverter inv262(interconnections[261], interconnections[262]);
	inverter inv263(interconnections[262], interconnections[263]);
	inverter inv264(interconnections[263], interconnections[264]);
	inverter inv265(interconnections[264], interconnections[265]);
	inverter inv266(interconnections[265], interconnections[266]);
	inverter inv267(interconnections[266], interconnections[267]);
	inverter inv268(interconnections[267], interconnections[268]);
	inverter inv269(interconnections[268], interconnections[269]);
	inverter inv270(interconnections[269], interconnections[270]);
	inverter inv271(interconnections[270], interconnections[271]);
	inverter inv272(interconnections[271], interconnections[272]);
	inverter inv273(interconnections[272], interconnections[273]);
	inverter inv274(interconnections[273], interconnections[274]);
	inverter inv275(interconnections[274], interconnections[275]);
	inverter inv276(interconnections[275], interconnections[276]);
	inverter inv277(interconnections[276], interconnections[277]);
	inverter inv278(interconnections[277], interconnections[278]);
	inverter inv279(interconnections[278], interconnections[279]);
	inverter inv280(interconnections[279], interconnections[280]);
	inverter inv281(interconnections[280], interconnections[281]);
	inverter inv282(interconnections[281], interconnections[282]);
	inverter inv283(interconnections[282], interconnections[283]);
	inverter inv284(interconnections[283], interconnections[284]);
	inverter inv285(interconnections[284], interconnections[285]);
	inverter inv286(interconnections[285], interconnections[286]);
	inverter inv287(interconnections[286], interconnections[287]);
	inverter inv288(interconnections[287], interconnections[288]);
	inverter inv289(interconnections[288], interconnections[289]);
	inverter inv290(interconnections[289], interconnections[290]);
	inverter inv291(interconnections[290], interconnections[291]);
	inverter inv292(interconnections[291], interconnections[292]);
	inverter inv293(interconnections[292], interconnections[293]);
	inverter inv294(interconnections[293], interconnections[294]);
	inverter inv295(interconnections[294], interconnections[295]);
	inverter inv296(interconnections[295], interconnections[296]);
	inverter inv297(interconnections[296], interconnections[297]);
	inverter inv298(interconnections[297], interconnections[298]);
	inverter inv299(interconnections[298], interconnections[299]);
	inverter inv300(interconnections[299], interconnections[300]);
	inverter inv301(interconnections[300], interconnections[301]);
	inverter inv302(interconnections[301], interconnections[302]);
	inverter inv303(interconnections[302], interconnections[303]);
	inverter inv304(interconnections[303], interconnections[304]);
	inverter inv305(interconnections[304], interconnections[305]);
	inverter inv306(interconnections[305], interconnections[306]);
	inverter inv307(interconnections[306], interconnections[307]);
	inverter inv308(interconnections[307], interconnections[308]);
	inverter inv309(interconnections[308], interconnections[309]);
	inverter inv310(interconnections[309], interconnections[310]);
	inverter inv311(interconnections[310], interconnections[311]);
	inverter inv312(interconnections[311], interconnections[312]);
	inverter inv313(interconnections[312], interconnections[313]);
	inverter inv314(interconnections[313], interconnections[314]);
	inverter inv315(interconnections[314], interconnections[315]);
	inverter inv316(interconnections[315], interconnections[316]);
	inverter inv317(interconnections[316], interconnections[317]);
	inverter inv318(interconnections[317], interconnections[318]);
	inverter inv319(interconnections[318], interconnections[319]);
	inverter inv320(interconnections[319], interconnections[320]);
	inverter inv321(interconnections[320], interconnections[321]);
	inverter inv322(interconnections[321], interconnections[322]);
	inverter inv323(interconnections[322], interconnections[323]);
	inverter inv324(interconnections[323], interconnections[324]);
	inverter inv325(interconnections[324], interconnections[325]);
	inverter inv326(interconnections[325], interconnections[326]);
	inverter inv327(interconnections[326], interconnections[327]);
	inverter inv328(interconnections[327], interconnections[328]);
	inverter inv329(interconnections[328], interconnections[329]);
	inverter inv330(interconnections[329], interconnections[330]);
	inverter inv331(interconnections[330], interconnections[331]);
	inverter inv332(interconnections[331], interconnections[332]);
	inverter inv333(interconnections[332], interconnections[333]);
	inverter inv334(interconnections[333], interconnections[334]);
	inverter inv335(interconnections[334], interconnections[335]);
	inverter inv336(interconnections[335], interconnections[336]);
	inverter inv337(interconnections[336], interconnections[337]);
	inverter inv338(interconnections[337], interconnections[338]);
	inverter inv339(interconnections[338], interconnections[339]);
	inverter inv340(interconnections[339], interconnections[340]);
	inverter inv341(interconnections[340], interconnections[341]);
	inverter inv342(interconnections[341], interconnections[342]);
	inverter inv343(interconnections[342], interconnections[343]);
	inverter inv344(interconnections[343], interconnections[344]);
	inverter inv345(interconnections[344], interconnections[345]);
	inverter inv346(interconnections[345], interconnections[346]);
	inverter inv347(interconnections[346], interconnections[347]);
	inverter inv348(interconnections[347], interconnections[348]);
	inverter inv349(interconnections[348], interconnections[349]);
	inverter inv350(interconnections[349], interconnections[350]);
	inverter inv351(interconnections[350], interconnections[351]);
	inverter inv352(interconnections[351], interconnections[352]);
	inverter inv353(interconnections[352], interconnections[353]);
	inverter inv354(interconnections[353], interconnections[354]);
	inverter inv355(interconnections[354], interconnections[355]);
	inverter inv356(interconnections[355], interconnections[356]);
	inverter inv357(interconnections[356], interconnections[357]);
	inverter inv358(interconnections[357], interconnections[358]);
	inverter inv359(interconnections[358], interconnections[359]);
	inverter inv360(interconnections[359], interconnections[360]);
	inverter inv361(interconnections[360], interconnections[361]);
	inverter inv362(interconnections[361], interconnections[362]);
	inverter inv363(interconnections[362], interconnections[363]);
	inverter inv364(interconnections[363], interconnections[364]);
	inverter inv365(interconnections[364], interconnections[365]);
	inverter inv366(interconnections[365], interconnections[366]);
	inverter inv367(interconnections[366], interconnections[367]);
	inverter inv368(interconnections[367], interconnections[368]);
	inverter inv369(interconnections[368], interconnections[369]);
	inverter inv370(interconnections[369], interconnections[370]);
	inverter inv371(interconnections[370], interconnections[371]);
	inverter inv372(interconnections[371], interconnections[372]);
	inverter inv373(interconnections[372], interconnections[373]);
	inverter inv374(interconnections[373], interconnections[374]);
	inverter inv375(interconnections[374], interconnections[375]);
	inverter inv376(interconnections[375], interconnections[376]);
	inverter inv377(interconnections[376], interconnections[377]);
	inverter inv378(interconnections[377], interconnections[378]);
	inverter inv379(interconnections[378], interconnections[379]);
	inverter inv380(interconnections[379], interconnections[380]);
	inverter inv381(interconnections[380], interconnections[381]);
	inverter inv382(interconnections[381], interconnections[382]);
	inverter inv383(interconnections[382], interconnections[383]);
	inverter inv384(interconnections[383], interconnections[384]);
	inverter inv385(interconnections[384], interconnections[385]);
	inverter inv386(interconnections[385], interconnections[386]);
	inverter inv387(interconnections[386], interconnections[387]);
	inverter inv388(interconnections[387], interconnections[388]);
	inverter inv389(interconnections[388], interconnections[389]);
	inverter inv390(interconnections[389], interconnections[390]);
	inverter inv391(interconnections[390], interconnections[391]);
	inverter inv392(interconnections[391], interconnections[392]);
	inverter inv393(interconnections[392], interconnections[393]);
	inverter inv394(interconnections[393], interconnections[394]);
	inverter inv395(interconnections[394], interconnections[395]);
	inverter inv396(interconnections[395], interconnections[396]);
	inverter inv397(interconnections[396], interconnections[397]);
	inverter inv398(interconnections[397], interconnections[398]);
	inverter inv399(interconnections[398], interconnections[399]);
	inverter inv400(interconnections[399], interconnections[400]);
	inverter inv401(interconnections[400], interconnections[401]);
	inverter inv402(interconnections[401], interconnections[402]);
	inverter inv403(interconnections[402], interconnections[403]);
	inverter inv404(interconnections[403], interconnections[404]);
	inverter inv405(interconnections[404], interconnections[405]);
	inverter inv406(interconnections[405], interconnections[406]);
	inverter inv407(interconnections[406], interconnections[407]);
	inverter inv408(interconnections[407], interconnections[408]);
	inverter inv409(interconnections[408], interconnections[409]);
	inverter inv410(interconnections[409], interconnections[410]);
	inverter inv411(interconnections[410], interconnections[411]);
	inverter inv412(interconnections[411], interconnections[412]);
	inverter inv413(interconnections[412], interconnections[413]);
	inverter inv414(interconnections[413], interconnections[414]);
	inverter inv415(interconnections[414], interconnections[415]);
	inverter inv416(interconnections[415], interconnections[416]);
	inverter inv417(interconnections[416], interconnections[417]);
	inverter inv418(interconnections[417], interconnections[418]);
	inverter inv419(interconnections[418], interconnections[419]);
	inverter inv420(interconnections[419], interconnections[420]);
	inverter inv421(interconnections[420], interconnections[421]);
	inverter inv422(interconnections[421], interconnections[422]);
	inverter inv423(interconnections[422], interconnections[423]);
	inverter inv424(interconnections[423], interconnections[424]);
	inverter inv425(interconnections[424], interconnections[425]);
	inverter inv426(interconnections[425], interconnections[426]);
	inverter inv427(interconnections[426], interconnections[427]);
	inverter inv428(interconnections[427], interconnections[428]);
	inverter inv429(interconnections[428], interconnections[429]);
	inverter inv430(interconnections[429], interconnections[430]);
	inverter inv431(interconnections[430], interconnections[431]);
	inverter inv432(interconnections[431], interconnections[432]);
	inverter inv433(interconnections[432], interconnections[433]);
	inverter inv434(interconnections[433], interconnections[434]);
	inverter inv435(interconnections[434], interconnections[435]);
	inverter inv436(interconnections[435], interconnections[436]);
	inverter inv437(interconnections[436], interconnections[437]);
	inverter inv438(interconnections[437], interconnections[438]);
	inverter inv439(interconnections[438], interconnections[439]);
	inverter inv440(interconnections[439], interconnections[440]);
	inverter inv441(interconnections[440], interconnections[441]);
	inverter inv442(interconnections[441], interconnections[442]);
	inverter inv443(interconnections[442], interconnections[443]);
	inverter inv444(interconnections[443], interconnections[444]);
	inverter inv445(interconnections[444], interconnections[445]);
	inverter inv446(interconnections[445], interconnections[446]);
	inverter inv447(interconnections[446], interconnections[447]);
	inverter inv448(interconnections[447], interconnections[448]);
	inverter inv449(interconnections[448], interconnections[449]);
	inverter inv450(interconnections[449], interconnections[450]);
	inverter inv451(interconnections[450], interconnections[451]);
	inverter inv452(interconnections[451], interconnections[452]);
	inverter inv453(interconnections[452], interconnections[453]);
	inverter inv454(interconnections[453], interconnections[454]);
	inverter inv455(interconnections[454], interconnections[455]);
	inverter inv456(interconnections[455], interconnections[456]);
	inverter inv457(interconnections[456], interconnections[457]);
	inverter inv458(interconnections[457], interconnections[458]);
	inverter inv459(interconnections[458], interconnections[459]);
	inverter inv460(interconnections[459], interconnections[460]);
	inverter inv461(interconnections[460], interconnections[461]);
	inverter inv462(interconnections[461], interconnections[462]);
	inverter inv463(interconnections[462], interconnections[463]);
	inverter inv464(interconnections[463], interconnections[464]);
	inverter inv465(interconnections[464], interconnections[465]);
	inverter inv466(interconnections[465], interconnections[466]);
	inverter inv467(interconnections[466], interconnections[467]);
	inverter inv468(interconnections[467], interconnections[468]);
	inverter inv469(interconnections[468], interconnections[469]);
	inverter inv470(interconnections[469], interconnections[470]);
	inverter inv471(interconnections[470], interconnections[471]);
	inverter inv472(interconnections[471], interconnections[472]);
	inverter inv473(interconnections[472], interconnections[473]);
	inverter inv474(interconnections[473], interconnections[474]);
	inverter inv475(interconnections[474], interconnections[475]);
	inverter inv476(interconnections[475], interconnections[476]);
	inverter inv477(interconnections[476], interconnections[477]);
	inverter inv478(interconnections[477], interconnections[478]);
	inverter inv479(interconnections[478], interconnections[479]);
	inverter inv480(interconnections[479], interconnections[480]);
	inverter inv481(interconnections[480], interconnections[481]);
	inverter inv482(interconnections[481], interconnections[482]);
	inverter inv483(interconnections[482], interconnections[483]);
	inverter inv484(interconnections[483], interconnections[484]);
	inverter inv485(interconnections[484], interconnections[485]);
	inverter inv486(interconnections[485], interconnections[486]);
	inverter inv487(interconnections[486], interconnections[487]);
	inverter inv488(interconnections[487], interconnections[488]);
	inverter inv489(interconnections[488], interconnections[489]);
	inverter inv490(interconnections[489], interconnections[490]);
	inverter inv491(interconnections[490], interconnections[491]);
	inverter inv492(interconnections[491], interconnections[492]);
	inverter inv493(interconnections[492], interconnections[493]);
	inverter inv494(interconnections[493], interconnections[494]);
	inverter inv495(interconnections[494], interconnections[495]);
	inverter inv496(interconnections[495], interconnections[496]);
	inverter inv497(interconnections[496], interconnections[497]);
	inverter inv498(interconnections[497], interconnections[498]);
	inverter inv499(interconnections[498], interconnections[499]);
	inverter inv500(interconnections[499], interconnections[500]);
	inverter inv501(interconnections[500], interconnections[501]);
	inverter inv502(interconnections[501], interconnections[502]);
	inverter inv503(interconnections[502], interconnections[503]);
	inverter inv504(interconnections[503], interconnections[504]);
	inverter inv505(interconnections[504], interconnections[505]);
	inverter inv506(interconnections[505], interconnections[506]);
	inverter inv507(interconnections[506], interconnections[507]);
	inverter inv508(interconnections[507], interconnections[508]);
	inverter inv509(interconnections[508], interconnections[509]);
	inverter inv510(interconnections[509], interconnections[510]);
	inverter inv511(interconnections[510], interconnections[511]);
	inverter inv512(interconnections[511], interconnections[512]);
	inverter inv513(interconnections[512], interconnections[513]);
	inverter inv514(interconnections[513], interconnections[514]);
	inverter inv515(interconnections[514], interconnections[515]);
	inverter inv516(interconnections[515], interconnections[516]);
	inverter inv517(interconnections[516], interconnections[517]);
	inverter inv518(interconnections[517], interconnections[518]);
	inverter inv519(interconnections[518], interconnections[519]);
	inverter inv520(interconnections[519], interconnections[520]);
	inverter inv521(interconnections[520], interconnections[521]);
	inverter inv522(interconnections[521], interconnections[522]);
	inverter inv523(interconnections[522], interconnections[523]);
	inverter inv524(interconnections[523], interconnections[524]);
	inverter inv525(interconnections[524], interconnections[525]);
	inverter inv526(interconnections[525], interconnections[526]);
	inverter inv527(interconnections[526], interconnections[527]);
	inverter inv528(interconnections[527], interconnections[528]);
	inverter inv529(interconnections[528], interconnections[529]);
	inverter inv530(interconnections[529], interconnections[530]);
	inverter inv531(interconnections[530], out);
endmodule