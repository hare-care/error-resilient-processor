magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 271 1326 582
rect -38 261 199 271
rect 524 261 1326 271
<< pwell >>
rect 279 176 487 229
rect 735 176 932 203
rect 279 157 932 176
rect 1103 157 1287 203
rect 1 40 1287 157
rect 1 21 271 40
rect 516 21 1287 40
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 366 119 396 203
rect 476 66 506 150
rect 621 47 651 125
rect 716 47 746 131
rect 824 47 854 177
rect 1012 47 1042 131
rect 1084 47 1114 131
rect 1179 47 1209 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 446 413 476 497
rect 570 413 600 497
rect 642 413 672 497
rect 832 297 862 497
rect 927 369 957 497
rect 1084 369 1114 497
rect 1179 297 1209 497
<< ndiff >>
rect 27 102 79 131
rect 27 68 35 102
rect 69 68 79 102
rect 27 47 79 68
rect 109 89 163 131
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 102 245 131
rect 193 68 203 102
rect 237 68 245 102
rect 193 47 245 68
rect 305 165 366 203
rect 305 131 313 165
rect 347 131 366 165
rect 305 119 366 131
rect 396 150 461 203
rect 396 119 476 150
rect 411 66 476 119
rect 506 125 556 150
rect 761 131 824 177
rect 666 125 716 131
rect 506 112 621 125
rect 506 78 574 112
rect 608 78 621 112
rect 506 66 621 78
rect 542 47 621 66
rect 651 47 716 125
rect 746 106 824 131
rect 746 72 780 106
rect 814 72 824 106
rect 746 47 824 72
rect 854 107 906 177
rect 1129 131 1179 177
rect 854 73 864 107
rect 898 73 906 107
rect 854 47 906 73
rect 960 108 1012 131
rect 960 74 968 108
rect 1002 74 1012 108
rect 960 47 1012 74
rect 1042 47 1084 131
rect 1114 93 1179 131
rect 1114 59 1134 93
rect 1168 59 1179 93
rect 1114 47 1179 59
rect 1209 101 1261 177
rect 1209 67 1219 101
rect 1253 67 1261 101
rect 1209 47 1261 67
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 369 351 451
rect 381 413 446 497
rect 476 485 570 497
rect 476 451 511 485
rect 545 451 570 485
rect 476 413 570 451
rect 600 413 642 497
rect 672 477 724 497
rect 672 443 682 477
rect 716 443 724 477
rect 672 413 724 443
rect 778 471 832 497
rect 778 437 788 471
rect 822 437 832 471
rect 381 369 431 413
rect 778 368 832 437
rect 778 334 788 368
rect 822 334 832 368
rect 778 297 832 334
rect 862 471 927 497
rect 862 437 875 471
rect 909 437 927 471
rect 862 369 927 437
rect 957 485 1084 497
rect 957 451 1017 485
rect 1051 451 1084 485
rect 957 417 1084 451
rect 957 383 1017 417
rect 1051 383 1084 417
rect 957 369 1084 383
rect 1114 476 1179 497
rect 1114 442 1135 476
rect 1169 442 1179 476
rect 1114 369 1179 442
rect 862 297 912 369
rect 1129 297 1179 369
rect 1209 475 1261 497
rect 1209 441 1219 475
rect 1253 441 1261 475
rect 1209 349 1261 441
rect 1209 315 1219 349
rect 1253 315 1261 349
rect 1209 297 1261 315
<< ndiffc >>
rect 35 68 69 102
rect 119 55 153 89
rect 203 68 237 102
rect 313 131 347 165
rect 574 78 608 112
rect 780 72 814 106
rect 864 73 898 107
rect 968 74 1002 108
rect 1134 59 1168 93
rect 1219 67 1253 101
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 451 341 485
rect 511 451 545 485
rect 682 443 716 477
rect 788 437 822 471
rect 788 334 822 368
rect 875 437 909 471
rect 1017 451 1051 485
rect 1017 383 1051 417
rect 1135 442 1169 476
rect 1219 441 1253 475
rect 1219 315 1253 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 446 497 476 523
rect 570 497 600 523
rect 642 497 672 523
rect 832 497 862 523
rect 927 497 957 523
rect 1084 497 1114 523
rect 1179 497 1209 523
rect 446 375 476 413
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 272 193 363
rect 351 337 381 369
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 262 193 272
rect 326 321 381 337
rect 446 365 528 375
rect 446 331 478 365
rect 512 331 528 365
rect 446 321 528 331
rect 326 287 336 321
rect 370 287 381 321
rect 326 271 381 287
rect 570 279 600 413
rect 642 373 672 413
rect 642 357 746 373
rect 642 323 686 357
rect 720 323 746 357
rect 642 307 746 323
rect 118 228 134 262
rect 168 228 193 262
rect 118 218 193 228
rect 351 248 381 271
rect 476 249 600 279
rect 351 218 396 248
rect 46 176 76 214
rect 163 176 193 218
rect 366 203 396 218
rect 46 146 109 176
rect 79 131 109 146
rect 163 146 290 176
rect 163 131 193 146
rect 260 51 290 146
rect 476 150 506 249
rect 578 197 651 207
rect 578 163 594 197
rect 628 163 651 197
rect 578 153 651 163
rect 366 93 396 119
rect 621 125 651 153
rect 716 131 746 307
rect 832 265 862 297
rect 927 265 957 369
rect 1084 287 1114 369
rect 1038 271 1114 287
rect 791 249 862 265
rect 791 215 801 249
rect 835 215 862 249
rect 791 199 862 215
rect 904 249 958 265
rect 904 215 914 249
rect 948 215 958 249
rect 1038 237 1048 271
rect 1082 237 1114 271
rect 1179 265 1209 297
rect 1038 221 1114 237
rect 904 199 958 215
rect 824 177 854 199
rect 476 51 506 66
rect 79 21 109 47
rect 163 21 193 47
rect 260 21 506 51
rect 928 176 958 199
rect 928 146 1042 176
rect 1012 131 1042 146
rect 1084 131 1114 221
rect 1156 249 1210 265
rect 1156 215 1166 249
rect 1200 215 1210 249
rect 1156 199 1210 215
rect 1179 177 1209 199
rect 621 21 651 47
rect 716 21 746 47
rect 824 21 854 47
rect 1012 21 1042 47
rect 1084 21 1114 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 478 331 512 365
rect 336 287 370 321
rect 686 323 720 357
rect 134 228 168 262
rect 594 163 628 197
rect 801 215 835 249
rect 914 215 948 249
rect 1048 237 1082 271
rect 1166 215 1200 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 203 409 248 443
rect 290 485 363 527
rect 290 451 307 485
rect 341 451 363 485
rect 495 451 511 485
rect 545 451 645 485
rect 290 439 363 451
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 255 32 264
rect 17 221 29 255
rect 63 221 66 230
rect 17 197 66 221
rect 122 278 156 359
rect 237 405 248 409
rect 237 375 518 405
rect 203 371 518 375
rect 122 262 168 278
rect 122 228 134 262
rect 122 212 168 228
rect 122 157 156 212
rect 35 123 156 157
rect 35 102 69 123
rect 203 102 256 371
rect 478 365 518 371
rect 305 321 437 337
rect 305 287 336 321
rect 370 287 437 321
rect 35 52 69 68
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 237 68 256 102
rect 203 52 256 68
rect 296 165 362 181
rect 296 131 313 165
rect 347 131 362 165
rect 296 17 362 131
rect 397 77 437 287
rect 512 331 518 365
rect 478 197 518 331
rect 611 265 645 451
rect 679 477 739 527
rect 679 443 682 477
rect 716 443 739 477
rect 679 427 739 443
rect 782 471 826 487
rect 782 437 788 471
rect 822 437 826 471
rect 782 373 826 437
rect 862 471 919 527
rect 862 437 875 471
rect 909 437 919 471
rect 862 402 919 437
rect 1001 485 1067 493
rect 1001 451 1017 485
rect 1051 451 1067 485
rect 1001 417 1067 451
rect 1114 476 1184 527
rect 1114 442 1135 476
rect 1169 442 1184 476
rect 1114 426 1184 442
rect 1218 475 1271 491
rect 1218 441 1219 475
rect 1253 441 1271 475
rect 686 368 826 373
rect 1001 383 1017 417
rect 1051 383 1067 417
rect 1001 379 1067 383
rect 686 357 788 368
rect 720 334 788 357
rect 822 334 942 368
rect 1001 345 1184 379
rect 720 323 942 334
rect 686 307 942 323
rect 869 265 942 307
rect 1038 271 1102 287
rect 611 249 835 265
rect 611 231 801 249
rect 711 215 801 231
rect 711 199 835 215
rect 869 249 948 265
rect 869 215 914 249
rect 1038 255 1048 271
rect 1038 221 1042 255
rect 1082 237 1102 271
rect 1076 221 1102 237
rect 1150 265 1184 345
rect 1218 349 1271 441
rect 1218 315 1219 349
rect 1253 315 1271 349
rect 1218 299 1271 315
rect 1150 249 1200 265
rect 869 199 948 215
rect 1150 215 1166 249
rect 478 163 594 197
rect 628 163 644 197
rect 711 112 745 199
rect 869 123 916 199
rect 1150 187 1200 215
rect 987 153 1200 187
rect 987 124 1031 153
rect 558 78 574 112
rect 608 78 745 112
rect 779 106 829 122
rect 779 72 780 106
rect 814 72 829 106
rect 779 17 829 72
rect 864 107 916 123
rect 898 73 916 107
rect 864 51 916 73
rect 968 108 1031 124
rect 1234 119 1271 299
rect 1002 74 1031 108
rect 968 58 1031 74
rect 1134 93 1168 109
rect 1134 17 1168 59
rect 1211 101 1271 119
rect 1211 67 1219 101
rect 1253 67 1271 101
rect 1211 51 1271 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 230 32 255
rect 32 230 63 255
rect 29 221 63 230
rect 1042 237 1048 255
rect 1048 237 1076 255
rect 1042 221 1076 237
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 17 255 76 261
rect 17 221 29 255
rect 63 252 76 255
rect 1030 255 1088 261
rect 1030 252 1042 255
rect 63 224 1042 252
rect 63 221 76 224
rect 17 215 76 221
rect 1030 221 1042 224
rect 1076 221 1088 255
rect 1030 215 1088 221
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 305 289 339 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1225 85 1259 119 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1225 425 1259 459 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1225 357 1259 391 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_1
rlabel locali s 1038 221 1102 287 1 CLK
port 1 nsew clock input
rlabel metal1 s 1030 252 1088 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 1030 215 1088 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 17 252 76 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 17 224 1088 252 1 CLK
port 1 nsew clock input
rlabel metal1 s 17 215 76 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 0 -48 1288 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 2647380
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2637414
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 32.200 13.600 
<< end >>
