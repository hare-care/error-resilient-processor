magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< metal1 >>
rect 17258 3312 17458 3318
rect 17310 3260 17332 3312
rect 17384 3260 17406 3312
rect 4955 3087 5065 3249
rect 17258 3244 17458 3260
rect 17310 3192 17332 3244
rect 17384 3192 17406 3244
tri 17458 3236 17492 3270 sw
rect 18288 3223 18388 3267
rect 17258 3176 17458 3192
rect 17310 3124 17332 3176
rect 17384 3124 17406 3176
rect 17258 3118 17458 3124
rect 19567 3087 19677 3249
rect 18610 3058 18726 3064
rect 18610 2936 18726 2942
tri 18718 2928 18726 2936 nw
rect 18438 2842 18444 2894
rect 18496 2842 18508 2894
rect 18560 2842 18566 2894
rect 18516 1553 18568 1559
rect 18516 1489 18568 1501
tri 18379 1431 18412 1464 se
rect 18516 1431 18568 1437
tri 18378 1430 18379 1431 se
rect 18379 1430 18412 1431
rect 18336 1378 18342 1430
rect 18394 1378 18406 1430
rect 18458 1378 18464 1430
rect 7030 1199 7127 1232
rect 15261 1201 15381 1230
rect 1892 908 2026 1038
rect 1689 350 1715 444
rect 15961 178 16026 230
rect 16078 178 16091 230
rect 16143 178 16156 230
rect 16208 178 16214 230
rect 18780 213 18836 298
rect 15961 158 16214 178
tri 15919 84 15961 126 se
rect 15961 106 16026 158
rect 16078 106 16091 158
rect 16143 106 16156 158
rect 16208 106 16214 158
rect 15961 86 16214 106
tri 15957 34 15961 38 ne
rect 15961 34 16026 86
rect 16078 34 16091 86
rect 16143 34 16156 86
rect 16208 34 16214 86
<< via1 >>
rect 17258 3260 17310 3312
rect 17332 3260 17384 3312
rect 17406 3260 17458 3312
rect 17258 3192 17310 3244
rect 17332 3192 17384 3244
rect 17406 3192 17458 3244
rect 17258 3124 17310 3176
rect 17332 3124 17384 3176
rect 17406 3124 17458 3176
rect 18610 2942 18726 3058
rect 18444 2842 18496 2894
rect 18508 2842 18560 2894
rect 18516 1501 18568 1553
rect 18516 1437 18568 1489
rect 18342 1378 18394 1430
rect 18406 1378 18458 1430
rect 16026 178 16078 230
rect 16091 178 16143 230
rect 16156 178 16208 230
rect 16026 106 16078 158
rect 16091 106 16143 158
rect 16156 106 16208 158
rect 16026 34 16078 86
rect 16091 34 16143 86
rect 16156 34 16208 86
<< metal2 >>
rect 15928 3312 17458 3318
rect 152 3162 402 3292
rect 15928 3260 17258 3312
rect 17310 3260 17332 3312
rect 17384 3260 17406 3312
rect 15928 3244 17458 3260
rect 15928 3192 17258 3244
rect 17310 3192 17332 3244
rect 17384 3192 17406 3244
rect 15928 3176 17458 3192
rect 15928 3124 17258 3176
rect 17310 3124 17332 3176
rect 17384 3124 17406 3176
rect 15928 3118 17458 3124
rect 18610 3058 18961 3064
rect 4338 2922 4472 3010
rect 18726 2942 18961 3058
rect 18610 2936 18961 2942
tri 18839 2922 18853 2936 ne
rect 18853 2922 18961 2936
tri 18853 2894 18881 2922 ne
rect 18881 2894 18961 2922
rect 18438 2842 18444 2894
rect 18496 2842 18508 2894
rect 18560 2866 18710 2894
tri 18710 2866 18738 2894 sw
tri 18881 2866 18909 2894 ne
rect 18560 2842 18738 2866
tri 18738 2842 18762 2866 sw
tri 18688 2821 18709 2842 ne
rect 18709 2821 18762 2842
tri 18762 2821 18783 2842 sw
tri 18709 2820 18710 2821 ne
rect 18710 2820 18783 2821
tri 18710 2799 18731 2820 ne
rect 15949 2235 16017 2342
rect 93 2032 163 2076
rect 89 1953 180 1995
rect 94 1840 193 1878
rect 131 1741 213 1779
tri 17139 1701 17173 1735 se
tri 17225 1701 17259 1735 sw
rect 9870 1649 17899 1701
tri 17899 1649 17951 1701 sw
tri 17877 1621 17905 1649 ne
rect 17905 1621 17951 1649
rect 9870 1575 17725 1621
tri 17725 1575 17771 1621 sw
tri 17905 1575 17951 1621 ne
tri 17951 1581 18019 1649 sw
rect 17951 1575 18019 1581
tri 18019 1575 18025 1581 sw
rect 9870 1569 17771 1575
tri 17771 1569 17777 1575 sw
tri 17951 1569 17957 1575 ne
rect 17957 1569 18025 1575
tri 17703 1553 17719 1569 ne
rect 17719 1553 17777 1569
tri 17777 1553 17793 1569 sw
tri 17957 1553 17973 1569 ne
rect 17973 1559 18025 1569
tri 18025 1559 18041 1575 sw
rect 17973 1553 18568 1559
tri 17719 1533 17739 1553 ne
rect 17739 1533 17793 1553
rect 136 1493 256 1533
tri 17739 1507 17765 1533 ne
rect 17765 1507 17793 1533
tri 17793 1507 17839 1553 sw
tri 17973 1507 18019 1553 ne
rect 18019 1507 18516 1553
tri 17765 1501 17771 1507 ne
rect 17771 1501 17839 1507
tri 17839 1501 17845 1507 sw
tri 18482 1501 18488 1507 ne
rect 18488 1501 18516 1507
tri 17771 1495 17777 1501 ne
rect 17777 1495 17845 1501
tri 17845 1495 17851 1501 sw
tri 18488 1495 18494 1501 ne
rect 18494 1495 18568 1501
tri 17777 1493 17779 1495 ne
rect 17779 1493 17851 1495
tri 17779 1489 17783 1493 ne
rect 17783 1489 17851 1493
tri 17851 1489 17857 1495 sw
tri 18494 1489 18500 1495 ne
rect 18500 1489 18568 1495
tri 17783 1455 17817 1489 ne
rect 17817 1455 17857 1489
rect 132 1413 224 1455
tri 17817 1437 17835 1455 ne
rect 17835 1437 17857 1455
tri 17857 1437 17909 1489 sw
tri 18500 1473 18516 1489 ne
rect 18731 1486 18783 2820
tri 17835 1431 17841 1437 ne
rect 17841 1431 17909 1437
tri 17909 1431 17915 1437 sw
rect 18516 1431 18568 1437
tri 17841 1430 17842 1431 ne
rect 17842 1430 17915 1431
tri 17915 1430 17916 1431 sw
tri 17842 1421 17851 1430 ne
rect 17851 1421 18342 1430
tri 17851 1413 17859 1421 ne
rect 17859 1413 18342 1421
tri 17859 1378 17894 1413 ne
rect 17894 1378 18342 1413
rect 18394 1378 18406 1430
rect 18458 1378 18464 1430
tri 18835 885 18909 959 se
rect 18909 937 18961 2894
tri 18909 885 18961 937 nw
tri 18833 883 18835 885 se
rect 18835 883 18907 885
tri 18907 883 18909 885 nw
rect 18596 831 18855 883
tri 18855 831 18907 883 nw
rect 18251 539 18336 585
tri 16013 230 16047 264 sw
rect 3547 53 3842 215
rect 15947 178 16026 230
rect 16078 178 16091 230
rect 16143 178 16156 230
rect 16208 178 16214 230
rect 15947 158 16214 178
rect 15947 106 16026 158
rect 16078 106 16091 158
rect 16143 106 16156 158
rect 16208 106 16214 158
rect 15947 86 16214 106
rect 15947 34 16026 86
rect 16078 34 16091 86
rect 16143 34 16156 86
rect 16208 34 16214 86
use sky130_fd_io__gpio_ovtv2_in_buf  sky130_fd_io__gpio_ovtv2_in_buf_0
timestamp 1694700623
transform 1 0 0 0 1 0
box -2286 -894 17248 3318
use sky130_fd_io__gpio_ovtv2_ipath_hvls  sky130_fd_io__gpio_ovtv2_ipath_hvls_0
timestamp 1694700623
transform 0 -1 19756 1 0 1415
box -457 10 1903 2559
use sky130_fd_io__gpio_ovtv2_ipath_lvls  sky130_fd_io__gpio_ovtv2_ipath_lvls_0
timestamp 1694700623
transform 0 1 16241 1 0 -240
box -7 -228 1518 2676
<< labels >>
flabel metal2 s 136 1493 256 1533 3 FreeSans 200 0 0 0 IN_H
port 2 nsew
flabel metal2 s 132 1413 224 1455 3 FreeSans 200 0 0 0 IN_VT
port 3 nsew
flabel metal2 s 89 1953 180 1995 3 FreeSans 200 0 0 0 MODE_NORMAL_N
port 4 nsew
flabel metal2 s 93 2032 163 2076 3 FreeSans 200 0 0 0 MODE_VCCD_N
port 5 nsew
flabel metal2 s 94 1840 193 1878 3 FreeSans 200 0 0 0 MODE_REF_3V_N
port 6 nsew
flabel metal2 s 152 3162 402 3292 3 FreeSans 200 0 0 0 VDDIO_Q
port 7 nsew
flabel metal2 s 3547 53 3842 215 3 FreeSans 200 0 0 0 VSSD
port 8 nsew
flabel metal2 s 15949 2235 16017 2342 3 FreeSans 200 0 0 0 VREFIN
port 9 nsew
flabel metal2 s 18251 539 18336 585 3 FreeSans 200 0 0 0 IBUFMUX_OUT
port 10 nsew
flabel metal2 s 131 1741 213 1779 3 FreeSans 200 0 0 0 MODE_REF_N
port 11 nsew
flabel metal2 s 4338 2922 4472 3010 3 FreeSans 200 0 0 0 VCCHIB
port 12 nsew
flabel metal1 s 15261 1201 15381 1230 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 14 nsew
flabel metal1 s 7030 1199 7127 1232 3 FreeSans 200 0 0 0 EN_H_N
port 15 nsew
flabel metal1 s 1689 350 1715 444 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 16 nsew
flabel metal1 s 18780 213 18836 298 3 FreeSans 200 0 0 0 VCCHIB
port 12 nsew
flabel metal1 s 1892 908 2026 1038 3 FreeSans 200 0 0 0 VDDIO_Q
port 7 nsew
flabel metal1 s 4955 3087 5065 3249 3 FreeSans 200 0 0 0 VSSD
port 8 nsew
flabel metal1 s 19567 3087 19677 3249 3 FreeSans 200 0 0 0 VSSD
port 8 nsew
flabel metal1 s 18288 3223 18388 3267 3 FreeSans 200 0 0 0 IBUFMUX_OUT_H
port 17 nsew
<< properties >>
string GDS_END 36518896
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36512312
<< end >>
