magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal4 >>
rect 0 41065 1000 45908
rect 0 19915 1000 24908
rect 0 18725 1000 19615
rect 0 17555 1000 18445
rect 0 17189 1000 17255
rect 0 16533 1000 17129
rect 0 16237 1000 16473
rect 0 15581 1000 16177
rect 0 15455 1000 15521
rect 0 14225 1000 15155
rect 0 13255 1000 13945
rect 0 12285 1000 12975
rect 0 11075 1000 12005
rect 0 9865 1000 10795
rect 0 8895 1000 9585
rect 0 7685 1000 8615
rect 0 6315 1000 7405
<< properties >>
string GDS_END 12450
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11358
<< end >>
