magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 67 397 203
rect 30 17 63 67
rect 29 -17 63 17
<< scnmos >>
rect 108 93 138 177
rect 192 93 222 177
rect 289 93 319 177
<< scpmoshvt >>
rect 120 355 150 439
rect 192 355 222 439
rect 289 355 319 483
<< ndiff >>
rect 56 149 108 177
rect 56 115 64 149
rect 98 115 108 149
rect 56 93 108 115
rect 138 149 192 177
rect 138 115 148 149
rect 182 115 192 149
rect 138 93 192 115
rect 222 149 289 177
rect 222 115 244 149
rect 278 115 289 149
rect 222 93 289 115
rect 319 154 371 177
rect 319 120 329 154
rect 363 120 371 154
rect 319 93 371 120
<< pdiff >>
rect 237 459 289 483
rect 237 439 245 459
rect 68 407 120 439
rect 68 373 76 407
rect 110 373 120 407
rect 68 355 120 373
rect 150 355 192 439
rect 222 425 245 439
rect 279 425 289 459
rect 222 355 289 425
rect 319 461 387 483
rect 319 427 345 461
rect 379 427 387 461
rect 319 355 387 427
<< ndiffc >>
rect 64 115 98 149
rect 148 115 182 149
rect 244 115 278 149
rect 329 120 363 154
<< pdiffc >>
rect 76 373 110 407
rect 245 425 279 459
rect 345 427 379 461
<< poly >>
rect 289 483 319 509
rect 120 439 150 465
rect 192 439 222 465
rect 120 265 150 355
rect 50 249 150 265
rect 50 215 66 249
rect 100 215 150 249
rect 50 199 150 215
rect 192 265 222 355
rect 289 265 319 355
rect 192 249 246 265
rect 192 215 202 249
rect 236 215 246 249
rect 192 199 246 215
rect 289 249 355 265
rect 289 215 305 249
rect 339 215 355 249
rect 289 199 355 215
rect 108 177 138 199
rect 192 177 222 199
rect 289 177 319 199
rect 108 67 138 93
rect 192 67 222 93
rect 289 67 319 93
<< polycont >>
rect 66 215 100 249
rect 202 215 236 249
rect 305 215 339 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 229 459 295 527
rect 54 407 132 426
rect 229 425 245 459
rect 279 425 295 459
rect 329 461 436 493
rect 329 427 345 461
rect 379 427 436 461
rect 54 373 76 407
rect 110 391 132 407
rect 110 373 339 391
rect 54 357 339 373
rect 29 249 100 323
rect 29 215 66 249
rect 29 199 100 215
rect 134 165 168 357
rect 202 249 267 323
rect 236 215 267 249
rect 202 199 267 215
rect 305 249 339 357
rect 305 199 339 215
rect 373 165 436 427
rect 50 149 98 165
rect 50 115 64 149
rect 50 17 98 115
rect 134 149 190 165
rect 134 115 148 149
rect 182 115 190 149
rect 134 85 190 115
rect 236 149 279 165
rect 236 115 244 149
rect 278 115 279 149
rect 236 17 279 115
rect 313 154 436 165
rect 313 120 329 154
rect 363 120 436 154
rect 313 105 436 120
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or2_0
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 980036
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 976142
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.300 0.000 
<< end >>
