magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 54 43 476 283
rect -26 -43 506 43
<< mvnmos >>
rect 137 107 237 257
rect 293 107 393 257
<< mvpmos >>
rect 151 443 251 743
rect 293 443 393 743
<< mvndiff >>
rect 80 249 137 257
rect 80 215 92 249
rect 126 215 137 249
rect 80 149 137 215
rect 80 115 92 149
rect 126 115 137 149
rect 80 107 137 115
rect 237 249 293 257
rect 237 215 248 249
rect 282 215 293 249
rect 237 149 293 215
rect 237 115 248 149
rect 282 115 293 149
rect 237 107 293 115
rect 393 249 450 257
rect 393 215 404 249
rect 438 215 450 249
rect 393 149 450 215
rect 393 115 404 149
rect 438 115 450 149
rect 393 107 450 115
<< mvpdiff >>
rect 94 735 151 743
rect 94 701 106 735
rect 140 701 151 735
rect 94 655 151 701
rect 94 621 106 655
rect 140 621 151 655
rect 94 574 151 621
rect 94 540 106 574
rect 140 540 151 574
rect 94 494 151 540
rect 94 460 106 494
rect 140 460 151 494
rect 94 443 151 460
rect 251 443 293 743
rect 393 735 450 743
rect 393 701 404 735
rect 438 701 450 735
rect 393 652 450 701
rect 393 618 404 652
rect 438 618 450 652
rect 393 568 450 618
rect 393 534 404 568
rect 438 534 450 568
rect 393 485 450 534
rect 393 451 404 485
rect 438 451 450 485
rect 393 443 450 451
<< mvndiffc >>
rect 92 215 126 249
rect 92 115 126 149
rect 248 215 282 249
rect 248 115 282 149
rect 404 215 438 249
rect 404 115 438 149
<< mvpdiffc >>
rect 106 701 140 735
rect 106 621 140 655
rect 106 540 140 574
rect 106 460 140 494
rect 404 701 438 735
rect 404 618 438 652
rect 404 534 438 568
rect 404 451 438 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
<< poly >>
rect 151 743 251 769
rect 293 743 393 769
rect 151 417 251 443
rect 137 395 251 417
rect 137 361 165 395
rect 199 361 251 395
rect 137 283 251 361
rect 293 395 393 443
rect 293 361 315 395
rect 349 361 393 395
rect 137 257 237 283
rect 293 257 393 361
rect 137 81 237 107
rect 293 81 393 107
<< polycont >>
rect 165 361 199 395
rect 315 361 349 395
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 18 735 352 751
rect 18 701 24 735
rect 58 701 96 735
rect 140 701 168 735
rect 202 701 240 735
rect 274 701 312 735
rect 346 701 352 735
rect 18 655 352 701
rect 18 621 106 655
rect 140 621 352 655
rect 18 574 352 621
rect 18 540 106 574
rect 140 540 352 574
rect 18 494 352 540
rect 18 460 106 494
rect 140 460 352 494
rect 404 735 455 751
rect 438 701 455 735
rect 404 652 455 701
rect 438 618 455 652
rect 404 568 455 618
rect 438 534 455 568
rect 404 485 455 534
rect 438 451 455 485
rect 25 395 263 424
rect 25 361 165 395
rect 199 361 263 395
rect 25 355 263 361
rect 299 395 365 424
rect 299 361 315 395
rect 349 361 365 395
rect 299 355 365 361
rect 404 319 455 451
rect 240 285 455 319
rect 18 249 204 265
rect 18 215 92 249
rect 126 215 204 249
rect 18 149 204 215
rect 18 115 92 149
rect 126 115 204 149
rect 18 113 204 115
rect 18 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 204 113
rect 240 249 306 285
rect 240 215 248 249
rect 282 215 306 249
rect 240 149 306 215
rect 240 115 248 149
rect 282 115 306 149
rect 240 99 306 115
rect 344 215 404 249
rect 438 215 462 249
rect 344 149 462 215
rect 344 115 404 149
rect 438 115 462 149
rect 344 113 462 115
rect 18 73 204 79
rect 344 79 350 113
rect 384 79 422 113
rect 456 79 462 113
rect 344 73 462 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 24 701 58 735
rect 96 701 106 735
rect 106 701 130 735
rect 168 701 202 735
rect 240 701 274 735
rect 312 701 346 735
rect 22 79 56 113
rect 94 79 128 113
rect 166 79 200 113
rect 350 79 384 113
rect 422 79 456 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 240 735
rect 274 701 312 735
rect 346 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 350 113
rect 384 79 422 113
rect 456 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor2_1
flabel metal1 s 0 51 480 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 480 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 480 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 480 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 612 449 646 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 480 814
string GDS_END 195320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 187998
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
