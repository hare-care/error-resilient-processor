magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< metal1 >>
rect 101889 69433 101895 69485
rect 101947 69473 101953 69485
rect 103955 69473 103961 69485
rect 101947 69445 103961 69473
rect 101947 69433 101953 69445
rect 103955 69433 103961 69445
rect 104013 69433 104019 69485
rect 101765 69331 101771 69383
rect 101823 69371 101829 69383
rect 102787 69371 102793 69383
rect 101823 69343 102793 69371
rect 101823 69331 101829 69343
rect 102787 69331 102793 69343
rect 102845 69331 102851 69383
rect 101889 68532 101895 68584
rect 101947 68532 101953 68584
rect 101765 67042 101771 67094
rect 101823 67042 101829 67094
<< via1 >>
rect 101895 69433 101947 69485
rect 103961 69433 104013 69485
rect 101771 69331 101823 69383
rect 102793 69331 102845 69383
rect 101895 68532 101947 68584
rect 101771 67042 101823 67094
<< metal2 >>
rect 101895 69485 101947 69491
rect 101895 69427 101947 69433
rect 101771 69383 101823 69389
rect 101771 69325 101823 69331
rect 101783 67100 101811 69325
rect 101907 68590 101935 69427
rect 102805 69389 102833 70732
rect 103973 69491 104001 70732
rect 103961 69485 104013 69491
rect 103961 69427 104013 69433
rect 102793 69383 102845 69389
rect 102793 69325 102845 69331
rect 101895 68584 101947 68590
rect 101895 68526 101947 68532
rect 101771 67094 101823 67100
rect 101771 67036 101823 67042
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1694700623
transform 1 0 103955 0 1 69427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1694700623
transform 1 0 101889 0 1 68526
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1694700623
transform 1 0 101889 0 1 69427
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1694700623
transform 1 0 102787 0 1 69325
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1694700623
transform 1 0 101765 0 1 67036
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1694700623
transform 1 0 101765 0 1 69325
box 0 0 1 1
<< properties >>
string FIXED_BBOX 101765 67036 104019 70732
string GDS_END 12234198
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 12233110
<< end >>
