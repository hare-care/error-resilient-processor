magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 170 157 735 203
rect 69 21 735 157
rect 29 -17 63 17
<< locali >>
rect 21 65 67 333
rect 350 199 435 323
rect 474 199 526 323
rect 660 53 716 491
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 21 409 69 487
rect 103 445 173 527
rect 21 369 171 409
rect 103 233 171 369
rect 207 269 273 491
rect 307 397 343 491
rect 377 431 443 527
rect 478 397 512 491
rect 307 357 512 397
rect 103 53 149 233
rect 207 209 316 269
rect 189 17 238 173
rect 272 163 316 209
rect 565 299 622 527
rect 568 163 620 265
rect 272 125 620 163
rect 272 53 358 125
rect 474 17 620 91
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 350 199 435 323 6 A1
port 1 nsew signal input
rlabel locali s 474 199 526 323 6 A2
port 2 nsew signal input
rlabel locali s 21 65 67 333 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 660 53 716 491 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3983636
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3976090
<< end >>
