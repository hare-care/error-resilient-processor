magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 347 21 1863 157
rect 29 -17 63 17
<< locali >>
rect 123 333 157 493
rect 295 333 329 493
rect 467 333 501 493
rect 639 333 673 493
rect 811 333 845 493
rect 1016 333 1050 493
rect 1193 333 1227 493
rect 1365 333 1399 493
rect 1537 333 1571 493
rect 1709 333 1743 493
rect 1881 333 1915 493
rect 2053 333 2087 493
rect 123 291 2096 333
rect 465 283 1751 291
rect 465 56 510 283
rect 631 56 682 283
rect 803 56 851 283
rect 981 56 1051 283
rect 1185 56 1235 283
rect 1357 56 1407 283
rect 1529 56 1579 283
rect 1701 56 1751 283
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 22 459 88 493
rect 22 425 26 459
rect 60 425 88 459
rect 22 299 88 425
rect 193 459 259 493
rect 193 425 198 459
rect 232 425 259 459
rect 193 367 259 425
rect 365 459 431 493
rect 365 425 378 459
rect 412 425 431 459
rect 365 367 431 425
rect 537 459 603 493
rect 537 425 554 459
rect 588 425 603 459
rect 537 367 603 425
rect 709 459 775 493
rect 709 425 738 459
rect 772 425 775 459
rect 709 367 775 425
rect 885 459 951 493
rect 885 425 910 459
rect 944 425 951 459
rect 885 367 951 425
rect 1090 459 1156 493
rect 1124 425 1156 459
rect 1090 367 1156 425
rect 1263 459 1329 493
rect 1263 425 1274 459
rect 1308 425 1329 459
rect 1263 367 1329 425
rect 1435 459 1501 493
rect 1435 425 1446 459
rect 1480 425 1501 459
rect 1435 367 1501 425
rect 1607 459 1673 493
rect 1607 425 1626 459
rect 1660 425 1673 459
rect 1607 367 1673 425
rect 1779 459 1845 493
rect 1779 425 1792 459
rect 1826 425 1845 459
rect 1779 367 1845 425
rect 1951 459 2017 493
rect 1951 425 1964 459
rect 1998 425 2017 459
rect 1951 367 2017 425
rect 2122 459 2188 493
rect 2122 425 2144 459
rect 2178 425 2188 459
rect 2122 367 2188 425
rect 69 221 305 255
rect 339 221 397 255
rect 69 179 431 221
rect 371 17 425 122
rect 544 17 597 122
rect 716 17 769 122
rect 893 17 946 122
rect 1098 17 1151 122
rect 1270 17 1315 122
rect 1442 17 1495 122
rect 1614 17 1667 122
rect 1786 221 1869 255
rect 1903 221 1961 255
rect 1995 221 2142 255
rect 1786 179 2142 221
rect 1786 17 1839 122
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 26 425 60 459
rect 198 425 232 459
rect 378 425 412 459
rect 554 425 588 459
rect 738 425 772 459
rect 910 425 944 459
rect 1090 425 1124 459
rect 1274 425 1308 459
rect 1446 425 1480 459
rect 1626 425 1660 459
rect 1792 425 1826 459
rect 1964 425 1998 459
rect 2144 425 2178 459
rect 305 221 339 255
rect 397 221 431 255
rect 1869 221 1903 255
rect 1961 221 1995 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 14 459 2194 468
rect 14 425 26 459
rect 60 428 198 459
rect 60 425 72 428
rect 14 416 72 425
rect 186 425 198 428
rect 232 428 378 459
rect 232 425 244 428
rect 186 416 244 425
rect 366 425 378 428
rect 412 428 554 459
rect 412 425 424 428
rect 366 416 424 425
rect 542 425 554 428
rect 588 428 738 459
rect 588 425 600 428
rect 542 416 600 425
rect 726 425 738 428
rect 772 428 910 459
rect 772 425 784 428
rect 726 416 784 425
rect 898 425 910 428
rect 944 428 1090 459
rect 944 425 956 428
rect 898 416 956 425
rect 1078 425 1090 428
rect 1124 428 1274 459
rect 1124 425 1136 428
rect 1078 416 1136 425
rect 1262 425 1274 428
rect 1308 428 1446 459
rect 1308 425 1320 428
rect 1262 416 1320 425
rect 1434 425 1446 428
rect 1480 428 1626 459
rect 1480 425 1492 428
rect 1434 416 1492 425
rect 1614 425 1626 428
rect 1660 428 1792 459
rect 1660 425 1672 428
rect 1614 416 1672 425
rect 1780 425 1792 428
rect 1826 428 1964 459
rect 1826 425 1838 428
rect 1780 416 1838 425
rect 1952 425 1964 428
rect 1998 428 2144 459
rect 1998 425 2010 428
rect 1952 416 2010 425
rect 2132 425 2144 428
rect 2178 428 2194 459
rect 2178 425 2190 428
rect 2132 416 2190 425
rect 293 255 443 261
rect 293 221 305 255
rect 339 221 397 255
rect 431 252 443 255
rect 1857 255 2007 261
rect 1857 252 1869 255
rect 431 224 1869 252
rect 431 221 443 224
rect 293 215 443 221
rect 1857 221 1869 224
rect 1903 221 1961 255
rect 1995 221 2007 255
rect 1857 215 2007 221
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
rlabel metal1 s 1857 215 2007 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 215 443 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 224 2007 252 6 A
port 1 nsew signal input
rlabel metal1 s 1857 252 2007 261 6 A
port 1 nsew signal input
rlabel metal1 s 293 252 443 261 6 A
port 1 nsew signal input
rlabel metal1 s 2132 416 2190 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1952 416 2010 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1780 416 1838 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1614 416 1672 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1434 416 1492 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1262 416 1320 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1078 416 1136 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 898 416 956 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 726 416 784 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 542 416 600 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 186 416 244 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 416 72 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 2194 468 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 2208 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1701 56 1751 283 6 Y
port 7 nsew signal output
rlabel locali s 1529 56 1579 283 6 Y
port 7 nsew signal output
rlabel locali s 1357 56 1407 283 6 Y
port 7 nsew signal output
rlabel locali s 1185 56 1235 283 6 Y
port 7 nsew signal output
rlabel locali s 981 56 1051 283 6 Y
port 7 nsew signal output
rlabel locali s 803 56 851 283 6 Y
port 7 nsew signal output
rlabel locali s 631 56 682 283 6 Y
port 7 nsew signal output
rlabel locali s 465 56 510 283 6 Y
port 7 nsew signal output
rlabel locali s 465 283 1751 291 6 Y
port 7 nsew signal output
rlabel locali s 123 291 2096 333 6 Y
port 7 nsew signal output
rlabel locali s 2053 333 2087 493 6 Y
port 7 nsew signal output
rlabel locali s 1881 333 1915 493 6 Y
port 7 nsew signal output
rlabel locali s 1709 333 1743 493 6 Y
port 7 nsew signal output
rlabel locali s 1537 333 1571 493 6 Y
port 7 nsew signal output
rlabel locali s 1365 333 1399 493 6 Y
port 7 nsew signal output
rlabel locali s 1193 333 1227 493 6 Y
port 7 nsew signal output
rlabel locali s 1016 333 1050 493 6 Y
port 7 nsew signal output
rlabel locali s 811 333 845 493 6 Y
port 7 nsew signal output
rlabel locali s 639 333 673 493 6 Y
port 7 nsew signal output
rlabel locali s 467 333 501 493 6 Y
port 7 nsew signal output
rlabel locali s 295 333 329 493 6 Y
port 7 nsew signal output
rlabel locali s 123 333 157 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2318066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2302824
<< end >>
