magic
tech sky130B
magscale 1 2
timestamp 1694700623
use sky130_fd_pr__dfm1sd__example_55959141808173  sky130_fd_pr__dfm1sd__example_55959141808173_0
timestamp 1694700623
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808173  sky130_fd_pr__dfm1sd__example_55959141808173_1
timestamp 1694700623
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_0
timestamp 1694700623
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_1
timestamp 1694700623
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_2
timestamp 1694700623
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_3
timestamp 1694700623
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180831  sky130_fd_pr__hvdfm1sd2__example_5595914180831_4
timestamp 1694700623
transform 1 0 724 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 39450600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39446970
<< end >>
