magic
tech sky130B
magscale 1 2
timestamp 1694700623
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1694700623
transform 1 0 1452 0 1 0
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1694700623
transform -1 0 820 0 1 0
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1694700623
transform 1 0 2922 0 1 0
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1694700623
transform -1 0 2287 0 1 0
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1694700623
transform 1 0 2105 0 1 0
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1694700623
transform -1 0 1634 0 1 0
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1694700623
transform 1 0 638 0 1 0
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2v2  sky130_fd_io__hvsbt_nand2v2_0
timestamp 1694700623
transform 1 0 0 0 1 0
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1694700623
transform -1 0 3104 0 1 0
box 107 226 460 873
<< properties >>
string GDS_END 3199754
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3176790
<< end >>
