magic
tech sky130A
magscale 1 2
timestamp 1694700623
<< obsli1 >>
rect 137 1789 1813 1813
rect 137 1755 259 1789
rect 293 1755 332 1789
rect 366 1755 405 1789
rect 439 1755 478 1789
rect 512 1755 551 1789
rect 585 1755 625 1789
rect 659 1755 699 1789
rect 733 1755 773 1789
rect 807 1755 847 1789
rect 881 1755 921 1789
rect 955 1755 995 1789
rect 1029 1755 1069 1789
rect 1103 1755 1143 1789
rect 1177 1755 1217 1789
rect 1251 1755 1291 1789
rect 1325 1755 1365 1789
rect 1399 1755 1439 1789
rect 1473 1755 1513 1789
rect 1547 1755 1587 1789
rect 1621 1755 1661 1789
rect 1695 1755 1813 1789
rect 137 1731 1813 1755
rect 137 1696 219 1731
rect 137 1662 161 1696
rect 195 1662 219 1696
rect 137 1622 219 1662
rect 137 1588 161 1622
rect 195 1588 219 1622
rect 1731 1696 1813 1731
rect 1731 1662 1755 1696
rect 1789 1662 1813 1696
rect 1731 1622 1813 1662
rect 137 1548 219 1588
rect 137 1514 161 1548
rect 195 1514 219 1548
rect 137 1474 219 1514
rect 137 1440 161 1474
rect 195 1440 219 1474
rect 137 1400 219 1440
rect 137 1366 161 1400
rect 195 1366 219 1400
rect 137 1326 219 1366
rect 137 1292 161 1326
rect 195 1292 219 1326
rect 137 1252 219 1292
rect 137 1218 161 1252
rect 195 1218 219 1252
rect 137 1178 219 1218
rect 137 1144 161 1178
rect 195 1144 219 1178
rect 137 1104 219 1144
rect 332 1593 1616 1616
rect 332 1559 414 1593
rect 448 1559 487 1593
rect 521 1559 560 1593
rect 594 1559 633 1593
rect 667 1559 706 1593
rect 740 1559 779 1593
rect 813 1559 852 1593
rect 886 1559 924 1593
rect 958 1559 996 1593
rect 1030 1559 1068 1593
rect 1102 1559 1140 1593
rect 1174 1559 1212 1593
rect 1246 1559 1284 1593
rect 1318 1559 1356 1593
rect 1390 1559 1428 1593
rect 1462 1559 1616 1593
rect 332 1536 1616 1559
rect 332 1522 414 1536
rect 332 1488 355 1522
rect 389 1488 414 1522
rect 332 1437 414 1488
rect 332 1403 355 1437
rect 389 1403 414 1437
rect 332 1352 414 1403
rect 332 1318 355 1352
rect 389 1318 414 1352
rect 332 1267 414 1318
rect 332 1233 355 1267
rect 389 1233 414 1267
rect 332 1182 414 1233
rect 332 1148 355 1182
rect 389 1148 414 1182
rect 332 1136 414 1148
rect 1536 1534 1616 1536
rect 1536 1500 1559 1534
rect 1593 1500 1616 1534
rect 1536 1461 1616 1500
rect 1536 1427 1559 1461
rect 1593 1427 1616 1461
rect 1536 1388 1616 1427
rect 1536 1354 1559 1388
rect 1593 1354 1616 1388
rect 1536 1315 1616 1354
rect 1536 1281 1559 1315
rect 1593 1281 1616 1315
rect 1536 1242 1616 1281
rect 1536 1208 1559 1242
rect 1593 1208 1616 1242
rect 1536 1170 1616 1208
rect 1536 1136 1559 1170
rect 1593 1136 1616 1170
rect 137 1070 161 1104
rect 195 1070 219 1104
rect 1536 1098 1616 1136
rect 137 1030 219 1070
rect 137 996 161 1030
rect 195 996 219 1030
rect 137 956 219 996
rect 137 922 161 956
rect 195 922 219 956
rect 137 882 219 922
rect 137 848 161 882
rect 195 848 219 882
rect 261 1042 295 1076
rect 329 1042 367 1076
rect 401 1042 439 1076
rect 473 1042 1076 1076
rect 261 992 1076 1042
rect 261 958 295 992
rect 329 958 367 992
rect 401 958 439 992
rect 473 958 1076 992
rect 261 908 1076 958
rect 261 874 295 908
rect 329 874 367 908
rect 401 874 439 908
rect 473 874 1076 908
rect 1536 1064 1559 1098
rect 1593 1064 1616 1098
rect 1536 1026 1616 1064
rect 1536 992 1559 1026
rect 1593 992 1616 1026
rect 1536 954 1616 992
rect 1536 920 1559 954
rect 1593 920 1616 954
rect 1536 882 1616 920
rect 137 808 219 848
rect 1536 848 1559 882
rect 1593 848 1616 882
rect 137 774 161 808
rect 195 774 219 808
rect 137 734 219 774
rect 137 700 161 734
rect 195 700 219 734
rect 137 660 219 700
rect 137 626 161 660
rect 195 626 219 660
rect 137 586 219 626
rect 137 552 161 586
rect 195 552 219 586
rect 137 512 219 552
rect 137 478 161 512
rect 195 478 219 512
rect 137 439 219 478
rect 137 405 161 439
rect 195 405 219 439
rect 137 366 219 405
rect 137 332 161 366
rect 195 332 219 366
rect 332 801 414 813
rect 332 767 355 801
rect 389 767 414 801
rect 332 714 414 767
rect 332 680 355 714
rect 389 680 414 714
rect 332 626 414 680
rect 332 592 355 626
rect 389 592 414 626
rect 332 538 414 592
rect 332 504 355 538
rect 389 504 414 538
rect 332 450 414 504
rect 332 416 355 450
rect 389 416 414 450
rect 332 414 414 416
rect 1536 810 1616 848
rect 1536 776 1559 810
rect 1593 776 1616 810
rect 1536 738 1616 776
rect 1536 704 1559 738
rect 1593 704 1616 738
rect 1536 666 1616 704
rect 1536 632 1559 666
rect 1593 632 1616 666
rect 1536 594 1616 632
rect 1536 560 1559 594
rect 1593 560 1616 594
rect 1536 522 1616 560
rect 1536 488 1559 522
rect 1593 488 1616 522
rect 1536 414 1616 488
rect 332 391 1616 414
rect 332 357 486 391
rect 520 357 558 391
rect 592 357 630 391
rect 664 357 702 391
rect 736 357 774 391
rect 808 357 846 391
rect 880 357 918 391
rect 952 357 990 391
rect 1024 357 1062 391
rect 1096 357 1135 391
rect 1169 357 1208 391
rect 1242 357 1281 391
rect 1315 357 1354 391
rect 1388 357 1427 391
rect 1461 357 1500 391
rect 1534 357 1616 391
rect 332 334 1616 357
rect 1731 1588 1755 1622
rect 1789 1588 1813 1622
rect 1731 1548 1813 1588
rect 1731 1514 1755 1548
rect 1789 1514 1813 1548
rect 1731 1474 1813 1514
rect 1731 1440 1755 1474
rect 1789 1440 1813 1474
rect 1731 1400 1813 1440
rect 1731 1366 1755 1400
rect 1789 1366 1813 1400
rect 1731 1326 1813 1366
rect 1731 1292 1755 1326
rect 1789 1292 1813 1326
rect 1731 1252 1813 1292
rect 1731 1218 1755 1252
rect 1789 1218 1813 1252
rect 1731 1178 1813 1218
rect 1731 1144 1755 1178
rect 1789 1144 1813 1178
rect 1731 1104 1813 1144
rect 1731 1070 1755 1104
rect 1789 1070 1813 1104
rect 1731 1030 1813 1070
rect 1731 996 1755 1030
rect 1789 996 1813 1030
rect 1731 956 1813 996
rect 1731 922 1755 956
rect 1789 922 1813 956
rect 1731 882 1813 922
rect 1731 848 1755 882
rect 1789 848 1813 882
rect 1731 808 1813 848
rect 1731 774 1755 808
rect 1789 774 1813 808
rect 1731 734 1813 774
rect 1731 700 1755 734
rect 1789 700 1813 734
rect 1731 660 1813 700
rect 1731 626 1755 660
rect 1789 626 1813 660
rect 1731 586 1813 626
rect 1731 552 1755 586
rect 1789 552 1813 586
rect 1731 512 1813 552
rect 1731 478 1755 512
rect 1789 478 1813 512
rect 1731 439 1813 478
rect 1731 405 1755 439
rect 1789 405 1813 439
rect 1731 366 1813 405
rect 137 293 219 332
rect 137 259 161 293
rect 195 259 219 293
rect 137 219 219 259
rect 1731 332 1755 366
rect 1789 332 1813 366
rect 1731 293 1813 332
rect 1731 259 1755 293
rect 1789 259 1813 293
rect 1731 219 1813 259
rect 137 195 1813 219
rect 137 161 259 195
rect 293 161 332 195
rect 366 161 405 195
rect 439 161 478 195
rect 512 161 551 195
rect 585 161 625 195
rect 659 161 699 195
rect 733 161 773 195
rect 807 161 847 195
rect 881 161 921 195
rect 955 161 995 195
rect 1029 161 1069 195
rect 1103 161 1143 195
rect 1177 161 1217 195
rect 1251 161 1291 195
rect 1325 161 1365 195
rect 1399 161 1439 195
rect 1473 161 1513 195
rect 1547 161 1587 195
rect 1621 161 1661 195
rect 1695 161 1813 195
rect 137 137 1813 161
<< obsli1c >>
rect 259 1755 293 1789
rect 332 1755 366 1789
rect 405 1755 439 1789
rect 478 1755 512 1789
rect 551 1755 585 1789
rect 625 1755 659 1789
rect 699 1755 733 1789
rect 773 1755 807 1789
rect 847 1755 881 1789
rect 921 1755 955 1789
rect 995 1755 1029 1789
rect 1069 1755 1103 1789
rect 1143 1755 1177 1789
rect 1217 1755 1251 1789
rect 1291 1755 1325 1789
rect 1365 1755 1399 1789
rect 1439 1755 1473 1789
rect 1513 1755 1547 1789
rect 1587 1755 1621 1789
rect 1661 1755 1695 1789
rect 161 1662 195 1696
rect 161 1588 195 1622
rect 1755 1662 1789 1696
rect 161 1514 195 1548
rect 161 1440 195 1474
rect 161 1366 195 1400
rect 161 1292 195 1326
rect 161 1218 195 1252
rect 161 1144 195 1178
rect 414 1559 448 1593
rect 487 1559 521 1593
rect 560 1559 594 1593
rect 633 1559 667 1593
rect 706 1559 740 1593
rect 779 1559 813 1593
rect 852 1559 886 1593
rect 924 1559 958 1593
rect 996 1559 1030 1593
rect 1068 1559 1102 1593
rect 1140 1559 1174 1593
rect 1212 1559 1246 1593
rect 1284 1559 1318 1593
rect 1356 1559 1390 1593
rect 1428 1559 1462 1593
rect 355 1488 389 1522
rect 355 1403 389 1437
rect 355 1318 389 1352
rect 355 1233 389 1267
rect 355 1148 389 1182
rect 1559 1500 1593 1534
rect 1559 1427 1593 1461
rect 1559 1354 1593 1388
rect 1559 1281 1593 1315
rect 1559 1208 1593 1242
rect 1559 1136 1593 1170
rect 161 1070 195 1104
rect 161 996 195 1030
rect 161 922 195 956
rect 161 848 195 882
rect 295 1042 329 1076
rect 367 1042 401 1076
rect 439 1042 473 1076
rect 295 958 329 992
rect 367 958 401 992
rect 439 958 473 992
rect 295 874 329 908
rect 367 874 401 908
rect 439 874 473 908
rect 1559 1064 1593 1098
rect 1559 992 1593 1026
rect 1559 920 1593 954
rect 1559 848 1593 882
rect 161 774 195 808
rect 161 700 195 734
rect 161 626 195 660
rect 161 552 195 586
rect 161 478 195 512
rect 161 405 195 439
rect 161 332 195 366
rect 355 767 389 801
rect 355 680 389 714
rect 355 592 389 626
rect 355 504 389 538
rect 355 416 389 450
rect 1559 776 1593 810
rect 1559 704 1593 738
rect 1559 632 1593 666
rect 1559 560 1593 594
rect 1559 488 1593 522
rect 486 357 520 391
rect 558 357 592 391
rect 630 357 664 391
rect 702 357 736 391
rect 774 357 808 391
rect 846 357 880 391
rect 918 357 952 391
rect 990 357 1024 391
rect 1062 357 1096 391
rect 1135 357 1169 391
rect 1208 357 1242 391
rect 1281 357 1315 391
rect 1354 357 1388 391
rect 1427 357 1461 391
rect 1500 357 1534 391
rect 1755 1588 1789 1622
rect 1755 1514 1789 1548
rect 1755 1440 1789 1474
rect 1755 1366 1789 1400
rect 1755 1292 1789 1326
rect 1755 1218 1789 1252
rect 1755 1144 1789 1178
rect 1755 1070 1789 1104
rect 1755 996 1789 1030
rect 1755 922 1789 956
rect 1755 848 1789 882
rect 1755 774 1789 808
rect 1755 700 1789 734
rect 1755 626 1789 660
rect 1755 552 1789 586
rect 1755 478 1789 512
rect 1755 405 1789 439
rect 161 259 195 293
rect 1755 332 1789 366
rect 1755 259 1789 293
rect 259 161 293 195
rect 332 161 366 195
rect 405 161 439 195
rect 478 161 512 195
rect 551 161 585 195
rect 625 161 659 195
rect 699 161 733 195
rect 773 161 807 195
rect 847 161 881 195
rect 921 161 955 195
rect 995 161 1029 195
rect 1069 161 1103 195
rect 1143 161 1177 195
rect 1217 161 1251 195
rect 1291 161 1325 195
rect 1365 161 1399 195
rect 1439 161 1473 195
rect 1513 161 1547 195
rect 1587 161 1621 195
rect 1661 161 1695 195
<< metal1 >>
rect 142 1789 1808 1809
rect 142 1755 259 1789
rect 293 1755 332 1789
rect 366 1755 405 1789
rect 439 1755 478 1789
rect 512 1755 551 1789
rect 585 1755 625 1789
rect 659 1755 699 1789
rect 733 1755 773 1789
rect 807 1755 847 1789
rect 881 1755 921 1789
rect 955 1755 995 1789
rect 1029 1755 1069 1789
rect 1103 1755 1143 1789
rect 1177 1755 1217 1789
rect 1251 1755 1291 1789
rect 1325 1755 1365 1789
rect 1399 1755 1439 1789
rect 1473 1755 1513 1789
rect 1547 1755 1587 1789
rect 1621 1755 1661 1789
rect 1695 1755 1808 1789
rect 142 1737 1808 1755
rect 142 1696 214 1737
rect 142 1662 161 1696
rect 195 1662 214 1696
rect 142 1622 214 1662
rect 142 1588 161 1622
rect 195 1588 214 1622
rect 1736 1696 1808 1737
rect 1736 1662 1755 1696
rect 1789 1662 1808 1696
rect 1736 1622 1808 1662
rect 142 1548 214 1588
rect 142 1514 161 1548
rect 195 1514 214 1548
rect 142 1474 214 1514
rect 142 1440 161 1474
rect 195 1440 214 1474
rect 142 1400 214 1440
rect 142 1366 161 1400
rect 195 1366 214 1400
rect 142 1326 214 1366
rect 142 1292 161 1326
rect 195 1292 214 1326
rect 142 1252 214 1292
rect 142 1218 161 1252
rect 195 1218 214 1252
rect 142 1178 214 1218
rect 142 1144 161 1178
rect 195 1144 214 1178
rect 142 1104 214 1144
rect 336 1593 1612 1612
rect 336 1559 414 1593
rect 448 1559 487 1593
rect 521 1559 560 1593
rect 594 1559 633 1593
rect 667 1559 706 1593
rect 740 1559 779 1593
rect 813 1559 852 1593
rect 886 1559 924 1593
rect 958 1559 996 1593
rect 1030 1559 1068 1593
rect 1102 1559 1140 1593
rect 1174 1559 1212 1593
rect 1246 1559 1284 1593
rect 1318 1559 1356 1593
rect 1390 1559 1428 1593
rect 1462 1559 1612 1593
rect 336 1540 1612 1559
rect 336 1522 408 1540
rect 336 1488 355 1522
rect 389 1488 408 1522
rect 336 1437 408 1488
rect 336 1403 355 1437
rect 389 1403 408 1437
rect 336 1352 408 1403
rect 336 1318 355 1352
rect 389 1318 408 1352
rect 336 1267 408 1318
rect 336 1233 355 1267
rect 389 1233 408 1267
rect 336 1182 408 1233
rect 336 1148 355 1182
rect 389 1148 408 1182
rect 336 1136 408 1148
rect 1540 1534 1612 1540
rect 1540 1500 1559 1534
rect 1593 1500 1612 1534
rect 1540 1461 1612 1500
rect 1540 1427 1559 1461
rect 1593 1427 1612 1461
rect 1540 1388 1612 1427
rect 1540 1354 1559 1388
rect 1593 1354 1612 1388
rect 1540 1315 1612 1354
rect 1540 1281 1559 1315
rect 1593 1281 1612 1315
rect 1540 1242 1612 1281
rect 1540 1208 1559 1242
rect 1593 1208 1612 1242
rect 1540 1170 1612 1208
rect 1540 1136 1559 1170
rect 1593 1136 1612 1170
rect 142 1070 161 1104
rect 195 1070 214 1104
rect 1540 1098 1612 1136
rect 142 1030 214 1070
rect 142 996 161 1030
rect 195 996 214 1030
rect 142 956 214 996
rect 142 922 161 956
rect 195 922 214 956
rect 142 882 214 922
rect 142 848 161 882
rect 195 848 214 882
rect 289 1076 479 1088
rect 289 1042 295 1076
rect 329 1042 367 1076
rect 401 1042 439 1076
rect 473 1042 479 1076
rect 289 992 479 1042
rect 289 958 295 992
rect 329 958 367 992
rect 401 958 439 992
rect 473 958 479 992
rect 289 908 479 958
rect 289 874 295 908
rect 329 874 367 908
rect 401 874 439 908
rect 473 874 479 908
rect 289 862 479 874
rect 1540 1064 1559 1098
rect 1593 1064 1612 1098
rect 1540 1026 1612 1064
rect 1540 992 1559 1026
rect 1593 992 1612 1026
rect 1540 954 1612 992
rect 1540 920 1559 954
rect 1593 920 1612 954
rect 1540 882 1612 920
rect 142 808 214 848
rect 1540 848 1559 882
rect 1593 848 1612 882
rect 142 774 161 808
rect 195 774 214 808
rect 142 734 214 774
rect 142 700 161 734
rect 195 700 214 734
rect 142 660 214 700
rect 142 626 161 660
rect 195 626 214 660
rect 142 586 214 626
rect 142 552 161 586
rect 195 552 214 586
rect 142 512 214 552
rect 142 478 161 512
rect 195 478 214 512
rect 142 439 214 478
rect 142 405 161 439
rect 195 405 214 439
rect 142 366 214 405
rect 142 332 161 366
rect 195 332 214 366
rect 336 801 408 813
rect 336 767 355 801
rect 389 767 408 801
rect 336 714 408 767
rect 336 680 355 714
rect 389 680 408 714
rect 336 626 408 680
rect 336 592 355 626
rect 389 592 408 626
rect 336 538 408 592
rect 336 504 355 538
rect 389 504 408 538
rect 336 450 408 504
rect 336 416 355 450
rect 389 416 408 450
rect 336 410 408 416
rect 1540 810 1612 848
rect 1540 776 1559 810
rect 1593 776 1612 810
rect 1540 738 1612 776
rect 1540 704 1559 738
rect 1593 704 1612 738
rect 1540 666 1612 704
rect 1540 632 1559 666
rect 1593 632 1612 666
rect 1540 594 1612 632
rect 1540 560 1559 594
rect 1593 560 1612 594
rect 1540 522 1612 560
rect 1540 488 1559 522
rect 1593 488 1612 522
rect 1540 410 1612 488
rect 336 391 1612 410
rect 336 357 486 391
rect 520 357 558 391
rect 592 357 630 391
rect 664 357 702 391
rect 736 357 774 391
rect 808 357 846 391
rect 880 357 918 391
rect 952 357 990 391
rect 1024 357 1062 391
rect 1096 357 1135 391
rect 1169 357 1208 391
rect 1242 357 1281 391
rect 1315 357 1354 391
rect 1388 357 1427 391
rect 1461 357 1500 391
rect 1534 357 1612 391
rect 336 338 1612 357
rect 1736 1588 1755 1622
rect 1789 1588 1808 1622
rect 1736 1548 1808 1588
rect 1736 1514 1755 1548
rect 1789 1514 1808 1548
rect 1736 1474 1808 1514
rect 1736 1440 1755 1474
rect 1789 1440 1808 1474
rect 1736 1400 1808 1440
rect 1736 1366 1755 1400
rect 1789 1366 1808 1400
rect 1736 1326 1808 1366
rect 1736 1292 1755 1326
rect 1789 1292 1808 1326
rect 1736 1252 1808 1292
rect 1736 1218 1755 1252
rect 1789 1218 1808 1252
rect 1736 1178 1808 1218
rect 1736 1144 1755 1178
rect 1789 1144 1808 1178
rect 1736 1104 1808 1144
rect 1736 1070 1755 1104
rect 1789 1070 1808 1104
rect 1736 1030 1808 1070
rect 1736 996 1755 1030
rect 1789 996 1808 1030
rect 1736 956 1808 996
rect 1736 922 1755 956
rect 1789 922 1808 956
rect 1736 882 1808 922
rect 1736 848 1755 882
rect 1789 848 1808 882
rect 1736 808 1808 848
rect 1736 774 1755 808
rect 1789 774 1808 808
rect 1736 734 1808 774
rect 1736 700 1755 734
rect 1789 700 1808 734
rect 1736 660 1808 700
rect 1736 626 1755 660
rect 1789 626 1808 660
rect 1736 586 1808 626
rect 1736 552 1755 586
rect 1789 552 1808 586
rect 1736 512 1808 552
rect 1736 478 1755 512
rect 1789 478 1808 512
rect 1736 439 1808 478
rect 1736 405 1755 439
rect 1789 405 1808 439
rect 1736 366 1808 405
rect 142 293 214 332
rect 142 259 161 293
rect 195 259 214 293
rect 142 214 214 259
rect 1736 332 1755 366
rect 1789 332 1808 366
rect 1736 293 1808 332
rect 1736 259 1755 293
rect 1789 259 1808 293
rect 1736 214 1808 259
rect 142 195 1808 214
rect 142 161 259 195
rect 293 161 332 195
rect 366 161 405 195
rect 439 161 478 195
rect 512 161 551 195
rect 585 161 625 195
rect 659 161 699 195
rect 733 161 773 195
rect 807 161 847 195
rect 881 161 921 195
rect 955 161 995 195
rect 1029 161 1069 195
rect 1103 161 1143 195
rect 1177 161 1217 195
rect 1251 161 1291 195
rect 1325 161 1365 195
rect 1399 161 1439 195
rect 1473 161 1513 195
rect 1547 161 1587 195
rect 1621 161 1661 195
rect 1695 161 1808 195
rect 142 142 1808 161
<< labels >>
rlabel metal1 s 1540 410 1612 1540 6 B
port 1 nsew
rlabel metal1 s 336 1540 1612 1612 6 B
port 1 nsew
rlabel metal1 s 336 1136 408 1540 6 B
port 1 nsew
rlabel metal1 s 336 410 408 813 6 B
port 1 nsew
rlabel metal1 s 336 338 1612 410 6 B
port 1 nsew
rlabel metal1 s 1736 214 1808 1737 6 C
port 2 nsew
rlabel metal1 s 142 1737 1808 1809 6 C
port 2 nsew
rlabel metal1 s 142 214 214 1737 6 C
port 2 nsew
rlabel metal1 s 142 142 1808 214 6 C
port 2 nsew
rlabel metal1 s 289 862 479 1088 6 E
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1950 1950
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__npn_11v0_W1p00L1p00
string library sky130
string parameter m=1
string GDS_END 9109982
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9086230
<< end >>
