magic
tech sky130B
magscale 1 2
timestamp 1694700623
<< nwell >>
rect 7397 350 11245 3602
<< pwell >>
rect 7207 3602 11425 3782
rect 7207 350 7397 3602
rect 11245 350 11425 3602
rect 7207 170 11425 350
<< mvpsubdiff >>
rect 7233 3732 11399 3756
rect 7233 3698 7353 3732
rect 7387 3698 7421 3732
rect 7455 3698 7489 3732
rect 7523 3698 7557 3732
rect 7591 3698 7625 3732
rect 7659 3698 7693 3732
rect 7727 3698 7761 3732
rect 7795 3698 7829 3732
rect 7863 3698 7897 3732
rect 7931 3698 7965 3732
rect 7999 3698 8033 3732
rect 8067 3698 8101 3732
rect 8135 3698 8169 3732
rect 8203 3698 8237 3732
rect 8271 3698 8305 3732
rect 8339 3698 8373 3732
rect 8407 3698 8441 3732
rect 8475 3698 8509 3732
rect 8543 3698 8577 3732
rect 8611 3698 8645 3732
rect 8679 3698 8713 3732
rect 8747 3698 8781 3732
rect 8815 3698 8849 3732
rect 8883 3698 8917 3732
rect 8951 3698 8985 3732
rect 9019 3698 9053 3732
rect 9087 3698 9121 3732
rect 9155 3698 9189 3732
rect 9223 3698 9257 3732
rect 9291 3698 9325 3732
rect 9359 3698 9393 3732
rect 9427 3698 9461 3732
rect 9495 3698 9529 3732
rect 9563 3698 9597 3732
rect 9631 3698 9665 3732
rect 9699 3698 9733 3732
rect 9767 3698 9801 3732
rect 9835 3698 9869 3732
rect 9903 3698 9937 3732
rect 9971 3698 10005 3732
rect 10039 3698 10073 3732
rect 10107 3698 10141 3732
rect 10175 3698 10209 3732
rect 10243 3698 10277 3732
rect 10311 3698 10345 3732
rect 10379 3698 10413 3732
rect 10447 3698 10481 3732
rect 10515 3698 10549 3732
rect 10583 3698 10617 3732
rect 10651 3698 10685 3732
rect 10719 3698 10753 3732
rect 10787 3698 10821 3732
rect 10855 3698 10889 3732
rect 10923 3698 10957 3732
rect 10991 3698 11025 3732
rect 11059 3698 11093 3732
rect 11127 3698 11161 3732
rect 11195 3698 11229 3732
rect 11263 3698 11399 3732
rect 7233 3628 11399 3698
rect 7233 3625 7371 3628
rect 7233 3591 7267 3625
rect 7301 3591 7371 3625
rect 7233 3557 7371 3591
rect 7233 3523 7267 3557
rect 7301 3523 7371 3557
rect 7233 3489 7371 3523
rect 7233 3455 7267 3489
rect 7301 3455 7371 3489
rect 11271 3625 11399 3628
rect 11271 3591 11341 3625
rect 11375 3591 11399 3625
rect 11271 3557 11399 3591
rect 11271 3523 11341 3557
rect 11375 3523 11399 3557
rect 11271 3489 11399 3523
rect 7233 3421 7371 3455
rect 7233 3387 7267 3421
rect 7301 3387 7371 3421
rect 7233 3353 7371 3387
rect 7233 3319 7267 3353
rect 7301 3319 7371 3353
rect 7233 3285 7371 3319
rect 7233 3251 7267 3285
rect 7301 3251 7371 3285
rect 7233 3217 7371 3251
rect 7233 3183 7267 3217
rect 7301 3183 7371 3217
rect 7233 3149 7371 3183
rect 7233 3115 7267 3149
rect 7301 3115 7371 3149
rect 7233 3081 7371 3115
rect 7233 3047 7267 3081
rect 7301 3047 7371 3081
rect 7233 3013 7371 3047
rect 7233 2979 7267 3013
rect 7301 2979 7371 3013
rect 7233 2945 7371 2979
rect 7233 2911 7267 2945
rect 7301 2911 7371 2945
rect 7233 2877 7371 2911
rect 7233 2843 7267 2877
rect 7301 2843 7371 2877
rect 7233 2809 7371 2843
rect 7233 2775 7267 2809
rect 7301 2775 7371 2809
rect 7233 2741 7371 2775
rect 7233 2707 7267 2741
rect 7301 2707 7371 2741
rect 7233 2673 7371 2707
rect 7233 2639 7267 2673
rect 7301 2639 7371 2673
rect 7233 2605 7371 2639
rect 7233 2571 7267 2605
rect 7301 2571 7371 2605
rect 7233 2537 7371 2571
rect 7233 2503 7267 2537
rect 7301 2503 7371 2537
rect 7233 2469 7371 2503
rect 7233 2435 7267 2469
rect 7301 2435 7371 2469
rect 7233 2401 7371 2435
rect 7233 2367 7267 2401
rect 7301 2367 7371 2401
rect 7233 2333 7371 2367
rect 7233 2299 7267 2333
rect 7301 2299 7371 2333
rect 7233 2265 7371 2299
rect 7233 2231 7267 2265
rect 7301 2231 7371 2265
rect 7233 2197 7371 2231
rect 7233 2163 7267 2197
rect 7301 2163 7371 2197
rect 7233 2129 7371 2163
rect 7233 2095 7267 2129
rect 7301 2095 7371 2129
rect 7233 2061 7371 2095
rect 7233 2027 7267 2061
rect 7301 2027 7371 2061
rect 7233 1993 7371 2027
rect 7233 1959 7267 1993
rect 7301 1959 7371 1993
rect 7233 1925 7371 1959
rect 7233 1891 7267 1925
rect 7301 1891 7371 1925
rect 7233 1857 7371 1891
rect 7233 1823 7267 1857
rect 7301 1823 7371 1857
rect 7233 1789 7371 1823
rect 7233 1755 7267 1789
rect 7301 1755 7371 1789
rect 7233 1721 7371 1755
rect 7233 1687 7267 1721
rect 7301 1687 7371 1721
rect 7233 1653 7371 1687
rect 7233 1619 7267 1653
rect 7301 1619 7371 1653
rect 7233 1585 7371 1619
rect 7233 1551 7267 1585
rect 7301 1551 7371 1585
rect 7233 1517 7371 1551
rect 7233 1483 7267 1517
rect 7301 1483 7371 1517
rect 7233 1449 7371 1483
rect 7233 1415 7267 1449
rect 7301 1415 7371 1449
rect 7233 1381 7371 1415
rect 7233 1347 7267 1381
rect 7301 1347 7371 1381
rect 7233 1313 7371 1347
rect 7233 1279 7267 1313
rect 7301 1279 7371 1313
rect 7233 1245 7371 1279
rect 7233 1211 7267 1245
rect 7301 1211 7371 1245
rect 7233 1177 7371 1211
rect 7233 1143 7267 1177
rect 7301 1143 7371 1177
rect 7233 1109 7371 1143
rect 7233 1075 7267 1109
rect 7301 1075 7371 1109
rect 7233 1041 7371 1075
rect 7233 1007 7267 1041
rect 7301 1007 7371 1041
rect 7233 973 7371 1007
rect 7233 939 7267 973
rect 7301 939 7371 973
rect 7233 905 7371 939
rect 7233 871 7267 905
rect 7301 871 7371 905
rect 7233 837 7371 871
rect 7233 803 7267 837
rect 7301 803 7371 837
rect 7233 769 7371 803
rect 7233 735 7267 769
rect 7301 735 7371 769
rect 7233 701 7371 735
rect 7233 667 7267 701
rect 7301 667 7371 701
rect 7233 633 7371 667
rect 7233 599 7267 633
rect 7301 599 7371 633
rect 7233 565 7371 599
rect 7233 531 7267 565
rect 7301 531 7371 565
rect 7233 497 7371 531
rect 7233 463 7267 497
rect 7301 463 7371 497
rect 11271 3455 11341 3489
rect 11375 3455 11399 3489
rect 11271 3421 11399 3455
rect 11271 3387 11341 3421
rect 11375 3387 11399 3421
rect 11271 3353 11399 3387
rect 11271 3319 11341 3353
rect 11375 3319 11399 3353
rect 11271 3285 11399 3319
rect 11271 3251 11341 3285
rect 11375 3251 11399 3285
rect 11271 3217 11399 3251
rect 11271 3183 11341 3217
rect 11375 3183 11399 3217
rect 11271 3149 11399 3183
rect 11271 3115 11341 3149
rect 11375 3115 11399 3149
rect 11271 3081 11399 3115
rect 11271 3047 11341 3081
rect 11375 3047 11399 3081
rect 11271 3013 11399 3047
rect 11271 2979 11341 3013
rect 11375 2979 11399 3013
rect 11271 2945 11399 2979
rect 11271 2911 11341 2945
rect 11375 2911 11399 2945
rect 11271 2877 11399 2911
rect 11271 2843 11341 2877
rect 11375 2843 11399 2877
rect 11271 2809 11399 2843
rect 11271 2775 11341 2809
rect 11375 2775 11399 2809
rect 11271 2741 11399 2775
rect 11271 2707 11341 2741
rect 11375 2707 11399 2741
rect 11271 2673 11399 2707
rect 11271 2639 11341 2673
rect 11375 2639 11399 2673
rect 11271 2605 11399 2639
rect 11271 2571 11341 2605
rect 11375 2571 11399 2605
rect 11271 2537 11399 2571
rect 11271 2503 11341 2537
rect 11375 2503 11399 2537
rect 11271 2469 11399 2503
rect 11271 2435 11341 2469
rect 11375 2435 11399 2469
rect 11271 2401 11399 2435
rect 11271 2367 11341 2401
rect 11375 2367 11399 2401
rect 11271 2333 11399 2367
rect 11271 2299 11341 2333
rect 11375 2299 11399 2333
rect 11271 2265 11399 2299
rect 11271 2231 11341 2265
rect 11375 2231 11399 2265
rect 11271 2197 11399 2231
rect 11271 2163 11341 2197
rect 11375 2163 11399 2197
rect 11271 2129 11399 2163
rect 11271 2095 11341 2129
rect 11375 2095 11399 2129
rect 11271 2061 11399 2095
rect 11271 2027 11341 2061
rect 11375 2027 11399 2061
rect 11271 1993 11399 2027
rect 11271 1959 11341 1993
rect 11375 1959 11399 1993
rect 11271 1925 11399 1959
rect 11271 1891 11341 1925
rect 11375 1891 11399 1925
rect 11271 1857 11399 1891
rect 11271 1823 11341 1857
rect 11375 1823 11399 1857
rect 11271 1789 11399 1823
rect 11271 1755 11341 1789
rect 11375 1755 11399 1789
rect 11271 1721 11399 1755
rect 11271 1687 11341 1721
rect 11375 1687 11399 1721
rect 11271 1653 11399 1687
rect 11271 1619 11341 1653
rect 11375 1619 11399 1653
rect 11271 1585 11399 1619
rect 11271 1551 11341 1585
rect 11375 1551 11399 1585
rect 11271 1517 11399 1551
rect 11271 1483 11341 1517
rect 11375 1483 11399 1517
rect 11271 1449 11399 1483
rect 11271 1415 11341 1449
rect 11375 1415 11399 1449
rect 11271 1381 11399 1415
rect 11271 1347 11341 1381
rect 11375 1347 11399 1381
rect 11271 1313 11399 1347
rect 11271 1279 11341 1313
rect 11375 1279 11399 1313
rect 11271 1245 11399 1279
rect 11271 1211 11341 1245
rect 11375 1211 11399 1245
rect 11271 1177 11399 1211
rect 11271 1143 11341 1177
rect 11375 1143 11399 1177
rect 11271 1109 11399 1143
rect 11271 1075 11341 1109
rect 11375 1075 11399 1109
rect 11271 1041 11399 1075
rect 11271 1007 11341 1041
rect 11375 1007 11399 1041
rect 11271 973 11399 1007
rect 11271 939 11341 973
rect 11375 939 11399 973
rect 11271 905 11399 939
rect 11271 871 11341 905
rect 11375 871 11399 905
rect 11271 837 11399 871
rect 11271 803 11341 837
rect 11375 803 11399 837
rect 11271 769 11399 803
rect 11271 735 11341 769
rect 11375 735 11399 769
rect 11271 701 11399 735
rect 11271 667 11341 701
rect 11375 667 11399 701
rect 11271 633 11399 667
rect 11271 599 11341 633
rect 11375 599 11399 633
rect 11271 565 11399 599
rect 11271 531 11341 565
rect 11375 531 11399 565
rect 11271 497 11399 531
rect 7233 429 7371 463
rect 7233 395 7267 429
rect 7301 395 7371 429
rect 7233 361 7371 395
rect 7233 327 7267 361
rect 7301 327 7371 361
rect 7233 324 7371 327
rect 11271 463 11341 497
rect 11375 463 11399 497
rect 11271 429 11399 463
rect 11271 395 11341 429
rect 11375 395 11399 429
rect 11271 361 11399 395
rect 11271 327 11341 361
rect 11375 327 11399 361
rect 11271 324 11399 327
rect 7233 254 11399 324
rect 7233 220 7343 254
rect 7377 220 7411 254
rect 7445 220 7479 254
rect 7513 220 7547 254
rect 7581 220 7615 254
rect 7649 220 7683 254
rect 7717 220 7751 254
rect 7785 220 7819 254
rect 7853 220 7887 254
rect 7921 220 7955 254
rect 7989 220 8023 254
rect 8057 220 8091 254
rect 8125 220 8159 254
rect 8193 220 8227 254
rect 8261 220 8295 254
rect 8329 220 8363 254
rect 8397 220 8431 254
rect 8465 220 8499 254
rect 8533 220 8567 254
rect 8601 220 8635 254
rect 8669 220 8703 254
rect 8737 220 8771 254
rect 8805 220 8839 254
rect 8873 220 8907 254
rect 8941 220 8975 254
rect 9009 220 9043 254
rect 9077 220 9111 254
rect 9145 220 9179 254
rect 9213 220 9247 254
rect 9281 220 9315 254
rect 9349 220 9383 254
rect 9417 220 9451 254
rect 9485 220 9519 254
rect 9553 220 9587 254
rect 9621 220 9655 254
rect 9689 220 9723 254
rect 9757 220 9791 254
rect 9825 220 9859 254
rect 9893 220 9927 254
rect 9961 220 9995 254
rect 10029 220 10063 254
rect 10097 220 10131 254
rect 10165 220 10199 254
rect 10233 220 10267 254
rect 10301 220 10335 254
rect 10369 220 10403 254
rect 10437 220 10471 254
rect 10505 220 10539 254
rect 10573 220 10607 254
rect 10641 220 10675 254
rect 10709 220 10743 254
rect 10777 220 10811 254
rect 10845 220 10879 254
rect 10913 220 10947 254
rect 10981 220 11015 254
rect 11049 220 11083 254
rect 11117 220 11151 254
rect 11185 220 11219 254
rect 11253 220 11399 254
rect 7233 196 11399 220
<< mvnsubdiff >>
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
<< mvpsubdiffcont >>
rect 7353 3698 7387 3732
rect 7421 3698 7455 3732
rect 7489 3698 7523 3732
rect 7557 3698 7591 3732
rect 7625 3698 7659 3732
rect 7693 3698 7727 3732
rect 7761 3698 7795 3732
rect 7829 3698 7863 3732
rect 7897 3698 7931 3732
rect 7965 3698 7999 3732
rect 8033 3698 8067 3732
rect 8101 3698 8135 3732
rect 8169 3698 8203 3732
rect 8237 3698 8271 3732
rect 8305 3698 8339 3732
rect 8373 3698 8407 3732
rect 8441 3698 8475 3732
rect 8509 3698 8543 3732
rect 8577 3698 8611 3732
rect 8645 3698 8679 3732
rect 8713 3698 8747 3732
rect 8781 3698 8815 3732
rect 8849 3698 8883 3732
rect 8917 3698 8951 3732
rect 8985 3698 9019 3732
rect 9053 3698 9087 3732
rect 9121 3698 9155 3732
rect 9189 3698 9223 3732
rect 9257 3698 9291 3732
rect 9325 3698 9359 3732
rect 9393 3698 9427 3732
rect 9461 3698 9495 3732
rect 9529 3698 9563 3732
rect 9597 3698 9631 3732
rect 9665 3698 9699 3732
rect 9733 3698 9767 3732
rect 9801 3698 9835 3732
rect 9869 3698 9903 3732
rect 9937 3698 9971 3732
rect 10005 3698 10039 3732
rect 10073 3698 10107 3732
rect 10141 3698 10175 3732
rect 10209 3698 10243 3732
rect 10277 3698 10311 3732
rect 10345 3698 10379 3732
rect 10413 3698 10447 3732
rect 10481 3698 10515 3732
rect 10549 3698 10583 3732
rect 10617 3698 10651 3732
rect 10685 3698 10719 3732
rect 10753 3698 10787 3732
rect 10821 3698 10855 3732
rect 10889 3698 10923 3732
rect 10957 3698 10991 3732
rect 11025 3698 11059 3732
rect 11093 3698 11127 3732
rect 11161 3698 11195 3732
rect 11229 3698 11263 3732
rect 7267 3591 7301 3625
rect 7267 3523 7301 3557
rect 7267 3455 7301 3489
rect 11341 3591 11375 3625
rect 11341 3523 11375 3557
rect 7267 3387 7301 3421
rect 7267 3319 7301 3353
rect 7267 3251 7301 3285
rect 7267 3183 7301 3217
rect 7267 3115 7301 3149
rect 7267 3047 7301 3081
rect 7267 2979 7301 3013
rect 7267 2911 7301 2945
rect 7267 2843 7301 2877
rect 7267 2775 7301 2809
rect 7267 2707 7301 2741
rect 7267 2639 7301 2673
rect 7267 2571 7301 2605
rect 7267 2503 7301 2537
rect 7267 2435 7301 2469
rect 7267 2367 7301 2401
rect 7267 2299 7301 2333
rect 7267 2231 7301 2265
rect 7267 2163 7301 2197
rect 7267 2095 7301 2129
rect 7267 2027 7301 2061
rect 7267 1959 7301 1993
rect 7267 1891 7301 1925
rect 7267 1823 7301 1857
rect 7267 1755 7301 1789
rect 7267 1687 7301 1721
rect 7267 1619 7301 1653
rect 7267 1551 7301 1585
rect 7267 1483 7301 1517
rect 7267 1415 7301 1449
rect 7267 1347 7301 1381
rect 7267 1279 7301 1313
rect 7267 1211 7301 1245
rect 7267 1143 7301 1177
rect 7267 1075 7301 1109
rect 7267 1007 7301 1041
rect 7267 939 7301 973
rect 7267 871 7301 905
rect 7267 803 7301 837
rect 7267 735 7301 769
rect 7267 667 7301 701
rect 7267 599 7301 633
rect 7267 531 7301 565
rect 7267 463 7301 497
rect 11341 3455 11375 3489
rect 11341 3387 11375 3421
rect 11341 3319 11375 3353
rect 11341 3251 11375 3285
rect 11341 3183 11375 3217
rect 11341 3115 11375 3149
rect 11341 3047 11375 3081
rect 11341 2979 11375 3013
rect 11341 2911 11375 2945
rect 11341 2843 11375 2877
rect 11341 2775 11375 2809
rect 11341 2707 11375 2741
rect 11341 2639 11375 2673
rect 11341 2571 11375 2605
rect 11341 2503 11375 2537
rect 11341 2435 11375 2469
rect 11341 2367 11375 2401
rect 11341 2299 11375 2333
rect 11341 2231 11375 2265
rect 11341 2163 11375 2197
rect 11341 2095 11375 2129
rect 11341 2027 11375 2061
rect 11341 1959 11375 1993
rect 11341 1891 11375 1925
rect 11341 1823 11375 1857
rect 11341 1755 11375 1789
rect 11341 1687 11375 1721
rect 11341 1619 11375 1653
rect 11341 1551 11375 1585
rect 11341 1483 11375 1517
rect 11341 1415 11375 1449
rect 11341 1347 11375 1381
rect 11341 1279 11375 1313
rect 11341 1211 11375 1245
rect 11341 1143 11375 1177
rect 11341 1075 11375 1109
rect 11341 1007 11375 1041
rect 11341 939 11375 973
rect 11341 871 11375 905
rect 11341 803 11375 837
rect 11341 735 11375 769
rect 11341 667 11375 701
rect 11341 599 11375 633
rect 11341 531 11375 565
rect 7267 395 7301 429
rect 7267 327 7301 361
rect 11341 463 11375 497
rect 11341 395 11375 429
rect 11341 327 11375 361
rect 7343 220 7377 254
rect 7411 220 7445 254
rect 7479 220 7513 254
rect 7547 220 7581 254
rect 7615 220 7649 254
rect 7683 220 7717 254
rect 7751 220 7785 254
rect 7819 220 7853 254
rect 7887 220 7921 254
rect 7955 220 7989 254
rect 8023 220 8057 254
rect 8091 220 8125 254
rect 8159 220 8193 254
rect 8227 220 8261 254
rect 8295 220 8329 254
rect 8363 220 8397 254
rect 8431 220 8465 254
rect 8499 220 8533 254
rect 8567 220 8601 254
rect 8635 220 8669 254
rect 8703 220 8737 254
rect 8771 220 8805 254
rect 8839 220 8873 254
rect 8907 220 8941 254
rect 8975 220 9009 254
rect 9043 220 9077 254
rect 9111 220 9145 254
rect 9179 220 9213 254
rect 9247 220 9281 254
rect 9315 220 9349 254
rect 9383 220 9417 254
rect 9451 220 9485 254
rect 9519 220 9553 254
rect 9587 220 9621 254
rect 9655 220 9689 254
rect 9723 220 9757 254
rect 9791 220 9825 254
rect 9859 220 9893 254
rect 9927 220 9961 254
rect 9995 220 10029 254
rect 10063 220 10097 254
rect 10131 220 10165 254
rect 10199 220 10233 254
rect 10267 220 10301 254
rect 10335 220 10369 254
rect 10403 220 10437 254
rect 10471 220 10505 254
rect 10539 220 10573 254
rect 10607 220 10641 254
rect 10675 220 10709 254
rect 10743 220 10777 254
rect 10811 220 10845 254
rect 10879 220 10913 254
rect 10947 220 10981 254
rect 11015 220 11049 254
rect 11083 220 11117 254
rect 11151 220 11185 254
rect 11219 220 11253 254
<< mvnsubdiffcont >>
rect 7554 531 7792 3421
rect 8378 531 8616 3421
rect 9202 531 9440 3421
rect 10026 531 10264 3421
rect 10850 531 11088 3421
<< mvpdiode >>
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
<< mvpdiodec >>
rect 7966 531 8204 3421
rect 8790 531 9028 3421
rect 9614 531 9852 3421
rect 10438 531 10676 3421
<< locali >>
rect 7233 3750 11399 3756
rect 7233 3716 7342 3750
rect 7376 3732 7501 3750
rect 7535 3732 7574 3750
rect 7608 3732 7646 3750
rect 7680 3732 7718 3750
rect 7752 3732 7790 3750
rect 7824 3732 7862 3750
rect 7896 3732 7934 3750
rect 7968 3732 8006 3750
rect 8040 3732 8078 3750
rect 8112 3732 8150 3750
rect 8184 3732 8222 3750
rect 8256 3732 8294 3750
rect 8328 3732 8366 3750
rect 8400 3732 8438 3750
rect 8472 3732 8510 3750
rect 8544 3732 8582 3750
rect 8616 3732 8654 3750
rect 8688 3732 8726 3750
rect 8760 3732 8798 3750
rect 8832 3732 8870 3750
rect 8904 3732 8942 3750
rect 8976 3732 9014 3750
rect 9048 3732 9086 3750
rect 9120 3732 9158 3750
rect 9192 3732 9230 3750
rect 9264 3732 9302 3750
rect 9336 3732 9374 3750
rect 9408 3732 9446 3750
rect 9480 3732 9518 3750
rect 9552 3732 9590 3750
rect 9624 3732 9662 3750
rect 9696 3732 9734 3750
rect 9768 3732 9806 3750
rect 9840 3732 9878 3750
rect 9912 3732 9950 3750
rect 9984 3732 10022 3750
rect 10056 3732 10094 3750
rect 10128 3732 10166 3750
rect 10200 3732 10238 3750
rect 10272 3732 10310 3750
rect 10344 3732 10382 3750
rect 10416 3732 10454 3750
rect 10488 3732 10526 3750
rect 10560 3732 10598 3750
rect 10632 3732 10670 3750
rect 10704 3732 10742 3750
rect 10776 3732 10814 3750
rect 10848 3732 10886 3750
rect 10920 3732 10958 3750
rect 10992 3732 11030 3750
rect 11064 3732 11102 3750
rect 11136 3732 11260 3750
rect 7233 3698 7353 3716
rect 7387 3698 7421 3732
rect 7455 3698 7489 3732
rect 7535 3716 7557 3732
rect 7608 3716 7625 3732
rect 7680 3716 7693 3732
rect 7752 3716 7761 3732
rect 7824 3716 7829 3732
rect 7896 3716 7897 3732
rect 7523 3698 7557 3716
rect 7591 3698 7625 3716
rect 7659 3698 7693 3716
rect 7727 3698 7761 3716
rect 7795 3698 7829 3716
rect 7863 3698 7897 3716
rect 7931 3716 7934 3732
rect 7999 3716 8006 3732
rect 8067 3716 8078 3732
rect 8135 3716 8150 3732
rect 8203 3716 8222 3732
rect 8271 3716 8294 3732
rect 8339 3716 8366 3732
rect 8407 3716 8438 3732
rect 7931 3698 7965 3716
rect 7999 3698 8033 3716
rect 8067 3698 8101 3716
rect 8135 3698 8169 3716
rect 8203 3698 8237 3716
rect 8271 3698 8305 3716
rect 8339 3698 8373 3716
rect 8407 3698 8441 3716
rect 8475 3698 8509 3732
rect 8544 3716 8577 3732
rect 8616 3716 8645 3732
rect 8688 3716 8713 3732
rect 8760 3716 8781 3732
rect 8832 3716 8849 3732
rect 8904 3716 8917 3732
rect 8976 3716 8985 3732
rect 9048 3716 9053 3732
rect 9120 3716 9121 3732
rect 8543 3698 8577 3716
rect 8611 3698 8645 3716
rect 8679 3698 8713 3716
rect 8747 3698 8781 3716
rect 8815 3698 8849 3716
rect 8883 3698 8917 3716
rect 8951 3698 8985 3716
rect 9019 3698 9053 3716
rect 9087 3698 9121 3716
rect 9155 3716 9158 3732
rect 9223 3716 9230 3732
rect 9291 3716 9302 3732
rect 9359 3716 9374 3732
rect 9427 3716 9446 3732
rect 9495 3716 9518 3732
rect 9563 3716 9590 3732
rect 9631 3716 9662 3732
rect 9155 3698 9189 3716
rect 9223 3698 9257 3716
rect 9291 3698 9325 3716
rect 9359 3698 9393 3716
rect 9427 3698 9461 3716
rect 9495 3698 9529 3716
rect 9563 3698 9597 3716
rect 9631 3698 9665 3716
rect 9699 3698 9733 3732
rect 9768 3716 9801 3732
rect 9840 3716 9869 3732
rect 9912 3716 9937 3732
rect 9984 3716 10005 3732
rect 10056 3716 10073 3732
rect 10128 3716 10141 3732
rect 10200 3716 10209 3732
rect 10272 3716 10277 3732
rect 10344 3716 10345 3732
rect 9767 3698 9801 3716
rect 9835 3698 9869 3716
rect 9903 3698 9937 3716
rect 9971 3698 10005 3716
rect 10039 3698 10073 3716
rect 10107 3698 10141 3716
rect 10175 3698 10209 3716
rect 10243 3698 10277 3716
rect 10311 3698 10345 3716
rect 10379 3716 10382 3732
rect 10447 3716 10454 3732
rect 10515 3716 10526 3732
rect 10583 3716 10598 3732
rect 10651 3716 10670 3732
rect 10719 3716 10742 3732
rect 10787 3716 10814 3732
rect 10855 3716 10886 3732
rect 10379 3698 10413 3716
rect 10447 3698 10481 3716
rect 10515 3698 10549 3716
rect 10583 3698 10617 3716
rect 10651 3698 10685 3716
rect 10719 3698 10753 3716
rect 10787 3698 10821 3716
rect 10855 3698 10889 3716
rect 10923 3698 10957 3732
rect 10992 3716 11025 3732
rect 11064 3716 11093 3732
rect 11136 3716 11161 3732
rect 10991 3698 11025 3716
rect 11059 3698 11093 3716
rect 11127 3698 11161 3716
rect 11195 3698 11229 3732
rect 11294 3716 11399 3750
rect 11263 3698 11399 3716
rect 7233 3642 11399 3698
rect 7233 3625 7342 3642
rect 7233 3622 7267 3625
rect 7233 3588 7264 3622
rect 7301 3608 7342 3625
rect 7376 3608 7501 3642
rect 7535 3608 7574 3642
rect 7608 3608 7646 3642
rect 7680 3608 7718 3642
rect 7752 3608 7790 3642
rect 7824 3608 7862 3642
rect 7896 3608 7934 3642
rect 7968 3608 8006 3642
rect 8040 3608 8078 3642
rect 8112 3608 8150 3642
rect 8184 3608 8222 3642
rect 8256 3608 8294 3642
rect 8328 3608 8366 3642
rect 8400 3608 8438 3642
rect 8472 3608 8510 3642
rect 8544 3608 8582 3642
rect 8616 3608 8654 3642
rect 8688 3608 8726 3642
rect 8760 3608 8798 3642
rect 8832 3608 8870 3642
rect 8904 3608 8942 3642
rect 8976 3608 9014 3642
rect 9048 3608 9086 3642
rect 9120 3608 9158 3642
rect 9192 3608 9230 3642
rect 9264 3608 9302 3642
rect 9336 3608 9374 3642
rect 9408 3608 9446 3642
rect 9480 3608 9518 3642
rect 9552 3608 9590 3642
rect 9624 3608 9662 3642
rect 9696 3608 9734 3642
rect 9768 3608 9806 3642
rect 9840 3608 9878 3642
rect 9912 3608 9950 3642
rect 9984 3608 10022 3642
rect 10056 3608 10094 3642
rect 10128 3608 10166 3642
rect 10200 3608 10238 3642
rect 10272 3608 10310 3642
rect 10344 3608 10382 3642
rect 10416 3608 10454 3642
rect 10488 3608 10526 3642
rect 10560 3608 10598 3642
rect 10632 3608 10670 3642
rect 10704 3608 10742 3642
rect 10776 3608 10814 3642
rect 10848 3608 10886 3642
rect 10920 3608 10958 3642
rect 10992 3608 11030 3642
rect 11064 3608 11102 3642
rect 11136 3608 11260 3642
rect 11294 3625 11399 3642
rect 11294 3622 11341 3625
rect 11294 3608 11338 3622
rect 7301 3602 11338 3608
rect 7301 3591 7325 3602
rect 7298 3588 7325 3591
rect 7233 3557 7325 3588
rect 7233 3523 7267 3557
rect 7301 3523 7325 3557
rect 7233 3489 7325 3523
rect 7233 3464 7267 3489
rect 7233 3430 7264 3464
rect 7301 3455 7325 3489
rect 11317 3588 11338 3602
rect 11375 3591 11399 3625
rect 11372 3588 11399 3591
rect 11317 3557 11399 3588
rect 11317 3523 11341 3557
rect 11375 3523 11399 3557
rect 11317 3489 11399 3523
rect 7298 3430 7325 3455
rect 7233 3421 7325 3430
rect 7233 3392 7267 3421
rect 7233 3358 7264 3392
rect 7301 3387 7325 3421
rect 7298 3358 7325 3387
rect 7233 3353 7325 3358
rect 7233 3320 7267 3353
rect 7233 3286 7264 3320
rect 7301 3319 7325 3353
rect 7298 3286 7325 3319
rect 7233 3285 7325 3286
rect 7233 3251 7267 3285
rect 7301 3251 7325 3285
rect 7233 3248 7325 3251
rect 7233 3214 7264 3248
rect 7298 3217 7325 3248
rect 7233 3183 7267 3214
rect 7301 3183 7325 3217
rect 7233 3176 7325 3183
rect 7233 3142 7264 3176
rect 7298 3149 7325 3176
rect 7233 3115 7267 3142
rect 7301 3115 7325 3149
rect 7233 3104 7325 3115
rect 7233 3070 7264 3104
rect 7298 3081 7325 3104
rect 7233 3047 7267 3070
rect 7301 3047 7325 3081
rect 7233 3032 7325 3047
rect 7233 2998 7264 3032
rect 7298 3013 7325 3032
rect 7233 2979 7267 2998
rect 7301 2979 7325 3013
rect 7233 2960 7325 2979
rect 7233 2926 7264 2960
rect 7298 2945 7325 2960
rect 7233 2911 7267 2926
rect 7301 2911 7325 2945
rect 7233 2888 7325 2911
rect 7233 2854 7264 2888
rect 7298 2877 7325 2888
rect 7233 2843 7267 2854
rect 7301 2843 7325 2877
rect 7233 2816 7325 2843
rect 7233 2782 7264 2816
rect 7298 2809 7325 2816
rect 7233 2775 7267 2782
rect 7301 2775 7325 2809
rect 7233 2744 7325 2775
rect 7233 2710 7264 2744
rect 7298 2741 7325 2744
rect 7233 2707 7267 2710
rect 7301 2707 7325 2741
rect 7233 2673 7325 2707
rect 7233 2672 7267 2673
rect 7233 2638 7264 2672
rect 7301 2639 7325 2673
rect 7298 2638 7325 2639
rect 7233 2605 7325 2638
rect 7233 2600 7267 2605
rect 7233 2566 7264 2600
rect 7301 2571 7325 2605
rect 7298 2566 7325 2571
rect 7233 2537 7325 2566
rect 7233 2528 7267 2537
rect 7233 2494 7264 2528
rect 7301 2503 7325 2537
rect 7298 2494 7325 2503
rect 7233 2469 7325 2494
rect 7233 2456 7267 2469
rect 7233 2422 7264 2456
rect 7301 2435 7325 2469
rect 7298 2422 7325 2435
rect 7233 2401 7325 2422
rect 7233 2384 7267 2401
rect 7233 2350 7264 2384
rect 7301 2367 7325 2401
rect 7298 2350 7325 2367
rect 7233 2333 7325 2350
rect 7233 2312 7267 2333
rect 7233 2278 7264 2312
rect 7301 2299 7325 2333
rect 7298 2278 7325 2299
rect 7233 2265 7325 2278
rect 7233 2240 7267 2265
rect 7233 2206 7264 2240
rect 7301 2231 7325 2265
rect 7298 2206 7325 2231
rect 7233 2197 7325 2206
rect 7233 2168 7267 2197
rect 7233 2134 7264 2168
rect 7301 2163 7325 2197
rect 7298 2134 7325 2163
rect 7233 2129 7325 2134
rect 7233 2096 7267 2129
rect 7233 2062 7264 2096
rect 7301 2095 7325 2129
rect 7298 2062 7325 2095
rect 7233 2061 7325 2062
rect 7233 2027 7267 2061
rect 7301 2027 7325 2061
rect 7233 2024 7325 2027
rect 7233 1990 7264 2024
rect 7298 1993 7325 2024
rect 7233 1959 7267 1990
rect 7301 1959 7325 1993
rect 7233 1952 7325 1959
rect 7233 1918 7264 1952
rect 7298 1925 7325 1952
rect 7233 1891 7267 1918
rect 7301 1891 7325 1925
rect 7233 1880 7325 1891
rect 7233 1846 7264 1880
rect 7298 1857 7325 1880
rect 7233 1823 7267 1846
rect 7301 1823 7325 1857
rect 7233 1808 7325 1823
rect 7233 1774 7264 1808
rect 7298 1789 7325 1808
rect 7233 1755 7267 1774
rect 7301 1755 7325 1789
rect 7233 1736 7325 1755
rect 7233 1702 7264 1736
rect 7298 1721 7325 1736
rect 7233 1687 7267 1702
rect 7301 1687 7325 1721
rect 7233 1664 7325 1687
rect 7233 1630 7264 1664
rect 7298 1653 7325 1664
rect 7233 1619 7267 1630
rect 7301 1619 7325 1653
rect 7233 1592 7325 1619
rect 7233 1558 7264 1592
rect 7298 1585 7325 1592
rect 7233 1551 7267 1558
rect 7301 1551 7325 1585
rect 7233 1520 7325 1551
rect 7233 1486 7264 1520
rect 7298 1517 7325 1520
rect 7233 1483 7267 1486
rect 7301 1483 7325 1517
rect 7233 1449 7325 1483
rect 7233 1448 7267 1449
rect 7233 1414 7264 1448
rect 7301 1415 7325 1449
rect 7298 1414 7325 1415
rect 7233 1381 7325 1414
rect 7233 1376 7267 1381
rect 7233 1342 7264 1376
rect 7301 1347 7325 1381
rect 7298 1342 7325 1347
rect 7233 1313 7325 1342
rect 7233 1304 7267 1313
rect 7233 1270 7264 1304
rect 7301 1279 7325 1313
rect 7298 1270 7325 1279
rect 7233 1245 7325 1270
rect 7233 1232 7267 1245
rect 7233 1198 7264 1232
rect 7301 1211 7325 1245
rect 7298 1198 7325 1211
rect 7233 1177 7325 1198
rect 7233 1160 7267 1177
rect 7233 1126 7264 1160
rect 7301 1143 7325 1177
rect 7298 1126 7325 1143
rect 7233 1109 7325 1126
rect 7233 1088 7267 1109
rect 7233 1054 7264 1088
rect 7301 1075 7325 1109
rect 7298 1054 7325 1075
rect 7233 1041 7325 1054
rect 7233 1016 7267 1041
rect 7233 982 7264 1016
rect 7301 1007 7325 1041
rect 7298 982 7325 1007
rect 7233 973 7325 982
rect 7233 944 7267 973
rect 7233 910 7264 944
rect 7301 939 7325 973
rect 7298 910 7325 939
rect 7233 905 7325 910
rect 7233 872 7267 905
rect 7233 838 7264 872
rect 7301 871 7325 905
rect 7298 838 7325 871
rect 7233 837 7325 838
rect 7233 803 7267 837
rect 7301 803 7325 837
rect 7233 800 7325 803
rect 7233 766 7264 800
rect 7298 769 7325 800
rect 7233 735 7267 766
rect 7301 735 7325 769
rect 7233 728 7325 735
rect 7233 694 7264 728
rect 7298 701 7325 728
rect 7233 667 7267 694
rect 7301 667 7325 701
rect 7233 656 7325 667
rect 7233 622 7264 656
rect 7298 633 7325 656
rect 7233 599 7267 622
rect 7301 599 7325 633
rect 7233 565 7325 599
rect 7233 531 7267 565
rect 7301 531 7325 565
rect 7233 497 7325 531
rect 7233 463 7267 497
rect 7301 463 7325 497
rect 7523 3421 7823 3476
rect 7523 531 7554 3421
rect 7792 531 7823 3421
rect 7523 476 7823 531
rect 7935 3421 8235 3476
rect 7935 531 7966 3421
rect 8204 531 8235 3421
rect 7935 476 8235 531
rect 8347 3421 8647 3476
rect 8347 531 8378 3421
rect 8616 531 8647 3421
rect 8347 476 8647 531
rect 8759 3421 9059 3476
rect 8759 531 8790 3421
rect 9028 531 9059 3421
rect 8759 476 9059 531
rect 9171 3421 9471 3476
rect 9171 531 9202 3421
rect 9440 531 9471 3421
rect 9171 476 9471 531
rect 9583 3421 9883 3476
rect 9583 531 9614 3421
rect 9852 531 9883 3421
rect 9583 476 9883 531
rect 9995 3421 10295 3476
rect 9995 531 10026 3421
rect 10264 531 10295 3421
rect 9995 476 10295 531
rect 10407 3421 10707 3476
rect 10407 531 10438 3421
rect 10676 531 10707 3421
rect 10407 476 10707 531
rect 10819 3421 11119 3476
rect 10819 531 10850 3421
rect 11088 531 11119 3421
rect 10819 476 11119 531
rect 11317 3464 11341 3489
rect 11317 3430 11338 3464
rect 11375 3455 11399 3489
rect 11372 3430 11399 3455
rect 11317 3421 11399 3430
rect 11317 3392 11341 3421
rect 11317 3358 11338 3392
rect 11375 3387 11399 3421
rect 11372 3358 11399 3387
rect 11317 3353 11399 3358
rect 11317 3320 11341 3353
rect 11317 3286 11338 3320
rect 11375 3319 11399 3353
rect 11372 3286 11399 3319
rect 11317 3285 11399 3286
rect 11317 3251 11341 3285
rect 11375 3251 11399 3285
rect 11317 3248 11399 3251
rect 11317 3214 11338 3248
rect 11372 3217 11399 3248
rect 11317 3183 11341 3214
rect 11375 3183 11399 3217
rect 11317 3176 11399 3183
rect 11317 3142 11338 3176
rect 11372 3149 11399 3176
rect 11317 3115 11341 3142
rect 11375 3115 11399 3149
rect 11317 3104 11399 3115
rect 11317 3070 11338 3104
rect 11372 3081 11399 3104
rect 11317 3047 11341 3070
rect 11375 3047 11399 3081
rect 11317 3032 11399 3047
rect 11317 2998 11338 3032
rect 11372 3013 11399 3032
rect 11317 2979 11341 2998
rect 11375 2979 11399 3013
rect 11317 2960 11399 2979
rect 11317 2926 11338 2960
rect 11372 2945 11399 2960
rect 11317 2911 11341 2926
rect 11375 2911 11399 2945
rect 11317 2888 11399 2911
rect 11317 2854 11338 2888
rect 11372 2877 11399 2888
rect 11317 2843 11341 2854
rect 11375 2843 11399 2877
rect 11317 2816 11399 2843
rect 11317 2782 11338 2816
rect 11372 2809 11399 2816
rect 11317 2775 11341 2782
rect 11375 2775 11399 2809
rect 11317 2744 11399 2775
rect 11317 2710 11338 2744
rect 11372 2741 11399 2744
rect 11317 2707 11341 2710
rect 11375 2707 11399 2741
rect 11317 2673 11399 2707
rect 11317 2672 11341 2673
rect 11317 2638 11338 2672
rect 11375 2639 11399 2673
rect 11372 2638 11399 2639
rect 11317 2605 11399 2638
rect 11317 2600 11341 2605
rect 11317 2566 11338 2600
rect 11375 2571 11399 2605
rect 11372 2566 11399 2571
rect 11317 2537 11399 2566
rect 11317 2528 11341 2537
rect 11317 2494 11338 2528
rect 11375 2503 11399 2537
rect 11372 2494 11399 2503
rect 11317 2469 11399 2494
rect 11317 2456 11341 2469
rect 11317 2422 11338 2456
rect 11375 2435 11399 2469
rect 11372 2422 11399 2435
rect 11317 2401 11399 2422
rect 11317 2384 11341 2401
rect 11317 2350 11338 2384
rect 11375 2367 11399 2401
rect 11372 2350 11399 2367
rect 11317 2333 11399 2350
rect 11317 2312 11341 2333
rect 11317 2278 11338 2312
rect 11375 2299 11399 2333
rect 11372 2278 11399 2299
rect 11317 2265 11399 2278
rect 11317 2240 11341 2265
rect 11317 2206 11338 2240
rect 11375 2231 11399 2265
rect 11372 2206 11399 2231
rect 11317 2197 11399 2206
rect 11317 2168 11341 2197
rect 11317 2134 11338 2168
rect 11375 2163 11399 2197
rect 11372 2134 11399 2163
rect 11317 2129 11399 2134
rect 11317 2096 11341 2129
rect 11317 2062 11338 2096
rect 11375 2095 11399 2129
rect 11372 2062 11399 2095
rect 11317 2061 11399 2062
rect 11317 2027 11341 2061
rect 11375 2027 11399 2061
rect 11317 2024 11399 2027
rect 11317 1990 11338 2024
rect 11372 1993 11399 2024
rect 11317 1959 11341 1990
rect 11375 1959 11399 1993
rect 11317 1952 11399 1959
rect 11317 1918 11338 1952
rect 11372 1925 11399 1952
rect 11317 1891 11341 1918
rect 11375 1891 11399 1925
rect 11317 1880 11399 1891
rect 11317 1846 11338 1880
rect 11372 1857 11399 1880
rect 11317 1823 11341 1846
rect 11375 1823 11399 1857
rect 11317 1808 11399 1823
rect 11317 1774 11338 1808
rect 11372 1789 11399 1808
rect 11317 1755 11341 1774
rect 11375 1755 11399 1789
rect 11317 1736 11399 1755
rect 11317 1702 11338 1736
rect 11372 1721 11399 1736
rect 11317 1687 11341 1702
rect 11375 1687 11399 1721
rect 11317 1664 11399 1687
rect 11317 1630 11338 1664
rect 11372 1653 11399 1664
rect 11317 1619 11341 1630
rect 11375 1619 11399 1653
rect 11317 1592 11399 1619
rect 11317 1558 11338 1592
rect 11372 1585 11399 1592
rect 11317 1551 11341 1558
rect 11375 1551 11399 1585
rect 11317 1520 11399 1551
rect 11317 1486 11338 1520
rect 11372 1517 11399 1520
rect 11317 1483 11341 1486
rect 11375 1483 11399 1517
rect 11317 1449 11399 1483
rect 11317 1448 11341 1449
rect 11317 1414 11338 1448
rect 11375 1415 11399 1449
rect 11372 1414 11399 1415
rect 11317 1381 11399 1414
rect 11317 1376 11341 1381
rect 11317 1342 11338 1376
rect 11375 1347 11399 1381
rect 11372 1342 11399 1347
rect 11317 1313 11399 1342
rect 11317 1304 11341 1313
rect 11317 1270 11338 1304
rect 11375 1279 11399 1313
rect 11372 1270 11399 1279
rect 11317 1245 11399 1270
rect 11317 1232 11341 1245
rect 11317 1198 11338 1232
rect 11375 1211 11399 1245
rect 11372 1198 11399 1211
rect 11317 1177 11399 1198
rect 11317 1160 11341 1177
rect 11317 1126 11338 1160
rect 11375 1143 11399 1177
rect 11372 1126 11399 1143
rect 11317 1109 11399 1126
rect 11317 1088 11341 1109
rect 11317 1054 11338 1088
rect 11375 1075 11399 1109
rect 11372 1054 11399 1075
rect 11317 1041 11399 1054
rect 11317 1016 11341 1041
rect 11317 982 11338 1016
rect 11375 1007 11399 1041
rect 11372 982 11399 1007
rect 11317 973 11399 982
rect 11317 944 11341 973
rect 11317 910 11338 944
rect 11375 939 11399 973
rect 11372 910 11399 939
rect 11317 905 11399 910
rect 11317 872 11341 905
rect 11317 838 11338 872
rect 11375 871 11399 905
rect 11372 838 11399 871
rect 11317 837 11399 838
rect 11317 803 11341 837
rect 11375 803 11399 837
rect 11317 800 11399 803
rect 11317 766 11338 800
rect 11372 769 11399 800
rect 11317 735 11341 766
rect 11375 735 11399 769
rect 11317 728 11399 735
rect 11317 694 11338 728
rect 11372 701 11399 728
rect 11317 667 11341 694
rect 11375 667 11399 701
rect 11317 656 11399 667
rect 11317 622 11338 656
rect 11372 633 11399 656
rect 11317 599 11341 622
rect 11375 599 11399 633
rect 11317 565 11399 599
rect 11317 531 11341 565
rect 11375 531 11399 565
rect 11317 497 11399 531
rect 7233 429 7325 463
rect 7233 395 7267 429
rect 7301 395 7325 429
rect 7233 361 7325 395
rect 7233 327 7267 361
rect 7301 327 7325 361
rect 7233 278 7325 327
rect 11317 463 11341 497
rect 11375 463 11399 497
rect 11317 429 11399 463
rect 11317 395 11341 429
rect 11375 395 11399 429
rect 11317 361 11399 395
rect 11317 327 11341 361
rect 11375 327 11399 361
rect 11317 278 11399 327
rect 7233 254 11399 278
rect 7233 220 7343 254
rect 7377 220 7411 254
rect 7445 220 7479 254
rect 7513 220 7547 254
rect 7581 220 7615 254
rect 7649 220 7683 254
rect 7717 220 7751 254
rect 7785 220 7819 254
rect 7853 220 7887 254
rect 7921 220 7955 254
rect 7989 220 8023 254
rect 8057 220 8091 254
rect 8125 220 8159 254
rect 8193 220 8227 254
rect 8261 220 8295 254
rect 8329 220 8363 254
rect 8397 220 8431 254
rect 8465 220 8499 254
rect 8533 220 8567 254
rect 8601 220 8635 254
rect 8669 220 8703 254
rect 8737 220 8771 254
rect 8805 220 8839 254
rect 8873 220 8907 254
rect 8941 220 8975 254
rect 9009 220 9043 254
rect 9077 220 9111 254
rect 9145 220 9179 254
rect 9213 220 9247 254
rect 9281 220 9315 254
rect 9349 220 9383 254
rect 9417 220 9451 254
rect 9485 220 9519 254
rect 9553 220 9587 254
rect 9621 220 9655 254
rect 9689 220 9723 254
rect 9757 220 9791 254
rect 9825 220 9859 254
rect 9893 220 9927 254
rect 9961 220 9995 254
rect 10029 220 10063 254
rect 10097 220 10131 254
rect 10165 220 10199 254
rect 10233 220 10267 254
rect 10301 220 10335 254
rect 10369 220 10403 254
rect 10437 220 10471 254
rect 10505 220 10539 254
rect 10573 220 10607 254
rect 10641 220 10675 254
rect 10709 220 10743 254
rect 10777 220 10811 254
rect 10845 220 10879 254
rect 10913 220 10947 254
rect 10981 220 11015 254
rect 11049 220 11083 254
rect 11117 220 11151 254
rect 11185 220 11219 254
rect 11253 220 11399 254
rect 7233 196 11399 220
<< viali >>
rect 7342 3732 7376 3750
rect 7501 3732 7535 3750
rect 7574 3732 7608 3750
rect 7646 3732 7680 3750
rect 7718 3732 7752 3750
rect 7790 3732 7824 3750
rect 7862 3732 7896 3750
rect 7934 3732 7968 3750
rect 8006 3732 8040 3750
rect 8078 3732 8112 3750
rect 8150 3732 8184 3750
rect 8222 3732 8256 3750
rect 8294 3732 8328 3750
rect 8366 3732 8400 3750
rect 8438 3732 8472 3750
rect 8510 3732 8544 3750
rect 8582 3732 8616 3750
rect 8654 3732 8688 3750
rect 8726 3732 8760 3750
rect 8798 3732 8832 3750
rect 8870 3732 8904 3750
rect 8942 3732 8976 3750
rect 9014 3732 9048 3750
rect 9086 3732 9120 3750
rect 9158 3732 9192 3750
rect 9230 3732 9264 3750
rect 9302 3732 9336 3750
rect 9374 3732 9408 3750
rect 9446 3732 9480 3750
rect 9518 3732 9552 3750
rect 9590 3732 9624 3750
rect 9662 3732 9696 3750
rect 9734 3732 9768 3750
rect 9806 3732 9840 3750
rect 9878 3732 9912 3750
rect 9950 3732 9984 3750
rect 10022 3732 10056 3750
rect 10094 3732 10128 3750
rect 10166 3732 10200 3750
rect 10238 3732 10272 3750
rect 10310 3732 10344 3750
rect 10382 3732 10416 3750
rect 10454 3732 10488 3750
rect 10526 3732 10560 3750
rect 10598 3732 10632 3750
rect 10670 3732 10704 3750
rect 10742 3732 10776 3750
rect 10814 3732 10848 3750
rect 10886 3732 10920 3750
rect 10958 3732 10992 3750
rect 11030 3732 11064 3750
rect 11102 3732 11136 3750
rect 11260 3732 11294 3750
rect 7342 3716 7353 3732
rect 7353 3716 7376 3732
rect 7501 3716 7523 3732
rect 7523 3716 7535 3732
rect 7574 3716 7591 3732
rect 7591 3716 7608 3732
rect 7646 3716 7659 3732
rect 7659 3716 7680 3732
rect 7718 3716 7727 3732
rect 7727 3716 7752 3732
rect 7790 3716 7795 3732
rect 7795 3716 7824 3732
rect 7862 3716 7863 3732
rect 7863 3716 7896 3732
rect 7934 3716 7965 3732
rect 7965 3716 7968 3732
rect 8006 3716 8033 3732
rect 8033 3716 8040 3732
rect 8078 3716 8101 3732
rect 8101 3716 8112 3732
rect 8150 3716 8169 3732
rect 8169 3716 8184 3732
rect 8222 3716 8237 3732
rect 8237 3716 8256 3732
rect 8294 3716 8305 3732
rect 8305 3716 8328 3732
rect 8366 3716 8373 3732
rect 8373 3716 8400 3732
rect 8438 3716 8441 3732
rect 8441 3716 8472 3732
rect 8510 3716 8543 3732
rect 8543 3716 8544 3732
rect 8582 3716 8611 3732
rect 8611 3716 8616 3732
rect 8654 3716 8679 3732
rect 8679 3716 8688 3732
rect 8726 3716 8747 3732
rect 8747 3716 8760 3732
rect 8798 3716 8815 3732
rect 8815 3716 8832 3732
rect 8870 3716 8883 3732
rect 8883 3716 8904 3732
rect 8942 3716 8951 3732
rect 8951 3716 8976 3732
rect 9014 3716 9019 3732
rect 9019 3716 9048 3732
rect 9086 3716 9087 3732
rect 9087 3716 9120 3732
rect 9158 3716 9189 3732
rect 9189 3716 9192 3732
rect 9230 3716 9257 3732
rect 9257 3716 9264 3732
rect 9302 3716 9325 3732
rect 9325 3716 9336 3732
rect 9374 3716 9393 3732
rect 9393 3716 9408 3732
rect 9446 3716 9461 3732
rect 9461 3716 9480 3732
rect 9518 3716 9529 3732
rect 9529 3716 9552 3732
rect 9590 3716 9597 3732
rect 9597 3716 9624 3732
rect 9662 3716 9665 3732
rect 9665 3716 9696 3732
rect 9734 3716 9767 3732
rect 9767 3716 9768 3732
rect 9806 3716 9835 3732
rect 9835 3716 9840 3732
rect 9878 3716 9903 3732
rect 9903 3716 9912 3732
rect 9950 3716 9971 3732
rect 9971 3716 9984 3732
rect 10022 3716 10039 3732
rect 10039 3716 10056 3732
rect 10094 3716 10107 3732
rect 10107 3716 10128 3732
rect 10166 3716 10175 3732
rect 10175 3716 10200 3732
rect 10238 3716 10243 3732
rect 10243 3716 10272 3732
rect 10310 3716 10311 3732
rect 10311 3716 10344 3732
rect 10382 3716 10413 3732
rect 10413 3716 10416 3732
rect 10454 3716 10481 3732
rect 10481 3716 10488 3732
rect 10526 3716 10549 3732
rect 10549 3716 10560 3732
rect 10598 3716 10617 3732
rect 10617 3716 10632 3732
rect 10670 3716 10685 3732
rect 10685 3716 10704 3732
rect 10742 3716 10753 3732
rect 10753 3716 10776 3732
rect 10814 3716 10821 3732
rect 10821 3716 10848 3732
rect 10886 3716 10889 3732
rect 10889 3716 10920 3732
rect 10958 3716 10991 3732
rect 10991 3716 10992 3732
rect 11030 3716 11059 3732
rect 11059 3716 11064 3732
rect 11102 3716 11127 3732
rect 11127 3716 11136 3732
rect 11260 3716 11263 3732
rect 11263 3716 11294 3732
rect 7264 3591 7267 3622
rect 7267 3591 7298 3622
rect 7342 3608 7376 3642
rect 7501 3608 7535 3642
rect 7574 3608 7608 3642
rect 7646 3608 7680 3642
rect 7718 3608 7752 3642
rect 7790 3608 7824 3642
rect 7862 3608 7896 3642
rect 7934 3608 7968 3642
rect 8006 3608 8040 3642
rect 8078 3608 8112 3642
rect 8150 3608 8184 3642
rect 8222 3608 8256 3642
rect 8294 3608 8328 3642
rect 8366 3608 8400 3642
rect 8438 3608 8472 3642
rect 8510 3608 8544 3642
rect 8582 3608 8616 3642
rect 8654 3608 8688 3642
rect 8726 3608 8760 3642
rect 8798 3608 8832 3642
rect 8870 3608 8904 3642
rect 8942 3608 8976 3642
rect 9014 3608 9048 3642
rect 9086 3608 9120 3642
rect 9158 3608 9192 3642
rect 9230 3608 9264 3642
rect 9302 3608 9336 3642
rect 9374 3608 9408 3642
rect 9446 3608 9480 3642
rect 9518 3608 9552 3642
rect 9590 3608 9624 3642
rect 9662 3608 9696 3642
rect 9734 3608 9768 3642
rect 9806 3608 9840 3642
rect 9878 3608 9912 3642
rect 9950 3608 9984 3642
rect 10022 3608 10056 3642
rect 10094 3608 10128 3642
rect 10166 3608 10200 3642
rect 10238 3608 10272 3642
rect 10310 3608 10344 3642
rect 10382 3608 10416 3642
rect 10454 3608 10488 3642
rect 10526 3608 10560 3642
rect 10598 3608 10632 3642
rect 10670 3608 10704 3642
rect 10742 3608 10776 3642
rect 10814 3608 10848 3642
rect 10886 3608 10920 3642
rect 10958 3608 10992 3642
rect 11030 3608 11064 3642
rect 11102 3608 11136 3642
rect 11260 3608 11294 3642
rect 7264 3588 7298 3591
rect 7264 3455 7267 3464
rect 7267 3455 7298 3464
rect 11338 3591 11341 3622
rect 11341 3591 11372 3622
rect 11338 3588 11372 3591
rect 7264 3430 7298 3455
rect 7264 3387 7267 3392
rect 7267 3387 7298 3392
rect 7264 3358 7298 3387
rect 7264 3319 7267 3320
rect 7267 3319 7298 3320
rect 7264 3286 7298 3319
rect 7264 3217 7298 3248
rect 7264 3214 7267 3217
rect 7267 3214 7298 3217
rect 7264 3149 7298 3176
rect 7264 3142 7267 3149
rect 7267 3142 7298 3149
rect 7264 3081 7298 3104
rect 7264 3070 7267 3081
rect 7267 3070 7298 3081
rect 7264 3013 7298 3032
rect 7264 2998 7267 3013
rect 7267 2998 7298 3013
rect 7264 2945 7298 2960
rect 7264 2926 7267 2945
rect 7267 2926 7298 2945
rect 7264 2877 7298 2888
rect 7264 2854 7267 2877
rect 7267 2854 7298 2877
rect 7264 2809 7298 2816
rect 7264 2782 7267 2809
rect 7267 2782 7298 2809
rect 7264 2741 7298 2744
rect 7264 2710 7267 2741
rect 7267 2710 7298 2741
rect 7264 2639 7267 2672
rect 7267 2639 7298 2672
rect 7264 2638 7298 2639
rect 7264 2571 7267 2600
rect 7267 2571 7298 2600
rect 7264 2566 7298 2571
rect 7264 2503 7267 2528
rect 7267 2503 7298 2528
rect 7264 2494 7298 2503
rect 7264 2435 7267 2456
rect 7267 2435 7298 2456
rect 7264 2422 7298 2435
rect 7264 2367 7267 2384
rect 7267 2367 7298 2384
rect 7264 2350 7298 2367
rect 7264 2299 7267 2312
rect 7267 2299 7298 2312
rect 7264 2278 7298 2299
rect 7264 2231 7267 2240
rect 7267 2231 7298 2240
rect 7264 2206 7298 2231
rect 7264 2163 7267 2168
rect 7267 2163 7298 2168
rect 7264 2134 7298 2163
rect 7264 2095 7267 2096
rect 7267 2095 7298 2096
rect 7264 2062 7298 2095
rect 7264 1993 7298 2024
rect 7264 1990 7267 1993
rect 7267 1990 7298 1993
rect 7264 1925 7298 1952
rect 7264 1918 7267 1925
rect 7267 1918 7298 1925
rect 7264 1857 7298 1880
rect 7264 1846 7267 1857
rect 7267 1846 7298 1857
rect 7264 1789 7298 1808
rect 7264 1774 7267 1789
rect 7267 1774 7298 1789
rect 7264 1721 7298 1736
rect 7264 1702 7267 1721
rect 7267 1702 7298 1721
rect 7264 1653 7298 1664
rect 7264 1630 7267 1653
rect 7267 1630 7298 1653
rect 7264 1585 7298 1592
rect 7264 1558 7267 1585
rect 7267 1558 7298 1585
rect 7264 1517 7298 1520
rect 7264 1486 7267 1517
rect 7267 1486 7298 1517
rect 7264 1415 7267 1448
rect 7267 1415 7298 1448
rect 7264 1414 7298 1415
rect 7264 1347 7267 1376
rect 7267 1347 7298 1376
rect 7264 1342 7298 1347
rect 7264 1279 7267 1304
rect 7267 1279 7298 1304
rect 7264 1270 7298 1279
rect 7264 1211 7267 1232
rect 7267 1211 7298 1232
rect 7264 1198 7298 1211
rect 7264 1143 7267 1160
rect 7267 1143 7298 1160
rect 7264 1126 7298 1143
rect 7264 1075 7267 1088
rect 7267 1075 7298 1088
rect 7264 1054 7298 1075
rect 7264 1007 7267 1016
rect 7267 1007 7298 1016
rect 7264 982 7298 1007
rect 7264 939 7267 944
rect 7267 939 7298 944
rect 7264 910 7298 939
rect 7264 871 7267 872
rect 7267 871 7298 872
rect 7264 838 7298 871
rect 7264 769 7298 800
rect 7264 766 7267 769
rect 7267 766 7298 769
rect 7264 701 7298 728
rect 7264 694 7267 701
rect 7267 694 7298 701
rect 7264 633 7298 656
rect 7264 622 7267 633
rect 7267 622 7298 633
rect 7584 3303 7618 3337
rect 7656 3303 7690 3337
rect 7728 3303 7762 3337
rect 7584 3207 7618 3241
rect 7656 3207 7690 3241
rect 7728 3207 7762 3241
rect 7584 3111 7618 3145
rect 7656 3111 7690 3145
rect 7728 3111 7762 3145
rect 7584 3015 7618 3049
rect 7656 3015 7690 3049
rect 7728 3015 7762 3049
rect 7584 2919 7618 2953
rect 7656 2919 7690 2953
rect 7728 2919 7762 2953
rect 7584 2823 7618 2857
rect 7656 2823 7690 2857
rect 7728 2823 7762 2857
rect 7584 2727 7618 2761
rect 7656 2727 7690 2761
rect 7728 2727 7762 2761
rect 7584 2631 7618 2665
rect 7656 2631 7690 2665
rect 7728 2631 7762 2665
rect 7584 2535 7618 2569
rect 7656 2535 7690 2569
rect 7728 2535 7762 2569
rect 7584 2439 7618 2473
rect 7656 2439 7690 2473
rect 7728 2439 7762 2473
rect 7584 2343 7618 2377
rect 7656 2343 7690 2377
rect 7728 2343 7762 2377
rect 7584 2247 7618 2281
rect 7656 2247 7690 2281
rect 7728 2247 7762 2281
rect 7584 2151 7618 2185
rect 7656 2151 7690 2185
rect 7728 2151 7762 2185
rect 7584 2055 7618 2089
rect 7656 2055 7690 2089
rect 7728 2055 7762 2089
rect 7584 1959 7618 1993
rect 7656 1959 7690 1993
rect 7728 1959 7762 1993
rect 7584 1863 7618 1897
rect 7656 1863 7690 1897
rect 7728 1863 7762 1897
rect 7584 1767 7618 1801
rect 7656 1767 7690 1801
rect 7728 1767 7762 1801
rect 7584 1671 7618 1705
rect 7656 1671 7690 1705
rect 7728 1671 7762 1705
rect 7584 1575 7618 1609
rect 7656 1575 7690 1609
rect 7728 1575 7762 1609
rect 7584 1479 7618 1513
rect 7656 1479 7690 1513
rect 7728 1479 7762 1513
rect 7584 1383 7618 1417
rect 7656 1383 7690 1417
rect 7728 1383 7762 1417
rect 7584 1287 7618 1321
rect 7656 1287 7690 1321
rect 7728 1287 7762 1321
rect 7584 1191 7618 1225
rect 7656 1191 7690 1225
rect 7728 1191 7762 1225
rect 7584 1095 7618 1129
rect 7656 1095 7690 1129
rect 7728 1095 7762 1129
rect 7584 999 7618 1033
rect 7656 999 7690 1033
rect 7728 999 7762 1033
rect 7584 903 7618 937
rect 7656 903 7690 937
rect 7728 903 7762 937
rect 7584 807 7618 841
rect 7656 807 7690 841
rect 7728 807 7762 841
rect 7584 711 7618 745
rect 7656 711 7690 745
rect 7728 711 7762 745
rect 7584 615 7618 649
rect 7656 615 7690 649
rect 7728 615 7762 649
rect 7996 3303 8030 3337
rect 8068 3303 8102 3337
rect 8140 3303 8174 3337
rect 7996 3207 8030 3241
rect 8068 3207 8102 3241
rect 8140 3207 8174 3241
rect 7996 3111 8030 3145
rect 8068 3111 8102 3145
rect 8140 3111 8174 3145
rect 7996 3015 8030 3049
rect 8068 3015 8102 3049
rect 8140 3015 8174 3049
rect 7996 2919 8030 2953
rect 8068 2919 8102 2953
rect 8140 2919 8174 2953
rect 7996 2823 8030 2857
rect 8068 2823 8102 2857
rect 8140 2823 8174 2857
rect 7996 2727 8030 2761
rect 8068 2727 8102 2761
rect 8140 2727 8174 2761
rect 7996 2631 8030 2665
rect 8068 2631 8102 2665
rect 8140 2631 8174 2665
rect 7996 2535 8030 2569
rect 8068 2535 8102 2569
rect 8140 2535 8174 2569
rect 7996 2439 8030 2473
rect 8068 2439 8102 2473
rect 8140 2439 8174 2473
rect 7996 2343 8030 2377
rect 8068 2343 8102 2377
rect 8140 2343 8174 2377
rect 7996 2247 8030 2281
rect 8068 2247 8102 2281
rect 8140 2247 8174 2281
rect 7996 2151 8030 2185
rect 8068 2151 8102 2185
rect 8140 2151 8174 2185
rect 7996 2055 8030 2089
rect 8068 2055 8102 2089
rect 8140 2055 8174 2089
rect 7996 1959 8030 1993
rect 8068 1959 8102 1993
rect 8140 1959 8174 1993
rect 7996 1863 8030 1897
rect 8068 1863 8102 1897
rect 8140 1863 8174 1897
rect 7996 1767 8030 1801
rect 8068 1767 8102 1801
rect 8140 1767 8174 1801
rect 7996 1671 8030 1705
rect 8068 1671 8102 1705
rect 8140 1671 8174 1705
rect 7996 1575 8030 1609
rect 8068 1575 8102 1609
rect 8140 1575 8174 1609
rect 7996 1479 8030 1513
rect 8068 1479 8102 1513
rect 8140 1479 8174 1513
rect 7996 1383 8030 1417
rect 8068 1383 8102 1417
rect 8140 1383 8174 1417
rect 7996 1287 8030 1321
rect 8068 1287 8102 1321
rect 8140 1287 8174 1321
rect 7996 1191 8030 1225
rect 8068 1191 8102 1225
rect 8140 1191 8174 1225
rect 7996 1095 8030 1129
rect 8068 1095 8102 1129
rect 8140 1095 8174 1129
rect 7996 999 8030 1033
rect 8068 999 8102 1033
rect 8140 999 8174 1033
rect 7996 903 8030 937
rect 8068 903 8102 937
rect 8140 903 8174 937
rect 7996 807 8030 841
rect 8068 807 8102 841
rect 8140 807 8174 841
rect 7996 711 8030 745
rect 8068 711 8102 745
rect 8140 711 8174 745
rect 7996 615 8030 649
rect 8068 615 8102 649
rect 8140 615 8174 649
rect 8408 3303 8442 3337
rect 8480 3303 8514 3337
rect 8552 3303 8586 3337
rect 8408 3207 8442 3241
rect 8480 3207 8514 3241
rect 8552 3207 8586 3241
rect 8408 3111 8442 3145
rect 8480 3111 8514 3145
rect 8552 3111 8586 3145
rect 8408 3015 8442 3049
rect 8480 3015 8514 3049
rect 8552 3015 8586 3049
rect 8408 2919 8442 2953
rect 8480 2919 8514 2953
rect 8552 2919 8586 2953
rect 8408 2823 8442 2857
rect 8480 2823 8514 2857
rect 8552 2823 8586 2857
rect 8408 2727 8442 2761
rect 8480 2727 8514 2761
rect 8552 2727 8586 2761
rect 8408 2631 8442 2665
rect 8480 2631 8514 2665
rect 8552 2631 8586 2665
rect 8408 2535 8442 2569
rect 8480 2535 8514 2569
rect 8552 2535 8586 2569
rect 8408 2439 8442 2473
rect 8480 2439 8514 2473
rect 8552 2439 8586 2473
rect 8408 2343 8442 2377
rect 8480 2343 8514 2377
rect 8552 2343 8586 2377
rect 8408 2247 8442 2281
rect 8480 2247 8514 2281
rect 8552 2247 8586 2281
rect 8408 2151 8442 2185
rect 8480 2151 8514 2185
rect 8552 2151 8586 2185
rect 8408 2055 8442 2089
rect 8480 2055 8514 2089
rect 8552 2055 8586 2089
rect 8408 1959 8442 1993
rect 8480 1959 8514 1993
rect 8552 1959 8586 1993
rect 8408 1863 8442 1897
rect 8480 1863 8514 1897
rect 8552 1863 8586 1897
rect 8408 1767 8442 1801
rect 8480 1767 8514 1801
rect 8552 1767 8586 1801
rect 8408 1671 8442 1705
rect 8480 1671 8514 1705
rect 8552 1671 8586 1705
rect 8408 1575 8442 1609
rect 8480 1575 8514 1609
rect 8552 1575 8586 1609
rect 8408 1479 8442 1513
rect 8480 1479 8514 1513
rect 8552 1479 8586 1513
rect 8408 1383 8442 1417
rect 8480 1383 8514 1417
rect 8552 1383 8586 1417
rect 8408 1287 8442 1321
rect 8480 1287 8514 1321
rect 8552 1287 8586 1321
rect 8408 1191 8442 1225
rect 8480 1191 8514 1225
rect 8552 1191 8586 1225
rect 8408 1095 8442 1129
rect 8480 1095 8514 1129
rect 8552 1095 8586 1129
rect 8408 999 8442 1033
rect 8480 999 8514 1033
rect 8552 999 8586 1033
rect 8408 903 8442 937
rect 8480 903 8514 937
rect 8552 903 8586 937
rect 8408 807 8442 841
rect 8480 807 8514 841
rect 8552 807 8586 841
rect 8408 711 8442 745
rect 8480 711 8514 745
rect 8552 711 8586 745
rect 8408 615 8442 649
rect 8480 615 8514 649
rect 8552 615 8586 649
rect 8820 3303 8854 3337
rect 8892 3303 8926 3337
rect 8964 3303 8998 3337
rect 8820 3207 8854 3241
rect 8892 3207 8926 3241
rect 8964 3207 8998 3241
rect 8820 3111 8854 3145
rect 8892 3111 8926 3145
rect 8964 3111 8998 3145
rect 8820 3015 8854 3049
rect 8892 3015 8926 3049
rect 8964 3015 8998 3049
rect 8820 2919 8854 2953
rect 8892 2919 8926 2953
rect 8964 2919 8998 2953
rect 8820 2823 8854 2857
rect 8892 2823 8926 2857
rect 8964 2823 8998 2857
rect 8820 2727 8854 2761
rect 8892 2727 8926 2761
rect 8964 2727 8998 2761
rect 8820 2631 8854 2665
rect 8892 2631 8926 2665
rect 8964 2631 8998 2665
rect 8820 2535 8854 2569
rect 8892 2535 8926 2569
rect 8964 2535 8998 2569
rect 8820 2439 8854 2473
rect 8892 2439 8926 2473
rect 8964 2439 8998 2473
rect 8820 2343 8854 2377
rect 8892 2343 8926 2377
rect 8964 2343 8998 2377
rect 8820 2247 8854 2281
rect 8892 2247 8926 2281
rect 8964 2247 8998 2281
rect 8820 2151 8854 2185
rect 8892 2151 8926 2185
rect 8964 2151 8998 2185
rect 8820 2055 8854 2089
rect 8892 2055 8926 2089
rect 8964 2055 8998 2089
rect 8820 1959 8854 1993
rect 8892 1959 8926 1993
rect 8964 1959 8998 1993
rect 8820 1863 8854 1897
rect 8892 1863 8926 1897
rect 8964 1863 8998 1897
rect 8820 1767 8854 1801
rect 8892 1767 8926 1801
rect 8964 1767 8998 1801
rect 8820 1671 8854 1705
rect 8892 1671 8926 1705
rect 8964 1671 8998 1705
rect 8820 1575 8854 1609
rect 8892 1575 8926 1609
rect 8964 1575 8998 1609
rect 8820 1479 8854 1513
rect 8892 1479 8926 1513
rect 8964 1479 8998 1513
rect 8820 1383 8854 1417
rect 8892 1383 8926 1417
rect 8964 1383 8998 1417
rect 8820 1287 8854 1321
rect 8892 1287 8926 1321
rect 8964 1287 8998 1321
rect 8820 1191 8854 1225
rect 8892 1191 8926 1225
rect 8964 1191 8998 1225
rect 8820 1095 8854 1129
rect 8892 1095 8926 1129
rect 8964 1095 8998 1129
rect 8820 999 8854 1033
rect 8892 999 8926 1033
rect 8964 999 8998 1033
rect 8820 903 8854 937
rect 8892 903 8926 937
rect 8964 903 8998 937
rect 8820 807 8854 841
rect 8892 807 8926 841
rect 8964 807 8998 841
rect 8820 711 8854 745
rect 8892 711 8926 745
rect 8964 711 8998 745
rect 8820 615 8854 649
rect 8892 615 8926 649
rect 8964 615 8998 649
rect 9232 3303 9266 3337
rect 9304 3303 9338 3337
rect 9376 3303 9410 3337
rect 9232 3207 9266 3241
rect 9304 3207 9338 3241
rect 9376 3207 9410 3241
rect 9232 3111 9266 3145
rect 9304 3111 9338 3145
rect 9376 3111 9410 3145
rect 9232 3015 9266 3049
rect 9304 3015 9338 3049
rect 9376 3015 9410 3049
rect 9232 2919 9266 2953
rect 9304 2919 9338 2953
rect 9376 2919 9410 2953
rect 9232 2823 9266 2857
rect 9304 2823 9338 2857
rect 9376 2823 9410 2857
rect 9232 2727 9266 2761
rect 9304 2727 9338 2761
rect 9376 2727 9410 2761
rect 9232 2631 9266 2665
rect 9304 2631 9338 2665
rect 9376 2631 9410 2665
rect 9232 2535 9266 2569
rect 9304 2535 9338 2569
rect 9376 2535 9410 2569
rect 9232 2439 9266 2473
rect 9304 2439 9338 2473
rect 9376 2439 9410 2473
rect 9232 2343 9266 2377
rect 9304 2343 9338 2377
rect 9376 2343 9410 2377
rect 9232 2247 9266 2281
rect 9304 2247 9338 2281
rect 9376 2247 9410 2281
rect 9232 2151 9266 2185
rect 9304 2151 9338 2185
rect 9376 2151 9410 2185
rect 9232 2055 9266 2089
rect 9304 2055 9338 2089
rect 9376 2055 9410 2089
rect 9232 1959 9266 1993
rect 9304 1959 9338 1993
rect 9376 1959 9410 1993
rect 9232 1863 9266 1897
rect 9304 1863 9338 1897
rect 9376 1863 9410 1897
rect 9232 1767 9266 1801
rect 9304 1767 9338 1801
rect 9376 1767 9410 1801
rect 9232 1671 9266 1705
rect 9304 1671 9338 1705
rect 9376 1671 9410 1705
rect 9232 1575 9266 1609
rect 9304 1575 9338 1609
rect 9376 1575 9410 1609
rect 9232 1479 9266 1513
rect 9304 1479 9338 1513
rect 9376 1479 9410 1513
rect 9232 1383 9266 1417
rect 9304 1383 9338 1417
rect 9376 1383 9410 1417
rect 9232 1287 9266 1321
rect 9304 1287 9338 1321
rect 9376 1287 9410 1321
rect 9232 1191 9266 1225
rect 9304 1191 9338 1225
rect 9376 1191 9410 1225
rect 9232 1095 9266 1129
rect 9304 1095 9338 1129
rect 9376 1095 9410 1129
rect 9232 999 9266 1033
rect 9304 999 9338 1033
rect 9376 999 9410 1033
rect 9232 903 9266 937
rect 9304 903 9338 937
rect 9376 903 9410 937
rect 9232 807 9266 841
rect 9304 807 9338 841
rect 9376 807 9410 841
rect 9232 711 9266 745
rect 9304 711 9338 745
rect 9376 711 9410 745
rect 9232 615 9266 649
rect 9304 615 9338 649
rect 9376 615 9410 649
rect 9644 3303 9678 3337
rect 9716 3303 9750 3337
rect 9788 3303 9822 3337
rect 9644 3207 9678 3241
rect 9716 3207 9750 3241
rect 9788 3207 9822 3241
rect 9644 3111 9678 3145
rect 9716 3111 9750 3145
rect 9788 3111 9822 3145
rect 9644 3015 9678 3049
rect 9716 3015 9750 3049
rect 9788 3015 9822 3049
rect 9644 2919 9678 2953
rect 9716 2919 9750 2953
rect 9788 2919 9822 2953
rect 9644 2823 9678 2857
rect 9716 2823 9750 2857
rect 9788 2823 9822 2857
rect 9644 2727 9678 2761
rect 9716 2727 9750 2761
rect 9788 2727 9822 2761
rect 9644 2631 9678 2665
rect 9716 2631 9750 2665
rect 9788 2631 9822 2665
rect 9644 2535 9678 2569
rect 9716 2535 9750 2569
rect 9788 2535 9822 2569
rect 9644 2439 9678 2473
rect 9716 2439 9750 2473
rect 9788 2439 9822 2473
rect 9644 2343 9678 2377
rect 9716 2343 9750 2377
rect 9788 2343 9822 2377
rect 9644 2247 9678 2281
rect 9716 2247 9750 2281
rect 9788 2247 9822 2281
rect 9644 2151 9678 2185
rect 9716 2151 9750 2185
rect 9788 2151 9822 2185
rect 9644 2055 9678 2089
rect 9716 2055 9750 2089
rect 9788 2055 9822 2089
rect 9644 1959 9678 1993
rect 9716 1959 9750 1993
rect 9788 1959 9822 1993
rect 9644 1863 9678 1897
rect 9716 1863 9750 1897
rect 9788 1863 9822 1897
rect 9644 1767 9678 1801
rect 9716 1767 9750 1801
rect 9788 1767 9822 1801
rect 9644 1671 9678 1705
rect 9716 1671 9750 1705
rect 9788 1671 9822 1705
rect 9644 1575 9678 1609
rect 9716 1575 9750 1609
rect 9788 1575 9822 1609
rect 9644 1479 9678 1513
rect 9716 1479 9750 1513
rect 9788 1479 9822 1513
rect 9644 1383 9678 1417
rect 9716 1383 9750 1417
rect 9788 1383 9822 1417
rect 9644 1287 9678 1321
rect 9716 1287 9750 1321
rect 9788 1287 9822 1321
rect 9644 1191 9678 1225
rect 9716 1191 9750 1225
rect 9788 1191 9822 1225
rect 9644 1095 9678 1129
rect 9716 1095 9750 1129
rect 9788 1095 9822 1129
rect 9644 999 9678 1033
rect 9716 999 9750 1033
rect 9788 999 9822 1033
rect 9644 903 9678 937
rect 9716 903 9750 937
rect 9788 903 9822 937
rect 9644 807 9678 841
rect 9716 807 9750 841
rect 9788 807 9822 841
rect 9644 711 9678 745
rect 9716 711 9750 745
rect 9788 711 9822 745
rect 9644 615 9678 649
rect 9716 615 9750 649
rect 9788 615 9822 649
rect 10056 3303 10090 3337
rect 10128 3303 10162 3337
rect 10200 3303 10234 3337
rect 10056 3207 10090 3241
rect 10128 3207 10162 3241
rect 10200 3207 10234 3241
rect 10056 3111 10090 3145
rect 10128 3111 10162 3145
rect 10200 3111 10234 3145
rect 10056 3015 10090 3049
rect 10128 3015 10162 3049
rect 10200 3015 10234 3049
rect 10056 2919 10090 2953
rect 10128 2919 10162 2953
rect 10200 2919 10234 2953
rect 10056 2823 10090 2857
rect 10128 2823 10162 2857
rect 10200 2823 10234 2857
rect 10056 2727 10090 2761
rect 10128 2727 10162 2761
rect 10200 2727 10234 2761
rect 10056 2631 10090 2665
rect 10128 2631 10162 2665
rect 10200 2631 10234 2665
rect 10056 2535 10090 2569
rect 10128 2535 10162 2569
rect 10200 2535 10234 2569
rect 10056 2439 10090 2473
rect 10128 2439 10162 2473
rect 10200 2439 10234 2473
rect 10056 2343 10090 2377
rect 10128 2343 10162 2377
rect 10200 2343 10234 2377
rect 10056 2247 10090 2281
rect 10128 2247 10162 2281
rect 10200 2247 10234 2281
rect 10056 2151 10090 2185
rect 10128 2151 10162 2185
rect 10200 2151 10234 2185
rect 10056 2055 10090 2089
rect 10128 2055 10162 2089
rect 10200 2055 10234 2089
rect 10056 1959 10090 1993
rect 10128 1959 10162 1993
rect 10200 1959 10234 1993
rect 10056 1863 10090 1897
rect 10128 1863 10162 1897
rect 10200 1863 10234 1897
rect 10056 1767 10090 1801
rect 10128 1767 10162 1801
rect 10200 1767 10234 1801
rect 10056 1671 10090 1705
rect 10128 1671 10162 1705
rect 10200 1671 10234 1705
rect 10056 1575 10090 1609
rect 10128 1575 10162 1609
rect 10200 1575 10234 1609
rect 10056 1479 10090 1513
rect 10128 1479 10162 1513
rect 10200 1479 10234 1513
rect 10056 1383 10090 1417
rect 10128 1383 10162 1417
rect 10200 1383 10234 1417
rect 10056 1287 10090 1321
rect 10128 1287 10162 1321
rect 10200 1287 10234 1321
rect 10056 1191 10090 1225
rect 10128 1191 10162 1225
rect 10200 1191 10234 1225
rect 10056 1095 10090 1129
rect 10128 1095 10162 1129
rect 10200 1095 10234 1129
rect 10056 999 10090 1033
rect 10128 999 10162 1033
rect 10200 999 10234 1033
rect 10056 903 10090 937
rect 10128 903 10162 937
rect 10200 903 10234 937
rect 10056 807 10090 841
rect 10128 807 10162 841
rect 10200 807 10234 841
rect 10056 711 10090 745
rect 10128 711 10162 745
rect 10200 711 10234 745
rect 10056 615 10090 649
rect 10128 615 10162 649
rect 10200 615 10234 649
rect 10468 3303 10502 3337
rect 10540 3303 10574 3337
rect 10612 3303 10646 3337
rect 10468 3207 10502 3241
rect 10540 3207 10574 3241
rect 10612 3207 10646 3241
rect 10468 3111 10502 3145
rect 10540 3111 10574 3145
rect 10612 3111 10646 3145
rect 10468 3015 10502 3049
rect 10540 3015 10574 3049
rect 10612 3015 10646 3049
rect 10468 2919 10502 2953
rect 10540 2919 10574 2953
rect 10612 2919 10646 2953
rect 10468 2823 10502 2857
rect 10540 2823 10574 2857
rect 10612 2823 10646 2857
rect 10468 2727 10502 2761
rect 10540 2727 10574 2761
rect 10612 2727 10646 2761
rect 10468 2631 10502 2665
rect 10540 2631 10574 2665
rect 10612 2631 10646 2665
rect 10468 2535 10502 2569
rect 10540 2535 10574 2569
rect 10612 2535 10646 2569
rect 10468 2439 10502 2473
rect 10540 2439 10574 2473
rect 10612 2439 10646 2473
rect 10468 2343 10502 2377
rect 10540 2343 10574 2377
rect 10612 2343 10646 2377
rect 10468 2247 10502 2281
rect 10540 2247 10574 2281
rect 10612 2247 10646 2281
rect 10468 2151 10502 2185
rect 10540 2151 10574 2185
rect 10612 2151 10646 2185
rect 10468 2055 10502 2089
rect 10540 2055 10574 2089
rect 10612 2055 10646 2089
rect 10468 1959 10502 1993
rect 10540 1959 10574 1993
rect 10612 1959 10646 1993
rect 10468 1863 10502 1897
rect 10540 1863 10574 1897
rect 10612 1863 10646 1897
rect 10468 1767 10502 1801
rect 10540 1767 10574 1801
rect 10612 1767 10646 1801
rect 10468 1671 10502 1705
rect 10540 1671 10574 1705
rect 10612 1671 10646 1705
rect 10468 1575 10502 1609
rect 10540 1575 10574 1609
rect 10612 1575 10646 1609
rect 10468 1479 10502 1513
rect 10540 1479 10574 1513
rect 10612 1479 10646 1513
rect 10468 1383 10502 1417
rect 10540 1383 10574 1417
rect 10612 1383 10646 1417
rect 10468 1287 10502 1321
rect 10540 1287 10574 1321
rect 10612 1287 10646 1321
rect 10468 1191 10502 1225
rect 10540 1191 10574 1225
rect 10612 1191 10646 1225
rect 10468 1095 10502 1129
rect 10540 1095 10574 1129
rect 10612 1095 10646 1129
rect 10468 999 10502 1033
rect 10540 999 10574 1033
rect 10612 999 10646 1033
rect 10468 903 10502 937
rect 10540 903 10574 937
rect 10612 903 10646 937
rect 10468 807 10502 841
rect 10540 807 10574 841
rect 10612 807 10646 841
rect 10468 711 10502 745
rect 10540 711 10574 745
rect 10612 711 10646 745
rect 10468 615 10502 649
rect 10540 615 10574 649
rect 10612 615 10646 649
rect 10880 3303 10914 3337
rect 10952 3303 10986 3337
rect 11024 3303 11058 3337
rect 10880 3207 10914 3241
rect 10952 3207 10986 3241
rect 11024 3207 11058 3241
rect 10880 3111 10914 3145
rect 10952 3111 10986 3145
rect 11024 3111 11058 3145
rect 10880 3015 10914 3049
rect 10952 3015 10986 3049
rect 11024 3015 11058 3049
rect 10880 2919 10914 2953
rect 10952 2919 10986 2953
rect 11024 2919 11058 2953
rect 10880 2823 10914 2857
rect 10952 2823 10986 2857
rect 11024 2823 11058 2857
rect 10880 2727 10914 2761
rect 10952 2727 10986 2761
rect 11024 2727 11058 2761
rect 10880 2631 10914 2665
rect 10952 2631 10986 2665
rect 11024 2631 11058 2665
rect 10880 2535 10914 2569
rect 10952 2535 10986 2569
rect 11024 2535 11058 2569
rect 10880 2439 10914 2473
rect 10952 2439 10986 2473
rect 11024 2439 11058 2473
rect 10880 2343 10914 2377
rect 10952 2343 10986 2377
rect 11024 2343 11058 2377
rect 10880 2247 10914 2281
rect 10952 2247 10986 2281
rect 11024 2247 11058 2281
rect 10880 2151 10914 2185
rect 10952 2151 10986 2185
rect 11024 2151 11058 2185
rect 10880 2055 10914 2089
rect 10952 2055 10986 2089
rect 11024 2055 11058 2089
rect 10880 1959 10914 1993
rect 10952 1959 10986 1993
rect 11024 1959 11058 1993
rect 10880 1863 10914 1897
rect 10952 1863 10986 1897
rect 11024 1863 11058 1897
rect 10880 1767 10914 1801
rect 10952 1767 10986 1801
rect 11024 1767 11058 1801
rect 10880 1671 10914 1705
rect 10952 1671 10986 1705
rect 11024 1671 11058 1705
rect 10880 1575 10914 1609
rect 10952 1575 10986 1609
rect 11024 1575 11058 1609
rect 10880 1479 10914 1513
rect 10952 1479 10986 1513
rect 11024 1479 11058 1513
rect 10880 1383 10914 1417
rect 10952 1383 10986 1417
rect 11024 1383 11058 1417
rect 10880 1287 10914 1321
rect 10952 1287 10986 1321
rect 11024 1287 11058 1321
rect 10880 1191 10914 1225
rect 10952 1191 10986 1225
rect 11024 1191 11058 1225
rect 10880 1095 10914 1129
rect 10952 1095 10986 1129
rect 11024 1095 11058 1129
rect 10880 999 10914 1033
rect 10952 999 10986 1033
rect 11024 999 11058 1033
rect 10880 903 10914 937
rect 10952 903 10986 937
rect 11024 903 11058 937
rect 10880 807 10914 841
rect 10952 807 10986 841
rect 11024 807 11058 841
rect 10880 711 10914 745
rect 10952 711 10986 745
rect 11024 711 11058 745
rect 10880 615 10914 649
rect 10952 615 10986 649
rect 11024 615 11058 649
rect 11338 3455 11341 3464
rect 11341 3455 11372 3464
rect 11338 3430 11372 3455
rect 11338 3387 11341 3392
rect 11341 3387 11372 3392
rect 11338 3358 11372 3387
rect 11338 3319 11341 3320
rect 11341 3319 11372 3320
rect 11338 3286 11372 3319
rect 11338 3217 11372 3248
rect 11338 3214 11341 3217
rect 11341 3214 11372 3217
rect 11338 3149 11372 3176
rect 11338 3142 11341 3149
rect 11341 3142 11372 3149
rect 11338 3081 11372 3104
rect 11338 3070 11341 3081
rect 11341 3070 11372 3081
rect 11338 3013 11372 3032
rect 11338 2998 11341 3013
rect 11341 2998 11372 3013
rect 11338 2945 11372 2960
rect 11338 2926 11341 2945
rect 11341 2926 11372 2945
rect 11338 2877 11372 2888
rect 11338 2854 11341 2877
rect 11341 2854 11372 2877
rect 11338 2809 11372 2816
rect 11338 2782 11341 2809
rect 11341 2782 11372 2809
rect 11338 2741 11372 2744
rect 11338 2710 11341 2741
rect 11341 2710 11372 2741
rect 11338 2639 11341 2672
rect 11341 2639 11372 2672
rect 11338 2638 11372 2639
rect 11338 2571 11341 2600
rect 11341 2571 11372 2600
rect 11338 2566 11372 2571
rect 11338 2503 11341 2528
rect 11341 2503 11372 2528
rect 11338 2494 11372 2503
rect 11338 2435 11341 2456
rect 11341 2435 11372 2456
rect 11338 2422 11372 2435
rect 11338 2367 11341 2384
rect 11341 2367 11372 2384
rect 11338 2350 11372 2367
rect 11338 2299 11341 2312
rect 11341 2299 11372 2312
rect 11338 2278 11372 2299
rect 11338 2231 11341 2240
rect 11341 2231 11372 2240
rect 11338 2206 11372 2231
rect 11338 2163 11341 2168
rect 11341 2163 11372 2168
rect 11338 2134 11372 2163
rect 11338 2095 11341 2096
rect 11341 2095 11372 2096
rect 11338 2062 11372 2095
rect 11338 1993 11372 2024
rect 11338 1990 11341 1993
rect 11341 1990 11372 1993
rect 11338 1925 11372 1952
rect 11338 1918 11341 1925
rect 11341 1918 11372 1925
rect 11338 1857 11372 1880
rect 11338 1846 11341 1857
rect 11341 1846 11372 1857
rect 11338 1789 11372 1808
rect 11338 1774 11341 1789
rect 11341 1774 11372 1789
rect 11338 1721 11372 1736
rect 11338 1702 11341 1721
rect 11341 1702 11372 1721
rect 11338 1653 11372 1664
rect 11338 1630 11341 1653
rect 11341 1630 11372 1653
rect 11338 1585 11372 1592
rect 11338 1558 11341 1585
rect 11341 1558 11372 1585
rect 11338 1517 11372 1520
rect 11338 1486 11341 1517
rect 11341 1486 11372 1517
rect 11338 1415 11341 1448
rect 11341 1415 11372 1448
rect 11338 1414 11372 1415
rect 11338 1347 11341 1376
rect 11341 1347 11372 1376
rect 11338 1342 11372 1347
rect 11338 1279 11341 1304
rect 11341 1279 11372 1304
rect 11338 1270 11372 1279
rect 11338 1211 11341 1232
rect 11341 1211 11372 1232
rect 11338 1198 11372 1211
rect 11338 1143 11341 1160
rect 11341 1143 11372 1160
rect 11338 1126 11372 1143
rect 11338 1075 11341 1088
rect 11341 1075 11372 1088
rect 11338 1054 11372 1075
rect 11338 1007 11341 1016
rect 11341 1007 11372 1016
rect 11338 982 11372 1007
rect 11338 939 11341 944
rect 11341 939 11372 944
rect 11338 910 11372 939
rect 11338 871 11341 872
rect 11341 871 11372 872
rect 11338 838 11372 871
rect 11338 769 11372 800
rect 11338 766 11341 769
rect 11341 766 11372 769
rect 11338 701 11372 728
rect 11338 694 11341 701
rect 11341 694 11372 701
rect 11338 633 11372 656
rect 11338 622 11341 633
rect 11341 622 11372 633
<< metal1 >>
rect 7147 3750 11399 3756
rect 7147 3740 7342 3750
rect 7376 3740 7501 3750
rect 7535 3740 7574 3750
rect 7608 3740 7646 3750
rect 7680 3740 7718 3750
rect 7752 3740 7790 3750
rect 7824 3740 7862 3750
rect 7896 3740 7934 3750
rect 7968 3740 8006 3750
rect 8040 3740 8078 3750
rect 8112 3740 8150 3750
rect 8184 3740 8222 3750
rect 8256 3740 8294 3750
rect 8328 3740 8366 3750
rect 8400 3740 8438 3750
rect 8472 3740 8510 3750
rect 8544 3740 8582 3750
rect 8616 3740 8654 3750
rect 8688 3740 8726 3750
rect 8760 3740 8798 3750
rect 8832 3740 8870 3750
rect 8904 3740 8942 3750
rect 8976 3740 9014 3750
rect 9048 3740 9086 3750
rect 9120 3740 9158 3750
rect 9192 3740 9230 3750
rect 9264 3740 9302 3750
rect 9336 3740 9374 3750
rect 9408 3740 9446 3750
rect 9480 3740 9518 3750
rect 9552 3740 9590 3750
rect 9624 3740 9662 3750
rect 9696 3740 9734 3750
rect 9768 3740 9806 3750
rect 9840 3740 9878 3750
rect 9912 3740 9950 3750
rect 9984 3740 10022 3750
rect 10056 3740 10094 3750
rect 10128 3740 10166 3750
rect 10200 3740 10238 3750
rect 10272 3740 10310 3750
rect 10344 3740 10382 3750
rect 10416 3740 10454 3750
rect 10488 3740 10526 3750
rect 10560 3740 10598 3750
rect 10632 3740 10670 3750
rect 10704 3740 10742 3750
rect 10776 3740 10814 3750
rect 10848 3740 10886 3750
rect 7147 3624 7215 3740
rect 10851 3716 10886 3740
rect 10920 3716 10958 3750
rect 10992 3716 11030 3750
rect 11064 3716 11102 3750
rect 11136 3716 11260 3750
rect 11294 3716 11399 3750
rect 10851 3642 11399 3716
rect 10851 3624 10886 3642
rect 7147 3622 7342 3624
rect 7147 3588 7264 3622
rect 7298 3608 7342 3622
rect 7376 3608 7501 3624
rect 7535 3608 7574 3624
rect 7608 3608 7646 3624
rect 7680 3608 7718 3624
rect 7752 3608 7790 3624
rect 7824 3608 7862 3624
rect 7896 3608 7934 3624
rect 7968 3608 8006 3624
rect 8040 3608 8078 3624
rect 8112 3608 8150 3624
rect 8184 3608 8222 3624
rect 8256 3608 8294 3624
rect 8328 3608 8366 3624
rect 8400 3608 8438 3624
rect 8472 3608 8510 3624
rect 8544 3608 8582 3624
rect 8616 3608 8654 3624
rect 8688 3608 8726 3624
rect 8760 3608 8798 3624
rect 8832 3608 8870 3624
rect 8904 3608 8942 3624
rect 8976 3608 9014 3624
rect 9048 3608 9086 3624
rect 9120 3608 9158 3624
rect 9192 3608 9230 3624
rect 9264 3608 9302 3624
rect 9336 3608 9374 3624
rect 9408 3608 9446 3624
rect 9480 3608 9518 3624
rect 9552 3608 9590 3624
rect 9624 3608 9662 3624
rect 9696 3608 9734 3624
rect 9768 3608 9806 3624
rect 9840 3608 9878 3624
rect 9912 3608 9950 3624
rect 9984 3608 10022 3624
rect 10056 3608 10094 3624
rect 10128 3608 10166 3624
rect 10200 3608 10238 3624
rect 10272 3608 10310 3624
rect 10344 3608 10382 3624
rect 10416 3608 10454 3624
rect 10488 3608 10526 3624
rect 10560 3608 10598 3624
rect 10632 3608 10670 3624
rect 10704 3608 10742 3624
rect 10776 3608 10814 3624
rect 10848 3608 10886 3624
rect 10920 3608 10958 3642
rect 10992 3608 11030 3642
rect 11064 3608 11102 3642
rect 11136 3608 11260 3642
rect 11294 3622 11399 3642
rect 11294 3608 11338 3622
rect 7298 3602 11338 3608
rect 7298 3588 7359 3602
tri 7359 3588 7373 3602 nw
tri 11283 3588 11297 3602 ne
rect 11297 3588 11338 3602
rect 11372 3588 11399 3622
rect 7147 3464 7325 3588
tri 7325 3554 7359 3588 nw
tri 11297 3568 11317 3588 ne
tri 7571 3464 7583 3476 se
rect 7583 3464 7763 3476
tri 7763 3464 7775 3476 sw
tri 7983 3464 7995 3476 se
rect 7995 3464 8175 3476
tri 8175 3464 8187 3476 sw
tri 8395 3464 8407 3476 se
rect 8407 3464 8587 3476
tri 8587 3464 8599 3476 sw
tri 8807 3464 8819 3476 se
rect 8819 3464 8999 3476
tri 8999 3464 9011 3476 sw
tri 9219 3464 9231 3476 se
rect 9231 3464 9411 3476
tri 9411 3464 9423 3476 sw
tri 9631 3464 9643 3476 se
rect 9643 3464 9823 3476
tri 9823 3464 9835 3476 sw
tri 10043 3464 10055 3476 se
rect 10055 3464 10235 3476
tri 10235 3464 10247 3476 sw
tri 10455 3464 10467 3476 se
rect 10467 3464 10647 3476
tri 10647 3464 10659 3476 sw
tri 10867 3464 10879 3476 se
rect 10879 3464 11059 3476
tri 11059 3464 11071 3476 sw
rect 11317 3464 11399 3588
rect 7147 3430 7264 3464
rect 7298 3430 7325 3464
tri 7537 3430 7571 3464 se
rect 7571 3430 7775 3464
tri 7775 3430 7809 3464 sw
tri 7949 3430 7983 3464 se
rect 7983 3430 8187 3464
tri 8187 3430 8221 3464 sw
tri 8361 3430 8395 3464 se
rect 8395 3430 8599 3464
tri 8599 3430 8633 3464 sw
tri 8773 3430 8807 3464 se
rect 8807 3430 9011 3464
tri 9011 3430 9045 3464 sw
tri 9185 3430 9219 3464 se
rect 9219 3430 9423 3464
tri 9423 3430 9457 3464 sw
tri 9597 3430 9631 3464 se
rect 9631 3430 9835 3464
tri 9835 3430 9869 3464 sw
tri 10009 3430 10043 3464 se
rect 10043 3430 10247 3464
tri 10247 3430 10281 3464 sw
tri 10421 3430 10455 3464 se
rect 10455 3430 10659 3464
tri 10659 3430 10693 3464 sw
tri 10833 3430 10867 3464 se
rect 10867 3430 11071 3464
tri 11071 3430 11105 3464 sw
rect 11317 3430 11338 3464
rect 11372 3430 11399 3464
rect 7147 3392 7325 3430
rect 7147 3358 7264 3392
rect 7298 3358 7325 3392
rect 7147 3320 7325 3358
rect 7147 3286 7264 3320
rect 7298 3286 7325 3320
rect 7147 3248 7325 3286
rect 7147 3214 7264 3248
rect 7298 3214 7325 3248
rect 7147 3176 7325 3214
rect 7147 3142 7264 3176
rect 7298 3142 7325 3176
rect 7147 3104 7325 3142
rect 7147 3070 7264 3104
rect 7298 3070 7325 3104
rect 7147 3032 7325 3070
rect 7147 2998 7264 3032
rect 7298 2998 7325 3032
rect 7147 2960 7325 2998
rect 7147 2926 7264 2960
rect 7298 2926 7325 2960
rect 7147 2888 7325 2926
rect 7147 2854 7264 2888
rect 7298 2854 7325 2888
rect 7147 2816 7325 2854
rect 7147 2782 7264 2816
rect 7298 2782 7325 2816
rect 7147 2744 7325 2782
rect 7147 2710 7264 2744
rect 7298 2710 7325 2744
rect 7147 2672 7325 2710
rect 7147 2638 7264 2672
rect 7298 2638 7325 2672
rect 7147 2600 7325 2638
rect 7147 2566 7264 2600
rect 7298 2566 7325 2600
rect 7147 2528 7325 2566
rect 7147 2494 7264 2528
rect 7298 2494 7325 2528
rect 7147 2456 7325 2494
rect 7147 2422 7264 2456
rect 7298 2422 7325 2456
rect 7147 2384 7325 2422
rect 7147 2350 7264 2384
rect 7298 2350 7325 2384
rect 7147 2312 7325 2350
rect 7147 2278 7264 2312
rect 7298 2278 7325 2312
rect 7147 2240 7325 2278
rect 7147 2206 7264 2240
rect 7298 2206 7325 2240
rect 7147 2168 7325 2206
rect 7147 2134 7264 2168
rect 7298 2134 7325 2168
rect 7147 2096 7325 2134
rect 7147 2062 7264 2096
rect 7298 2062 7325 2096
rect 7147 2024 7325 2062
rect 7147 1990 7264 2024
rect 7298 1990 7325 2024
rect 7147 1952 7325 1990
rect 7147 1918 7264 1952
rect 7298 1918 7325 1952
rect 7147 1880 7325 1918
rect 7147 1846 7264 1880
rect 7298 1846 7325 1880
rect 7147 1808 7325 1846
rect 7147 1774 7264 1808
rect 7298 1774 7325 1808
rect 7147 1736 7325 1774
rect 7147 1702 7264 1736
rect 7298 1702 7325 1736
rect 7147 1664 7325 1702
rect 7147 1630 7264 1664
rect 7298 1630 7325 1664
rect 7147 1592 7325 1630
rect 7147 1558 7264 1592
rect 7298 1558 7325 1592
rect 7147 1520 7325 1558
rect 7147 1486 7264 1520
rect 7298 1486 7325 1520
rect 7147 1448 7325 1486
rect 7147 1414 7264 1448
rect 7298 1414 7325 1448
rect 7147 1376 7325 1414
rect 7147 1342 7264 1376
rect 7298 1342 7325 1376
rect 7147 1304 7325 1342
rect 7147 1270 7264 1304
rect 7298 1270 7325 1304
rect 7147 1232 7325 1270
rect 7147 1198 7264 1232
rect 7298 1198 7325 1232
rect 7147 1160 7325 1198
rect 7147 1126 7264 1160
rect 7298 1126 7325 1160
rect 7147 1088 7325 1126
rect 7147 1054 7264 1088
rect 7298 1054 7325 1088
rect 7147 1016 7325 1054
rect 7147 982 7264 1016
rect 7298 982 7325 1016
rect 7147 944 7325 982
rect 7147 910 7264 944
rect 7298 910 7325 944
rect 7147 872 7325 910
rect 7147 838 7264 872
rect 7298 838 7325 872
rect 7147 800 7325 838
rect 7147 766 7264 800
rect 7298 766 7325 800
rect 7147 728 7325 766
rect 7147 694 7264 728
rect 7298 694 7325 728
rect 7147 656 7325 694
rect 7147 622 7264 656
rect 7298 622 7325 656
rect 7147 609 7325 622
tri 7523 3416 7537 3430 se
rect 7537 3416 7809 3430
tri 7809 3416 7823 3430 sw
rect 7523 3382 7823 3416
rect 7523 2050 7551 3382
rect 7795 2050 7823 3382
rect 7523 1993 7823 2050
rect 7523 1959 7584 1993
rect 7618 1959 7656 1993
rect 7690 1959 7728 1993
rect 7762 1959 7823 1993
rect 7523 1897 7823 1959
rect 7523 1863 7584 1897
rect 7618 1863 7656 1897
rect 7690 1863 7728 1897
rect 7762 1863 7823 1897
rect 7523 1801 7823 1863
rect 7523 1767 7584 1801
rect 7618 1767 7656 1801
rect 7690 1767 7728 1801
rect 7762 1767 7823 1801
rect 7523 1705 7823 1767
rect 7523 1671 7584 1705
rect 7618 1671 7656 1705
rect 7690 1671 7728 1705
rect 7762 1671 7823 1705
rect 7523 1609 7823 1671
rect 7523 1575 7584 1609
rect 7618 1575 7656 1609
rect 7690 1575 7728 1609
rect 7762 1575 7823 1609
rect 7523 1513 7823 1575
rect 7523 1479 7584 1513
rect 7618 1479 7656 1513
rect 7690 1479 7728 1513
rect 7762 1479 7823 1513
rect 7523 1417 7823 1479
rect 7523 1383 7584 1417
rect 7618 1383 7656 1417
rect 7690 1383 7728 1417
rect 7762 1383 7823 1417
rect 7523 1321 7823 1383
rect 7523 1287 7584 1321
rect 7618 1287 7656 1321
rect 7690 1287 7728 1321
rect 7762 1287 7823 1321
rect 7523 1225 7823 1287
rect 7523 1191 7584 1225
rect 7618 1191 7656 1225
rect 7690 1191 7728 1225
rect 7762 1191 7823 1225
rect 7523 1129 7823 1191
rect 7523 1095 7584 1129
rect 7618 1095 7656 1129
rect 7690 1095 7728 1129
rect 7762 1095 7823 1129
rect 7523 1033 7823 1095
rect 7523 999 7584 1033
rect 7618 999 7656 1033
rect 7690 999 7728 1033
rect 7762 999 7823 1033
rect 7523 937 7823 999
rect 7523 903 7584 937
rect 7618 903 7656 937
rect 7690 903 7728 937
rect 7762 903 7823 937
rect 7523 841 7823 903
rect 7523 807 7584 841
rect 7618 807 7656 841
rect 7690 807 7728 841
rect 7762 807 7823 841
rect 7523 745 7823 807
rect 7523 711 7584 745
rect 7618 711 7656 745
rect 7690 711 7728 745
rect 7762 711 7823 745
rect 7523 649 7823 711
rect 7523 615 7584 649
rect 7618 615 7656 649
rect 7690 615 7728 649
rect 7762 615 7823 649
rect 7523 536 7823 615
tri 7523 476 7583 536 ne
rect 7583 476 7763 536
tri 7763 476 7823 536 nw
tri 7935 3416 7949 3430 se
rect 7949 3416 8221 3430
tri 8221 3416 8235 3430 sw
rect 7935 3337 8235 3416
rect 7935 3303 7996 3337
rect 8030 3303 8068 3337
rect 8102 3303 8140 3337
rect 8174 3303 8235 3337
rect 7935 3241 8235 3303
rect 7935 3207 7996 3241
rect 8030 3207 8068 3241
rect 8102 3207 8140 3241
rect 8174 3207 8235 3241
rect 7935 3145 8235 3207
rect 7935 3111 7996 3145
rect 8030 3111 8068 3145
rect 8102 3111 8140 3145
rect 8174 3111 8235 3145
rect 7935 3049 8235 3111
rect 7935 3015 7996 3049
rect 8030 3015 8068 3049
rect 8102 3015 8140 3049
rect 8174 3015 8235 3049
rect 7935 2953 8235 3015
rect 7935 2919 7996 2953
rect 8030 2919 8068 2953
rect 8102 2919 8140 2953
rect 8174 2919 8235 2953
rect 7935 2857 8235 2919
rect 7935 2823 7996 2857
rect 8030 2823 8068 2857
rect 8102 2823 8140 2857
rect 8174 2823 8235 2857
rect 7935 2761 8235 2823
rect 7935 2727 7996 2761
rect 8030 2727 8068 2761
rect 8102 2727 8140 2761
rect 8174 2727 8235 2761
rect 7935 2665 8235 2727
rect 7935 2631 7996 2665
rect 8030 2631 8068 2665
rect 8102 2631 8140 2665
rect 8174 2631 8235 2665
rect 7935 2569 8235 2631
rect 7935 2535 7996 2569
rect 8030 2535 8068 2569
rect 8102 2535 8140 2569
rect 8174 2535 8235 2569
rect 7935 2473 8235 2535
rect 7935 2439 7996 2473
rect 8030 2439 8068 2473
rect 8102 2439 8140 2473
rect 8174 2439 8235 2473
rect 7935 2377 8235 2439
rect 7935 2343 7996 2377
rect 8030 2343 8068 2377
rect 8102 2343 8140 2377
rect 8174 2343 8235 2377
rect 7935 2281 8235 2343
rect 7935 2247 7996 2281
rect 8030 2247 8068 2281
rect 8102 2247 8140 2281
rect 8174 2247 8235 2281
rect 7935 2185 8235 2247
rect 7935 2151 7996 2185
rect 8030 2151 8068 2185
rect 8102 2151 8140 2185
rect 8174 2151 8235 2185
rect 7935 2089 8235 2151
rect 7935 2055 7996 2089
rect 8030 2055 8068 2089
rect 8102 2055 8140 2089
rect 8174 2055 8235 2089
rect 7935 1993 8235 2055
rect 7935 1959 7996 1993
rect 8030 1959 8068 1993
rect 8102 1959 8140 1993
rect 8174 1959 8235 1993
rect 7935 1897 8235 1959
rect 7935 1888 7996 1897
rect 8030 1888 8068 1897
rect 8102 1888 8140 1897
rect 8174 1888 8235 1897
tri 7793 278 7935 420 se
rect 7935 300 7963 1888
rect 8207 300 8235 1888
tri 8347 3416 8361 3430 se
rect 8361 3416 8633 3430
tri 8633 3416 8647 3430 sw
rect 8347 3382 8647 3416
rect 8347 2050 8375 3382
rect 8619 2050 8647 3382
rect 8347 1993 8647 2050
rect 8347 1959 8408 1993
rect 8442 1959 8480 1993
rect 8514 1959 8552 1993
rect 8586 1959 8647 1993
rect 8347 1897 8647 1959
rect 8347 1863 8408 1897
rect 8442 1863 8480 1897
rect 8514 1863 8552 1897
rect 8586 1863 8647 1897
rect 8347 1801 8647 1863
rect 8347 1767 8408 1801
rect 8442 1767 8480 1801
rect 8514 1767 8552 1801
rect 8586 1767 8647 1801
rect 8347 1705 8647 1767
rect 8347 1671 8408 1705
rect 8442 1671 8480 1705
rect 8514 1671 8552 1705
rect 8586 1671 8647 1705
rect 8347 1609 8647 1671
rect 8347 1575 8408 1609
rect 8442 1575 8480 1609
rect 8514 1575 8552 1609
rect 8586 1575 8647 1609
rect 8347 1513 8647 1575
rect 8347 1479 8408 1513
rect 8442 1479 8480 1513
rect 8514 1479 8552 1513
rect 8586 1479 8647 1513
rect 8347 1417 8647 1479
rect 8347 1383 8408 1417
rect 8442 1383 8480 1417
rect 8514 1383 8552 1417
rect 8586 1383 8647 1417
rect 8347 1321 8647 1383
rect 8347 1287 8408 1321
rect 8442 1287 8480 1321
rect 8514 1287 8552 1321
rect 8586 1287 8647 1321
rect 8347 1225 8647 1287
rect 8347 1191 8408 1225
rect 8442 1191 8480 1225
rect 8514 1191 8552 1225
rect 8586 1191 8647 1225
rect 8347 1129 8647 1191
rect 8347 1095 8408 1129
rect 8442 1095 8480 1129
rect 8514 1095 8552 1129
rect 8586 1095 8647 1129
rect 8347 1033 8647 1095
rect 8347 999 8408 1033
rect 8442 999 8480 1033
rect 8514 999 8552 1033
rect 8586 999 8647 1033
rect 8347 937 8647 999
rect 8347 903 8408 937
rect 8442 903 8480 937
rect 8514 903 8552 937
rect 8586 903 8647 937
rect 8347 841 8647 903
rect 8347 807 8408 841
rect 8442 807 8480 841
rect 8514 807 8552 841
rect 8586 807 8647 841
rect 8347 745 8647 807
rect 8347 711 8408 745
rect 8442 711 8480 745
rect 8514 711 8552 745
rect 8586 711 8647 745
rect 8347 649 8647 711
rect 8347 615 8408 649
rect 8442 615 8480 649
rect 8514 615 8552 649
rect 8586 615 8647 649
rect 8347 536 8647 615
tri 8347 476 8407 536 ne
rect 8407 476 8587 536
tri 8587 476 8647 536 nw
tri 8759 3416 8773 3430 se
rect 8773 3416 9045 3430
tri 9045 3416 9059 3430 sw
rect 8759 3337 9059 3416
rect 8759 3303 8820 3337
rect 8854 3303 8892 3337
rect 8926 3303 8964 3337
rect 8998 3303 9059 3337
rect 8759 3241 9059 3303
rect 8759 3207 8820 3241
rect 8854 3207 8892 3241
rect 8926 3207 8964 3241
rect 8998 3207 9059 3241
rect 8759 3145 9059 3207
rect 8759 3111 8820 3145
rect 8854 3111 8892 3145
rect 8926 3111 8964 3145
rect 8998 3111 9059 3145
rect 8759 3049 9059 3111
rect 8759 3015 8820 3049
rect 8854 3015 8892 3049
rect 8926 3015 8964 3049
rect 8998 3015 9059 3049
rect 8759 2953 9059 3015
rect 8759 2919 8820 2953
rect 8854 2919 8892 2953
rect 8926 2919 8964 2953
rect 8998 2919 9059 2953
rect 8759 2857 9059 2919
rect 8759 2823 8820 2857
rect 8854 2823 8892 2857
rect 8926 2823 8964 2857
rect 8998 2823 9059 2857
rect 8759 2761 9059 2823
rect 8759 2727 8820 2761
rect 8854 2727 8892 2761
rect 8926 2727 8964 2761
rect 8998 2727 9059 2761
rect 8759 2665 9059 2727
rect 8759 2631 8820 2665
rect 8854 2631 8892 2665
rect 8926 2631 8964 2665
rect 8998 2631 9059 2665
rect 8759 2569 9059 2631
rect 8759 2535 8820 2569
rect 8854 2535 8892 2569
rect 8926 2535 8964 2569
rect 8998 2535 9059 2569
rect 8759 2473 9059 2535
rect 8759 2439 8820 2473
rect 8854 2439 8892 2473
rect 8926 2439 8964 2473
rect 8998 2439 9059 2473
rect 8759 2377 9059 2439
rect 8759 2343 8820 2377
rect 8854 2343 8892 2377
rect 8926 2343 8964 2377
rect 8998 2343 9059 2377
rect 8759 2281 9059 2343
rect 8759 2247 8820 2281
rect 8854 2247 8892 2281
rect 8926 2247 8964 2281
rect 8998 2247 9059 2281
rect 8759 2185 9059 2247
rect 8759 2151 8820 2185
rect 8854 2151 8892 2185
rect 8926 2151 8964 2185
rect 8998 2151 9059 2185
rect 8759 2089 9059 2151
rect 8759 2055 8820 2089
rect 8854 2055 8892 2089
rect 8926 2055 8964 2089
rect 8998 2055 9059 2089
rect 8759 1993 9059 2055
rect 8759 1959 8820 1993
rect 8854 1959 8892 1993
rect 8926 1959 8964 1993
rect 8998 1959 9059 1993
rect 8759 1897 9059 1959
rect 8759 1888 8820 1897
rect 8854 1888 8892 1897
rect 8926 1888 8964 1897
rect 8998 1888 9059 1897
rect 7935 278 8235 300
tri 8235 278 8377 420 sw
tri 8617 278 8759 420 se
rect 8759 300 8787 1888
rect 9031 300 9059 1888
tri 9171 3416 9185 3430 se
rect 9185 3416 9457 3430
tri 9457 3416 9471 3430 sw
rect 9171 3382 9471 3416
rect 9171 2050 9199 3382
rect 9443 2050 9471 3382
rect 9171 1993 9471 2050
rect 9171 1959 9232 1993
rect 9266 1959 9304 1993
rect 9338 1959 9376 1993
rect 9410 1959 9471 1993
rect 9171 1897 9471 1959
rect 9171 1863 9232 1897
rect 9266 1863 9304 1897
rect 9338 1863 9376 1897
rect 9410 1863 9471 1897
rect 9171 1801 9471 1863
rect 9171 1767 9232 1801
rect 9266 1767 9304 1801
rect 9338 1767 9376 1801
rect 9410 1767 9471 1801
rect 9171 1705 9471 1767
rect 9171 1671 9232 1705
rect 9266 1671 9304 1705
rect 9338 1671 9376 1705
rect 9410 1671 9471 1705
rect 9171 1609 9471 1671
rect 9171 1575 9232 1609
rect 9266 1575 9304 1609
rect 9338 1575 9376 1609
rect 9410 1575 9471 1609
rect 9171 1513 9471 1575
rect 9171 1479 9232 1513
rect 9266 1479 9304 1513
rect 9338 1479 9376 1513
rect 9410 1479 9471 1513
rect 9171 1417 9471 1479
rect 9171 1383 9232 1417
rect 9266 1383 9304 1417
rect 9338 1383 9376 1417
rect 9410 1383 9471 1417
rect 9171 1321 9471 1383
rect 9171 1287 9232 1321
rect 9266 1287 9304 1321
rect 9338 1287 9376 1321
rect 9410 1287 9471 1321
rect 9171 1225 9471 1287
rect 9171 1191 9232 1225
rect 9266 1191 9304 1225
rect 9338 1191 9376 1225
rect 9410 1191 9471 1225
rect 9171 1129 9471 1191
rect 9171 1095 9232 1129
rect 9266 1095 9304 1129
rect 9338 1095 9376 1129
rect 9410 1095 9471 1129
rect 9171 1033 9471 1095
rect 9171 999 9232 1033
rect 9266 999 9304 1033
rect 9338 999 9376 1033
rect 9410 999 9471 1033
rect 9171 937 9471 999
rect 9171 903 9232 937
rect 9266 903 9304 937
rect 9338 903 9376 937
rect 9410 903 9471 937
rect 9171 841 9471 903
rect 9171 807 9232 841
rect 9266 807 9304 841
rect 9338 807 9376 841
rect 9410 807 9471 841
rect 9171 745 9471 807
rect 9171 711 9232 745
rect 9266 711 9304 745
rect 9338 711 9376 745
rect 9410 711 9471 745
rect 9171 649 9471 711
rect 9171 615 9232 649
rect 9266 615 9304 649
rect 9338 615 9376 649
rect 9410 615 9471 649
rect 9171 536 9471 615
tri 9171 476 9231 536 ne
rect 9231 476 9411 536
tri 9411 476 9471 536 nw
tri 9583 3416 9597 3430 se
rect 9597 3416 9869 3430
tri 9869 3416 9883 3430 sw
rect 9583 3337 9883 3416
rect 9583 3303 9644 3337
rect 9678 3303 9716 3337
rect 9750 3303 9788 3337
rect 9822 3303 9883 3337
rect 9583 3241 9883 3303
rect 9583 3207 9644 3241
rect 9678 3207 9716 3241
rect 9750 3207 9788 3241
rect 9822 3207 9883 3241
rect 9583 3145 9883 3207
rect 9583 3111 9644 3145
rect 9678 3111 9716 3145
rect 9750 3111 9788 3145
rect 9822 3111 9883 3145
rect 9583 3049 9883 3111
rect 9583 3015 9644 3049
rect 9678 3015 9716 3049
rect 9750 3015 9788 3049
rect 9822 3015 9883 3049
rect 9583 2953 9883 3015
rect 9583 2919 9644 2953
rect 9678 2919 9716 2953
rect 9750 2919 9788 2953
rect 9822 2919 9883 2953
rect 9583 2857 9883 2919
rect 9583 2823 9644 2857
rect 9678 2823 9716 2857
rect 9750 2823 9788 2857
rect 9822 2823 9883 2857
rect 9583 2761 9883 2823
rect 9583 2727 9644 2761
rect 9678 2727 9716 2761
rect 9750 2727 9788 2761
rect 9822 2727 9883 2761
rect 9583 2665 9883 2727
rect 9583 2631 9644 2665
rect 9678 2631 9716 2665
rect 9750 2631 9788 2665
rect 9822 2631 9883 2665
rect 9583 2569 9883 2631
rect 9583 2535 9644 2569
rect 9678 2535 9716 2569
rect 9750 2535 9788 2569
rect 9822 2535 9883 2569
rect 9583 2473 9883 2535
rect 9583 2439 9644 2473
rect 9678 2439 9716 2473
rect 9750 2439 9788 2473
rect 9822 2439 9883 2473
rect 9583 2377 9883 2439
rect 9583 2343 9644 2377
rect 9678 2343 9716 2377
rect 9750 2343 9788 2377
rect 9822 2343 9883 2377
rect 9583 2281 9883 2343
rect 9583 2247 9644 2281
rect 9678 2247 9716 2281
rect 9750 2247 9788 2281
rect 9822 2247 9883 2281
rect 9583 2185 9883 2247
rect 9583 2151 9644 2185
rect 9678 2151 9716 2185
rect 9750 2151 9788 2185
rect 9822 2151 9883 2185
rect 9583 2089 9883 2151
rect 9583 2055 9644 2089
rect 9678 2055 9716 2089
rect 9750 2055 9788 2089
rect 9822 2055 9883 2089
rect 9583 1993 9883 2055
rect 9583 1959 9644 1993
rect 9678 1959 9716 1993
rect 9750 1959 9788 1993
rect 9822 1959 9883 1993
rect 9583 1897 9883 1959
rect 9583 1888 9644 1897
rect 9678 1888 9716 1897
rect 9750 1888 9788 1897
rect 9822 1888 9883 1897
rect 8759 278 9059 300
tri 9059 278 9201 420 sw
tri 9441 278 9583 420 se
rect 9583 300 9611 1888
rect 9855 300 9883 1888
tri 9995 3416 10009 3430 se
rect 10009 3416 10281 3430
tri 10281 3416 10295 3430 sw
rect 9995 3382 10295 3416
rect 9995 2050 10023 3382
rect 10267 2050 10295 3382
rect 9995 1993 10295 2050
rect 9995 1959 10056 1993
rect 10090 1959 10128 1993
rect 10162 1959 10200 1993
rect 10234 1959 10295 1993
rect 9995 1897 10295 1959
rect 9995 1863 10056 1897
rect 10090 1863 10128 1897
rect 10162 1863 10200 1897
rect 10234 1863 10295 1897
rect 9995 1801 10295 1863
rect 9995 1767 10056 1801
rect 10090 1767 10128 1801
rect 10162 1767 10200 1801
rect 10234 1767 10295 1801
rect 9995 1705 10295 1767
rect 9995 1671 10056 1705
rect 10090 1671 10128 1705
rect 10162 1671 10200 1705
rect 10234 1671 10295 1705
rect 9995 1609 10295 1671
rect 9995 1575 10056 1609
rect 10090 1575 10128 1609
rect 10162 1575 10200 1609
rect 10234 1575 10295 1609
rect 9995 1513 10295 1575
rect 9995 1479 10056 1513
rect 10090 1479 10128 1513
rect 10162 1479 10200 1513
rect 10234 1479 10295 1513
rect 9995 1417 10295 1479
rect 9995 1383 10056 1417
rect 10090 1383 10128 1417
rect 10162 1383 10200 1417
rect 10234 1383 10295 1417
rect 9995 1321 10295 1383
rect 9995 1287 10056 1321
rect 10090 1287 10128 1321
rect 10162 1287 10200 1321
rect 10234 1287 10295 1321
rect 9995 1225 10295 1287
rect 9995 1191 10056 1225
rect 10090 1191 10128 1225
rect 10162 1191 10200 1225
rect 10234 1191 10295 1225
rect 9995 1129 10295 1191
rect 9995 1095 10056 1129
rect 10090 1095 10128 1129
rect 10162 1095 10200 1129
rect 10234 1095 10295 1129
rect 9995 1033 10295 1095
rect 9995 999 10056 1033
rect 10090 999 10128 1033
rect 10162 999 10200 1033
rect 10234 999 10295 1033
rect 9995 937 10295 999
rect 9995 903 10056 937
rect 10090 903 10128 937
rect 10162 903 10200 937
rect 10234 903 10295 937
rect 9995 841 10295 903
rect 9995 807 10056 841
rect 10090 807 10128 841
rect 10162 807 10200 841
rect 10234 807 10295 841
rect 9995 745 10295 807
rect 9995 711 10056 745
rect 10090 711 10128 745
rect 10162 711 10200 745
rect 10234 711 10295 745
rect 9995 649 10295 711
rect 9995 615 10056 649
rect 10090 615 10128 649
rect 10162 615 10200 649
rect 10234 615 10295 649
rect 9995 536 10295 615
tri 9995 476 10055 536 ne
rect 10055 476 10235 536
tri 10235 476 10295 536 nw
tri 10407 3416 10421 3430 se
rect 10421 3416 10693 3430
tri 10693 3416 10707 3430 sw
rect 10407 3337 10707 3416
rect 10407 3303 10468 3337
rect 10502 3303 10540 3337
rect 10574 3303 10612 3337
rect 10646 3303 10707 3337
rect 10407 3241 10707 3303
rect 10407 3207 10468 3241
rect 10502 3207 10540 3241
rect 10574 3207 10612 3241
rect 10646 3207 10707 3241
rect 10407 3145 10707 3207
rect 10407 3111 10468 3145
rect 10502 3111 10540 3145
rect 10574 3111 10612 3145
rect 10646 3111 10707 3145
rect 10407 3049 10707 3111
rect 10407 3015 10468 3049
rect 10502 3015 10540 3049
rect 10574 3015 10612 3049
rect 10646 3015 10707 3049
rect 10407 2953 10707 3015
rect 10407 2919 10468 2953
rect 10502 2919 10540 2953
rect 10574 2919 10612 2953
rect 10646 2919 10707 2953
rect 10407 2857 10707 2919
rect 10407 2823 10468 2857
rect 10502 2823 10540 2857
rect 10574 2823 10612 2857
rect 10646 2823 10707 2857
rect 10407 2761 10707 2823
rect 10407 2727 10468 2761
rect 10502 2727 10540 2761
rect 10574 2727 10612 2761
rect 10646 2727 10707 2761
rect 10407 2665 10707 2727
rect 10407 2631 10468 2665
rect 10502 2631 10540 2665
rect 10574 2631 10612 2665
rect 10646 2631 10707 2665
rect 10407 2569 10707 2631
rect 10407 2535 10468 2569
rect 10502 2535 10540 2569
rect 10574 2535 10612 2569
rect 10646 2535 10707 2569
rect 10407 2473 10707 2535
rect 10407 2439 10468 2473
rect 10502 2439 10540 2473
rect 10574 2439 10612 2473
rect 10646 2439 10707 2473
rect 10407 2377 10707 2439
rect 10407 2343 10468 2377
rect 10502 2343 10540 2377
rect 10574 2343 10612 2377
rect 10646 2343 10707 2377
rect 10407 2281 10707 2343
rect 10407 2247 10468 2281
rect 10502 2247 10540 2281
rect 10574 2247 10612 2281
rect 10646 2247 10707 2281
rect 10407 2185 10707 2247
rect 10407 2151 10468 2185
rect 10502 2151 10540 2185
rect 10574 2151 10612 2185
rect 10646 2151 10707 2185
rect 10407 2089 10707 2151
rect 10407 2055 10468 2089
rect 10502 2055 10540 2089
rect 10574 2055 10612 2089
rect 10646 2055 10707 2089
rect 10407 1993 10707 2055
rect 10407 1959 10468 1993
rect 10502 1959 10540 1993
rect 10574 1959 10612 1993
rect 10646 1959 10707 1993
rect 10407 1897 10707 1959
rect 10407 1888 10468 1897
rect 10502 1888 10540 1897
rect 10574 1888 10612 1897
rect 10646 1888 10707 1897
rect 9583 278 9883 300
tri 9883 278 10025 420 sw
tri 10265 278 10407 420 se
rect 10407 300 10435 1888
rect 10679 300 10707 1888
tri 10819 3416 10833 3430 se
rect 10833 3416 11105 3430
tri 11105 3416 11119 3430 sw
rect 10819 3382 11119 3416
rect 10819 2050 10847 3382
rect 11091 2050 11119 3382
rect 10819 1993 11119 2050
rect 10819 1959 10880 1993
rect 10914 1959 10952 1993
rect 10986 1959 11024 1993
rect 11058 1959 11119 1993
rect 10819 1897 11119 1959
rect 10819 1863 10880 1897
rect 10914 1863 10952 1897
rect 10986 1863 11024 1897
rect 11058 1863 11119 1897
rect 10819 1801 11119 1863
rect 10819 1767 10880 1801
rect 10914 1767 10952 1801
rect 10986 1767 11024 1801
rect 11058 1767 11119 1801
rect 10819 1705 11119 1767
rect 10819 1671 10880 1705
rect 10914 1671 10952 1705
rect 10986 1671 11024 1705
rect 11058 1671 11119 1705
rect 10819 1609 11119 1671
rect 10819 1575 10880 1609
rect 10914 1575 10952 1609
rect 10986 1575 11024 1609
rect 11058 1575 11119 1609
rect 10819 1513 11119 1575
rect 10819 1479 10880 1513
rect 10914 1479 10952 1513
rect 10986 1479 11024 1513
rect 11058 1479 11119 1513
rect 10819 1417 11119 1479
rect 10819 1383 10880 1417
rect 10914 1383 10952 1417
rect 10986 1383 11024 1417
rect 11058 1383 11119 1417
rect 10819 1321 11119 1383
rect 10819 1287 10880 1321
rect 10914 1287 10952 1321
rect 10986 1287 11024 1321
rect 11058 1287 11119 1321
rect 10819 1225 11119 1287
rect 10819 1191 10880 1225
rect 10914 1191 10952 1225
rect 10986 1191 11024 1225
rect 11058 1191 11119 1225
rect 10819 1129 11119 1191
rect 10819 1095 10880 1129
rect 10914 1095 10952 1129
rect 10986 1095 11024 1129
rect 11058 1095 11119 1129
rect 10819 1033 11119 1095
rect 10819 999 10880 1033
rect 10914 999 10952 1033
rect 10986 999 11024 1033
rect 11058 999 11119 1033
rect 10819 937 11119 999
rect 10819 903 10880 937
rect 10914 903 10952 937
rect 10986 903 11024 937
rect 11058 903 11119 937
rect 10819 841 11119 903
rect 10819 807 10880 841
rect 10914 807 10952 841
rect 10986 807 11024 841
rect 11058 807 11119 841
rect 10819 745 11119 807
rect 10819 711 10880 745
rect 10914 711 10952 745
rect 10986 711 11024 745
rect 11058 711 11119 745
rect 10819 649 11119 711
rect 10819 615 10880 649
rect 10914 615 10952 649
rect 10986 615 11024 649
rect 11058 615 11119 649
rect 10819 536 11119 615
rect 11317 3392 11399 3430
rect 11317 3358 11338 3392
rect 11372 3358 11399 3392
rect 11317 3320 11399 3358
rect 11317 3286 11338 3320
rect 11372 3286 11399 3320
rect 11317 3248 11399 3286
rect 11317 3214 11338 3248
rect 11372 3214 11399 3248
rect 11317 3176 11399 3214
rect 11317 3142 11338 3176
rect 11372 3142 11399 3176
rect 11317 3104 11399 3142
rect 11317 3070 11338 3104
rect 11372 3070 11399 3104
rect 11317 3032 11399 3070
rect 11317 2998 11338 3032
rect 11372 2998 11399 3032
rect 11317 2960 11399 2998
rect 11317 2926 11338 2960
rect 11372 2926 11399 2960
rect 11317 2888 11399 2926
rect 11317 2854 11338 2888
rect 11372 2854 11399 2888
rect 11317 2816 11399 2854
rect 11317 2782 11338 2816
rect 11372 2782 11399 2816
rect 11317 2744 11399 2782
rect 11317 2710 11338 2744
rect 11372 2710 11399 2744
rect 11317 2672 11399 2710
rect 11317 2638 11338 2672
rect 11372 2638 11399 2672
rect 11317 2600 11399 2638
rect 11317 2566 11338 2600
rect 11372 2566 11399 2600
rect 11317 2528 11399 2566
rect 11317 2494 11338 2528
rect 11372 2494 11399 2528
rect 11317 2456 11399 2494
rect 11317 2422 11338 2456
rect 11372 2422 11399 2456
rect 11317 2384 11399 2422
rect 11317 2350 11338 2384
rect 11372 2350 11399 2384
rect 11317 2312 11399 2350
rect 11317 2278 11338 2312
rect 11372 2278 11399 2312
rect 11317 2240 11399 2278
rect 11317 2206 11338 2240
rect 11372 2206 11399 2240
rect 11317 2168 11399 2206
rect 11317 2134 11338 2168
rect 11372 2134 11399 2168
rect 11317 2096 11399 2134
rect 11317 2062 11338 2096
rect 11372 2062 11399 2096
rect 11317 2024 11399 2062
rect 11317 1990 11338 2024
rect 11372 1990 11399 2024
rect 11317 1952 11399 1990
rect 11317 1918 11338 1952
rect 11372 1918 11399 1952
rect 11317 1880 11399 1918
rect 11317 1846 11338 1880
rect 11372 1846 11399 1880
rect 11317 1808 11399 1846
rect 11317 1774 11338 1808
rect 11372 1774 11399 1808
rect 11317 1736 11399 1774
rect 11317 1702 11338 1736
rect 11372 1702 11399 1736
rect 11317 1664 11399 1702
rect 11317 1630 11338 1664
rect 11372 1630 11399 1664
rect 11317 1592 11399 1630
rect 11317 1558 11338 1592
rect 11372 1558 11399 1592
rect 11317 1520 11399 1558
rect 11317 1486 11338 1520
rect 11372 1486 11399 1520
rect 11317 1448 11399 1486
rect 11317 1414 11338 1448
rect 11372 1414 11399 1448
rect 11317 1376 11399 1414
rect 11317 1342 11338 1376
rect 11372 1342 11399 1376
rect 11317 1304 11399 1342
rect 11317 1270 11338 1304
rect 11372 1270 11399 1304
rect 11317 1232 11399 1270
rect 11317 1198 11338 1232
rect 11372 1198 11399 1232
rect 11317 1160 11399 1198
rect 11317 1126 11338 1160
rect 11372 1126 11399 1160
rect 11317 1088 11399 1126
rect 11317 1054 11338 1088
rect 11372 1054 11399 1088
rect 11317 1016 11399 1054
rect 11317 982 11338 1016
rect 11372 982 11399 1016
rect 11317 944 11399 982
rect 11317 910 11338 944
rect 11372 910 11399 944
rect 11317 872 11399 910
rect 11317 838 11338 872
rect 11372 838 11399 872
rect 11317 800 11399 838
rect 11317 766 11338 800
rect 11372 766 11399 800
rect 11317 728 11399 766
rect 11317 694 11338 728
rect 11372 694 11399 728
rect 11317 656 11399 694
rect 11317 622 11338 656
rect 11372 622 11399 656
rect 11317 609 11399 622
tri 10819 476 10879 536 ne
rect 10879 476 11059 536
tri 11059 476 11119 536 nw
rect 10407 278 10707 300
tri 10707 278 10849 420 sw
tri 11175 278 11317 420 se
rect 11317 278 11399 506
rect 7147 250 11399 278
rect 7147 -58 7227 250
rect 10671 -58 11399 250
rect 7147 -86 11399 -58
<< via1 >>
rect 7215 3716 7342 3740
rect 7342 3716 7376 3740
rect 7376 3716 7501 3740
rect 7501 3716 7535 3740
rect 7535 3716 7574 3740
rect 7574 3716 7608 3740
rect 7608 3716 7646 3740
rect 7646 3716 7680 3740
rect 7680 3716 7718 3740
rect 7718 3716 7752 3740
rect 7752 3716 7790 3740
rect 7790 3716 7824 3740
rect 7824 3716 7862 3740
rect 7862 3716 7896 3740
rect 7896 3716 7934 3740
rect 7934 3716 7968 3740
rect 7968 3716 8006 3740
rect 8006 3716 8040 3740
rect 8040 3716 8078 3740
rect 8078 3716 8112 3740
rect 8112 3716 8150 3740
rect 8150 3716 8184 3740
rect 8184 3716 8222 3740
rect 8222 3716 8256 3740
rect 8256 3716 8294 3740
rect 8294 3716 8328 3740
rect 8328 3716 8366 3740
rect 8366 3716 8400 3740
rect 8400 3716 8438 3740
rect 8438 3716 8472 3740
rect 8472 3716 8510 3740
rect 8510 3716 8544 3740
rect 8544 3716 8582 3740
rect 8582 3716 8616 3740
rect 8616 3716 8654 3740
rect 8654 3716 8688 3740
rect 8688 3716 8726 3740
rect 8726 3716 8760 3740
rect 8760 3716 8798 3740
rect 8798 3716 8832 3740
rect 8832 3716 8870 3740
rect 8870 3716 8904 3740
rect 8904 3716 8942 3740
rect 8942 3716 8976 3740
rect 8976 3716 9014 3740
rect 9014 3716 9048 3740
rect 9048 3716 9086 3740
rect 9086 3716 9120 3740
rect 9120 3716 9158 3740
rect 9158 3716 9192 3740
rect 9192 3716 9230 3740
rect 9230 3716 9264 3740
rect 9264 3716 9302 3740
rect 9302 3716 9336 3740
rect 9336 3716 9374 3740
rect 9374 3716 9408 3740
rect 9408 3716 9446 3740
rect 9446 3716 9480 3740
rect 9480 3716 9518 3740
rect 9518 3716 9552 3740
rect 9552 3716 9590 3740
rect 9590 3716 9624 3740
rect 9624 3716 9662 3740
rect 9662 3716 9696 3740
rect 9696 3716 9734 3740
rect 9734 3716 9768 3740
rect 9768 3716 9806 3740
rect 9806 3716 9840 3740
rect 9840 3716 9878 3740
rect 9878 3716 9912 3740
rect 9912 3716 9950 3740
rect 9950 3716 9984 3740
rect 9984 3716 10022 3740
rect 10022 3716 10056 3740
rect 10056 3716 10094 3740
rect 10094 3716 10128 3740
rect 10128 3716 10166 3740
rect 10166 3716 10200 3740
rect 10200 3716 10238 3740
rect 10238 3716 10272 3740
rect 10272 3716 10310 3740
rect 10310 3716 10344 3740
rect 10344 3716 10382 3740
rect 10382 3716 10416 3740
rect 10416 3716 10454 3740
rect 10454 3716 10488 3740
rect 10488 3716 10526 3740
rect 10526 3716 10560 3740
rect 10560 3716 10598 3740
rect 10598 3716 10632 3740
rect 10632 3716 10670 3740
rect 10670 3716 10704 3740
rect 10704 3716 10742 3740
rect 10742 3716 10776 3740
rect 10776 3716 10814 3740
rect 10814 3716 10848 3740
rect 10848 3716 10851 3740
rect 7215 3642 10851 3716
rect 7215 3624 7342 3642
rect 7342 3624 7376 3642
rect 7376 3624 7501 3642
rect 7501 3624 7535 3642
rect 7535 3624 7574 3642
rect 7574 3624 7608 3642
rect 7608 3624 7646 3642
rect 7646 3624 7680 3642
rect 7680 3624 7718 3642
rect 7718 3624 7752 3642
rect 7752 3624 7790 3642
rect 7790 3624 7824 3642
rect 7824 3624 7862 3642
rect 7862 3624 7896 3642
rect 7896 3624 7934 3642
rect 7934 3624 7968 3642
rect 7968 3624 8006 3642
rect 8006 3624 8040 3642
rect 8040 3624 8078 3642
rect 8078 3624 8112 3642
rect 8112 3624 8150 3642
rect 8150 3624 8184 3642
rect 8184 3624 8222 3642
rect 8222 3624 8256 3642
rect 8256 3624 8294 3642
rect 8294 3624 8328 3642
rect 8328 3624 8366 3642
rect 8366 3624 8400 3642
rect 8400 3624 8438 3642
rect 8438 3624 8472 3642
rect 8472 3624 8510 3642
rect 8510 3624 8544 3642
rect 8544 3624 8582 3642
rect 8582 3624 8616 3642
rect 8616 3624 8654 3642
rect 8654 3624 8688 3642
rect 8688 3624 8726 3642
rect 8726 3624 8760 3642
rect 8760 3624 8798 3642
rect 8798 3624 8832 3642
rect 8832 3624 8870 3642
rect 8870 3624 8904 3642
rect 8904 3624 8942 3642
rect 8942 3624 8976 3642
rect 8976 3624 9014 3642
rect 9014 3624 9048 3642
rect 9048 3624 9086 3642
rect 9086 3624 9120 3642
rect 9120 3624 9158 3642
rect 9158 3624 9192 3642
rect 9192 3624 9230 3642
rect 9230 3624 9264 3642
rect 9264 3624 9302 3642
rect 9302 3624 9336 3642
rect 9336 3624 9374 3642
rect 9374 3624 9408 3642
rect 9408 3624 9446 3642
rect 9446 3624 9480 3642
rect 9480 3624 9518 3642
rect 9518 3624 9552 3642
rect 9552 3624 9590 3642
rect 9590 3624 9624 3642
rect 9624 3624 9662 3642
rect 9662 3624 9696 3642
rect 9696 3624 9734 3642
rect 9734 3624 9768 3642
rect 9768 3624 9806 3642
rect 9806 3624 9840 3642
rect 9840 3624 9878 3642
rect 9878 3624 9912 3642
rect 9912 3624 9950 3642
rect 9950 3624 9984 3642
rect 9984 3624 10022 3642
rect 10022 3624 10056 3642
rect 10056 3624 10094 3642
rect 10094 3624 10128 3642
rect 10128 3624 10166 3642
rect 10166 3624 10200 3642
rect 10200 3624 10238 3642
rect 10238 3624 10272 3642
rect 10272 3624 10310 3642
rect 10310 3624 10344 3642
rect 10344 3624 10382 3642
rect 10382 3624 10416 3642
rect 10416 3624 10454 3642
rect 10454 3624 10488 3642
rect 10488 3624 10526 3642
rect 10526 3624 10560 3642
rect 10560 3624 10598 3642
rect 10598 3624 10632 3642
rect 10632 3624 10670 3642
rect 10670 3624 10704 3642
rect 10704 3624 10742 3642
rect 10742 3624 10776 3642
rect 10776 3624 10814 3642
rect 10814 3624 10848 3642
rect 10848 3624 10851 3642
rect 7551 3337 7795 3382
rect 7551 3303 7584 3337
rect 7584 3303 7618 3337
rect 7618 3303 7656 3337
rect 7656 3303 7690 3337
rect 7690 3303 7728 3337
rect 7728 3303 7762 3337
rect 7762 3303 7795 3337
rect 7551 3241 7795 3303
rect 7551 3207 7584 3241
rect 7584 3207 7618 3241
rect 7618 3207 7656 3241
rect 7656 3207 7690 3241
rect 7690 3207 7728 3241
rect 7728 3207 7762 3241
rect 7762 3207 7795 3241
rect 7551 3145 7795 3207
rect 7551 3111 7584 3145
rect 7584 3111 7618 3145
rect 7618 3111 7656 3145
rect 7656 3111 7690 3145
rect 7690 3111 7728 3145
rect 7728 3111 7762 3145
rect 7762 3111 7795 3145
rect 7551 3049 7795 3111
rect 7551 3015 7584 3049
rect 7584 3015 7618 3049
rect 7618 3015 7656 3049
rect 7656 3015 7690 3049
rect 7690 3015 7728 3049
rect 7728 3015 7762 3049
rect 7762 3015 7795 3049
rect 7551 2953 7795 3015
rect 7551 2919 7584 2953
rect 7584 2919 7618 2953
rect 7618 2919 7656 2953
rect 7656 2919 7690 2953
rect 7690 2919 7728 2953
rect 7728 2919 7762 2953
rect 7762 2919 7795 2953
rect 7551 2857 7795 2919
rect 7551 2823 7584 2857
rect 7584 2823 7618 2857
rect 7618 2823 7656 2857
rect 7656 2823 7690 2857
rect 7690 2823 7728 2857
rect 7728 2823 7762 2857
rect 7762 2823 7795 2857
rect 7551 2761 7795 2823
rect 7551 2727 7584 2761
rect 7584 2727 7618 2761
rect 7618 2727 7656 2761
rect 7656 2727 7690 2761
rect 7690 2727 7728 2761
rect 7728 2727 7762 2761
rect 7762 2727 7795 2761
rect 7551 2665 7795 2727
rect 7551 2631 7584 2665
rect 7584 2631 7618 2665
rect 7618 2631 7656 2665
rect 7656 2631 7690 2665
rect 7690 2631 7728 2665
rect 7728 2631 7762 2665
rect 7762 2631 7795 2665
rect 7551 2569 7795 2631
rect 7551 2535 7584 2569
rect 7584 2535 7618 2569
rect 7618 2535 7656 2569
rect 7656 2535 7690 2569
rect 7690 2535 7728 2569
rect 7728 2535 7762 2569
rect 7762 2535 7795 2569
rect 7551 2473 7795 2535
rect 7551 2439 7584 2473
rect 7584 2439 7618 2473
rect 7618 2439 7656 2473
rect 7656 2439 7690 2473
rect 7690 2439 7728 2473
rect 7728 2439 7762 2473
rect 7762 2439 7795 2473
rect 7551 2377 7795 2439
rect 7551 2343 7584 2377
rect 7584 2343 7618 2377
rect 7618 2343 7656 2377
rect 7656 2343 7690 2377
rect 7690 2343 7728 2377
rect 7728 2343 7762 2377
rect 7762 2343 7795 2377
rect 7551 2281 7795 2343
rect 7551 2247 7584 2281
rect 7584 2247 7618 2281
rect 7618 2247 7656 2281
rect 7656 2247 7690 2281
rect 7690 2247 7728 2281
rect 7728 2247 7762 2281
rect 7762 2247 7795 2281
rect 7551 2185 7795 2247
rect 7551 2151 7584 2185
rect 7584 2151 7618 2185
rect 7618 2151 7656 2185
rect 7656 2151 7690 2185
rect 7690 2151 7728 2185
rect 7728 2151 7762 2185
rect 7762 2151 7795 2185
rect 7551 2089 7795 2151
rect 7551 2055 7584 2089
rect 7584 2055 7618 2089
rect 7618 2055 7656 2089
rect 7656 2055 7690 2089
rect 7690 2055 7728 2089
rect 7728 2055 7762 2089
rect 7762 2055 7795 2089
rect 7551 2050 7795 2055
rect 7963 1863 7996 1888
rect 7996 1863 8030 1888
rect 8030 1863 8068 1888
rect 8068 1863 8102 1888
rect 8102 1863 8140 1888
rect 8140 1863 8174 1888
rect 8174 1863 8207 1888
rect 7963 1801 8207 1863
rect 7963 1767 7996 1801
rect 7996 1767 8030 1801
rect 8030 1767 8068 1801
rect 8068 1767 8102 1801
rect 8102 1767 8140 1801
rect 8140 1767 8174 1801
rect 8174 1767 8207 1801
rect 7963 1705 8207 1767
rect 7963 1671 7996 1705
rect 7996 1671 8030 1705
rect 8030 1671 8068 1705
rect 8068 1671 8102 1705
rect 8102 1671 8140 1705
rect 8140 1671 8174 1705
rect 8174 1671 8207 1705
rect 7963 1609 8207 1671
rect 7963 1575 7996 1609
rect 7996 1575 8030 1609
rect 8030 1575 8068 1609
rect 8068 1575 8102 1609
rect 8102 1575 8140 1609
rect 8140 1575 8174 1609
rect 8174 1575 8207 1609
rect 7963 1513 8207 1575
rect 7963 1479 7996 1513
rect 7996 1479 8030 1513
rect 8030 1479 8068 1513
rect 8068 1479 8102 1513
rect 8102 1479 8140 1513
rect 8140 1479 8174 1513
rect 8174 1479 8207 1513
rect 7963 1417 8207 1479
rect 7963 1383 7996 1417
rect 7996 1383 8030 1417
rect 8030 1383 8068 1417
rect 8068 1383 8102 1417
rect 8102 1383 8140 1417
rect 8140 1383 8174 1417
rect 8174 1383 8207 1417
rect 7963 1321 8207 1383
rect 7963 1287 7996 1321
rect 7996 1287 8030 1321
rect 8030 1287 8068 1321
rect 8068 1287 8102 1321
rect 8102 1287 8140 1321
rect 8140 1287 8174 1321
rect 8174 1287 8207 1321
rect 7963 1225 8207 1287
rect 7963 1191 7996 1225
rect 7996 1191 8030 1225
rect 8030 1191 8068 1225
rect 8068 1191 8102 1225
rect 8102 1191 8140 1225
rect 8140 1191 8174 1225
rect 8174 1191 8207 1225
rect 7963 1129 8207 1191
rect 7963 1095 7996 1129
rect 7996 1095 8030 1129
rect 8030 1095 8068 1129
rect 8068 1095 8102 1129
rect 8102 1095 8140 1129
rect 8140 1095 8174 1129
rect 8174 1095 8207 1129
rect 7963 1033 8207 1095
rect 7963 999 7996 1033
rect 7996 999 8030 1033
rect 8030 999 8068 1033
rect 8068 999 8102 1033
rect 8102 999 8140 1033
rect 8140 999 8174 1033
rect 8174 999 8207 1033
rect 7963 937 8207 999
rect 7963 903 7996 937
rect 7996 903 8030 937
rect 8030 903 8068 937
rect 8068 903 8102 937
rect 8102 903 8140 937
rect 8140 903 8174 937
rect 8174 903 8207 937
rect 7963 841 8207 903
rect 7963 807 7996 841
rect 7996 807 8030 841
rect 8030 807 8068 841
rect 8068 807 8102 841
rect 8102 807 8140 841
rect 8140 807 8174 841
rect 8174 807 8207 841
rect 7963 745 8207 807
rect 7963 711 7996 745
rect 7996 711 8030 745
rect 8030 711 8068 745
rect 8068 711 8102 745
rect 8102 711 8140 745
rect 8140 711 8174 745
rect 8174 711 8207 745
rect 7963 649 8207 711
rect 7963 615 7996 649
rect 7996 615 8030 649
rect 8030 615 8068 649
rect 8068 615 8102 649
rect 8102 615 8140 649
rect 8140 615 8174 649
rect 8174 615 8207 649
rect 7963 300 8207 615
rect 8375 3337 8619 3382
rect 8375 3303 8408 3337
rect 8408 3303 8442 3337
rect 8442 3303 8480 3337
rect 8480 3303 8514 3337
rect 8514 3303 8552 3337
rect 8552 3303 8586 3337
rect 8586 3303 8619 3337
rect 8375 3241 8619 3303
rect 8375 3207 8408 3241
rect 8408 3207 8442 3241
rect 8442 3207 8480 3241
rect 8480 3207 8514 3241
rect 8514 3207 8552 3241
rect 8552 3207 8586 3241
rect 8586 3207 8619 3241
rect 8375 3145 8619 3207
rect 8375 3111 8408 3145
rect 8408 3111 8442 3145
rect 8442 3111 8480 3145
rect 8480 3111 8514 3145
rect 8514 3111 8552 3145
rect 8552 3111 8586 3145
rect 8586 3111 8619 3145
rect 8375 3049 8619 3111
rect 8375 3015 8408 3049
rect 8408 3015 8442 3049
rect 8442 3015 8480 3049
rect 8480 3015 8514 3049
rect 8514 3015 8552 3049
rect 8552 3015 8586 3049
rect 8586 3015 8619 3049
rect 8375 2953 8619 3015
rect 8375 2919 8408 2953
rect 8408 2919 8442 2953
rect 8442 2919 8480 2953
rect 8480 2919 8514 2953
rect 8514 2919 8552 2953
rect 8552 2919 8586 2953
rect 8586 2919 8619 2953
rect 8375 2857 8619 2919
rect 8375 2823 8408 2857
rect 8408 2823 8442 2857
rect 8442 2823 8480 2857
rect 8480 2823 8514 2857
rect 8514 2823 8552 2857
rect 8552 2823 8586 2857
rect 8586 2823 8619 2857
rect 8375 2761 8619 2823
rect 8375 2727 8408 2761
rect 8408 2727 8442 2761
rect 8442 2727 8480 2761
rect 8480 2727 8514 2761
rect 8514 2727 8552 2761
rect 8552 2727 8586 2761
rect 8586 2727 8619 2761
rect 8375 2665 8619 2727
rect 8375 2631 8408 2665
rect 8408 2631 8442 2665
rect 8442 2631 8480 2665
rect 8480 2631 8514 2665
rect 8514 2631 8552 2665
rect 8552 2631 8586 2665
rect 8586 2631 8619 2665
rect 8375 2569 8619 2631
rect 8375 2535 8408 2569
rect 8408 2535 8442 2569
rect 8442 2535 8480 2569
rect 8480 2535 8514 2569
rect 8514 2535 8552 2569
rect 8552 2535 8586 2569
rect 8586 2535 8619 2569
rect 8375 2473 8619 2535
rect 8375 2439 8408 2473
rect 8408 2439 8442 2473
rect 8442 2439 8480 2473
rect 8480 2439 8514 2473
rect 8514 2439 8552 2473
rect 8552 2439 8586 2473
rect 8586 2439 8619 2473
rect 8375 2377 8619 2439
rect 8375 2343 8408 2377
rect 8408 2343 8442 2377
rect 8442 2343 8480 2377
rect 8480 2343 8514 2377
rect 8514 2343 8552 2377
rect 8552 2343 8586 2377
rect 8586 2343 8619 2377
rect 8375 2281 8619 2343
rect 8375 2247 8408 2281
rect 8408 2247 8442 2281
rect 8442 2247 8480 2281
rect 8480 2247 8514 2281
rect 8514 2247 8552 2281
rect 8552 2247 8586 2281
rect 8586 2247 8619 2281
rect 8375 2185 8619 2247
rect 8375 2151 8408 2185
rect 8408 2151 8442 2185
rect 8442 2151 8480 2185
rect 8480 2151 8514 2185
rect 8514 2151 8552 2185
rect 8552 2151 8586 2185
rect 8586 2151 8619 2185
rect 8375 2089 8619 2151
rect 8375 2055 8408 2089
rect 8408 2055 8442 2089
rect 8442 2055 8480 2089
rect 8480 2055 8514 2089
rect 8514 2055 8552 2089
rect 8552 2055 8586 2089
rect 8586 2055 8619 2089
rect 8375 2050 8619 2055
rect 8787 1863 8820 1888
rect 8820 1863 8854 1888
rect 8854 1863 8892 1888
rect 8892 1863 8926 1888
rect 8926 1863 8964 1888
rect 8964 1863 8998 1888
rect 8998 1863 9031 1888
rect 8787 1801 9031 1863
rect 8787 1767 8820 1801
rect 8820 1767 8854 1801
rect 8854 1767 8892 1801
rect 8892 1767 8926 1801
rect 8926 1767 8964 1801
rect 8964 1767 8998 1801
rect 8998 1767 9031 1801
rect 8787 1705 9031 1767
rect 8787 1671 8820 1705
rect 8820 1671 8854 1705
rect 8854 1671 8892 1705
rect 8892 1671 8926 1705
rect 8926 1671 8964 1705
rect 8964 1671 8998 1705
rect 8998 1671 9031 1705
rect 8787 1609 9031 1671
rect 8787 1575 8820 1609
rect 8820 1575 8854 1609
rect 8854 1575 8892 1609
rect 8892 1575 8926 1609
rect 8926 1575 8964 1609
rect 8964 1575 8998 1609
rect 8998 1575 9031 1609
rect 8787 1513 9031 1575
rect 8787 1479 8820 1513
rect 8820 1479 8854 1513
rect 8854 1479 8892 1513
rect 8892 1479 8926 1513
rect 8926 1479 8964 1513
rect 8964 1479 8998 1513
rect 8998 1479 9031 1513
rect 8787 1417 9031 1479
rect 8787 1383 8820 1417
rect 8820 1383 8854 1417
rect 8854 1383 8892 1417
rect 8892 1383 8926 1417
rect 8926 1383 8964 1417
rect 8964 1383 8998 1417
rect 8998 1383 9031 1417
rect 8787 1321 9031 1383
rect 8787 1287 8820 1321
rect 8820 1287 8854 1321
rect 8854 1287 8892 1321
rect 8892 1287 8926 1321
rect 8926 1287 8964 1321
rect 8964 1287 8998 1321
rect 8998 1287 9031 1321
rect 8787 1225 9031 1287
rect 8787 1191 8820 1225
rect 8820 1191 8854 1225
rect 8854 1191 8892 1225
rect 8892 1191 8926 1225
rect 8926 1191 8964 1225
rect 8964 1191 8998 1225
rect 8998 1191 9031 1225
rect 8787 1129 9031 1191
rect 8787 1095 8820 1129
rect 8820 1095 8854 1129
rect 8854 1095 8892 1129
rect 8892 1095 8926 1129
rect 8926 1095 8964 1129
rect 8964 1095 8998 1129
rect 8998 1095 9031 1129
rect 8787 1033 9031 1095
rect 8787 999 8820 1033
rect 8820 999 8854 1033
rect 8854 999 8892 1033
rect 8892 999 8926 1033
rect 8926 999 8964 1033
rect 8964 999 8998 1033
rect 8998 999 9031 1033
rect 8787 937 9031 999
rect 8787 903 8820 937
rect 8820 903 8854 937
rect 8854 903 8892 937
rect 8892 903 8926 937
rect 8926 903 8964 937
rect 8964 903 8998 937
rect 8998 903 9031 937
rect 8787 841 9031 903
rect 8787 807 8820 841
rect 8820 807 8854 841
rect 8854 807 8892 841
rect 8892 807 8926 841
rect 8926 807 8964 841
rect 8964 807 8998 841
rect 8998 807 9031 841
rect 8787 745 9031 807
rect 8787 711 8820 745
rect 8820 711 8854 745
rect 8854 711 8892 745
rect 8892 711 8926 745
rect 8926 711 8964 745
rect 8964 711 8998 745
rect 8998 711 9031 745
rect 8787 649 9031 711
rect 8787 615 8820 649
rect 8820 615 8854 649
rect 8854 615 8892 649
rect 8892 615 8926 649
rect 8926 615 8964 649
rect 8964 615 8998 649
rect 8998 615 9031 649
rect 8787 300 9031 615
rect 9199 3337 9443 3382
rect 9199 3303 9232 3337
rect 9232 3303 9266 3337
rect 9266 3303 9304 3337
rect 9304 3303 9338 3337
rect 9338 3303 9376 3337
rect 9376 3303 9410 3337
rect 9410 3303 9443 3337
rect 9199 3241 9443 3303
rect 9199 3207 9232 3241
rect 9232 3207 9266 3241
rect 9266 3207 9304 3241
rect 9304 3207 9338 3241
rect 9338 3207 9376 3241
rect 9376 3207 9410 3241
rect 9410 3207 9443 3241
rect 9199 3145 9443 3207
rect 9199 3111 9232 3145
rect 9232 3111 9266 3145
rect 9266 3111 9304 3145
rect 9304 3111 9338 3145
rect 9338 3111 9376 3145
rect 9376 3111 9410 3145
rect 9410 3111 9443 3145
rect 9199 3049 9443 3111
rect 9199 3015 9232 3049
rect 9232 3015 9266 3049
rect 9266 3015 9304 3049
rect 9304 3015 9338 3049
rect 9338 3015 9376 3049
rect 9376 3015 9410 3049
rect 9410 3015 9443 3049
rect 9199 2953 9443 3015
rect 9199 2919 9232 2953
rect 9232 2919 9266 2953
rect 9266 2919 9304 2953
rect 9304 2919 9338 2953
rect 9338 2919 9376 2953
rect 9376 2919 9410 2953
rect 9410 2919 9443 2953
rect 9199 2857 9443 2919
rect 9199 2823 9232 2857
rect 9232 2823 9266 2857
rect 9266 2823 9304 2857
rect 9304 2823 9338 2857
rect 9338 2823 9376 2857
rect 9376 2823 9410 2857
rect 9410 2823 9443 2857
rect 9199 2761 9443 2823
rect 9199 2727 9232 2761
rect 9232 2727 9266 2761
rect 9266 2727 9304 2761
rect 9304 2727 9338 2761
rect 9338 2727 9376 2761
rect 9376 2727 9410 2761
rect 9410 2727 9443 2761
rect 9199 2665 9443 2727
rect 9199 2631 9232 2665
rect 9232 2631 9266 2665
rect 9266 2631 9304 2665
rect 9304 2631 9338 2665
rect 9338 2631 9376 2665
rect 9376 2631 9410 2665
rect 9410 2631 9443 2665
rect 9199 2569 9443 2631
rect 9199 2535 9232 2569
rect 9232 2535 9266 2569
rect 9266 2535 9304 2569
rect 9304 2535 9338 2569
rect 9338 2535 9376 2569
rect 9376 2535 9410 2569
rect 9410 2535 9443 2569
rect 9199 2473 9443 2535
rect 9199 2439 9232 2473
rect 9232 2439 9266 2473
rect 9266 2439 9304 2473
rect 9304 2439 9338 2473
rect 9338 2439 9376 2473
rect 9376 2439 9410 2473
rect 9410 2439 9443 2473
rect 9199 2377 9443 2439
rect 9199 2343 9232 2377
rect 9232 2343 9266 2377
rect 9266 2343 9304 2377
rect 9304 2343 9338 2377
rect 9338 2343 9376 2377
rect 9376 2343 9410 2377
rect 9410 2343 9443 2377
rect 9199 2281 9443 2343
rect 9199 2247 9232 2281
rect 9232 2247 9266 2281
rect 9266 2247 9304 2281
rect 9304 2247 9338 2281
rect 9338 2247 9376 2281
rect 9376 2247 9410 2281
rect 9410 2247 9443 2281
rect 9199 2185 9443 2247
rect 9199 2151 9232 2185
rect 9232 2151 9266 2185
rect 9266 2151 9304 2185
rect 9304 2151 9338 2185
rect 9338 2151 9376 2185
rect 9376 2151 9410 2185
rect 9410 2151 9443 2185
rect 9199 2089 9443 2151
rect 9199 2055 9232 2089
rect 9232 2055 9266 2089
rect 9266 2055 9304 2089
rect 9304 2055 9338 2089
rect 9338 2055 9376 2089
rect 9376 2055 9410 2089
rect 9410 2055 9443 2089
rect 9199 2050 9443 2055
rect 9611 1863 9644 1888
rect 9644 1863 9678 1888
rect 9678 1863 9716 1888
rect 9716 1863 9750 1888
rect 9750 1863 9788 1888
rect 9788 1863 9822 1888
rect 9822 1863 9855 1888
rect 9611 1801 9855 1863
rect 9611 1767 9644 1801
rect 9644 1767 9678 1801
rect 9678 1767 9716 1801
rect 9716 1767 9750 1801
rect 9750 1767 9788 1801
rect 9788 1767 9822 1801
rect 9822 1767 9855 1801
rect 9611 1705 9855 1767
rect 9611 1671 9644 1705
rect 9644 1671 9678 1705
rect 9678 1671 9716 1705
rect 9716 1671 9750 1705
rect 9750 1671 9788 1705
rect 9788 1671 9822 1705
rect 9822 1671 9855 1705
rect 9611 1609 9855 1671
rect 9611 1575 9644 1609
rect 9644 1575 9678 1609
rect 9678 1575 9716 1609
rect 9716 1575 9750 1609
rect 9750 1575 9788 1609
rect 9788 1575 9822 1609
rect 9822 1575 9855 1609
rect 9611 1513 9855 1575
rect 9611 1479 9644 1513
rect 9644 1479 9678 1513
rect 9678 1479 9716 1513
rect 9716 1479 9750 1513
rect 9750 1479 9788 1513
rect 9788 1479 9822 1513
rect 9822 1479 9855 1513
rect 9611 1417 9855 1479
rect 9611 1383 9644 1417
rect 9644 1383 9678 1417
rect 9678 1383 9716 1417
rect 9716 1383 9750 1417
rect 9750 1383 9788 1417
rect 9788 1383 9822 1417
rect 9822 1383 9855 1417
rect 9611 1321 9855 1383
rect 9611 1287 9644 1321
rect 9644 1287 9678 1321
rect 9678 1287 9716 1321
rect 9716 1287 9750 1321
rect 9750 1287 9788 1321
rect 9788 1287 9822 1321
rect 9822 1287 9855 1321
rect 9611 1225 9855 1287
rect 9611 1191 9644 1225
rect 9644 1191 9678 1225
rect 9678 1191 9716 1225
rect 9716 1191 9750 1225
rect 9750 1191 9788 1225
rect 9788 1191 9822 1225
rect 9822 1191 9855 1225
rect 9611 1129 9855 1191
rect 9611 1095 9644 1129
rect 9644 1095 9678 1129
rect 9678 1095 9716 1129
rect 9716 1095 9750 1129
rect 9750 1095 9788 1129
rect 9788 1095 9822 1129
rect 9822 1095 9855 1129
rect 9611 1033 9855 1095
rect 9611 999 9644 1033
rect 9644 999 9678 1033
rect 9678 999 9716 1033
rect 9716 999 9750 1033
rect 9750 999 9788 1033
rect 9788 999 9822 1033
rect 9822 999 9855 1033
rect 9611 937 9855 999
rect 9611 903 9644 937
rect 9644 903 9678 937
rect 9678 903 9716 937
rect 9716 903 9750 937
rect 9750 903 9788 937
rect 9788 903 9822 937
rect 9822 903 9855 937
rect 9611 841 9855 903
rect 9611 807 9644 841
rect 9644 807 9678 841
rect 9678 807 9716 841
rect 9716 807 9750 841
rect 9750 807 9788 841
rect 9788 807 9822 841
rect 9822 807 9855 841
rect 9611 745 9855 807
rect 9611 711 9644 745
rect 9644 711 9678 745
rect 9678 711 9716 745
rect 9716 711 9750 745
rect 9750 711 9788 745
rect 9788 711 9822 745
rect 9822 711 9855 745
rect 9611 649 9855 711
rect 9611 615 9644 649
rect 9644 615 9678 649
rect 9678 615 9716 649
rect 9716 615 9750 649
rect 9750 615 9788 649
rect 9788 615 9822 649
rect 9822 615 9855 649
rect 9611 300 9855 615
rect 10023 3337 10267 3382
rect 10023 3303 10056 3337
rect 10056 3303 10090 3337
rect 10090 3303 10128 3337
rect 10128 3303 10162 3337
rect 10162 3303 10200 3337
rect 10200 3303 10234 3337
rect 10234 3303 10267 3337
rect 10023 3241 10267 3303
rect 10023 3207 10056 3241
rect 10056 3207 10090 3241
rect 10090 3207 10128 3241
rect 10128 3207 10162 3241
rect 10162 3207 10200 3241
rect 10200 3207 10234 3241
rect 10234 3207 10267 3241
rect 10023 3145 10267 3207
rect 10023 3111 10056 3145
rect 10056 3111 10090 3145
rect 10090 3111 10128 3145
rect 10128 3111 10162 3145
rect 10162 3111 10200 3145
rect 10200 3111 10234 3145
rect 10234 3111 10267 3145
rect 10023 3049 10267 3111
rect 10023 3015 10056 3049
rect 10056 3015 10090 3049
rect 10090 3015 10128 3049
rect 10128 3015 10162 3049
rect 10162 3015 10200 3049
rect 10200 3015 10234 3049
rect 10234 3015 10267 3049
rect 10023 2953 10267 3015
rect 10023 2919 10056 2953
rect 10056 2919 10090 2953
rect 10090 2919 10128 2953
rect 10128 2919 10162 2953
rect 10162 2919 10200 2953
rect 10200 2919 10234 2953
rect 10234 2919 10267 2953
rect 10023 2857 10267 2919
rect 10023 2823 10056 2857
rect 10056 2823 10090 2857
rect 10090 2823 10128 2857
rect 10128 2823 10162 2857
rect 10162 2823 10200 2857
rect 10200 2823 10234 2857
rect 10234 2823 10267 2857
rect 10023 2761 10267 2823
rect 10023 2727 10056 2761
rect 10056 2727 10090 2761
rect 10090 2727 10128 2761
rect 10128 2727 10162 2761
rect 10162 2727 10200 2761
rect 10200 2727 10234 2761
rect 10234 2727 10267 2761
rect 10023 2665 10267 2727
rect 10023 2631 10056 2665
rect 10056 2631 10090 2665
rect 10090 2631 10128 2665
rect 10128 2631 10162 2665
rect 10162 2631 10200 2665
rect 10200 2631 10234 2665
rect 10234 2631 10267 2665
rect 10023 2569 10267 2631
rect 10023 2535 10056 2569
rect 10056 2535 10090 2569
rect 10090 2535 10128 2569
rect 10128 2535 10162 2569
rect 10162 2535 10200 2569
rect 10200 2535 10234 2569
rect 10234 2535 10267 2569
rect 10023 2473 10267 2535
rect 10023 2439 10056 2473
rect 10056 2439 10090 2473
rect 10090 2439 10128 2473
rect 10128 2439 10162 2473
rect 10162 2439 10200 2473
rect 10200 2439 10234 2473
rect 10234 2439 10267 2473
rect 10023 2377 10267 2439
rect 10023 2343 10056 2377
rect 10056 2343 10090 2377
rect 10090 2343 10128 2377
rect 10128 2343 10162 2377
rect 10162 2343 10200 2377
rect 10200 2343 10234 2377
rect 10234 2343 10267 2377
rect 10023 2281 10267 2343
rect 10023 2247 10056 2281
rect 10056 2247 10090 2281
rect 10090 2247 10128 2281
rect 10128 2247 10162 2281
rect 10162 2247 10200 2281
rect 10200 2247 10234 2281
rect 10234 2247 10267 2281
rect 10023 2185 10267 2247
rect 10023 2151 10056 2185
rect 10056 2151 10090 2185
rect 10090 2151 10128 2185
rect 10128 2151 10162 2185
rect 10162 2151 10200 2185
rect 10200 2151 10234 2185
rect 10234 2151 10267 2185
rect 10023 2089 10267 2151
rect 10023 2055 10056 2089
rect 10056 2055 10090 2089
rect 10090 2055 10128 2089
rect 10128 2055 10162 2089
rect 10162 2055 10200 2089
rect 10200 2055 10234 2089
rect 10234 2055 10267 2089
rect 10023 2050 10267 2055
rect 10435 1863 10468 1888
rect 10468 1863 10502 1888
rect 10502 1863 10540 1888
rect 10540 1863 10574 1888
rect 10574 1863 10612 1888
rect 10612 1863 10646 1888
rect 10646 1863 10679 1888
rect 10435 1801 10679 1863
rect 10435 1767 10468 1801
rect 10468 1767 10502 1801
rect 10502 1767 10540 1801
rect 10540 1767 10574 1801
rect 10574 1767 10612 1801
rect 10612 1767 10646 1801
rect 10646 1767 10679 1801
rect 10435 1705 10679 1767
rect 10435 1671 10468 1705
rect 10468 1671 10502 1705
rect 10502 1671 10540 1705
rect 10540 1671 10574 1705
rect 10574 1671 10612 1705
rect 10612 1671 10646 1705
rect 10646 1671 10679 1705
rect 10435 1609 10679 1671
rect 10435 1575 10468 1609
rect 10468 1575 10502 1609
rect 10502 1575 10540 1609
rect 10540 1575 10574 1609
rect 10574 1575 10612 1609
rect 10612 1575 10646 1609
rect 10646 1575 10679 1609
rect 10435 1513 10679 1575
rect 10435 1479 10468 1513
rect 10468 1479 10502 1513
rect 10502 1479 10540 1513
rect 10540 1479 10574 1513
rect 10574 1479 10612 1513
rect 10612 1479 10646 1513
rect 10646 1479 10679 1513
rect 10435 1417 10679 1479
rect 10435 1383 10468 1417
rect 10468 1383 10502 1417
rect 10502 1383 10540 1417
rect 10540 1383 10574 1417
rect 10574 1383 10612 1417
rect 10612 1383 10646 1417
rect 10646 1383 10679 1417
rect 10435 1321 10679 1383
rect 10435 1287 10468 1321
rect 10468 1287 10502 1321
rect 10502 1287 10540 1321
rect 10540 1287 10574 1321
rect 10574 1287 10612 1321
rect 10612 1287 10646 1321
rect 10646 1287 10679 1321
rect 10435 1225 10679 1287
rect 10435 1191 10468 1225
rect 10468 1191 10502 1225
rect 10502 1191 10540 1225
rect 10540 1191 10574 1225
rect 10574 1191 10612 1225
rect 10612 1191 10646 1225
rect 10646 1191 10679 1225
rect 10435 1129 10679 1191
rect 10435 1095 10468 1129
rect 10468 1095 10502 1129
rect 10502 1095 10540 1129
rect 10540 1095 10574 1129
rect 10574 1095 10612 1129
rect 10612 1095 10646 1129
rect 10646 1095 10679 1129
rect 10435 1033 10679 1095
rect 10435 999 10468 1033
rect 10468 999 10502 1033
rect 10502 999 10540 1033
rect 10540 999 10574 1033
rect 10574 999 10612 1033
rect 10612 999 10646 1033
rect 10646 999 10679 1033
rect 10435 937 10679 999
rect 10435 903 10468 937
rect 10468 903 10502 937
rect 10502 903 10540 937
rect 10540 903 10574 937
rect 10574 903 10612 937
rect 10612 903 10646 937
rect 10646 903 10679 937
rect 10435 841 10679 903
rect 10435 807 10468 841
rect 10468 807 10502 841
rect 10502 807 10540 841
rect 10540 807 10574 841
rect 10574 807 10612 841
rect 10612 807 10646 841
rect 10646 807 10679 841
rect 10435 745 10679 807
rect 10435 711 10468 745
rect 10468 711 10502 745
rect 10502 711 10540 745
rect 10540 711 10574 745
rect 10574 711 10612 745
rect 10612 711 10646 745
rect 10646 711 10679 745
rect 10435 649 10679 711
rect 10435 615 10468 649
rect 10468 615 10502 649
rect 10502 615 10540 649
rect 10540 615 10574 649
rect 10574 615 10612 649
rect 10612 615 10646 649
rect 10646 615 10679 649
rect 10435 300 10679 615
rect 10847 3337 11091 3382
rect 10847 3303 10880 3337
rect 10880 3303 10914 3337
rect 10914 3303 10952 3337
rect 10952 3303 10986 3337
rect 10986 3303 11024 3337
rect 11024 3303 11058 3337
rect 11058 3303 11091 3337
rect 10847 3241 11091 3303
rect 10847 3207 10880 3241
rect 10880 3207 10914 3241
rect 10914 3207 10952 3241
rect 10952 3207 10986 3241
rect 10986 3207 11024 3241
rect 11024 3207 11058 3241
rect 11058 3207 11091 3241
rect 10847 3145 11091 3207
rect 10847 3111 10880 3145
rect 10880 3111 10914 3145
rect 10914 3111 10952 3145
rect 10952 3111 10986 3145
rect 10986 3111 11024 3145
rect 11024 3111 11058 3145
rect 11058 3111 11091 3145
rect 10847 3049 11091 3111
rect 10847 3015 10880 3049
rect 10880 3015 10914 3049
rect 10914 3015 10952 3049
rect 10952 3015 10986 3049
rect 10986 3015 11024 3049
rect 11024 3015 11058 3049
rect 11058 3015 11091 3049
rect 10847 2953 11091 3015
rect 10847 2919 10880 2953
rect 10880 2919 10914 2953
rect 10914 2919 10952 2953
rect 10952 2919 10986 2953
rect 10986 2919 11024 2953
rect 11024 2919 11058 2953
rect 11058 2919 11091 2953
rect 10847 2857 11091 2919
rect 10847 2823 10880 2857
rect 10880 2823 10914 2857
rect 10914 2823 10952 2857
rect 10952 2823 10986 2857
rect 10986 2823 11024 2857
rect 11024 2823 11058 2857
rect 11058 2823 11091 2857
rect 10847 2761 11091 2823
rect 10847 2727 10880 2761
rect 10880 2727 10914 2761
rect 10914 2727 10952 2761
rect 10952 2727 10986 2761
rect 10986 2727 11024 2761
rect 11024 2727 11058 2761
rect 11058 2727 11091 2761
rect 10847 2665 11091 2727
rect 10847 2631 10880 2665
rect 10880 2631 10914 2665
rect 10914 2631 10952 2665
rect 10952 2631 10986 2665
rect 10986 2631 11024 2665
rect 11024 2631 11058 2665
rect 11058 2631 11091 2665
rect 10847 2569 11091 2631
rect 10847 2535 10880 2569
rect 10880 2535 10914 2569
rect 10914 2535 10952 2569
rect 10952 2535 10986 2569
rect 10986 2535 11024 2569
rect 11024 2535 11058 2569
rect 11058 2535 11091 2569
rect 10847 2473 11091 2535
rect 10847 2439 10880 2473
rect 10880 2439 10914 2473
rect 10914 2439 10952 2473
rect 10952 2439 10986 2473
rect 10986 2439 11024 2473
rect 11024 2439 11058 2473
rect 11058 2439 11091 2473
rect 10847 2377 11091 2439
rect 10847 2343 10880 2377
rect 10880 2343 10914 2377
rect 10914 2343 10952 2377
rect 10952 2343 10986 2377
rect 10986 2343 11024 2377
rect 11024 2343 11058 2377
rect 11058 2343 11091 2377
rect 10847 2281 11091 2343
rect 10847 2247 10880 2281
rect 10880 2247 10914 2281
rect 10914 2247 10952 2281
rect 10952 2247 10986 2281
rect 10986 2247 11024 2281
rect 11024 2247 11058 2281
rect 11058 2247 11091 2281
rect 10847 2185 11091 2247
rect 10847 2151 10880 2185
rect 10880 2151 10914 2185
rect 10914 2151 10952 2185
rect 10952 2151 10986 2185
rect 10986 2151 11024 2185
rect 11024 2151 11058 2185
rect 11058 2151 11091 2185
rect 10847 2089 11091 2151
rect 10847 2055 10880 2089
rect 10880 2055 10914 2089
rect 10914 2055 10952 2089
rect 10952 2055 10986 2089
rect 10986 2055 11024 2089
rect 11024 2055 11058 2089
rect 11058 2055 11091 2089
rect 10847 2050 11091 2055
rect 7227 -58 10671 250
<< metal2 >>
rect 7075 3740 10869 3752
rect 7075 3624 7215 3740
rect 10851 3624 10869 3740
rect 7075 3612 10869 3624
rect 7075 3382 11119 3416
rect 7075 2050 7551 3382
rect 7795 2050 8375 3382
rect 8619 2050 9199 3382
rect 9443 2050 10023 3382
rect 10267 2050 10847 3382
rect 11091 2050 11119 3382
rect 7075 2016 11119 2050
rect 7075 1888 11141 1908
rect 7075 300 7963 1888
rect 8207 300 8787 1888
rect 9031 300 9611 1888
rect 9855 300 10435 1888
rect 10679 300 11141 1888
rect 7075 250 11141 300
rect 7075 -58 7227 250
rect 10671 -58 11141 250
rect 7075 -86 11141 -58
<< properties >>
string GDS_END 4448810
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 4186382
<< end >>
